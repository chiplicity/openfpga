magic
tech EFS8A
magscale 1 2
timestamp 1602530918
<< locali >>
rect 11563 24225 11598 24259
rect 16991 22049 17026 22083
rect 18331 20009 18337 20043
rect 18331 19941 18365 20009
rect 6227 19873 6262 19907
rect 11839 19873 11874 19907
rect 20855 19873 20982 19907
rect 4123 19465 4169 19499
rect 19533 19227 19567 19465
rect 10919 19193 10964 19227
rect 14651 19159 14685 19227
rect 14651 19125 14657 19159
rect 9631 18785 9758 18819
rect 18337 18615 18371 18785
rect 4807 17833 4813 17867
rect 4807 17765 4841 17833
rect 21281 17051 21315 17289
rect 5083 16983 5117 17051
rect 5083 16949 5089 16983
rect 9631 16609 9758 16643
rect 4629 15963 4663 16133
rect 13179 14569 13185 14603
rect 18331 14569 18337 14603
rect 13179 14501 13213 14569
rect 18331 14501 18365 14569
rect 25087 13345 25122 13379
rect 1443 12733 1570 12767
rect 3433 12631 3467 12733
rect 22511 12257 22546 12291
rect 6929 11543 6963 11645
rect 18699 11543 18733 11611
rect 18699 11509 18705 11543
rect 18153 11169 18314 11203
rect 18153 10999 18187 11169
rect 18981 10999 19015 11237
rect 22511 10081 22546 10115
rect 24627 10081 24662 10115
rect 19751 8993 19786 9027
rect 10051 6953 10057 6987
rect 10051 6885 10085 6953
rect 23811 6409 23949 6443
rect 1443 3553 1478 3587
rect 20223 2601 20361 2635
<< viali >>
rect 7481 24361 7515 24395
rect 7297 24225 7331 24259
rect 11529 24225 11563 24259
rect 11667 24021 11701 24055
rect 8033 23817 8067 23851
rect 10793 23817 10827 23851
rect 11621 23817 11655 23851
rect 18337 23817 18371 23851
rect 20729 23817 20763 23851
rect 21741 23817 21775 23851
rect 25237 23817 25271 23851
rect 11253 23749 11287 23783
rect 24823 23749 24857 23783
rect 1869 23681 1903 23715
rect 1476 23613 1510 23647
rect 7849 23613 7883 23647
rect 8401 23613 8435 23647
rect 10609 23613 10643 23647
rect 15996 23613 16030 23647
rect 16083 23613 16117 23647
rect 16497 23613 16531 23647
rect 18153 23613 18187 23647
rect 18705 23613 18739 23647
rect 20244 23613 20278 23647
rect 21240 23613 21274 23647
rect 23740 23613 23774 23647
rect 24752 23613 24786 23647
rect 21327 23545 21361 23579
rect 24225 23545 24259 23579
rect 1547 23477 1581 23511
rect 7389 23477 7423 23511
rect 20315 23477 20349 23511
rect 23811 23477 23845 23511
rect 15669 23205 15703 23239
rect 1476 23137 1510 23171
rect 8620 23137 8654 23171
rect 13645 23137 13679 23171
rect 14105 23137 14139 23171
rect 17084 23137 17118 23171
rect 20980 23137 21014 23171
rect 14289 23069 14323 23103
rect 15577 23069 15611 23103
rect 8723 23001 8757 23035
rect 16129 23001 16163 23035
rect 1547 22933 1581 22967
rect 12725 22933 12759 22967
rect 14657 22933 14691 22967
rect 17187 22933 17221 22967
rect 21051 22933 21085 22967
rect 2237 22729 2271 22763
rect 14105 22729 14139 22763
rect 14473 22729 14507 22763
rect 16405 22729 16439 22763
rect 21005 22729 21039 22763
rect 13277 22593 13311 22627
rect 15485 22593 15519 22627
rect 16773 22593 16807 22627
rect 17095 22593 17129 22627
rect 1444 22525 1478 22559
rect 1869 22525 1903 22559
rect 12725 22525 12759 22559
rect 13185 22525 13219 22559
rect 14289 22525 14323 22559
rect 17008 22525 17042 22559
rect 17417 22525 17451 22559
rect 17785 22525 17819 22559
rect 18096 22525 18130 22559
rect 14933 22457 14967 22491
rect 15301 22457 15335 22491
rect 15577 22457 15611 22491
rect 16129 22457 16163 22491
rect 18521 22457 18555 22491
rect 1547 22389 1581 22423
rect 8585 22389 8619 22423
rect 12265 22389 12299 22423
rect 13737 22389 13771 22423
rect 18199 22389 18233 22423
rect 13461 22185 13495 22219
rect 13737 22117 13771 22151
rect 13829 22117 13863 22151
rect 15577 22117 15611 22151
rect 18429 22117 18463 22151
rect 18521 22117 18555 22151
rect 12668 22049 12702 22083
rect 14381 22049 14415 22083
rect 16957 22049 16991 22083
rect 15485 21981 15519 22015
rect 16129 21981 16163 22015
rect 19073 21981 19107 22015
rect 17095 21913 17129 21947
rect 12771 21845 12805 21879
rect 12173 21641 12207 21675
rect 16957 21641 16991 21675
rect 17417 21641 17451 21675
rect 24777 21641 24811 21675
rect 14473 21505 14507 21539
rect 16037 21505 16071 21539
rect 18613 21505 18647 21539
rect 19533 21505 19567 21539
rect 12633 21437 12667 21471
rect 13093 21437 13127 21471
rect 24593 21437 24627 21471
rect 25145 21437 25179 21471
rect 11897 21369 11931 21403
rect 13369 21369 13403 21403
rect 14565 21369 14599 21403
rect 15117 21369 15151 21403
rect 16129 21369 16163 21403
rect 16681 21369 16715 21403
rect 18429 21369 18463 21403
rect 18705 21369 18739 21403
rect 19257 21369 19291 21403
rect 13737 21301 13771 21335
rect 14197 21301 14231 21335
rect 15393 21301 15427 21335
rect 15761 21301 15795 21335
rect 17877 21301 17911 21335
rect 13277 21097 13311 21131
rect 15117 21097 15151 21131
rect 17003 21097 17037 21131
rect 11529 21029 11563 21063
rect 13737 21029 13771 21063
rect 13829 21029 13863 21063
rect 15485 21029 15519 21063
rect 18521 21029 18555 21063
rect 19073 21029 19107 21063
rect 1476 20961 1510 20995
rect 9724 20961 9758 20995
rect 16932 20961 16966 20995
rect 24660 20961 24694 20995
rect 8309 20893 8343 20927
rect 11437 20893 11471 20927
rect 12081 20893 12115 20927
rect 15393 20893 15427 20927
rect 15669 20893 15703 20927
rect 18429 20893 18463 20927
rect 14289 20825 14323 20859
rect 1547 20757 1581 20791
rect 8861 20757 8895 20791
rect 9827 20757 9861 20791
rect 10333 20757 10367 20791
rect 12633 20757 12667 20791
rect 14657 20757 14691 20791
rect 16405 20757 16439 20791
rect 24731 20757 24765 20791
rect 1593 20553 1627 20587
rect 4077 20553 4111 20587
rect 11437 20553 11471 20587
rect 14749 20553 14783 20587
rect 15393 20553 15427 20587
rect 17785 20553 17819 20587
rect 18797 20553 18831 20587
rect 24685 20553 24719 20587
rect 10149 20485 10183 20519
rect 14105 20485 14139 20519
rect 14473 20485 14507 20519
rect 19993 20485 20027 20519
rect 21557 20485 21591 20519
rect 4445 20417 4479 20451
rect 11805 20417 11839 20451
rect 13185 20417 13219 20451
rect 14933 20417 14967 20451
rect 20453 20417 20487 20451
rect 21005 20417 21039 20451
rect 3893 20349 3927 20383
rect 7700 20349 7734 20383
rect 8125 20349 8159 20383
rect 8585 20349 8619 20383
rect 8677 20349 8711 20383
rect 9229 20349 9263 20383
rect 10241 20349 10275 20383
rect 10793 20349 10827 20383
rect 17141 20349 17175 20383
rect 7803 20281 7837 20315
rect 13547 20281 13581 20315
rect 16497 20281 16531 20315
rect 16589 20281 16623 20315
rect 18337 20281 18371 20315
rect 19165 20281 19199 20315
rect 19441 20281 19475 20315
rect 19533 20281 19567 20315
rect 21097 20281 21131 20315
rect 8953 20213 8987 20247
rect 9689 20213 9723 20247
rect 10333 20213 10367 20247
rect 13001 20213 13035 20247
rect 15761 20213 15795 20247
rect 16313 20213 16347 20247
rect 17417 20213 17451 20247
rect 20729 20213 20763 20247
rect 7757 20009 7791 20043
rect 14197 20009 14231 20043
rect 14473 20009 14507 20043
rect 17003 20009 17037 20043
rect 18337 20009 18371 20043
rect 18889 20009 18923 20043
rect 19349 20009 19383 20043
rect 24777 20009 24811 20043
rect 4813 19941 4847 19975
rect 8033 19941 8067 19975
rect 8125 19941 8159 19975
rect 10378 19941 10412 19975
rect 13598 19941 13632 19975
rect 15485 19941 15519 19975
rect 6193 19873 6227 19907
rect 10057 19873 10091 19907
rect 11805 19873 11839 19907
rect 13277 19873 13311 19907
rect 16932 19873 16966 19907
rect 19752 19873 19786 19907
rect 20821 19873 20855 19907
rect 24593 19873 24627 19907
rect 4721 19805 4755 19839
rect 4997 19805 5031 19839
rect 8677 19805 8711 19839
rect 15393 19805 15427 19839
rect 16037 19805 16071 19839
rect 17969 19805 18003 19839
rect 16497 19737 16531 19771
rect 19855 19737 19889 19771
rect 5641 19669 5675 19703
rect 6331 19669 6365 19703
rect 10977 19669 11011 19703
rect 11345 19669 11379 19703
rect 11943 19669 11977 19703
rect 12449 19669 12483 19703
rect 20269 19669 20303 19703
rect 21051 19669 21085 19703
rect 21373 19669 21407 19703
rect 21833 19669 21867 19703
rect 1593 19465 1627 19499
rect 3893 19465 3927 19499
rect 4169 19465 4203 19499
rect 6285 19465 6319 19499
rect 8309 19465 8343 19499
rect 9781 19465 9815 19499
rect 11529 19465 11563 19499
rect 18981 19465 19015 19499
rect 19257 19465 19291 19499
rect 19533 19465 19567 19499
rect 11897 19397 11931 19431
rect 17141 19397 17175 19431
rect 5089 19329 5123 19363
rect 5365 19329 5399 19363
rect 8585 19329 8619 19363
rect 8861 19329 8895 19363
rect 12541 19329 12575 19363
rect 12817 19329 12851 19363
rect 13461 19329 13495 19363
rect 14289 19329 14323 19363
rect 16405 19329 16439 19363
rect 1409 19261 1443 19295
rect 4052 19261 4086 19295
rect 6653 19261 6687 19295
rect 7205 19261 7239 19295
rect 7481 19261 7515 19295
rect 10609 19261 10643 19295
rect 18061 19261 18095 19295
rect 19625 19329 19659 19363
rect 19901 19329 19935 19363
rect 24593 19329 24627 19363
rect 21649 19261 21683 19295
rect 21833 19261 21867 19295
rect 3525 19193 3559 19227
rect 5181 19193 5215 19227
rect 7665 19193 7699 19227
rect 8677 19193 8711 19227
rect 10885 19193 10919 19227
rect 12265 19193 12299 19227
rect 12633 19193 12667 19227
rect 15577 19193 15611 19227
rect 16129 19193 16163 19227
rect 16221 19193 16255 19227
rect 18382 19193 18416 19227
rect 19533 19193 19567 19227
rect 19993 19193 20027 19227
rect 20545 19193 20579 19227
rect 1961 19125 1995 19159
rect 4629 19125 4663 19159
rect 8033 19125 8067 19159
rect 10149 19125 10183 19159
rect 10425 19125 10459 19159
rect 14197 19125 14231 19159
rect 14657 19125 14691 19159
rect 15209 19125 15243 19159
rect 15853 19125 15887 19159
rect 17417 19125 17451 19159
rect 17785 19125 17819 19159
rect 21005 19125 21039 19159
rect 21465 19125 21499 19159
rect 2973 18921 3007 18955
rect 7021 18921 7055 18955
rect 8585 18921 8619 18955
rect 8953 18921 8987 18955
rect 12449 18921 12483 18955
rect 13369 18921 13403 18955
rect 14151 18921 14185 18955
rect 15117 18921 15151 18955
rect 16681 18921 16715 18955
rect 18613 18921 18647 18955
rect 5733 18853 5767 18887
rect 6285 18853 6319 18887
rect 7665 18853 7699 18887
rect 10701 18853 10735 18887
rect 10977 18853 11011 18887
rect 15485 18853 15519 18887
rect 16037 18853 16071 18887
rect 19441 18853 19475 18887
rect 4604 18785 4638 18819
rect 9597 18785 9631 18819
rect 12357 18785 12391 18819
rect 12909 18785 12943 18819
rect 14080 18785 14114 18819
rect 17233 18785 17267 18819
rect 17693 18785 17727 18819
rect 18337 18785 18371 18819
rect 20913 18785 20947 18819
rect 21373 18785 21407 18819
rect 5641 18717 5675 18751
rect 7573 18717 7607 18751
rect 7849 18717 7883 18751
rect 9827 18717 9861 18751
rect 10333 18717 10367 18751
rect 10885 18717 10919 18751
rect 11161 18717 11195 18751
rect 15393 18717 15427 18751
rect 17877 18717 17911 18751
rect 4675 18649 4709 18683
rect 5365 18649 5399 18683
rect 7389 18649 7423 18683
rect 19349 18717 19383 18751
rect 19993 18717 20027 18751
rect 21465 18717 21499 18751
rect 5089 18581 5123 18615
rect 14565 18581 14599 18615
rect 16405 18581 16439 18615
rect 18153 18581 18187 18615
rect 18337 18581 18371 18615
rect 6193 18377 6227 18411
rect 8309 18377 8343 18411
rect 9781 18377 9815 18411
rect 10517 18377 10551 18411
rect 16865 18377 16899 18411
rect 18981 18377 19015 18411
rect 19717 18377 19751 18411
rect 20913 18377 20947 18411
rect 24777 18377 24811 18411
rect 10149 18309 10183 18343
rect 20545 18309 20579 18343
rect 4353 18241 4387 18275
rect 5273 18241 5307 18275
rect 5549 18241 5583 18275
rect 7389 18241 7423 18275
rect 7849 18241 7883 18275
rect 8861 18241 8895 18275
rect 10701 18241 10735 18275
rect 11345 18241 11379 18275
rect 14933 18241 14967 18275
rect 15853 18241 15887 18275
rect 16497 18241 16531 18275
rect 18061 18241 18095 18275
rect 3525 18173 3559 18207
rect 4261 18173 4295 18207
rect 12265 18173 12299 18207
rect 12725 18173 12759 18207
rect 13001 18173 13035 18207
rect 14197 18173 14231 18207
rect 14749 18173 14783 18207
rect 24593 18173 24627 18207
rect 25145 18173 25179 18207
rect 5089 18105 5123 18139
rect 5365 18105 5399 18139
rect 7205 18105 7239 18139
rect 7481 18105 7515 18139
rect 8769 18105 8803 18139
rect 9223 18105 9257 18139
rect 10793 18105 10827 18139
rect 15669 18105 15703 18139
rect 15945 18105 15979 18139
rect 18382 18105 18416 18139
rect 19993 18105 20027 18139
rect 20085 18105 20119 18139
rect 4721 18037 4755 18071
rect 11805 18037 11839 18071
rect 12541 18037 12575 18071
rect 13645 18037 13679 18071
rect 14105 18037 14139 18071
rect 15301 18037 15335 18071
rect 17233 18037 17267 18071
rect 17785 18037 17819 18071
rect 19257 18037 19291 18071
rect 21281 18037 21315 18071
rect 4813 17833 4847 17867
rect 5733 17833 5767 17867
rect 10701 17833 10735 17867
rect 11345 17833 11379 17867
rect 15025 17833 15059 17867
rect 16221 17833 16255 17867
rect 18061 17833 18095 17867
rect 19257 17833 19291 17867
rect 6193 17765 6227 17799
rect 8217 17765 8251 17799
rect 9873 17765 9907 17799
rect 11758 17765 11792 17799
rect 15622 17765 15656 17799
rect 18658 17765 18692 17799
rect 20545 17765 20579 17799
rect 21005 17765 21039 17799
rect 21097 17765 21131 17799
rect 6285 17697 6319 17731
rect 11437 17697 11471 17731
rect 13645 17697 13679 17731
rect 14197 17697 14231 17731
rect 4445 17629 4479 17663
rect 7481 17629 7515 17663
rect 8125 17629 8159 17663
rect 8401 17629 8435 17663
rect 9781 17629 9815 17663
rect 10057 17629 10091 17663
rect 14381 17629 14415 17663
rect 15301 17629 15335 17663
rect 18337 17629 18371 17663
rect 21281 17629 21315 17663
rect 5365 17561 5399 17595
rect 12357 17493 12391 17527
rect 12725 17493 12759 17527
rect 13093 17493 13127 17527
rect 19533 17493 19567 17527
rect 19993 17493 20027 17527
rect 2835 17289 2869 17323
rect 5641 17289 5675 17323
rect 6193 17289 6227 17323
rect 9137 17289 9171 17323
rect 10609 17289 10643 17323
rect 11805 17289 11839 17323
rect 12265 17289 12299 17323
rect 14565 17289 14599 17323
rect 15669 17289 15703 17323
rect 21281 17289 21315 17323
rect 21465 17289 21499 17323
rect 23811 17289 23845 17323
rect 8861 17221 8895 17255
rect 9597 17221 9631 17255
rect 9873 17221 9907 17255
rect 16405 17221 16439 17255
rect 7941 17153 7975 17187
rect 10885 17153 10919 17187
rect 11161 17153 11195 17187
rect 12817 17153 12851 17187
rect 14105 17153 14139 17187
rect 20821 17153 20855 17187
rect 2764 17085 2798 17119
rect 3709 17085 3743 17119
rect 4721 17085 4755 17119
rect 6904 17085 6938 17119
rect 9689 17085 9723 17119
rect 10149 17085 10183 17119
rect 14749 17085 14783 17119
rect 16497 17085 16531 17119
rect 16957 17085 16991 17119
rect 18705 17085 18739 17119
rect 22569 17153 22603 17187
rect 22017 17085 22051 17119
rect 22477 17085 22511 17119
rect 23740 17085 23774 17119
rect 24133 17085 24167 17119
rect 3617 17017 3651 17051
rect 7849 17017 7883 17051
rect 8303 17017 8337 17051
rect 10977 17017 11011 17051
rect 12541 17017 12575 17051
rect 12633 17017 12667 17051
rect 15070 17017 15104 17051
rect 15945 17017 15979 17051
rect 19026 17017 19060 17051
rect 20545 17017 20579 17051
rect 20637 17017 20671 17051
rect 21281 17017 21315 17051
rect 21833 17017 21867 17051
rect 3249 16949 3283 16983
rect 4537 16949 4571 16983
rect 5089 16949 5123 16983
rect 6975 16949 7009 16983
rect 7389 16949 7423 16983
rect 13645 16949 13679 16983
rect 16681 16949 16715 16983
rect 17509 16949 17543 16983
rect 17785 16949 17819 16983
rect 18521 16949 18555 16983
rect 19625 16949 19659 16983
rect 20269 16949 20303 16983
rect 4813 16745 4847 16779
rect 8217 16745 8251 16779
rect 10517 16745 10551 16779
rect 12449 16745 12483 16779
rect 14749 16745 14783 16779
rect 16221 16745 16255 16779
rect 16497 16745 16531 16779
rect 18981 16745 19015 16779
rect 19349 16745 19383 16779
rect 21005 16745 21039 16779
rect 22017 16745 22051 16779
rect 5181 16677 5215 16711
rect 8585 16677 8619 16711
rect 11523 16677 11557 16711
rect 15622 16677 15656 16711
rect 18382 16677 18416 16711
rect 20729 16677 20763 16711
rect 1752 16609 1786 16643
rect 7297 16609 7331 16643
rect 9597 16609 9631 16643
rect 10885 16609 10919 16643
rect 12081 16609 12115 16643
rect 12909 16609 12943 16643
rect 13369 16609 13403 16643
rect 15301 16609 15335 16643
rect 19876 16609 19910 16643
rect 21097 16609 21131 16643
rect 21465 16609 21499 16643
rect 22477 16609 22511 16643
rect 22937 16609 22971 16643
rect 2973 16541 3007 16575
rect 5089 16541 5123 16575
rect 5549 16541 5583 16575
rect 11161 16541 11195 16575
rect 13461 16541 13495 16575
rect 18061 16541 18095 16575
rect 23029 16541 23063 16575
rect 1823 16405 1857 16439
rect 4445 16405 4479 16439
rect 7481 16405 7515 16439
rect 9827 16405 9861 16439
rect 13921 16405 13955 16439
rect 16957 16405 16991 16439
rect 19625 16405 19659 16439
rect 19947 16405 19981 16439
rect 2053 16201 2087 16235
rect 4445 16201 4479 16235
rect 4813 16201 4847 16235
rect 7113 16201 7147 16235
rect 7481 16201 7515 16235
rect 10241 16201 10275 16235
rect 11805 16201 11839 16235
rect 12633 16201 12667 16235
rect 15025 16201 15059 16235
rect 15945 16201 15979 16235
rect 17509 16201 17543 16235
rect 18981 16201 19015 16235
rect 20177 16201 20211 16235
rect 21373 16201 21407 16235
rect 22661 16201 22695 16235
rect 23029 16201 23063 16235
rect 4629 16133 4663 16167
rect 5549 16133 5583 16167
rect 9873 16133 9907 16167
rect 11437 16133 11471 16167
rect 19809 16133 19843 16167
rect 4077 16065 4111 16099
rect 1409 15997 1443 16031
rect 3249 15997 3283 16031
rect 3985 15997 4019 16031
rect 4997 16065 5031 16099
rect 5917 16065 5951 16099
rect 7757 16065 7791 16099
rect 9321 16065 9355 16099
rect 10885 16065 10919 16099
rect 12265 16065 12299 16099
rect 17141 16065 17175 16099
rect 18291 16065 18325 16099
rect 19257 16065 19291 16099
rect 21741 16065 21775 16099
rect 12449 15997 12483 16031
rect 12909 15997 12943 16031
rect 15152 15997 15186 16031
rect 15577 15997 15611 16031
rect 16405 15997 16439 16031
rect 16957 15997 16991 16031
rect 18204 15997 18238 16031
rect 18613 15997 18647 16031
rect 4629 15929 4663 15963
rect 5089 15929 5123 15963
rect 7849 15929 7883 15963
rect 8401 15929 8435 15963
rect 9413 15929 9447 15963
rect 10977 15929 11011 15963
rect 13277 15929 13311 15963
rect 13645 15929 13679 15963
rect 13737 15929 13771 15963
rect 14289 15929 14323 15963
rect 19349 15929 19383 15963
rect 21833 15929 21867 15963
rect 22385 15929 22419 15963
rect 1593 15861 1627 15895
rect 9137 15861 9171 15895
rect 10701 15861 10735 15895
rect 14565 15861 14599 15895
rect 15255 15861 15289 15895
rect 17785 15861 17819 15895
rect 21005 15861 21039 15895
rect 1593 15657 1627 15691
rect 5273 15657 5307 15691
rect 7297 15657 7331 15691
rect 9229 15657 9263 15691
rect 11253 15657 11287 15691
rect 17693 15657 17727 15691
rect 21925 15657 21959 15691
rect 22293 15657 22327 15691
rect 4445 15589 4479 15623
rect 4997 15589 5031 15623
rect 6377 15589 6411 15623
rect 7941 15589 7975 15623
rect 8493 15589 8527 15623
rect 10149 15589 10183 15623
rect 10241 15589 10275 15623
rect 11529 15589 11563 15623
rect 13185 15589 13219 15623
rect 16174 15589 16208 15623
rect 19441 15589 19475 15623
rect 21097 15589 21131 15623
rect 22569 15589 22603 15623
rect 22661 15589 22695 15623
rect 2973 15521 3007 15555
rect 12024 15521 12058 15555
rect 15853 15521 15887 15555
rect 16773 15521 16807 15555
rect 17877 15521 17911 15555
rect 18153 15521 18187 15555
rect 24593 15521 24627 15555
rect 4353 15453 4387 15487
rect 6285 15453 6319 15487
rect 6929 15453 6963 15487
rect 7849 15453 7883 15487
rect 10425 15453 10459 15487
rect 12127 15453 12161 15487
rect 13093 15453 13127 15487
rect 13369 15453 13403 15487
rect 18797 15453 18831 15487
rect 19349 15453 19383 15487
rect 21005 15453 21039 15487
rect 21281 15453 21315 15487
rect 22845 15453 22879 15487
rect 19901 15385 19935 15419
rect 24777 15385 24811 15419
rect 3157 15317 3191 15351
rect 3801 15317 3835 15351
rect 6009 15317 6043 15351
rect 7573 15317 7607 15351
rect 14013 15317 14047 15351
rect 15669 15317 15703 15351
rect 19073 15317 19107 15351
rect 5549 15113 5583 15147
rect 7849 15113 7883 15147
rect 8125 15113 8159 15147
rect 10793 15113 10827 15147
rect 11989 15113 12023 15147
rect 14565 15113 14599 15147
rect 14933 15113 14967 15147
rect 15255 15113 15289 15147
rect 15945 15113 15979 15147
rect 17233 15113 17267 15147
rect 17693 15113 17727 15147
rect 18199 15113 18233 15147
rect 22845 15113 22879 15147
rect 5273 15045 5307 15079
rect 8493 15045 8527 15079
rect 14197 15045 14231 15079
rect 19993 15045 20027 15079
rect 20453 15045 20487 15079
rect 20821 15045 20855 15079
rect 21925 15045 21959 15079
rect 6929 14977 6963 15011
rect 10149 14977 10183 15011
rect 13093 14977 13127 15011
rect 13369 14977 13403 15011
rect 13645 14977 13679 15011
rect 16221 14977 16255 15011
rect 16865 14977 16899 15011
rect 22569 14977 22603 15011
rect 24685 14977 24719 15011
rect 3376 14909 3410 14943
rect 3801 14909 3835 14943
rect 4353 14909 4387 14943
rect 10977 14909 11011 14943
rect 11437 14909 11471 14943
rect 15152 14909 15186 14943
rect 15577 14909 15611 14943
rect 18128 14909 18162 14943
rect 18521 14909 18555 14943
rect 19073 14909 19107 14943
rect 23673 14909 23707 14943
rect 24133 14909 24167 14943
rect 4261 14841 4295 14875
rect 4715 14841 4749 14875
rect 6653 14841 6687 14875
rect 7291 14841 7325 14875
rect 9505 14841 9539 14875
rect 9597 14841 9631 14875
rect 13737 14841 13771 14875
rect 16313 14841 16347 14875
rect 19394 14841 19428 14875
rect 21373 14841 21407 14875
rect 21465 14841 21499 14875
rect 23489 14841 23523 14875
rect 1593 14773 1627 14807
rect 2973 14773 3007 14807
rect 3479 14773 3513 14807
rect 6193 14773 6227 14807
rect 9321 14773 9355 14807
rect 10517 14773 10551 14807
rect 11161 14773 11195 14807
rect 12541 14773 12575 14807
rect 18889 14773 18923 14807
rect 21097 14773 21131 14807
rect 23765 14773 23799 14807
rect 1593 14569 1627 14603
rect 3111 14569 3145 14603
rect 3525 14569 3559 14603
rect 6653 14569 6687 14603
rect 8447 14569 8481 14603
rect 9505 14569 9539 14603
rect 13185 14569 13219 14603
rect 13737 14569 13771 14603
rect 16221 14569 16255 14603
rect 18337 14569 18371 14603
rect 18889 14569 18923 14603
rect 19947 14569 19981 14603
rect 20729 14569 20763 14603
rect 22569 14569 22603 14603
rect 23765 14569 23799 14603
rect 4353 14501 4387 14535
rect 4445 14501 4479 14535
rect 4997 14501 5031 14535
rect 6837 14501 6871 14535
rect 6929 14501 6963 14535
rect 7481 14501 7515 14535
rect 10517 14501 10551 14535
rect 16589 14501 16623 14535
rect 19533 14501 19567 14535
rect 21097 14501 21131 14535
rect 1409 14433 1443 14467
rect 3040 14433 3074 14467
rect 8344 14433 8378 14467
rect 15301 14433 15335 14467
rect 19876 14433 19910 14467
rect 22477 14433 22511 14467
rect 22937 14433 22971 14467
rect 24108 14433 24142 14467
rect 10425 14365 10459 14399
rect 12817 14365 12851 14399
rect 16497 14365 16531 14399
rect 17969 14365 18003 14399
rect 21005 14365 21039 14399
rect 21281 14365 21315 14399
rect 10977 14297 11011 14331
rect 17049 14297 17083 14331
rect 2053 14229 2087 14263
rect 3893 14229 3927 14263
rect 6285 14229 6319 14263
rect 9873 14229 9907 14263
rect 12541 14229 12575 14263
rect 14289 14229 14323 14263
rect 15485 14229 15519 14263
rect 15853 14229 15887 14263
rect 19165 14229 19199 14263
rect 22109 14229 22143 14263
rect 24179 14229 24213 14263
rect 1547 14025 1581 14059
rect 4813 14025 4847 14059
rect 5089 14025 5123 14059
rect 7757 14025 7791 14059
rect 8309 14025 8343 14059
rect 8907 14025 8941 14059
rect 11345 14025 11379 14059
rect 12173 14025 12207 14059
rect 14013 14025 14047 14059
rect 15853 14025 15887 14059
rect 16865 14025 16899 14059
rect 19993 14025 20027 14059
rect 21465 14025 21499 14059
rect 23397 14025 23431 14059
rect 25421 14025 25455 14059
rect 1961 13957 1995 13991
rect 6653 13957 6687 13991
rect 9597 13957 9631 13991
rect 10701 13957 10735 13991
rect 10977 13957 11011 13991
rect 13369 13957 13403 13991
rect 23029 13957 23063 13991
rect 2237 13889 2271 13923
rect 6837 13889 6871 13923
rect 14289 13889 14323 13923
rect 14565 13889 14599 13923
rect 15945 13889 15979 13923
rect 24225 13889 24259 13923
rect 1444 13821 1478 13855
rect 2789 13821 2823 13855
rect 2881 13821 2915 13855
rect 3893 13821 3927 13855
rect 5733 13821 5767 13855
rect 6193 13821 6227 13855
rect 8836 13821 8870 13855
rect 9229 13821 9263 13855
rect 9777 13821 9811 13855
rect 12449 13821 12483 13855
rect 18705 13821 18739 13855
rect 22753 13821 22787 13855
rect 23673 13821 23707 13855
rect 24133 13821 24167 13855
rect 25237 13821 25271 13855
rect 25789 13821 25823 13855
rect 4255 13753 4289 13787
rect 7158 13753 7192 13787
rect 10143 13753 10177 13787
rect 12770 13753 12804 13787
rect 14381 13753 14415 13787
rect 16266 13753 16300 13787
rect 17509 13753 17543 13787
rect 19026 13753 19060 13787
rect 20545 13753 20579 13787
rect 20637 13753 20671 13787
rect 21189 13753 21223 13787
rect 22109 13753 22143 13787
rect 22201 13753 22235 13787
rect 24685 13753 24719 13787
rect 3065 13685 3099 13719
rect 3433 13685 3467 13719
rect 3801 13685 3835 13719
rect 5457 13685 5491 13719
rect 5917 13685 5951 13719
rect 13645 13685 13679 13719
rect 15393 13685 15427 13719
rect 17785 13685 17819 13719
rect 18245 13685 18279 13719
rect 19625 13685 19659 13719
rect 20269 13685 20303 13719
rect 21833 13685 21867 13719
rect 3433 13481 3467 13515
rect 5089 13481 5123 13515
rect 6101 13481 6135 13515
rect 12817 13481 12851 13515
rect 14289 13481 14323 13515
rect 15393 13481 15427 13515
rect 16681 13481 16715 13515
rect 17325 13481 17359 13515
rect 19165 13481 19199 13515
rect 20361 13481 20395 13515
rect 20913 13481 20947 13515
rect 22937 13481 22971 13515
rect 4813 13413 4847 13447
rect 6193 13413 6227 13447
rect 10051 13413 10085 13447
rect 12173 13413 12207 13447
rect 12449 13413 12483 13447
rect 13414 13413 13448 13447
rect 18566 13413 18600 13447
rect 22109 13413 22143 13447
rect 22661 13413 22695 13447
rect 1476 13345 1510 13379
rect 2513 13345 2547 13379
rect 4721 13345 4755 13379
rect 6469 13345 6503 13379
rect 8309 13345 8343 13379
rect 8585 13345 8619 13379
rect 11437 13345 11471 13379
rect 11897 13345 11931 13379
rect 15301 13345 15335 13379
rect 15853 13345 15887 13379
rect 16932 13345 16966 13379
rect 23489 13345 23523 13379
rect 23949 13345 23983 13379
rect 24501 13345 24535 13379
rect 25053 13345 25087 13379
rect 8769 13277 8803 13311
rect 9689 13277 9723 13311
rect 13093 13277 13127 13311
rect 18245 13277 18279 13311
rect 22017 13277 22051 13311
rect 24041 13277 24075 13311
rect 1547 13209 1581 13243
rect 17003 13209 17037 13243
rect 20729 13209 20763 13243
rect 1869 13141 1903 13175
rect 2237 13141 2271 13175
rect 2697 13141 2731 13175
rect 3893 13141 3927 13175
rect 7481 13141 7515 13175
rect 10609 13141 10643 13175
rect 14013 13141 14047 13175
rect 16313 13141 16347 13175
rect 18153 13141 18187 13175
rect 19993 13141 20027 13175
rect 21557 13141 21591 13175
rect 25191 13141 25225 13175
rect 1639 12937 1673 12971
rect 2145 12937 2179 12971
rect 2421 12937 2455 12971
rect 8861 12937 8895 12971
rect 9321 12937 9355 12971
rect 9689 12937 9723 12971
rect 10793 12937 10827 12971
rect 12265 12937 12299 12971
rect 13645 12937 13679 12971
rect 14013 12937 14047 12971
rect 15301 12937 15335 12971
rect 16865 12937 16899 12971
rect 22477 12937 22511 12971
rect 23857 12937 23891 12971
rect 24225 12937 24259 12971
rect 25145 12937 25179 12971
rect 2697 12869 2731 12903
rect 6561 12869 6595 12903
rect 7481 12869 7515 12903
rect 10425 12869 10459 12903
rect 17785 12869 17819 12903
rect 19073 12869 19107 12903
rect 20545 12869 20579 12903
rect 24777 12869 24811 12903
rect 3341 12801 3375 12835
rect 8125 12801 8159 12835
rect 9873 12801 9907 12835
rect 11483 12801 11517 12835
rect 14289 12801 14323 12835
rect 18613 12801 18647 12835
rect 21833 12801 21867 12835
rect 1409 12733 1443 12767
rect 2605 12733 2639 12767
rect 2881 12733 2915 12767
rect 3433 12733 3467 12767
rect 4169 12733 4203 12767
rect 4629 12733 4663 12767
rect 5181 12733 5215 12767
rect 5365 12733 5399 12767
rect 7389 12733 7423 12767
rect 7665 12733 7699 12767
rect 11380 12733 11414 12767
rect 12449 12733 12483 12767
rect 15761 12733 15795 12767
rect 16313 12733 16347 12767
rect 18061 12733 18095 12767
rect 18521 12733 18555 12767
rect 24593 12733 24627 12767
rect 3985 12665 4019 12699
rect 9965 12665 9999 12699
rect 11805 12665 11839 12699
rect 12770 12665 12804 12699
rect 14381 12665 14415 12699
rect 14933 12665 14967 12699
rect 17509 12665 17543 12699
rect 19993 12665 20027 12699
rect 20085 12665 20119 12699
rect 21557 12665 21591 12699
rect 21649 12665 21683 12699
rect 3433 12597 3467 12631
rect 3709 12597 3743 12631
rect 4261 12597 4295 12631
rect 6009 12597 6043 12631
rect 7205 12597 7239 12631
rect 8493 12597 8527 12631
rect 11253 12597 11287 12631
rect 13369 12597 13403 12631
rect 15853 12597 15887 12631
rect 19809 12597 19843 12631
rect 21281 12597 21315 12631
rect 1593 12393 1627 12427
rect 1961 12393 1995 12427
rect 3801 12393 3835 12427
rect 4629 12393 4663 12427
rect 6469 12393 6503 12427
rect 6837 12393 6871 12427
rect 9505 12393 9539 12427
rect 9781 12393 9815 12427
rect 11529 12393 11563 12427
rect 17049 12393 17083 12427
rect 18337 12393 18371 12427
rect 20637 12393 20671 12427
rect 23627 12393 23661 12427
rect 24685 12393 24719 12427
rect 3525 12325 3559 12359
rect 7205 12325 7239 12359
rect 8125 12325 8159 12359
rect 12541 12325 12575 12359
rect 13093 12325 13127 12359
rect 13553 12325 13587 12359
rect 14105 12325 14139 12359
rect 19441 12325 19475 12359
rect 19993 12325 20027 12359
rect 21005 12325 21039 12359
rect 21097 12325 21131 12359
rect 1409 12257 1443 12291
rect 2421 12257 2455 12291
rect 2697 12257 2731 12291
rect 4353 12257 4387 12291
rect 4813 12257 4847 12291
rect 5365 12257 5399 12291
rect 5733 12257 5767 12291
rect 7389 12257 7423 12291
rect 7481 12257 7515 12291
rect 7665 12257 7699 12291
rect 9965 12257 9999 12291
rect 10241 12257 10275 12291
rect 11897 12257 11931 12291
rect 12357 12257 12391 12291
rect 15577 12257 15611 12291
rect 16037 12257 16071 12291
rect 17233 12257 17267 12291
rect 17693 12257 17727 12291
rect 22477 12257 22511 12291
rect 23556 12257 23590 12291
rect 2329 12189 2363 12223
rect 2513 12189 2547 12223
rect 3157 12189 3191 12223
rect 6101 12189 6135 12223
rect 13461 12189 13495 12223
rect 16129 12189 16163 12223
rect 16681 12189 16715 12223
rect 17969 12189 18003 12223
rect 18705 12189 18739 12223
rect 19349 12189 19383 12223
rect 21281 12189 21315 12223
rect 22615 12121 22649 12155
rect 10701 12053 10735 12087
rect 21925 12053 21959 12087
rect 2881 11849 2915 11883
rect 5825 11849 5859 11883
rect 8585 11849 8619 11883
rect 9045 11849 9079 11883
rect 9321 11849 9355 11883
rect 12265 11849 12299 11883
rect 14473 11849 14507 11883
rect 15209 11849 15243 11883
rect 22753 11849 22787 11883
rect 23857 11849 23891 11883
rect 3893 11781 3927 11815
rect 7021 11781 7055 11815
rect 11345 11781 11379 11815
rect 17233 11781 17267 11815
rect 21189 11781 21223 11815
rect 1685 11713 1719 11747
rect 7297 11713 7331 11747
rect 7941 11713 7975 11747
rect 8309 11713 8343 11747
rect 10701 11713 10735 11747
rect 13553 11713 13587 11747
rect 16037 11713 16071 11747
rect 18337 11713 18371 11747
rect 20269 11713 20303 11747
rect 20913 11713 20947 11747
rect 21557 11713 21591 11747
rect 1869 11645 1903 11679
rect 3985 11645 4019 11679
rect 4537 11645 4571 11679
rect 4813 11645 4847 11679
rect 5365 11645 5399 11679
rect 6929 11645 6963 11679
rect 7205 11645 7239 11679
rect 7481 11645 7515 11679
rect 9137 11645 9171 11679
rect 9689 11645 9723 11679
rect 10241 11645 10275 11679
rect 10333 11645 10367 11679
rect 10517 11645 10551 11679
rect 12449 11645 12483 11679
rect 15025 11645 15059 11679
rect 15485 11645 15519 11679
rect 17693 11645 17727 11679
rect 21741 11645 21775 11679
rect 22201 11645 22235 11679
rect 3525 11577 3559 11611
rect 6193 11577 6227 11611
rect 12909 11577 12943 11611
rect 13645 11577 13679 11611
rect 14197 11577 14231 11611
rect 14933 11577 14967 11611
rect 16358 11577 16392 11611
rect 20361 11577 20395 11611
rect 2237 11509 2271 11543
rect 4077 11509 4111 11543
rect 6561 11509 6595 11543
rect 6929 11509 6963 11543
rect 10149 11509 10183 11543
rect 11897 11509 11931 11543
rect 12633 11509 12667 11543
rect 13277 11509 13311 11543
rect 15945 11509 15979 11543
rect 16957 11509 16991 11543
rect 18705 11509 18739 11543
rect 19257 11509 19291 11543
rect 19625 11509 19659 11543
rect 20085 11509 20119 11543
rect 21833 11509 21867 11543
rect 1869 11305 1903 11339
rect 3065 11305 3099 11339
rect 3893 11305 3927 11339
rect 5457 11305 5491 11339
rect 6653 11305 6687 11339
rect 6929 11305 6963 11339
rect 10241 11305 10275 11339
rect 13553 11305 13587 11339
rect 14197 11305 14231 11339
rect 15577 11305 15611 11339
rect 16129 11305 16163 11339
rect 18383 11305 18417 11339
rect 20361 11305 20395 11339
rect 22661 11305 22695 11339
rect 2145 11237 2179 11271
rect 2237 11237 2271 11271
rect 5825 11237 5859 11271
rect 12627 11237 12661 11271
rect 16313 11237 16347 11271
rect 16405 11237 16439 11271
rect 18981 11237 19015 11271
rect 19165 11237 19199 11271
rect 19441 11237 19475 11271
rect 21097 11237 21131 11271
rect 4169 11169 4203 11203
rect 4537 11169 4571 11203
rect 4905 11169 4939 11203
rect 5457 11169 5491 11203
rect 7389 11169 7423 11203
rect 7573 11169 7607 11203
rect 7941 11169 7975 11203
rect 8493 11169 8527 11203
rect 8861 11169 8895 11203
rect 9689 11169 9723 11203
rect 11345 11169 11379 11203
rect 13185 11169 13219 11203
rect 14013 11169 14047 11203
rect 18705 11169 18739 11203
rect 2421 11101 2455 11135
rect 3525 11101 3559 11135
rect 8585 11101 8619 11135
rect 12265 11101 12299 11135
rect 9873 11033 9907 11067
rect 11161 11033 11195 11067
rect 16865 11033 16899 11067
rect 6285 10965 6319 10999
rect 13829 10965 13863 10999
rect 18153 10965 18187 10999
rect 22477 11169 22511 11203
rect 19349 11101 19383 11135
rect 21005 11101 21039 11135
rect 19901 11033 19935 11067
rect 21557 11033 21591 11067
rect 18981 10965 19015 10999
rect 20637 10965 20671 10999
rect 3157 10761 3191 10795
rect 4997 10761 5031 10795
rect 6653 10761 6687 10795
rect 7021 10761 7055 10795
rect 11345 10761 11379 10795
rect 11805 10761 11839 10795
rect 12265 10761 12299 10795
rect 12725 10761 12759 10795
rect 14013 10761 14047 10795
rect 14749 10761 14783 10795
rect 17141 10761 17175 10795
rect 19809 10761 19843 10795
rect 21373 10761 21407 10795
rect 21741 10761 21775 10795
rect 22063 10761 22097 10795
rect 3433 10693 3467 10727
rect 5273 10693 5307 10727
rect 9137 10693 9171 10727
rect 2145 10625 2179 10659
rect 2421 10625 2455 10659
rect 4629 10625 4663 10659
rect 5917 10625 5951 10659
rect 8677 10625 8711 10659
rect 12817 10625 12851 10659
rect 15485 10625 15519 10659
rect 15945 10625 15979 10659
rect 17877 10625 17911 10659
rect 18613 10625 18647 10659
rect 20453 10625 20487 10659
rect 22477 10625 22511 10659
rect 3709 10557 3743 10591
rect 5181 10557 5215 10591
rect 5457 10557 5491 10591
rect 7389 10557 7423 10591
rect 7665 10557 7699 10591
rect 8217 10557 8251 10591
rect 8585 10557 8619 10591
rect 9965 10557 9999 10591
rect 10057 10557 10091 10591
rect 10241 10557 10275 10591
rect 14565 10557 14599 10591
rect 15025 10557 15059 10591
rect 19533 10557 19567 10591
rect 20177 10557 20211 10591
rect 21992 10557 22026 10591
rect 2237 10489 2271 10523
rect 9873 10489 9907 10523
rect 10701 10489 10735 10523
rect 13138 10489 13172 10523
rect 15761 10489 15795 10523
rect 16266 10489 16300 10523
rect 18934 10489 18968 10523
rect 20545 10489 20579 10523
rect 21097 10489 21131 10523
rect 1961 10421 1995 10455
rect 4077 10421 4111 10455
rect 6193 10421 6227 10455
rect 9413 10421 9447 10455
rect 11069 10421 11103 10455
rect 13737 10421 13771 10455
rect 16865 10421 16899 10455
rect 18245 10421 18279 10455
rect 22753 10421 22787 10455
rect 2789 10217 2823 10251
rect 4169 10217 4203 10251
rect 6837 10217 6871 10251
rect 8769 10217 8803 10251
rect 12633 10217 12667 10251
rect 12909 10217 12943 10251
rect 15485 10217 15519 10251
rect 16313 10217 16347 10251
rect 19349 10217 19383 10251
rect 20453 10217 20487 10251
rect 2190 10149 2224 10183
rect 3157 10149 3191 10183
rect 9965 10149 9999 10183
rect 12265 10149 12299 10183
rect 13737 10149 13771 10183
rect 14289 10149 14323 10183
rect 14565 10149 14599 10183
rect 16681 10149 16715 10183
rect 16773 10149 16807 10183
rect 18750 10149 18784 10183
rect 21097 10149 21131 10183
rect 1869 10081 1903 10115
rect 3433 10081 3467 10115
rect 4077 10081 4111 10115
rect 4629 10081 4663 10115
rect 4905 10081 4939 10115
rect 5365 10081 5399 10115
rect 6837 10081 6871 10115
rect 7297 10081 7331 10115
rect 7389 10081 7423 10115
rect 7941 10081 7975 10115
rect 10517 10081 10551 10115
rect 11529 10081 11563 10115
rect 11805 10081 11839 10115
rect 15301 10081 15335 10115
rect 17325 10081 17359 10115
rect 22477 10081 22511 10115
rect 24593 10081 24627 10115
rect 13645 10013 13679 10047
rect 18429 10013 18463 10047
rect 21005 10013 21039 10047
rect 21281 10013 21315 10047
rect 3893 9945 3927 9979
rect 11621 9945 11655 9979
rect 19717 9945 19751 9979
rect 22615 9945 22649 9979
rect 1777 9877 1811 9911
rect 6101 9877 6135 9911
rect 6377 9877 6411 9911
rect 8309 9877 8343 9911
rect 9137 9877 9171 9911
rect 10977 9877 11011 9911
rect 11345 9877 11379 9911
rect 15853 9877 15887 9911
rect 24731 9877 24765 9911
rect 9413 9673 9447 9707
rect 13553 9673 13587 9707
rect 16865 9673 16899 9707
rect 17877 9673 17911 9707
rect 21189 9673 21223 9707
rect 21557 9673 21591 9707
rect 24685 9673 24719 9707
rect 6653 9605 6687 9639
rect 10609 9605 10643 9639
rect 11529 9605 11563 9639
rect 11897 9605 11931 9639
rect 15209 9605 15243 9639
rect 17141 9605 17175 9639
rect 22477 9605 22511 9639
rect 2053 9537 2087 9571
rect 2329 9537 2363 9571
rect 8585 9537 8619 9571
rect 11253 9537 11287 9571
rect 14289 9537 14323 9571
rect 14933 9537 14967 9571
rect 16129 9537 16163 9571
rect 18245 9537 18279 9571
rect 18429 9537 18463 9571
rect 20269 9537 20303 9571
rect 20913 9537 20947 9571
rect 4261 9469 4295 9503
rect 4629 9469 4663 9503
rect 4813 9469 4847 9503
rect 5365 9469 5399 9503
rect 7113 9469 7147 9503
rect 7389 9469 7423 9503
rect 7665 9469 7699 9503
rect 8217 9469 8251 9503
rect 9505 9469 9539 9503
rect 10517 9469 10551 9503
rect 10793 9469 10827 9503
rect 12633 9469 12667 9503
rect 12909 9469 12943 9503
rect 2145 9401 2179 9435
rect 6285 9401 6319 9435
rect 14381 9401 14415 9435
rect 15853 9401 15887 9435
rect 15945 9401 15979 9435
rect 18750 9401 18784 9435
rect 20361 9401 20395 9435
rect 1869 9333 1903 9367
rect 2973 9333 3007 9367
rect 3525 9333 3559 9367
rect 3801 9333 3835 9367
rect 4077 9333 4111 9367
rect 5733 9333 5767 9367
rect 6929 9333 6963 9367
rect 9045 9333 9079 9367
rect 9689 9333 9723 9367
rect 10057 9333 10091 9367
rect 10425 9333 10459 9367
rect 12541 9333 12575 9367
rect 14013 9333 14047 9367
rect 15577 9333 15611 9367
rect 19349 9333 19383 9367
rect 19993 9333 20027 9367
rect 1777 9129 1811 9163
rect 3801 9129 3835 9163
rect 8677 9129 8711 9163
rect 11529 9129 11563 9163
rect 12817 9129 12851 9163
rect 18429 9129 18463 9163
rect 20177 9129 20211 9163
rect 20913 9129 20947 9163
rect 22477 9129 22511 9163
rect 2231 9061 2265 9095
rect 3433 9061 3467 9095
rect 4261 9061 4295 9095
rect 5825 9061 5859 9095
rect 10885 9061 10919 9095
rect 14381 9061 14415 9095
rect 18061 9061 18095 9095
rect 1869 8993 1903 9027
rect 5917 8993 5951 9027
rect 7205 8993 7239 9027
rect 7389 8993 7423 9027
rect 7757 8993 7791 9027
rect 8309 8993 8343 9027
rect 10793 8993 10827 9027
rect 11713 8993 11747 9027
rect 11989 8993 12023 9027
rect 13829 8993 13863 9027
rect 15393 8993 15427 9027
rect 17325 8993 17359 9027
rect 17785 8993 17819 9027
rect 19717 8993 19751 9027
rect 22293 8993 22327 9027
rect 4169 8925 4203 8959
rect 4445 8925 4479 8959
rect 8401 8925 8435 8959
rect 12449 8925 12483 8959
rect 3157 8857 3191 8891
rect 6561 8857 6595 8891
rect 11805 8857 11839 8891
rect 2789 8789 2823 8823
rect 5089 8789 5123 8823
rect 6101 8789 6135 8823
rect 9137 8789 9171 8823
rect 13553 8789 13587 8823
rect 15761 8789 15795 8823
rect 18797 8789 18831 8823
rect 19855 8789 19889 8823
rect 3617 8585 3651 8619
rect 6193 8585 6227 8619
rect 6561 8585 6595 8619
rect 7113 8585 7147 8619
rect 7481 8585 7515 8619
rect 10241 8585 10275 8619
rect 13461 8585 13495 8619
rect 14197 8585 14231 8619
rect 15393 8585 15427 8619
rect 15761 8585 15795 8619
rect 17325 8585 17359 8619
rect 22293 8585 22327 8619
rect 23811 8585 23845 8619
rect 3341 8517 3375 8551
rect 13829 8517 13863 8551
rect 17049 8517 17083 8551
rect 19809 8517 19843 8551
rect 2145 8449 2179 8483
rect 12541 8449 12575 8483
rect 15025 8449 15059 8483
rect 16221 8449 16255 8483
rect 18797 8449 18831 8483
rect 19441 8449 19475 8483
rect 19993 8449 20027 8483
rect 20269 8449 20303 8483
rect 3433 8381 3467 8415
rect 4721 8381 4755 8415
rect 5181 8381 5215 8415
rect 5273 8381 5307 8415
rect 5641 8381 5675 8415
rect 6929 8381 6963 8415
rect 7941 8381 7975 8415
rect 8401 8381 8435 8415
rect 8953 8381 8987 8415
rect 9137 8381 9171 8415
rect 11805 8381 11839 8415
rect 17785 8381 17819 8415
rect 18061 8381 18095 8415
rect 18521 8381 18555 8415
rect 23740 8381 23774 8415
rect 24133 8381 24167 8415
rect 1777 8313 1811 8347
rect 1869 8313 1903 8347
rect 5917 8313 5951 8347
rect 9413 8313 9447 8347
rect 10517 8313 10551 8347
rect 10609 8313 10643 8347
rect 11161 8313 11195 8347
rect 12903 8313 12937 8347
rect 14381 8313 14415 8347
rect 14473 8313 14507 8347
rect 15945 8313 15979 8347
rect 16037 8313 16071 8347
rect 20085 8313 20119 8347
rect 2789 8245 2823 8279
rect 4077 8245 4111 8279
rect 7849 8245 7883 8279
rect 9689 8245 9723 8279
rect 12265 8245 12299 8279
rect 2053 8041 2087 8075
rect 3525 8041 3559 8075
rect 3801 8041 3835 8075
rect 12725 8041 12759 8075
rect 14197 8041 14231 8075
rect 16405 8041 16439 8075
rect 18521 8041 18555 8075
rect 19993 8041 20027 8075
rect 1777 7973 1811 8007
rect 2421 7973 2455 8007
rect 2973 7973 3007 8007
rect 11161 7973 11195 8007
rect 11529 7973 11563 8007
rect 12449 7973 12483 8007
rect 13639 7973 13673 8007
rect 15393 7973 15427 8007
rect 15485 7973 15519 8007
rect 4537 7905 4571 7939
rect 5273 7905 5307 7939
rect 5733 7905 5767 7939
rect 6009 7905 6043 7939
rect 6193 7905 6227 7939
rect 7573 7905 7607 7939
rect 7757 7905 7791 7939
rect 8125 7905 8159 7939
rect 8493 7905 8527 7939
rect 10425 7905 10459 7939
rect 13277 7905 13311 7939
rect 16865 7905 16899 7939
rect 2329 7837 2363 7871
rect 4905 7837 4939 7871
rect 6469 7837 6503 7871
rect 11437 7837 11471 7871
rect 12081 7837 12115 7871
rect 17969 7837 18003 7871
rect 8677 7769 8711 7803
rect 14473 7769 14507 7803
rect 15945 7769 15979 7803
rect 6929 7701 6963 7735
rect 9137 7701 9171 7735
rect 9413 7701 9447 7735
rect 10057 7701 10091 7735
rect 10885 7701 10919 7735
rect 17049 7701 17083 7735
rect 2789 7497 2823 7531
rect 4629 7497 4663 7531
rect 5549 7497 5583 7531
rect 5917 7497 5951 7531
rect 6975 7497 7009 7531
rect 11345 7497 11379 7531
rect 11713 7497 11747 7531
rect 14151 7497 14185 7531
rect 16313 7497 16347 7531
rect 18613 7497 18647 7531
rect 3893 7429 3927 7463
rect 7665 7429 7699 7463
rect 13829 7429 13863 7463
rect 16911 7429 16945 7463
rect 17601 7429 17635 7463
rect 2421 7361 2455 7395
rect 7389 7361 7423 7395
rect 10149 7361 10183 7395
rect 12817 7361 12851 7395
rect 15301 7361 15335 7395
rect 15945 7361 15979 7395
rect 2329 7293 2363 7327
rect 3709 7293 3743 7327
rect 4721 7293 4755 7327
rect 5181 7293 5215 7327
rect 5733 7293 5767 7327
rect 6193 7293 6227 7327
rect 6904 7293 6938 7327
rect 8033 7293 8067 7327
rect 8401 7293 8435 7327
rect 8861 7293 8895 7327
rect 9137 7293 9171 7327
rect 11069 7293 11103 7327
rect 14080 7293 14114 7327
rect 14473 7293 14507 7327
rect 16808 7293 16842 7327
rect 17233 7293 17267 7327
rect 18112 7293 18146 7327
rect 24660 7293 24694 7327
rect 4261 7225 4295 7259
rect 9321 7225 9355 7259
rect 10470 7225 10504 7259
rect 12541 7225 12575 7259
rect 12633 7225 12667 7259
rect 15393 7225 15427 7259
rect 18199 7225 18233 7259
rect 3157 7157 3191 7191
rect 3525 7157 3559 7191
rect 4905 7157 4939 7191
rect 6561 7157 6595 7191
rect 9597 7157 9631 7191
rect 9965 7157 9999 7191
rect 12173 7157 12207 7191
rect 13461 7157 13495 7191
rect 15117 7157 15151 7191
rect 16589 7157 16623 7191
rect 24731 7157 24765 7191
rect 25145 7157 25179 7191
rect 1409 6953 1443 6987
rect 4261 6953 4295 6987
rect 6653 6953 6687 6987
rect 8493 6953 8527 6987
rect 8861 6953 8895 6987
rect 9229 6953 9263 6987
rect 10057 6953 10091 6987
rect 10609 6953 10643 6987
rect 12817 6953 12851 6987
rect 13461 6953 13495 6987
rect 15117 6953 15151 6987
rect 15577 6953 15611 6987
rect 24777 6953 24811 6987
rect 1869 6885 1903 6919
rect 2329 6885 2363 6919
rect 3157 6885 3191 6919
rect 5549 6885 5583 6919
rect 10885 6885 10919 6919
rect 12173 6885 12207 6919
rect 2421 6817 2455 6851
rect 2697 6817 2731 6851
rect 4905 6817 4939 6851
rect 6377 6817 6411 6851
rect 7113 6817 7147 6851
rect 7205 6817 7239 6851
rect 7665 6817 7699 6851
rect 8217 6817 8251 6851
rect 11529 6817 11563 6851
rect 13001 6817 13035 6851
rect 13277 6817 13311 6851
rect 15485 6817 15519 6851
rect 16900 6817 16934 6851
rect 24593 6817 24627 6851
rect 9689 6749 9723 6783
rect 13093 6749 13127 6783
rect 2513 6681 2547 6715
rect 3433 6613 3467 6647
rect 4629 6613 4663 6647
rect 5825 6613 5859 6647
rect 6193 6613 6227 6647
rect 11345 6613 11379 6647
rect 12449 6613 12483 6647
rect 14289 6613 14323 6647
rect 17003 6613 17037 6647
rect 1593 6409 1627 6443
rect 6101 6409 6135 6443
rect 10057 6409 10091 6443
rect 11253 6409 11287 6443
rect 14013 6409 14047 6443
rect 15393 6409 15427 6443
rect 16865 6409 16899 6443
rect 23949 6409 23983 6443
rect 5641 6341 5675 6375
rect 11805 6341 11839 6375
rect 5089 6273 5123 6307
rect 9045 6273 9079 6307
rect 10333 6273 10367 6307
rect 10977 6273 11011 6307
rect 12449 6273 12483 6307
rect 15761 6273 15795 6307
rect 1409 6205 1443 6239
rect 1961 6205 1995 6239
rect 3065 6205 3099 6239
rect 3157 6205 3191 6239
rect 3341 6205 3375 6239
rect 4629 6205 4663 6239
rect 4721 6205 4755 6239
rect 4905 6205 4939 6239
rect 7297 6205 7331 6239
rect 7757 6205 7791 6239
rect 8125 6205 8159 6239
rect 8677 6205 8711 6239
rect 13369 6205 13403 6239
rect 14473 6205 14507 6239
rect 18061 6205 18095 6239
rect 18613 6205 18647 6239
rect 23740 6205 23774 6239
rect 24133 6205 24167 6239
rect 2881 6137 2915 6171
rect 3801 6137 3835 6171
rect 7205 6137 7239 6171
rect 10425 6137 10459 6171
rect 12770 6137 12804 6171
rect 14197 6137 14231 6171
rect 24593 6137 24627 6171
rect 2513 6069 2547 6103
rect 4077 6069 4111 6103
rect 4445 6069 4479 6103
rect 6469 6069 6503 6103
rect 7573 6069 7607 6103
rect 9689 6069 9723 6103
rect 12265 6069 12299 6103
rect 13737 6069 13771 6103
rect 18245 6069 18279 6103
rect 3433 5865 3467 5899
rect 5089 5865 5123 5899
rect 6009 5865 6043 5899
rect 6469 5865 6503 5899
rect 7389 5865 7423 5899
rect 8769 5865 8803 5899
rect 11437 5865 11471 5899
rect 13093 5865 13127 5899
rect 14059 5865 14093 5899
rect 3157 5797 3191 5831
rect 4077 5797 4111 5831
rect 7665 5797 7699 5831
rect 8170 5797 8204 5831
rect 9873 5797 9907 5831
rect 12494 5797 12528 5831
rect 13369 5797 13403 5831
rect 15485 5797 15519 5831
rect 2789 5729 2823 5763
rect 4169 5729 4203 5763
rect 5825 5729 5859 5763
rect 6872 5729 6906 5763
rect 7849 5729 7883 5763
rect 12173 5729 12207 5763
rect 13956 5729 13990 5763
rect 2329 5661 2363 5695
rect 9781 5661 9815 5695
rect 10425 5661 10459 5695
rect 15393 5661 15427 5695
rect 16037 5661 16071 5695
rect 6975 5525 7009 5559
rect 10701 5525 10735 5559
rect 14473 5525 14507 5559
rect 4537 5321 4571 5355
rect 5917 5321 5951 5355
rect 12173 5321 12207 5355
rect 13921 5321 13955 5355
rect 16865 5321 16899 5355
rect 5641 5253 5675 5287
rect 6285 5253 6319 5287
rect 14933 5253 14967 5287
rect 15669 5253 15703 5287
rect 2881 5185 2915 5219
rect 4077 5185 4111 5219
rect 6837 5185 6871 5219
rect 10885 5185 10919 5219
rect 13461 5185 13495 5219
rect 15393 5185 15427 5219
rect 15853 5185 15887 5219
rect 2789 5117 2823 5151
rect 3065 5117 3099 5151
rect 4353 5117 4387 5151
rect 4813 5117 4847 5151
rect 5733 5117 5767 5151
rect 15945 5117 15979 5151
rect 3525 5049 3559 5083
rect 6561 5049 6595 5083
rect 7158 5049 7192 5083
rect 8033 5049 8067 5083
rect 8677 5049 8711 5083
rect 8769 5049 8803 5083
rect 9321 5049 9355 5083
rect 9689 5049 9723 5083
rect 10241 5049 10275 5083
rect 10333 5049 10367 5083
rect 11897 5049 11931 5083
rect 12817 5049 12851 5083
rect 12909 5049 12943 5083
rect 14381 5049 14415 5083
rect 14473 5049 14507 5083
rect 2053 4981 2087 5015
rect 2513 4981 2547 5015
rect 7757 4981 7791 5015
rect 8401 4981 8435 5015
rect 9965 4981 9999 5015
rect 11161 4981 11195 5015
rect 7297 4777 7331 4811
rect 8401 4777 8435 4811
rect 9965 4777 9999 4811
rect 11759 4777 11793 4811
rect 14657 4777 14691 4811
rect 2145 4709 2179 4743
rect 3157 4709 3191 4743
rect 7481 4709 7515 4743
rect 7573 4709 7607 4743
rect 8125 4709 8159 4743
rect 9413 4709 9447 4743
rect 12173 4709 12207 4743
rect 13838 4709 13872 4743
rect 15485 4709 15519 4743
rect 16037 4709 16071 4743
rect 1501 4641 1535 4675
rect 5768 4641 5802 4675
rect 10333 4641 10367 4675
rect 11656 4641 11690 4675
rect 12668 4641 12702 4675
rect 24660 4641 24694 4675
rect 5871 4573 5905 4607
rect 8769 4573 8803 4607
rect 12771 4573 12805 4607
rect 13737 4573 13771 4607
rect 14381 4573 14415 4607
rect 15393 4573 15427 4607
rect 6837 4505 6871 4539
rect 13185 4505 13219 4539
rect 2789 4437 2823 4471
rect 24731 4437 24765 4471
rect 5733 4233 5767 4267
rect 7941 4233 7975 4267
rect 9275 4233 9309 4267
rect 11805 4233 11839 4267
rect 12633 4233 12667 4267
rect 13737 4233 13771 4267
rect 15393 4233 15427 4267
rect 24685 4233 24719 4267
rect 9965 4165 9999 4199
rect 14105 4165 14139 4199
rect 7665 4097 7699 4131
rect 10149 4097 10183 4131
rect 11345 4097 11379 4131
rect 13185 4097 13219 4131
rect 14565 4097 14599 4131
rect 15669 4097 15703 4131
rect 6653 4029 6687 4063
rect 7573 4029 7607 4063
rect 9204 4029 9238 4063
rect 14289 3961 14323 3995
rect 14381 3961 14415 3995
rect 1593 3893 1627 3927
rect 9597 3893 9631 3927
rect 1547 3689 1581 3723
rect 7389 3689 7423 3723
rect 13737 3689 13771 3723
rect 1409 3553 1443 3587
rect 15368 3553 15402 3587
rect 24660 3553 24694 3587
rect 14289 3417 14323 3451
rect 24731 3417 24765 3451
rect 15439 3349 15473 3383
rect 9781 3145 9815 3179
rect 11437 3145 11471 3179
rect 15393 3145 15427 3179
rect 24685 3145 24719 3179
rect 1593 3077 1627 3111
rect 9321 3077 9355 3111
rect 10977 3077 11011 3111
rect 9137 2941 9171 2975
rect 10793 2941 10827 2975
rect 15669 2941 15703 2975
rect 16221 2941 16255 2975
rect 15853 2805 15887 2839
rect 14841 2601 14875 2635
rect 16267 2601 16301 2635
rect 20361 2601 20395 2635
rect 22799 2601 22833 2635
rect 23213 2533 23247 2567
rect 6929 2465 6963 2499
rect 7573 2465 7607 2499
rect 11161 2465 11195 2499
rect 11713 2465 11747 2499
rect 14289 2465 14323 2499
rect 16196 2465 16230 2499
rect 20152 2465 20186 2499
rect 21624 2465 21658 2499
rect 22728 2465 22762 2499
rect 24108 2465 24142 2499
rect 11345 2329 11379 2363
rect 20637 2329 20671 2363
rect 7113 2261 7147 2295
rect 14473 2261 14507 2295
rect 16681 2261 16715 2295
rect 21695 2261 21729 2295
rect 22109 2261 22143 2295
rect 24179 2261 24213 2295
rect 24593 2261 24627 2295
<< metal1 >>
rect 14 27480 20 27532
rect 72 27520 78 27532
rect 658 27520 664 27532
rect 72 27492 664 27520
rect 72 27480 78 27492
rect 658 27480 664 27492
rect 716 27480 722 27532
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 11606 24828 11612 24880
rect 11664 24868 11670 24880
rect 27614 24868 27620 24880
rect 11664 24840 27620 24868
rect 11664 24828 11670 24840
rect 27614 24828 27620 24840
rect 27672 24828 27678 24880
rect 11238 24556 11244 24608
rect 11296 24596 11302 24608
rect 13170 24596 13176 24608
rect 11296 24568 13176 24596
rect 11296 24556 11302 24568
rect 13170 24556 13176 24568
rect 13228 24556 13234 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 7466 24392 7472 24404
rect 7427 24364 7472 24392
rect 7466 24352 7472 24364
rect 7524 24352 7530 24404
rect 7282 24256 7288 24268
rect 7243 24228 7288 24256
rect 7282 24216 7288 24228
rect 7340 24216 7346 24268
rect 11517 24259 11575 24265
rect 11517 24225 11529 24259
rect 11563 24256 11575 24259
rect 11606 24256 11612 24268
rect 11563 24228 11612 24256
rect 11563 24225 11575 24228
rect 11517 24219 11575 24225
rect 11606 24216 11612 24228
rect 11664 24216 11670 24268
rect 10042 24012 10048 24064
rect 10100 24052 10106 24064
rect 11655 24055 11713 24061
rect 11655 24052 11667 24055
rect 10100 24024 11667 24052
rect 10100 24012 10106 24024
rect 11655 24021 11667 24024
rect 11701 24021 11713 24055
rect 11655 24015 11713 24021
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 8021 23851 8079 23857
rect 8021 23817 8033 23851
rect 8067 23848 8079 23851
rect 9030 23848 9036 23860
rect 8067 23820 9036 23848
rect 8067 23817 8079 23820
rect 8021 23811 8079 23817
rect 9030 23808 9036 23820
rect 9088 23808 9094 23860
rect 10781 23851 10839 23857
rect 10781 23817 10793 23851
rect 10827 23848 10839 23851
rect 11422 23848 11428 23860
rect 10827 23820 11428 23848
rect 10827 23817 10839 23820
rect 10781 23811 10839 23817
rect 11422 23808 11428 23820
rect 11480 23808 11486 23860
rect 11606 23848 11612 23860
rect 11567 23820 11612 23848
rect 11606 23808 11612 23820
rect 11664 23808 11670 23860
rect 18325 23851 18383 23857
rect 18325 23817 18337 23851
rect 18371 23848 18383 23851
rect 20162 23848 20168 23860
rect 18371 23820 20168 23848
rect 18371 23817 18383 23820
rect 18325 23811 18383 23817
rect 20162 23808 20168 23820
rect 20220 23808 20226 23860
rect 20717 23851 20775 23857
rect 20717 23817 20729 23851
rect 20763 23848 20775 23851
rect 21634 23848 21640 23860
rect 20763 23820 21640 23848
rect 20763 23817 20775 23820
rect 20717 23811 20775 23817
rect 11238 23780 11244 23792
rect 11199 23752 11244 23780
rect 11238 23740 11244 23752
rect 11296 23740 11302 23792
rect 1302 23672 1308 23724
rect 1360 23712 1366 23724
rect 1857 23715 1915 23721
rect 1857 23712 1869 23715
rect 1360 23684 1869 23712
rect 1360 23672 1366 23684
rect 1479 23653 1507 23684
rect 1857 23681 1869 23684
rect 1903 23681 1915 23715
rect 1857 23675 1915 23681
rect 1464 23647 1522 23653
rect 1464 23613 1476 23647
rect 1510 23613 1522 23647
rect 7834 23644 7840 23656
rect 7747 23616 7840 23644
rect 1464 23607 1522 23613
rect 7834 23604 7840 23616
rect 7892 23644 7898 23656
rect 8389 23647 8447 23653
rect 8389 23644 8401 23647
rect 7892 23616 8401 23644
rect 7892 23604 7898 23616
rect 8389 23613 8401 23616
rect 8435 23613 8447 23647
rect 8389 23607 8447 23613
rect 10597 23647 10655 23653
rect 10597 23613 10609 23647
rect 10643 23644 10655 23647
rect 11238 23644 11244 23656
rect 10643 23616 11244 23644
rect 10643 23613 10655 23616
rect 10597 23607 10655 23613
rect 11238 23604 11244 23616
rect 11296 23604 11302 23656
rect 15984 23647 16042 23653
rect 15984 23613 15996 23647
rect 16030 23644 16042 23647
rect 16071 23647 16129 23653
rect 16030 23613 16043 23644
rect 15984 23607 16043 23613
rect 16071 23613 16083 23647
rect 16117 23644 16129 23647
rect 16390 23644 16396 23656
rect 16117 23616 16396 23644
rect 16117 23613 16129 23616
rect 16071 23607 16129 23613
rect 16015 23576 16043 23607
rect 16390 23604 16396 23616
rect 16448 23604 16454 23656
rect 16482 23604 16488 23656
rect 16540 23644 16546 23656
rect 18138 23644 18144 23656
rect 16540 23616 16585 23644
rect 18051 23616 18144 23644
rect 16540 23604 16546 23616
rect 18138 23604 18144 23616
rect 18196 23644 18202 23656
rect 18693 23647 18751 23653
rect 18693 23644 18705 23647
rect 18196 23616 18705 23644
rect 18196 23604 18202 23616
rect 18693 23613 18705 23616
rect 18739 23613 18751 23647
rect 18693 23607 18751 23613
rect 20232 23647 20290 23653
rect 20232 23613 20244 23647
rect 20278 23644 20290 23647
rect 20732 23644 20760 23811
rect 21634 23808 21640 23820
rect 21692 23808 21698 23860
rect 21729 23851 21787 23857
rect 21729 23817 21741 23851
rect 21775 23848 21787 23851
rect 23014 23848 23020 23860
rect 21775 23820 23020 23848
rect 21775 23817 21787 23820
rect 21729 23811 21787 23817
rect 20278 23616 20760 23644
rect 21228 23647 21286 23653
rect 20278 23613 20290 23616
rect 20232 23607 20290 23613
rect 21228 23613 21240 23647
rect 21274 23644 21286 23647
rect 21744 23644 21772 23811
rect 23014 23808 23020 23820
rect 23072 23808 23078 23860
rect 25225 23851 25283 23857
rect 25225 23817 25237 23851
rect 25271 23848 25283 23851
rect 27154 23848 27160 23860
rect 25271 23820 27160 23848
rect 25271 23817 25283 23820
rect 25225 23811 25283 23817
rect 22278 23740 22284 23792
rect 22336 23780 22342 23792
rect 24811 23783 24869 23789
rect 24811 23780 24823 23783
rect 22336 23752 24823 23780
rect 22336 23740 22342 23752
rect 24811 23749 24823 23752
rect 24857 23749 24869 23783
rect 24811 23743 24869 23749
rect 21274 23616 21772 23644
rect 23728 23647 23786 23653
rect 21274 23613 21286 23616
rect 21228 23607 21286 23613
rect 23728 23613 23740 23647
rect 23774 23644 23786 23647
rect 24740 23647 24798 23653
rect 23774 23616 24256 23644
rect 23774 23613 23786 23616
rect 23728 23607 23786 23613
rect 16500 23576 16528 23604
rect 16015 23548 16528 23576
rect 19426 23536 19432 23588
rect 19484 23576 19490 23588
rect 24228 23585 24256 23616
rect 24740 23613 24752 23647
rect 24786 23644 24798 23647
rect 25240 23644 25268 23811
rect 27154 23808 27160 23820
rect 27212 23808 27218 23860
rect 24786 23616 25268 23644
rect 24786 23613 24798 23616
rect 24740 23607 24798 23613
rect 21315 23579 21373 23585
rect 21315 23576 21327 23579
rect 19484 23548 21327 23576
rect 19484 23536 19490 23548
rect 21315 23545 21327 23548
rect 21361 23545 21373 23579
rect 21315 23539 21373 23545
rect 24213 23579 24271 23585
rect 24213 23545 24225 23579
rect 24259 23576 24271 23579
rect 25774 23576 25780 23588
rect 24259 23548 25780 23576
rect 24259 23545 24271 23548
rect 24213 23539 24271 23545
rect 25774 23536 25780 23548
rect 25832 23536 25838 23588
rect 1535 23511 1593 23517
rect 1535 23477 1547 23511
rect 1581 23508 1593 23511
rect 1670 23508 1676 23520
rect 1581 23480 1676 23508
rect 1581 23477 1593 23480
rect 1535 23471 1593 23477
rect 1670 23468 1676 23480
rect 1728 23468 1734 23520
rect 7282 23468 7288 23520
rect 7340 23508 7346 23520
rect 7377 23511 7435 23517
rect 7377 23508 7389 23511
rect 7340 23480 7389 23508
rect 7340 23468 7346 23480
rect 7377 23477 7389 23480
rect 7423 23508 7435 23511
rect 7742 23508 7748 23520
rect 7423 23480 7748 23508
rect 7423 23477 7435 23480
rect 7377 23471 7435 23477
rect 7742 23468 7748 23480
rect 7800 23468 7806 23520
rect 19978 23468 19984 23520
rect 20036 23508 20042 23520
rect 20303 23511 20361 23517
rect 20303 23508 20315 23511
rect 20036 23480 20315 23508
rect 20036 23468 20042 23480
rect 20303 23477 20315 23480
rect 20349 23477 20361 23511
rect 20303 23471 20361 23477
rect 22554 23468 22560 23520
rect 22612 23508 22618 23520
rect 23799 23511 23857 23517
rect 23799 23508 23811 23511
rect 22612 23480 23811 23508
rect 22612 23468 22618 23480
rect 23799 23477 23811 23480
rect 23845 23477 23857 23511
rect 23799 23471 23857 23477
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 15654 23236 15660 23248
rect 15615 23208 15660 23236
rect 15654 23196 15660 23208
rect 15712 23196 15718 23248
rect 1210 23128 1216 23180
rect 1268 23168 1274 23180
rect 1464 23171 1522 23177
rect 1464 23168 1476 23171
rect 1268 23140 1476 23168
rect 1268 23128 1274 23140
rect 1464 23137 1476 23140
rect 1510 23168 1522 23171
rect 2222 23168 2228 23180
rect 1510 23140 2228 23168
rect 1510 23137 1522 23140
rect 1464 23131 1522 23137
rect 2222 23128 2228 23140
rect 2280 23128 2286 23180
rect 8478 23128 8484 23180
rect 8536 23168 8542 23180
rect 8608 23171 8666 23177
rect 8608 23168 8620 23171
rect 8536 23140 8620 23168
rect 8536 23128 8542 23140
rect 8608 23137 8620 23140
rect 8654 23137 8666 23171
rect 13630 23168 13636 23180
rect 13591 23140 13636 23168
rect 8608 23131 8666 23137
rect 13630 23128 13636 23140
rect 13688 23128 13694 23180
rect 14090 23168 14096 23180
rect 14051 23140 14096 23168
rect 14090 23128 14096 23140
rect 14148 23128 14154 23180
rect 16298 23128 16304 23180
rect 16356 23168 16362 23180
rect 17072 23171 17130 23177
rect 17072 23168 17084 23171
rect 16356 23140 17084 23168
rect 16356 23128 16362 23140
rect 17072 23137 17084 23140
rect 17118 23168 17130 23171
rect 17310 23168 17316 23180
rect 17118 23140 17316 23168
rect 17118 23137 17130 23140
rect 17072 23131 17130 23137
rect 17310 23128 17316 23140
rect 17368 23128 17374 23180
rect 20990 23177 20996 23180
rect 20968 23171 20996 23177
rect 20968 23168 20980 23171
rect 20903 23140 20980 23168
rect 20968 23137 20980 23140
rect 21048 23168 21054 23180
rect 24118 23168 24124 23180
rect 21048 23140 24124 23168
rect 20968 23131 20996 23137
rect 20990 23128 20996 23131
rect 21048 23128 21054 23140
rect 24118 23128 24124 23140
rect 24176 23128 24182 23180
rect 14274 23100 14280 23112
rect 14235 23072 14280 23100
rect 14274 23060 14280 23072
rect 14332 23060 14338 23112
rect 15565 23103 15623 23109
rect 15565 23069 15577 23103
rect 15611 23100 15623 23103
rect 16390 23100 16396 23112
rect 15611 23072 16396 23100
rect 15611 23069 15623 23072
rect 15565 23063 15623 23069
rect 16390 23060 16396 23072
rect 16448 23060 16454 23112
rect 8711 23035 8769 23041
rect 8711 23001 8723 23035
rect 8757 23032 8769 23035
rect 10962 23032 10968 23044
rect 8757 23004 10968 23032
rect 8757 23001 8769 23004
rect 8711 22995 8769 23001
rect 10962 22992 10968 23004
rect 11020 22992 11026 23044
rect 14366 22992 14372 23044
rect 14424 23032 14430 23044
rect 16117 23035 16175 23041
rect 16117 23032 16129 23035
rect 14424 23004 16129 23032
rect 14424 22992 14430 23004
rect 16117 23001 16129 23004
rect 16163 23001 16175 23035
rect 16117 22995 16175 23001
rect 1535 22967 1593 22973
rect 1535 22933 1547 22967
rect 1581 22964 1593 22967
rect 12434 22964 12440 22976
rect 1581 22936 12440 22964
rect 1581 22933 1593 22936
rect 1535 22927 1593 22933
rect 12434 22924 12440 22936
rect 12492 22924 12498 22976
rect 12710 22964 12716 22976
rect 12671 22936 12716 22964
rect 12710 22924 12716 22936
rect 12768 22924 12774 22976
rect 14642 22964 14648 22976
rect 14603 22936 14648 22964
rect 14642 22924 14648 22936
rect 14700 22924 14706 22976
rect 17175 22967 17233 22973
rect 17175 22933 17187 22967
rect 17221 22964 17233 22967
rect 17402 22964 17408 22976
rect 17221 22936 17408 22964
rect 17221 22933 17233 22936
rect 17175 22927 17233 22933
rect 17402 22924 17408 22936
rect 17460 22924 17466 22976
rect 21039 22967 21097 22973
rect 21039 22933 21051 22967
rect 21085 22964 21097 22967
rect 21174 22964 21180 22976
rect 21085 22936 21180 22964
rect 21085 22933 21097 22936
rect 21039 22927 21097 22933
rect 21174 22924 21180 22936
rect 21232 22924 21238 22976
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 2222 22760 2228 22772
rect 2183 22732 2228 22760
rect 2222 22720 2228 22732
rect 2280 22720 2286 22772
rect 14090 22760 14096 22772
rect 14051 22732 14096 22760
rect 14090 22720 14096 22732
rect 14148 22720 14154 22772
rect 14458 22760 14464 22772
rect 14419 22732 14464 22760
rect 14458 22720 14464 22732
rect 14516 22720 14522 22772
rect 16390 22760 16396 22772
rect 16351 22732 16396 22760
rect 16390 22720 16396 22732
rect 16448 22720 16454 22772
rect 20990 22760 20996 22772
rect 20951 22732 20996 22760
rect 20990 22720 20996 22732
rect 21048 22720 21054 22772
rect 13262 22624 13268 22636
rect 13223 22596 13268 22624
rect 13262 22584 13268 22596
rect 13320 22584 13326 22636
rect 15473 22627 15531 22633
rect 15473 22593 15485 22627
rect 15519 22624 15531 22627
rect 16761 22627 16819 22633
rect 16761 22624 16773 22627
rect 15519 22596 16773 22624
rect 15519 22593 15531 22596
rect 15473 22587 15531 22593
rect 16761 22593 16773 22596
rect 16807 22624 16819 22627
rect 17083 22627 17141 22633
rect 17083 22624 17095 22627
rect 16807 22596 17095 22624
rect 16807 22593 16819 22596
rect 16761 22587 16819 22593
rect 17083 22593 17095 22596
rect 17129 22593 17141 22627
rect 17083 22587 17141 22593
rect 106 22516 112 22568
rect 164 22556 170 22568
rect 1432 22559 1490 22565
rect 1432 22556 1444 22559
rect 164 22528 1444 22556
rect 164 22516 170 22528
rect 1432 22525 1444 22528
rect 1478 22556 1490 22559
rect 1857 22559 1915 22565
rect 1857 22556 1869 22559
rect 1478 22528 1869 22556
rect 1478 22525 1490 22528
rect 1432 22519 1490 22525
rect 1857 22525 1869 22528
rect 1903 22525 1915 22559
rect 12710 22556 12716 22568
rect 12671 22528 12716 22556
rect 1857 22519 1915 22525
rect 12710 22516 12716 22528
rect 12768 22516 12774 22568
rect 13173 22559 13231 22565
rect 13173 22525 13185 22559
rect 13219 22556 13231 22559
rect 14090 22556 14096 22568
rect 13219 22528 14096 22556
rect 13219 22525 13231 22528
rect 13173 22519 13231 22525
rect 13188 22488 13216 22519
rect 14090 22516 14096 22528
rect 14148 22516 14154 22568
rect 14277 22559 14335 22565
rect 14277 22525 14289 22559
rect 14323 22525 14335 22559
rect 14277 22519 14335 22525
rect 16996 22559 17054 22565
rect 16996 22525 17008 22559
rect 17042 22556 17054 22559
rect 17310 22556 17316 22568
rect 17042 22528 17316 22556
rect 17042 22525 17054 22528
rect 16996 22519 17054 22525
rect 12268 22460 13216 22488
rect 12268 22432 12296 22460
rect 1535 22423 1593 22429
rect 1535 22389 1547 22423
rect 1581 22420 1593 22423
rect 1762 22420 1768 22432
rect 1581 22392 1768 22420
rect 1581 22389 1593 22392
rect 1535 22383 1593 22389
rect 1762 22380 1768 22392
rect 1820 22380 1826 22432
rect 8478 22380 8484 22432
rect 8536 22420 8542 22432
rect 8573 22423 8631 22429
rect 8573 22420 8585 22423
rect 8536 22392 8585 22420
rect 8536 22380 8542 22392
rect 8573 22389 8585 22392
rect 8619 22389 8631 22423
rect 12250 22420 12256 22432
rect 12211 22392 12256 22420
rect 8573 22383 8631 22389
rect 12250 22380 12256 22392
rect 12308 22380 12314 22432
rect 13630 22380 13636 22432
rect 13688 22420 13694 22432
rect 13725 22423 13783 22429
rect 13725 22420 13737 22423
rect 13688 22392 13737 22420
rect 13688 22380 13694 22392
rect 13725 22389 13737 22392
rect 13771 22389 13783 22423
rect 14292 22420 14320 22519
rect 17310 22516 17316 22528
rect 17368 22556 17374 22568
rect 17405 22559 17463 22565
rect 17405 22556 17417 22559
rect 17368 22528 17417 22556
rect 17368 22516 17374 22528
rect 17405 22525 17417 22528
rect 17451 22556 17463 22559
rect 17773 22559 17831 22565
rect 17773 22556 17785 22559
rect 17451 22528 17785 22556
rect 17451 22525 17463 22528
rect 17405 22519 17463 22525
rect 17773 22525 17785 22528
rect 17819 22525 17831 22559
rect 17773 22519 17831 22525
rect 18084 22559 18142 22565
rect 18084 22525 18096 22559
rect 18130 22525 18142 22559
rect 18084 22519 18142 22525
rect 14458 22448 14464 22500
rect 14516 22488 14522 22500
rect 14921 22491 14979 22497
rect 14921 22488 14933 22491
rect 14516 22460 14933 22488
rect 14516 22448 14522 22460
rect 14921 22457 14933 22460
rect 14967 22488 14979 22491
rect 15289 22491 15347 22497
rect 15289 22488 15301 22491
rect 14967 22460 15301 22488
rect 14967 22457 14979 22460
rect 14921 22451 14979 22457
rect 15289 22457 15301 22460
rect 15335 22488 15347 22491
rect 15565 22491 15623 22497
rect 15565 22488 15577 22491
rect 15335 22460 15577 22488
rect 15335 22457 15347 22460
rect 15289 22451 15347 22457
rect 15565 22457 15577 22460
rect 15611 22488 15623 22491
rect 15654 22488 15660 22500
rect 15611 22460 15660 22488
rect 15611 22457 15623 22460
rect 15565 22451 15623 22457
rect 15654 22448 15660 22460
rect 15712 22448 15718 22500
rect 16114 22488 16120 22500
rect 16075 22460 16120 22488
rect 16114 22448 16120 22460
rect 16172 22448 16178 22500
rect 18099 22488 18127 22519
rect 18509 22491 18567 22497
rect 18509 22488 18521 22491
rect 18099 22460 18521 22488
rect 14642 22420 14648 22432
rect 14292 22392 14648 22420
rect 13725 22383 13783 22389
rect 14642 22380 14648 22392
rect 14700 22420 14706 22432
rect 15378 22420 15384 22432
rect 14700 22392 15384 22420
rect 14700 22380 14706 22392
rect 15378 22380 15384 22392
rect 15436 22380 15442 22432
rect 16942 22380 16948 22432
rect 17000 22420 17006 22432
rect 17770 22420 17776 22432
rect 17000 22392 17776 22420
rect 17000 22380 17006 22392
rect 17770 22380 17776 22392
rect 17828 22420 17834 22432
rect 18099 22420 18127 22460
rect 18509 22457 18521 22460
rect 18555 22457 18567 22491
rect 18509 22451 18567 22457
rect 17828 22392 18127 22420
rect 18187 22423 18245 22429
rect 17828 22380 17834 22392
rect 18187 22389 18199 22423
rect 18233 22420 18245 22423
rect 18414 22420 18420 22432
rect 18233 22392 18420 22420
rect 18233 22389 18245 22392
rect 18187 22383 18245 22389
rect 18414 22380 18420 22392
rect 18472 22380 18478 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 12434 22176 12440 22228
rect 12492 22216 12498 22228
rect 13449 22219 13507 22225
rect 13449 22216 13461 22219
rect 12492 22188 13461 22216
rect 12492 22176 12498 22188
rect 13449 22185 13461 22188
rect 13495 22216 13507 22219
rect 13495 22188 13768 22216
rect 13495 22185 13507 22188
rect 13449 22179 13507 22185
rect 13740 22157 13768 22188
rect 13725 22151 13783 22157
rect 13725 22117 13737 22151
rect 13771 22117 13783 22151
rect 13725 22111 13783 22117
rect 13814 22108 13820 22160
rect 13872 22148 13878 22160
rect 15565 22151 15623 22157
rect 15565 22148 15577 22151
rect 13872 22120 15577 22148
rect 13872 22108 13878 22120
rect 15565 22117 15577 22120
rect 15611 22117 15623 22151
rect 15565 22111 15623 22117
rect 17402 22108 17408 22160
rect 17460 22148 17466 22160
rect 18417 22151 18475 22157
rect 18417 22148 18429 22151
rect 17460 22120 18429 22148
rect 17460 22108 17466 22120
rect 18417 22117 18429 22120
rect 18463 22117 18475 22151
rect 18417 22111 18475 22117
rect 18506 22108 18512 22160
rect 18564 22148 18570 22160
rect 18564 22120 18609 22148
rect 18564 22108 18570 22120
rect 12158 22040 12164 22092
rect 12216 22080 12222 22092
rect 12656 22083 12714 22089
rect 12656 22080 12668 22083
rect 12216 22052 12668 22080
rect 12216 22040 12222 22052
rect 12656 22049 12668 22052
rect 12702 22049 12714 22083
rect 12656 22043 12714 22049
rect 14366 22040 14372 22092
rect 14424 22080 14430 22092
rect 16942 22080 16948 22092
rect 14424 22052 14469 22080
rect 16903 22052 16948 22080
rect 14424 22040 14430 22052
rect 16942 22040 16948 22052
rect 17000 22040 17006 22092
rect 15473 22015 15531 22021
rect 15473 21981 15485 22015
rect 15519 21981 15531 22015
rect 16114 22012 16120 22024
rect 16027 21984 16120 22012
rect 15473 21975 15531 21981
rect 15286 21904 15292 21956
rect 15344 21944 15350 21956
rect 15488 21944 15516 21975
rect 16114 21972 16120 21984
rect 16172 22012 16178 22024
rect 16666 22012 16672 22024
rect 16172 21984 16672 22012
rect 16172 21972 16178 21984
rect 16666 21972 16672 21984
rect 16724 21972 16730 22024
rect 19058 22012 19064 22024
rect 19019 21984 19064 22012
rect 19058 21972 19064 21984
rect 19116 21972 19122 22024
rect 17083 21947 17141 21953
rect 17083 21944 17095 21947
rect 15344 21916 17095 21944
rect 15344 21904 15350 21916
rect 17083 21913 17095 21916
rect 17129 21913 17141 21947
rect 17083 21907 17141 21913
rect 12759 21879 12817 21885
rect 12759 21845 12771 21879
rect 12805 21876 12817 21879
rect 13170 21876 13176 21888
rect 12805 21848 13176 21876
rect 12805 21845 12817 21848
rect 12759 21839 12817 21845
rect 13170 21836 13176 21848
rect 13228 21836 13234 21888
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 12158 21672 12164 21684
rect 12119 21644 12164 21672
rect 12158 21632 12164 21644
rect 12216 21632 12222 21684
rect 16942 21672 16948 21684
rect 16903 21644 16948 21672
rect 16942 21632 16948 21644
rect 17000 21632 17006 21684
rect 17402 21672 17408 21684
rect 17363 21644 17408 21672
rect 17402 21632 17408 21644
rect 17460 21632 17466 21684
rect 24762 21672 24768 21684
rect 24723 21644 24768 21672
rect 24762 21632 24768 21644
rect 24820 21632 24826 21684
rect 14461 21539 14519 21545
rect 14461 21505 14473 21539
rect 14507 21536 14519 21539
rect 14642 21536 14648 21548
rect 14507 21508 14648 21536
rect 14507 21505 14519 21508
rect 14461 21499 14519 21505
rect 14642 21496 14648 21508
rect 14700 21496 14706 21548
rect 16025 21539 16083 21545
rect 16025 21505 16037 21539
rect 16071 21536 16083 21539
rect 16390 21536 16396 21548
rect 16071 21508 16396 21536
rect 16071 21505 16083 21508
rect 16025 21499 16083 21505
rect 16390 21496 16396 21508
rect 16448 21496 16454 21548
rect 18414 21496 18420 21548
rect 18472 21536 18478 21548
rect 18601 21539 18659 21545
rect 18601 21536 18613 21539
rect 18472 21508 18613 21536
rect 18472 21496 18478 21508
rect 18601 21505 18613 21508
rect 18647 21536 18659 21539
rect 19521 21539 19579 21545
rect 19521 21536 19533 21539
rect 18647 21508 19533 21536
rect 18647 21505 18659 21508
rect 18601 21499 18659 21505
rect 19521 21505 19533 21508
rect 19567 21505 19579 21539
rect 19521 21499 19579 21505
rect 12618 21468 12624 21480
rect 12579 21440 12624 21468
rect 12618 21428 12624 21440
rect 12676 21428 12682 21480
rect 12894 21428 12900 21480
rect 12952 21468 12958 21480
rect 13081 21471 13139 21477
rect 13081 21468 13093 21471
rect 12952 21440 13093 21468
rect 12952 21428 12958 21440
rect 13081 21437 13093 21440
rect 13127 21437 13139 21471
rect 13081 21431 13139 21437
rect 23842 21428 23848 21480
rect 23900 21468 23906 21480
rect 24581 21471 24639 21477
rect 24581 21468 24593 21471
rect 23900 21440 24593 21468
rect 23900 21428 23906 21440
rect 24581 21437 24593 21440
rect 24627 21468 24639 21471
rect 25133 21471 25191 21477
rect 25133 21468 25145 21471
rect 24627 21440 25145 21468
rect 24627 21437 24639 21440
rect 24581 21431 24639 21437
rect 25133 21437 25145 21440
rect 25179 21437 25191 21471
rect 25133 21431 25191 21437
rect 11885 21403 11943 21409
rect 11885 21369 11897 21403
rect 11931 21400 11943 21403
rect 12250 21400 12256 21412
rect 11931 21372 12256 21400
rect 11931 21369 11943 21372
rect 11885 21363 11943 21369
rect 12250 21360 12256 21372
rect 12308 21400 12314 21412
rect 12912 21400 12940 21428
rect 13354 21400 13360 21412
rect 12308 21372 12940 21400
rect 13315 21372 13360 21400
rect 12308 21360 12314 21372
rect 13354 21360 13360 21372
rect 13412 21360 13418 21412
rect 14553 21403 14611 21409
rect 14553 21369 14565 21403
rect 14599 21369 14611 21403
rect 14553 21363 14611 21369
rect 15105 21403 15163 21409
rect 15105 21369 15117 21403
rect 15151 21400 15163 21403
rect 15194 21400 15200 21412
rect 15151 21372 15200 21400
rect 15151 21369 15163 21372
rect 15105 21363 15163 21369
rect 13725 21335 13783 21341
rect 13725 21301 13737 21335
rect 13771 21332 13783 21335
rect 13814 21332 13820 21344
rect 13771 21304 13820 21332
rect 13771 21301 13783 21304
rect 13725 21295 13783 21301
rect 13814 21292 13820 21304
rect 13872 21332 13878 21344
rect 14182 21332 14188 21344
rect 13872 21304 14188 21332
rect 13872 21292 13878 21304
rect 14182 21292 14188 21304
rect 14240 21332 14246 21344
rect 14568 21332 14596 21363
rect 15194 21360 15200 21372
rect 15252 21360 15258 21412
rect 16117 21403 16175 21409
rect 16117 21400 16129 21403
rect 15764 21372 16129 21400
rect 15381 21335 15439 21341
rect 15381 21332 15393 21335
rect 14240 21304 15393 21332
rect 14240 21292 14246 21304
rect 15381 21301 15393 21304
rect 15427 21301 15439 21335
rect 15381 21295 15439 21301
rect 15470 21292 15476 21344
rect 15528 21332 15534 21344
rect 15764 21341 15792 21372
rect 16117 21369 16129 21372
rect 16163 21369 16175 21403
rect 16666 21400 16672 21412
rect 16627 21372 16672 21400
rect 16117 21363 16175 21369
rect 16666 21360 16672 21372
rect 16724 21360 16730 21412
rect 18417 21403 18475 21409
rect 18417 21369 18429 21403
rect 18463 21400 18475 21403
rect 18693 21403 18751 21409
rect 18693 21400 18705 21403
rect 18463 21372 18705 21400
rect 18463 21369 18475 21372
rect 18417 21363 18475 21369
rect 18693 21369 18705 21372
rect 18739 21400 18751 21403
rect 18966 21400 18972 21412
rect 18739 21372 18972 21400
rect 18739 21369 18751 21372
rect 18693 21363 18751 21369
rect 18966 21360 18972 21372
rect 19024 21360 19030 21412
rect 19242 21400 19248 21412
rect 19203 21372 19248 21400
rect 19242 21360 19248 21372
rect 19300 21360 19306 21412
rect 15749 21335 15807 21341
rect 15749 21332 15761 21335
rect 15528 21304 15761 21332
rect 15528 21292 15534 21304
rect 15749 21301 15761 21304
rect 15795 21301 15807 21335
rect 17862 21332 17868 21344
rect 17823 21304 17868 21332
rect 15749 21295 15807 21301
rect 17862 21292 17868 21304
rect 17920 21292 17926 21344
rect 19426 21292 19432 21344
rect 19484 21332 19490 21344
rect 20346 21332 20352 21344
rect 19484 21304 20352 21332
rect 19484 21292 19490 21304
rect 20346 21292 20352 21304
rect 20404 21292 20410 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 13265 21131 13323 21137
rect 13265 21097 13277 21131
rect 13311 21128 13323 21131
rect 13354 21128 13360 21140
rect 13311 21100 13360 21128
rect 13311 21097 13323 21100
rect 13265 21091 13323 21097
rect 13354 21088 13360 21100
rect 13412 21088 13418 21140
rect 15105 21131 15163 21137
rect 15105 21097 15117 21131
rect 15151 21128 15163 21131
rect 15286 21128 15292 21140
rect 15151 21100 15292 21128
rect 15151 21097 15163 21100
rect 15105 21091 15163 21097
rect 15286 21088 15292 21100
rect 15344 21088 15350 21140
rect 15378 21088 15384 21140
rect 15436 21128 15442 21140
rect 16991 21131 17049 21137
rect 16991 21128 17003 21131
rect 15436 21100 17003 21128
rect 15436 21088 15442 21100
rect 16991 21097 17003 21100
rect 17037 21097 17049 21131
rect 16991 21091 17049 21097
rect 1210 21020 1216 21072
rect 1268 21060 1274 21072
rect 11514 21060 11520 21072
rect 1268 21032 1507 21060
rect 11475 21032 11520 21060
rect 1268 21020 1274 21032
rect 1479 21001 1507 21032
rect 11514 21020 11520 21032
rect 11572 21020 11578 21072
rect 13170 21020 13176 21072
rect 13228 21060 13234 21072
rect 13722 21060 13728 21072
rect 13228 21032 13728 21060
rect 13228 21020 13234 21032
rect 13722 21020 13728 21032
rect 13780 21020 13786 21072
rect 13817 21063 13875 21069
rect 13817 21029 13829 21063
rect 13863 21060 13875 21063
rect 14458 21060 14464 21072
rect 13863 21032 14464 21060
rect 13863 21029 13875 21032
rect 13817 21023 13875 21029
rect 14458 21020 14464 21032
rect 14516 21020 14522 21072
rect 15470 21060 15476 21072
rect 15431 21032 15476 21060
rect 15470 21020 15476 21032
rect 15528 21020 15534 21072
rect 17862 21020 17868 21072
rect 17920 21060 17926 21072
rect 18506 21060 18512 21072
rect 17920 21032 18512 21060
rect 17920 21020 17926 21032
rect 18506 21020 18512 21032
rect 18564 21020 18570 21072
rect 19061 21063 19119 21069
rect 19061 21029 19073 21063
rect 19107 21060 19119 21063
rect 19242 21060 19248 21072
rect 19107 21032 19248 21060
rect 19107 21029 19119 21032
rect 19061 21023 19119 21029
rect 19242 21020 19248 21032
rect 19300 21060 19306 21072
rect 20070 21060 20076 21072
rect 19300 21032 20076 21060
rect 19300 21020 19306 21032
rect 20070 21020 20076 21032
rect 20128 21020 20134 21072
rect 1464 20995 1522 21001
rect 1464 20961 1476 20995
rect 1510 20961 1522 20995
rect 1464 20955 1522 20961
rect 9582 20952 9588 21004
rect 9640 20992 9646 21004
rect 9712 20995 9770 21001
rect 9712 20992 9724 20995
rect 9640 20964 9724 20992
rect 9640 20952 9646 20964
rect 9712 20961 9724 20964
rect 9758 20961 9770 20995
rect 9712 20955 9770 20961
rect 16920 20995 16978 21001
rect 16920 20961 16932 20995
rect 16966 20992 16978 20995
rect 17402 20992 17408 21004
rect 16966 20964 17408 20992
rect 16966 20961 16978 20964
rect 16920 20955 16978 20961
rect 17402 20952 17408 20964
rect 17460 20952 17466 21004
rect 24670 21001 24676 21004
rect 24648 20995 24676 21001
rect 24648 20992 24660 20995
rect 24583 20964 24660 20992
rect 24648 20961 24660 20964
rect 24728 20992 24734 21004
rect 25130 20992 25136 21004
rect 24728 20964 25136 20992
rect 24648 20955 24676 20961
rect 24670 20952 24676 20955
rect 24728 20952 24734 20964
rect 25130 20952 25136 20964
rect 25188 20952 25194 21004
rect 8294 20924 8300 20936
rect 8255 20896 8300 20924
rect 8294 20884 8300 20896
rect 8352 20884 8358 20936
rect 10042 20884 10048 20936
rect 10100 20924 10106 20936
rect 11054 20924 11060 20936
rect 10100 20896 11060 20924
rect 10100 20884 10106 20896
rect 11054 20884 11060 20896
rect 11112 20884 11118 20936
rect 11425 20927 11483 20933
rect 11425 20893 11437 20927
rect 11471 20924 11483 20927
rect 11790 20924 11796 20936
rect 11471 20896 11796 20924
rect 11471 20893 11483 20896
rect 11425 20887 11483 20893
rect 11790 20884 11796 20896
rect 11848 20884 11854 20936
rect 12069 20927 12127 20933
rect 12069 20893 12081 20927
rect 12115 20924 12127 20927
rect 12802 20924 12808 20936
rect 12115 20896 12808 20924
rect 12115 20893 12127 20896
rect 12069 20887 12127 20893
rect 12802 20884 12808 20896
rect 12860 20884 12866 20936
rect 15378 20924 15384 20936
rect 15339 20896 15384 20924
rect 15378 20884 15384 20896
rect 15436 20884 15442 20936
rect 15657 20927 15715 20933
rect 15657 20893 15669 20927
rect 15703 20893 15715 20927
rect 15657 20887 15715 20893
rect 14277 20859 14335 20865
rect 14277 20825 14289 20859
rect 14323 20856 14335 20859
rect 15286 20856 15292 20868
rect 14323 20828 15292 20856
rect 14323 20825 14335 20828
rect 14277 20819 14335 20825
rect 15286 20816 15292 20828
rect 15344 20856 15350 20868
rect 15672 20856 15700 20887
rect 17770 20884 17776 20936
rect 17828 20924 17834 20936
rect 18417 20927 18475 20933
rect 18417 20924 18429 20927
rect 17828 20896 18429 20924
rect 17828 20884 17834 20896
rect 18417 20893 18429 20896
rect 18463 20893 18475 20927
rect 18417 20887 18475 20893
rect 15344 20828 15700 20856
rect 15344 20816 15350 20828
rect 18046 20816 18052 20868
rect 18104 20856 18110 20868
rect 19978 20856 19984 20868
rect 18104 20828 19984 20856
rect 18104 20816 18110 20828
rect 19978 20816 19984 20828
rect 20036 20816 20042 20868
rect 1535 20791 1593 20797
rect 1535 20757 1547 20791
rect 1581 20788 1593 20791
rect 7650 20788 7656 20800
rect 1581 20760 7656 20788
rect 1581 20757 1593 20760
rect 1535 20751 1593 20757
rect 7650 20748 7656 20760
rect 7708 20748 7714 20800
rect 8846 20788 8852 20800
rect 8807 20760 8852 20788
rect 8846 20748 8852 20760
rect 8904 20748 8910 20800
rect 9815 20791 9873 20797
rect 9815 20757 9827 20791
rect 9861 20788 9873 20791
rect 10042 20788 10048 20800
rect 9861 20760 10048 20788
rect 9861 20757 9873 20760
rect 9815 20751 9873 20757
rect 10042 20748 10048 20760
rect 10100 20748 10106 20800
rect 10318 20788 10324 20800
rect 10279 20760 10324 20788
rect 10318 20748 10324 20760
rect 10376 20748 10382 20800
rect 11606 20748 11612 20800
rect 11664 20788 11670 20800
rect 12618 20788 12624 20800
rect 11664 20760 12624 20788
rect 11664 20748 11670 20760
rect 12618 20748 12624 20760
rect 12676 20748 12682 20800
rect 14642 20788 14648 20800
rect 14603 20760 14648 20788
rect 14642 20748 14648 20760
rect 14700 20748 14706 20800
rect 16390 20788 16396 20800
rect 16351 20760 16396 20788
rect 16390 20748 16396 20760
rect 16448 20748 16454 20800
rect 18598 20748 18604 20800
rect 18656 20788 18662 20800
rect 24719 20791 24777 20797
rect 24719 20788 24731 20791
rect 18656 20760 24731 20788
rect 18656 20748 18662 20760
rect 24719 20757 24731 20760
rect 24765 20757 24777 20791
rect 24719 20751 24777 20757
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 1210 20544 1216 20596
rect 1268 20584 1274 20596
rect 1581 20587 1639 20593
rect 1581 20584 1593 20587
rect 1268 20556 1593 20584
rect 1268 20544 1274 20556
rect 1581 20553 1593 20556
rect 1627 20553 1639 20587
rect 4062 20584 4068 20596
rect 4023 20556 4068 20584
rect 1581 20547 1639 20553
rect 4062 20544 4068 20556
rect 4120 20544 4126 20596
rect 11425 20587 11483 20593
rect 11425 20553 11437 20587
rect 11471 20584 11483 20587
rect 11514 20584 11520 20596
rect 11471 20556 11520 20584
rect 11471 20553 11483 20556
rect 11425 20547 11483 20553
rect 11514 20544 11520 20556
rect 11572 20544 11578 20596
rect 13722 20544 13728 20596
rect 13780 20584 13786 20596
rect 14737 20587 14795 20593
rect 14737 20584 14749 20587
rect 13780 20556 14749 20584
rect 13780 20544 13786 20556
rect 14737 20553 14749 20556
rect 14783 20553 14795 20587
rect 15378 20584 15384 20596
rect 14737 20547 14795 20553
rect 14936 20556 15384 20584
rect 10137 20519 10195 20525
rect 10137 20485 10149 20519
rect 10183 20516 10195 20519
rect 10226 20516 10232 20528
rect 10183 20488 10232 20516
rect 10183 20485 10195 20488
rect 10137 20479 10195 20485
rect 10226 20476 10232 20488
rect 10284 20516 10290 20528
rect 12710 20516 12716 20528
rect 10284 20488 12716 20516
rect 10284 20476 10290 20488
rect 12710 20476 12716 20488
rect 12768 20516 12774 20528
rect 13538 20516 13544 20528
rect 12768 20488 13544 20516
rect 12768 20476 12774 20488
rect 13538 20476 13544 20488
rect 13596 20476 13602 20528
rect 14093 20519 14151 20525
rect 14093 20485 14105 20519
rect 14139 20516 14151 20519
rect 14458 20516 14464 20528
rect 14139 20488 14464 20516
rect 14139 20485 14151 20488
rect 14093 20479 14151 20485
rect 14458 20476 14464 20488
rect 14516 20476 14522 20528
rect 4154 20448 4160 20460
rect 3896 20420 4160 20448
rect 3896 20389 3924 20420
rect 4154 20408 4160 20420
rect 4212 20448 4218 20460
rect 4433 20451 4491 20457
rect 4433 20448 4445 20451
rect 4212 20420 4445 20448
rect 4212 20408 4218 20420
rect 4433 20417 4445 20420
rect 4479 20417 4491 20451
rect 4433 20411 4491 20417
rect 7834 20408 7840 20460
rect 7892 20408 7898 20460
rect 11606 20448 11612 20460
rect 8680 20420 11612 20448
rect 3881 20383 3939 20389
rect 3881 20349 3893 20383
rect 3927 20349 3939 20383
rect 3881 20343 3939 20349
rect 6362 20340 6368 20392
rect 6420 20380 6426 20392
rect 7688 20383 7746 20389
rect 7688 20380 7700 20383
rect 6420 20352 7700 20380
rect 6420 20340 6426 20352
rect 7688 20349 7700 20352
rect 7734 20380 7746 20383
rect 7852 20380 7880 20408
rect 8680 20389 8708 20420
rect 11606 20408 11612 20420
rect 11664 20408 11670 20460
rect 11790 20448 11796 20460
rect 11751 20420 11796 20448
rect 11790 20408 11796 20420
rect 11848 20408 11854 20460
rect 13173 20451 13231 20457
rect 13173 20417 13185 20451
rect 13219 20448 13231 20451
rect 13354 20448 13360 20460
rect 13219 20420 13360 20448
rect 13219 20417 13231 20420
rect 13173 20411 13231 20417
rect 13354 20408 13360 20420
rect 13412 20408 13418 20460
rect 14936 20457 14964 20556
rect 15378 20544 15384 20556
rect 15436 20544 15442 20596
rect 17770 20584 17776 20596
rect 17731 20556 17776 20584
rect 17770 20544 17776 20556
rect 17828 20544 17834 20596
rect 18506 20544 18512 20596
rect 18564 20584 18570 20596
rect 18785 20587 18843 20593
rect 18785 20584 18797 20587
rect 18564 20556 18797 20584
rect 18564 20544 18570 20556
rect 18785 20553 18797 20556
rect 18831 20553 18843 20587
rect 24670 20584 24676 20596
rect 24631 20556 24676 20584
rect 18785 20547 18843 20553
rect 24670 20544 24676 20556
rect 24728 20544 24734 20596
rect 19981 20519 20039 20525
rect 19981 20485 19993 20519
rect 20027 20516 20039 20519
rect 20530 20516 20536 20528
rect 20027 20488 20536 20516
rect 20027 20485 20039 20488
rect 19981 20479 20039 20485
rect 20530 20476 20536 20488
rect 20588 20516 20594 20528
rect 21545 20519 21603 20525
rect 21545 20516 21557 20519
rect 20588 20488 21557 20516
rect 20588 20476 20594 20488
rect 21545 20485 21557 20488
rect 21591 20485 21603 20519
rect 21545 20479 21603 20485
rect 14921 20451 14979 20457
rect 14921 20417 14933 20451
rect 14967 20417 14979 20451
rect 14921 20411 14979 20417
rect 20441 20451 20499 20457
rect 20441 20417 20453 20451
rect 20487 20448 20499 20451
rect 20993 20451 21051 20457
rect 20993 20448 21005 20451
rect 20487 20420 21005 20448
rect 20487 20417 20499 20420
rect 20441 20411 20499 20417
rect 20993 20417 21005 20420
rect 21039 20448 21051 20451
rect 21174 20448 21180 20460
rect 21039 20420 21180 20448
rect 21039 20417 21051 20420
rect 20993 20411 21051 20417
rect 21174 20408 21180 20420
rect 21232 20408 21238 20460
rect 8113 20383 8171 20389
rect 8113 20380 8125 20383
rect 7734 20352 8125 20380
rect 7734 20349 7746 20352
rect 7688 20343 7746 20349
rect 8113 20349 8125 20352
rect 8159 20349 8171 20383
rect 8113 20343 8171 20349
rect 8573 20383 8631 20389
rect 8573 20349 8585 20383
rect 8619 20380 8631 20383
rect 8665 20383 8723 20389
rect 8665 20380 8677 20383
rect 8619 20352 8677 20380
rect 8619 20349 8631 20352
rect 8573 20343 8631 20349
rect 8665 20349 8677 20352
rect 8711 20349 8723 20383
rect 8665 20343 8723 20349
rect 8846 20340 8852 20392
rect 8904 20380 8910 20392
rect 9217 20383 9275 20389
rect 9217 20380 9229 20383
rect 8904 20352 9229 20380
rect 8904 20340 8910 20352
rect 9217 20349 9229 20352
rect 9263 20380 9275 20383
rect 10226 20380 10232 20392
rect 9263 20352 9996 20380
rect 10187 20352 10232 20380
rect 9263 20349 9275 20352
rect 9217 20343 9275 20349
rect 7791 20315 7849 20321
rect 7791 20281 7803 20315
rect 7837 20312 7849 20315
rect 9766 20312 9772 20324
rect 7837 20284 9772 20312
rect 7837 20281 7849 20284
rect 7791 20275 7849 20281
rect 9766 20272 9772 20284
rect 9824 20272 9830 20324
rect 9968 20312 9996 20352
rect 10226 20340 10232 20352
rect 10284 20340 10290 20392
rect 10318 20340 10324 20392
rect 10376 20380 10382 20392
rect 10781 20383 10839 20389
rect 10781 20380 10793 20383
rect 10376 20352 10793 20380
rect 10376 20340 10382 20352
rect 10781 20349 10793 20352
rect 10827 20380 10839 20383
rect 11238 20380 11244 20392
rect 10827 20352 11244 20380
rect 10827 20349 10839 20352
rect 10781 20343 10839 20349
rect 11238 20340 11244 20352
rect 11296 20340 11302 20392
rect 12618 20340 12624 20392
rect 12676 20380 12682 20392
rect 16298 20380 16304 20392
rect 12676 20352 16304 20380
rect 12676 20340 12682 20352
rect 16298 20340 16304 20352
rect 16356 20340 16362 20392
rect 17129 20383 17187 20389
rect 17129 20349 17141 20383
rect 17175 20380 17187 20383
rect 19058 20380 19064 20392
rect 17175 20352 19064 20380
rect 17175 20349 17187 20352
rect 17129 20343 17187 20349
rect 19058 20340 19064 20352
rect 19116 20340 19122 20392
rect 10336 20312 10364 20340
rect 9968 20284 10364 20312
rect 13535 20315 13593 20321
rect 13535 20281 13547 20315
rect 13581 20312 13593 20315
rect 13722 20312 13728 20324
rect 13581 20284 13728 20312
rect 13581 20281 13593 20284
rect 13535 20275 13593 20281
rect 13722 20272 13728 20284
rect 13780 20272 13786 20324
rect 16482 20312 16488 20324
rect 16443 20284 16488 20312
rect 16482 20272 16488 20284
rect 16540 20272 16546 20324
rect 16577 20315 16635 20321
rect 16577 20281 16589 20315
rect 16623 20281 16635 20315
rect 16577 20275 16635 20281
rect 18325 20315 18383 20321
rect 18325 20281 18337 20315
rect 18371 20312 18383 20315
rect 19153 20315 19211 20321
rect 19153 20312 19165 20315
rect 18371 20284 19165 20312
rect 18371 20281 18383 20284
rect 18325 20275 18383 20281
rect 19153 20281 19165 20284
rect 19199 20312 19211 20315
rect 19429 20315 19487 20321
rect 19429 20312 19441 20315
rect 19199 20284 19441 20312
rect 19199 20281 19211 20284
rect 19153 20275 19211 20281
rect 19429 20281 19441 20284
rect 19475 20281 19487 20315
rect 19429 20275 19487 20281
rect 8938 20244 8944 20256
rect 8899 20216 8944 20244
rect 8938 20204 8944 20216
rect 8996 20204 9002 20256
rect 9582 20204 9588 20256
rect 9640 20244 9646 20256
rect 9677 20247 9735 20253
rect 9677 20244 9689 20247
rect 9640 20216 9689 20244
rect 9640 20204 9646 20216
rect 9677 20213 9689 20216
rect 9723 20213 9735 20247
rect 9677 20207 9735 20213
rect 10134 20204 10140 20256
rect 10192 20244 10198 20256
rect 10321 20247 10379 20253
rect 10321 20244 10333 20247
rect 10192 20216 10333 20244
rect 10192 20204 10198 20216
rect 10321 20213 10333 20216
rect 10367 20213 10379 20247
rect 10321 20207 10379 20213
rect 10870 20204 10876 20256
rect 10928 20244 10934 20256
rect 12989 20247 13047 20253
rect 12989 20244 13001 20247
rect 10928 20216 13001 20244
rect 10928 20204 10934 20216
rect 12989 20213 13001 20216
rect 13035 20244 13047 20247
rect 13354 20244 13360 20256
rect 13035 20216 13360 20244
rect 13035 20213 13047 20216
rect 12989 20207 13047 20213
rect 13354 20204 13360 20216
rect 13412 20204 13418 20256
rect 15470 20204 15476 20256
rect 15528 20244 15534 20256
rect 15749 20247 15807 20253
rect 15749 20244 15761 20247
rect 15528 20216 15761 20244
rect 15528 20204 15534 20216
rect 15749 20213 15761 20216
rect 15795 20213 15807 20247
rect 15749 20207 15807 20213
rect 16301 20247 16359 20253
rect 16301 20213 16313 20247
rect 16347 20244 16359 20247
rect 16592 20244 16620 20275
rect 19518 20272 19524 20324
rect 19576 20312 19582 20324
rect 21085 20315 21143 20321
rect 19576 20284 19621 20312
rect 19576 20272 19582 20284
rect 21085 20281 21097 20315
rect 21131 20281 21143 20315
rect 21085 20275 21143 20281
rect 17218 20244 17224 20256
rect 16347 20216 17224 20244
rect 16347 20213 16359 20216
rect 16301 20207 16359 20213
rect 17218 20204 17224 20216
rect 17276 20204 17282 20256
rect 17402 20244 17408 20256
rect 17363 20216 17408 20244
rect 17402 20204 17408 20216
rect 17460 20204 17466 20256
rect 19978 20204 19984 20256
rect 20036 20244 20042 20256
rect 20717 20247 20775 20253
rect 20717 20244 20729 20247
rect 20036 20216 20729 20244
rect 20036 20204 20042 20216
rect 20717 20213 20729 20216
rect 20763 20244 20775 20247
rect 21100 20244 21128 20275
rect 20763 20216 21128 20244
rect 20763 20213 20775 20216
rect 20717 20207 20775 20213
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 7650 20000 7656 20052
rect 7708 20040 7714 20052
rect 7745 20043 7803 20049
rect 7745 20040 7757 20043
rect 7708 20012 7757 20040
rect 7708 20000 7714 20012
rect 7745 20009 7757 20012
rect 7791 20009 7803 20043
rect 7745 20003 7803 20009
rect 4338 19932 4344 19984
rect 4396 19972 4402 19984
rect 4801 19975 4859 19981
rect 4801 19972 4813 19975
rect 4396 19944 4813 19972
rect 4396 19932 4402 19944
rect 4801 19941 4813 19944
rect 4847 19941 4859 19975
rect 7760 19972 7788 20003
rect 7834 20000 7840 20052
rect 7892 20040 7898 20052
rect 8846 20040 8852 20052
rect 7892 20012 8852 20040
rect 7892 20000 7898 20012
rect 8846 20000 8852 20012
rect 8904 20000 8910 20052
rect 14182 20040 14188 20052
rect 14143 20012 14188 20040
rect 14182 20000 14188 20012
rect 14240 20000 14246 20052
rect 14274 20000 14280 20052
rect 14332 20040 14338 20052
rect 14461 20043 14519 20049
rect 14461 20040 14473 20043
rect 14332 20012 14473 20040
rect 14332 20000 14338 20012
rect 14461 20009 14473 20012
rect 14507 20009 14519 20043
rect 14461 20003 14519 20009
rect 16390 20000 16396 20052
rect 16448 20040 16454 20052
rect 16991 20043 17049 20049
rect 16991 20040 17003 20043
rect 16448 20012 17003 20040
rect 16448 20000 16454 20012
rect 16991 20009 17003 20012
rect 17037 20009 17049 20043
rect 18322 20040 18328 20052
rect 18283 20012 18328 20040
rect 16991 20003 17049 20009
rect 18322 20000 18328 20012
rect 18380 20000 18386 20052
rect 18506 20000 18512 20052
rect 18564 20040 18570 20052
rect 18877 20043 18935 20049
rect 18877 20040 18889 20043
rect 18564 20012 18889 20040
rect 18564 20000 18570 20012
rect 18877 20009 18889 20012
rect 18923 20040 18935 20043
rect 19337 20043 19395 20049
rect 19337 20040 19349 20043
rect 18923 20012 19349 20040
rect 18923 20009 18935 20012
rect 18877 20003 18935 20009
rect 19337 20009 19349 20012
rect 19383 20040 19395 20043
rect 19518 20040 19524 20052
rect 19383 20012 19524 20040
rect 19383 20009 19395 20012
rect 19337 20003 19395 20009
rect 19518 20000 19524 20012
rect 19576 20000 19582 20052
rect 24762 20040 24768 20052
rect 24723 20012 24768 20040
rect 24762 20000 24768 20012
rect 24820 20000 24826 20052
rect 8021 19975 8079 19981
rect 8021 19972 8033 19975
rect 7760 19944 8033 19972
rect 4801 19935 4859 19941
rect 8021 19941 8033 19944
rect 8067 19941 8079 19975
rect 8021 19935 8079 19941
rect 8110 19932 8116 19984
rect 8168 19972 8174 19984
rect 8168 19944 8213 19972
rect 8168 19932 8174 19944
rect 10226 19932 10232 19984
rect 10284 19972 10290 19984
rect 10366 19975 10424 19981
rect 10366 19972 10378 19975
rect 10284 19944 10378 19972
rect 10284 19932 10290 19944
rect 10366 19941 10378 19944
rect 10412 19941 10424 19975
rect 10366 19935 10424 19941
rect 13354 19932 13360 19984
rect 13412 19972 13418 19984
rect 13586 19975 13644 19981
rect 13586 19972 13598 19975
rect 13412 19944 13598 19972
rect 13412 19932 13418 19944
rect 13586 19941 13598 19944
rect 13632 19972 13644 19975
rect 13722 19972 13728 19984
rect 13632 19944 13728 19972
rect 13632 19941 13644 19944
rect 13586 19935 13644 19941
rect 13722 19932 13728 19944
rect 13780 19932 13786 19984
rect 15473 19975 15531 19981
rect 15473 19941 15485 19975
rect 15519 19972 15531 19975
rect 15746 19972 15752 19984
rect 15519 19944 15752 19972
rect 15519 19941 15531 19944
rect 15473 19935 15531 19941
rect 15746 19932 15752 19944
rect 15804 19932 15810 19984
rect 6181 19907 6239 19913
rect 6181 19873 6193 19907
rect 6227 19904 6239 19907
rect 6270 19904 6276 19916
rect 6227 19876 6276 19904
rect 6227 19873 6239 19876
rect 6181 19867 6239 19873
rect 6270 19864 6276 19876
rect 6328 19864 6334 19916
rect 10045 19907 10103 19913
rect 10045 19873 10057 19907
rect 10091 19904 10103 19907
rect 10134 19904 10140 19916
rect 10091 19876 10140 19904
rect 10091 19873 10103 19876
rect 10045 19867 10103 19873
rect 10134 19864 10140 19876
rect 10192 19864 10198 19916
rect 11793 19907 11851 19913
rect 11793 19873 11805 19907
rect 11839 19904 11851 19907
rect 11882 19904 11888 19916
rect 11839 19876 11888 19904
rect 11839 19873 11851 19876
rect 11793 19867 11851 19873
rect 11882 19864 11888 19876
rect 11940 19864 11946 19916
rect 13262 19904 13268 19916
rect 13223 19876 13268 19904
rect 13262 19864 13268 19876
rect 13320 19864 13326 19916
rect 16920 19907 16978 19913
rect 16920 19873 16932 19907
rect 16966 19904 16978 19907
rect 17126 19904 17132 19916
rect 16966 19876 17132 19904
rect 16966 19873 16978 19876
rect 16920 19867 16978 19873
rect 17126 19864 17132 19876
rect 17184 19864 17190 19916
rect 19426 19864 19432 19916
rect 19484 19904 19490 19916
rect 19740 19907 19798 19913
rect 19740 19904 19752 19907
rect 19484 19876 19752 19904
rect 19484 19864 19490 19876
rect 19740 19873 19752 19876
rect 19786 19873 19798 19907
rect 19740 19867 19798 19873
rect 20809 19907 20867 19913
rect 20809 19873 20821 19907
rect 20855 19904 20867 19907
rect 20990 19904 20996 19916
rect 20855 19876 20996 19904
rect 20855 19873 20867 19876
rect 20809 19867 20867 19873
rect 20990 19864 20996 19876
rect 21048 19864 21054 19916
rect 24581 19907 24639 19913
rect 24581 19873 24593 19907
rect 24627 19904 24639 19907
rect 24670 19904 24676 19916
rect 24627 19876 24676 19904
rect 24627 19873 24639 19876
rect 24581 19867 24639 19873
rect 24670 19864 24676 19876
rect 24728 19864 24734 19916
rect 3970 19796 3976 19848
rect 4028 19836 4034 19848
rect 4709 19839 4767 19845
rect 4709 19836 4721 19839
rect 4028 19808 4721 19836
rect 4028 19796 4034 19808
rect 4709 19805 4721 19808
rect 4755 19805 4767 19839
rect 4709 19799 4767 19805
rect 4985 19839 5043 19845
rect 4985 19805 4997 19839
rect 5031 19805 5043 19839
rect 4985 19799 5043 19805
rect 3878 19728 3884 19780
rect 3936 19768 3942 19780
rect 5000 19768 5028 19799
rect 5442 19796 5448 19848
rect 5500 19836 5506 19848
rect 5994 19836 6000 19848
rect 5500 19808 6000 19836
rect 5500 19796 5506 19808
rect 5994 19796 6000 19808
rect 6052 19796 6058 19848
rect 8665 19839 8723 19845
rect 8665 19805 8677 19839
rect 8711 19836 8723 19839
rect 8846 19836 8852 19848
rect 8711 19808 8852 19836
rect 8711 19805 8723 19808
rect 8665 19799 8723 19805
rect 8846 19796 8852 19808
rect 8904 19796 8910 19848
rect 15381 19839 15439 19845
rect 15381 19805 15393 19839
rect 15427 19805 15439 19839
rect 15381 19799 15439 19805
rect 16025 19839 16083 19845
rect 16025 19805 16037 19839
rect 16071 19836 16083 19839
rect 16390 19836 16396 19848
rect 16071 19808 16396 19836
rect 16071 19805 16083 19808
rect 16025 19799 16083 19805
rect 5350 19768 5356 19780
rect 3936 19740 5356 19768
rect 3936 19728 3942 19740
rect 5350 19728 5356 19740
rect 5408 19728 5414 19780
rect 15286 19728 15292 19780
rect 15344 19768 15350 19780
rect 15396 19768 15424 19799
rect 16390 19796 16396 19808
rect 16448 19836 16454 19848
rect 17402 19836 17408 19848
rect 16448 19808 17408 19836
rect 16448 19796 16454 19808
rect 17402 19796 17408 19808
rect 17460 19796 17466 19848
rect 17954 19836 17960 19848
rect 17915 19808 17960 19836
rect 17954 19796 17960 19808
rect 18012 19796 18018 19848
rect 16482 19768 16488 19780
rect 15344 19740 15424 19768
rect 16395 19740 16488 19768
rect 15344 19728 15350 19740
rect 16482 19728 16488 19740
rect 16540 19768 16546 19780
rect 19843 19771 19901 19777
rect 19843 19768 19855 19771
rect 16540 19740 19855 19768
rect 16540 19728 16546 19740
rect 19843 19737 19855 19740
rect 19889 19737 19901 19771
rect 19843 19731 19901 19737
rect 5074 19660 5080 19712
rect 5132 19700 5138 19712
rect 5629 19703 5687 19709
rect 5629 19700 5641 19703
rect 5132 19672 5641 19700
rect 5132 19660 5138 19672
rect 5629 19669 5641 19672
rect 5675 19669 5687 19703
rect 5629 19663 5687 19669
rect 5994 19660 6000 19712
rect 6052 19700 6058 19712
rect 6319 19703 6377 19709
rect 6319 19700 6331 19703
rect 6052 19672 6331 19700
rect 6052 19660 6058 19672
rect 6319 19669 6331 19672
rect 6365 19669 6377 19703
rect 6319 19663 6377 19669
rect 10965 19703 11023 19709
rect 10965 19669 10977 19703
rect 11011 19700 11023 19703
rect 11146 19700 11152 19712
rect 11011 19672 11152 19700
rect 11011 19669 11023 19672
rect 10965 19663 11023 19669
rect 11146 19660 11152 19672
rect 11204 19660 11210 19712
rect 11330 19700 11336 19712
rect 11291 19672 11336 19700
rect 11330 19660 11336 19672
rect 11388 19660 11394 19712
rect 11931 19703 11989 19709
rect 11931 19669 11943 19703
rect 11977 19700 11989 19703
rect 12437 19703 12495 19709
rect 12437 19700 12449 19703
rect 11977 19672 12449 19700
rect 11977 19669 11989 19672
rect 11931 19663 11989 19669
rect 12437 19669 12449 19672
rect 12483 19700 12495 19703
rect 12526 19700 12532 19712
rect 12483 19672 12532 19700
rect 12483 19669 12495 19672
rect 12437 19663 12495 19669
rect 12526 19660 12532 19672
rect 12584 19660 12590 19712
rect 20254 19700 20260 19712
rect 20167 19672 20260 19700
rect 20254 19660 20260 19672
rect 20312 19700 20318 19712
rect 21039 19703 21097 19709
rect 21039 19700 21051 19703
rect 20312 19672 21051 19700
rect 20312 19660 20318 19672
rect 21039 19669 21051 19672
rect 21085 19669 21097 19703
rect 21358 19700 21364 19712
rect 21319 19672 21364 19700
rect 21039 19663 21097 19669
rect 21358 19660 21364 19672
rect 21416 19660 21422 19712
rect 21818 19700 21824 19712
rect 21779 19672 21824 19700
rect 21818 19660 21824 19672
rect 21876 19660 21882 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 1578 19496 1584 19508
rect 1539 19468 1584 19496
rect 1578 19456 1584 19468
rect 1636 19456 1642 19508
rect 3881 19499 3939 19505
rect 3881 19465 3893 19499
rect 3927 19496 3939 19499
rect 3970 19496 3976 19508
rect 3927 19468 3976 19496
rect 3927 19465 3939 19468
rect 3881 19459 3939 19465
rect 3970 19456 3976 19468
rect 4028 19456 4034 19508
rect 4154 19456 4160 19508
rect 4212 19496 4218 19508
rect 6270 19496 6276 19508
rect 4212 19468 4257 19496
rect 6231 19468 6276 19496
rect 4212 19456 4218 19468
rect 6270 19456 6276 19468
rect 6328 19456 6334 19508
rect 8294 19496 8300 19508
rect 8255 19468 8300 19496
rect 8294 19456 8300 19468
rect 8352 19456 8358 19508
rect 9769 19499 9827 19505
rect 9769 19465 9781 19499
rect 9815 19496 9827 19499
rect 10134 19496 10140 19508
rect 9815 19468 10140 19496
rect 9815 19465 9827 19468
rect 9769 19459 9827 19465
rect 10134 19456 10140 19468
rect 10192 19456 10198 19508
rect 11514 19496 11520 19508
rect 11475 19468 11520 19496
rect 11514 19456 11520 19468
rect 11572 19456 11578 19508
rect 17218 19456 17224 19508
rect 17276 19496 17282 19508
rect 18969 19499 19027 19505
rect 18969 19496 18981 19499
rect 17276 19468 18981 19496
rect 17276 19456 17282 19468
rect 18969 19465 18981 19468
rect 19015 19496 19027 19499
rect 19245 19499 19303 19505
rect 19245 19496 19257 19499
rect 19015 19468 19257 19496
rect 19015 19465 19027 19468
rect 18969 19459 19027 19465
rect 19245 19465 19257 19468
rect 19291 19496 19303 19499
rect 19521 19499 19579 19505
rect 19521 19496 19533 19499
rect 19291 19468 19533 19496
rect 19291 19465 19303 19468
rect 19245 19459 19303 19465
rect 19521 19465 19533 19468
rect 19567 19465 19579 19499
rect 19521 19459 19579 19465
rect 5074 19360 5080 19372
rect 5035 19332 5080 19360
rect 5074 19320 5080 19332
rect 5132 19320 5138 19372
rect 5350 19360 5356 19372
rect 5311 19332 5356 19360
rect 5350 19320 5356 19332
rect 5408 19320 5414 19372
rect 8312 19360 8340 19456
rect 10226 19388 10232 19440
rect 10284 19428 10290 19440
rect 10870 19428 10876 19440
rect 10284 19400 10876 19428
rect 10284 19388 10290 19400
rect 10870 19388 10876 19400
rect 10928 19388 10934 19440
rect 8573 19363 8631 19369
rect 8573 19360 8585 19363
rect 8312 19332 8585 19360
rect 8573 19329 8585 19332
rect 8619 19329 8631 19363
rect 8846 19360 8852 19372
rect 8807 19332 8852 19360
rect 8573 19323 8631 19329
rect 8846 19320 8852 19332
rect 8904 19320 8910 19372
rect 11532 19360 11560 19456
rect 11882 19428 11888 19440
rect 11795 19400 11888 19428
rect 11882 19388 11888 19400
rect 11940 19428 11946 19440
rect 17126 19428 17132 19440
rect 11940 19400 16620 19428
rect 17039 19400 17132 19428
rect 11940 19388 11946 19400
rect 12526 19360 12532 19372
rect 9416 19332 11560 19360
rect 12487 19332 12532 19360
rect 1397 19295 1455 19301
rect 1397 19261 1409 19295
rect 1443 19292 1455 19295
rect 4040 19295 4098 19301
rect 1443 19264 1992 19292
rect 1443 19261 1455 19264
rect 1397 19255 1455 19261
rect 1964 19168 1992 19264
rect 4040 19261 4052 19295
rect 4086 19292 4098 19295
rect 6641 19295 6699 19301
rect 4086 19264 4154 19292
rect 4086 19261 4098 19264
rect 4040 19255 4098 19261
rect 3513 19227 3571 19233
rect 3513 19193 3525 19227
rect 3559 19224 3571 19227
rect 3878 19224 3884 19236
rect 3559 19196 3884 19224
rect 3559 19193 3571 19196
rect 3513 19187 3571 19193
rect 3878 19184 3884 19196
rect 3936 19224 3942 19236
rect 4126 19224 4154 19264
rect 6641 19261 6653 19295
rect 6687 19292 6699 19295
rect 7190 19292 7196 19304
rect 6687 19264 7196 19292
rect 6687 19261 6699 19264
rect 6641 19255 6699 19261
rect 7190 19252 7196 19264
rect 7248 19252 7254 19304
rect 7466 19292 7472 19304
rect 7379 19264 7472 19292
rect 7466 19252 7472 19264
rect 7524 19292 7530 19304
rect 7834 19292 7840 19304
rect 7524 19264 7840 19292
rect 7524 19252 7530 19264
rect 7834 19252 7840 19264
rect 7892 19252 7898 19304
rect 5166 19224 5172 19236
rect 3936 19196 4154 19224
rect 5127 19196 5172 19224
rect 3936 19184 3942 19196
rect 5166 19184 5172 19196
rect 5224 19184 5230 19236
rect 7650 19224 7656 19236
rect 7611 19196 7656 19224
rect 7650 19184 7656 19196
rect 7708 19184 7714 19236
rect 8570 19184 8576 19236
rect 8628 19224 8634 19236
rect 8665 19227 8723 19233
rect 8665 19224 8677 19227
rect 8628 19196 8677 19224
rect 8628 19184 8634 19196
rect 8665 19193 8677 19196
rect 8711 19224 8723 19227
rect 9416 19224 9444 19332
rect 12526 19320 12532 19332
rect 12584 19320 12590 19372
rect 12802 19360 12808 19372
rect 12763 19332 12808 19360
rect 12802 19320 12808 19332
rect 12860 19320 12866 19372
rect 13446 19360 13452 19372
rect 13407 19332 13452 19360
rect 13446 19320 13452 19332
rect 13504 19320 13510 19372
rect 14274 19360 14280 19372
rect 14235 19332 14280 19360
rect 14274 19320 14280 19332
rect 14332 19320 14338 19372
rect 16390 19360 16396 19372
rect 16351 19332 16396 19360
rect 16390 19320 16396 19332
rect 16448 19320 16454 19372
rect 16592 19360 16620 19400
rect 17126 19388 17132 19400
rect 17184 19428 17190 19440
rect 20990 19428 20996 19440
rect 17184 19400 20996 19428
rect 17184 19388 17190 19400
rect 20990 19388 20996 19400
rect 21048 19388 21054 19440
rect 18782 19360 18788 19372
rect 16592 19332 18788 19360
rect 18782 19320 18788 19332
rect 18840 19320 18846 19372
rect 19426 19320 19432 19372
rect 19484 19360 19490 19372
rect 19613 19363 19671 19369
rect 19613 19360 19625 19363
rect 19484 19332 19625 19360
rect 19484 19320 19490 19332
rect 19613 19329 19625 19332
rect 19659 19329 19671 19363
rect 19613 19323 19671 19329
rect 19889 19363 19947 19369
rect 19889 19329 19901 19363
rect 19935 19360 19947 19363
rect 20254 19360 20260 19372
rect 19935 19332 20260 19360
rect 19935 19329 19947 19332
rect 19889 19323 19947 19329
rect 20254 19320 20260 19332
rect 20312 19320 20318 19372
rect 23382 19320 23388 19372
rect 23440 19360 23446 19372
rect 24581 19363 24639 19369
rect 24581 19360 24593 19363
rect 23440 19332 24593 19360
rect 23440 19320 23446 19332
rect 24581 19329 24593 19332
rect 24627 19360 24639 19363
rect 24670 19360 24676 19372
rect 24627 19332 24676 19360
rect 24627 19329 24639 19332
rect 24581 19323 24639 19329
rect 24670 19320 24676 19332
rect 24728 19320 24734 19372
rect 10597 19295 10655 19301
rect 10597 19261 10609 19295
rect 10643 19292 10655 19295
rect 11330 19292 11336 19304
rect 10643 19264 11336 19292
rect 10643 19261 10655 19264
rect 10597 19255 10655 19261
rect 11330 19252 11336 19264
rect 11388 19252 11394 19304
rect 18049 19295 18107 19301
rect 18049 19292 18061 19295
rect 17420 19264 18061 19292
rect 10870 19224 10876 19236
rect 8711 19196 9444 19224
rect 9692 19196 10548 19224
rect 10831 19196 10876 19224
rect 8711 19193 8723 19196
rect 8665 19187 8723 19193
rect 1946 19156 1952 19168
rect 1907 19128 1952 19156
rect 1946 19116 1952 19128
rect 2004 19116 2010 19168
rect 4338 19116 4344 19168
rect 4396 19156 4402 19168
rect 4617 19159 4675 19165
rect 4617 19156 4629 19159
rect 4396 19128 4629 19156
rect 4396 19116 4402 19128
rect 4617 19125 4629 19128
rect 4663 19125 4675 19159
rect 4617 19119 4675 19125
rect 8021 19159 8079 19165
rect 8021 19125 8033 19159
rect 8067 19156 8079 19159
rect 8110 19156 8116 19168
rect 8067 19128 8116 19156
rect 8067 19125 8079 19128
rect 8021 19119 8079 19125
rect 8110 19116 8116 19128
rect 8168 19156 8174 19168
rect 9692 19156 9720 19196
rect 10134 19156 10140 19168
rect 8168 19128 9720 19156
rect 10095 19128 10140 19156
rect 8168 19116 8174 19128
rect 10134 19116 10140 19128
rect 10192 19156 10198 19168
rect 10413 19159 10471 19165
rect 10413 19156 10425 19159
rect 10192 19128 10425 19156
rect 10192 19116 10198 19128
rect 10413 19125 10425 19128
rect 10459 19125 10471 19159
rect 10520 19156 10548 19196
rect 10870 19184 10876 19196
rect 10928 19184 10934 19236
rect 11146 19184 11152 19236
rect 11204 19224 11210 19236
rect 12253 19227 12311 19233
rect 12253 19224 12265 19227
rect 11204 19196 12265 19224
rect 11204 19184 11210 19196
rect 12253 19193 12265 19196
rect 12299 19224 12311 19227
rect 12621 19227 12679 19233
rect 12621 19224 12633 19227
rect 12299 19196 12633 19224
rect 12299 19193 12311 19196
rect 12253 19187 12311 19193
rect 12621 19193 12633 19196
rect 12667 19193 12679 19227
rect 12621 19187 12679 19193
rect 15565 19227 15623 19233
rect 15565 19193 15577 19227
rect 15611 19224 15623 19227
rect 15746 19224 15752 19236
rect 15611 19196 15752 19224
rect 15611 19193 15623 19196
rect 15565 19187 15623 19193
rect 15746 19184 15752 19196
rect 15804 19184 15810 19236
rect 16114 19224 16120 19236
rect 16075 19196 16120 19224
rect 16114 19184 16120 19196
rect 16172 19184 16178 19236
rect 16209 19227 16267 19233
rect 16209 19193 16221 19227
rect 16255 19193 16267 19227
rect 16209 19187 16267 19193
rect 11164 19156 11192 19184
rect 10520 19128 11192 19156
rect 10413 19119 10471 19125
rect 13446 19116 13452 19168
rect 13504 19156 13510 19168
rect 14185 19159 14243 19165
rect 14185 19156 14197 19159
rect 13504 19128 14197 19156
rect 13504 19116 13510 19128
rect 14185 19125 14197 19128
rect 14231 19156 14243 19159
rect 14645 19159 14703 19165
rect 14645 19156 14657 19159
rect 14231 19128 14657 19156
rect 14231 19125 14243 19128
rect 14185 19119 14243 19125
rect 14645 19125 14657 19128
rect 14691 19125 14703 19159
rect 14645 19119 14703 19125
rect 15197 19159 15255 19165
rect 15197 19125 15209 19159
rect 15243 19156 15255 19159
rect 15470 19156 15476 19168
rect 15243 19128 15476 19156
rect 15243 19125 15255 19128
rect 15197 19119 15255 19125
rect 15470 19116 15476 19128
rect 15528 19116 15534 19168
rect 15654 19116 15660 19168
rect 15712 19156 15718 19168
rect 15841 19159 15899 19165
rect 15841 19156 15853 19159
rect 15712 19128 15853 19156
rect 15712 19116 15718 19128
rect 15841 19125 15853 19128
rect 15887 19156 15899 19159
rect 16224 19156 16252 19187
rect 17420 19168 17448 19264
rect 18049 19261 18061 19264
rect 18095 19261 18107 19295
rect 18049 19255 18107 19261
rect 21358 19252 21364 19304
rect 21416 19292 21422 19304
rect 21637 19295 21695 19301
rect 21637 19292 21649 19295
rect 21416 19264 21649 19292
rect 21416 19252 21422 19264
rect 21637 19261 21649 19264
rect 21683 19261 21695 19295
rect 21818 19292 21824 19304
rect 21779 19264 21824 19292
rect 21637 19255 21695 19261
rect 18322 19224 18328 19236
rect 18280 19196 18328 19224
rect 18322 19184 18328 19196
rect 18380 19233 18386 19236
rect 18380 19227 18428 19233
rect 18380 19193 18382 19227
rect 18416 19193 18428 19227
rect 18380 19187 18428 19193
rect 19521 19227 19579 19233
rect 19521 19193 19533 19227
rect 19567 19224 19579 19227
rect 19978 19224 19984 19236
rect 19567 19196 19984 19224
rect 19567 19193 19579 19196
rect 19521 19187 19579 19193
rect 18380 19184 18413 19187
rect 19978 19184 19984 19196
rect 20036 19184 20042 19236
rect 20070 19184 20076 19236
rect 20128 19224 20134 19236
rect 20533 19227 20591 19233
rect 20533 19224 20545 19227
rect 20128 19196 20545 19224
rect 20128 19184 20134 19196
rect 20533 19193 20545 19196
rect 20579 19224 20591 19227
rect 20806 19224 20812 19236
rect 20579 19196 20812 19224
rect 20579 19193 20591 19196
rect 20533 19187 20591 19193
rect 20806 19184 20812 19196
rect 20864 19184 20870 19236
rect 21652 19224 21680 19255
rect 21818 19252 21824 19264
rect 21876 19252 21882 19304
rect 23474 19224 23480 19236
rect 21652 19196 23480 19224
rect 23474 19184 23480 19196
rect 23532 19184 23538 19236
rect 17402 19156 17408 19168
rect 15887 19128 16252 19156
rect 17363 19128 17408 19156
rect 15887 19125 15899 19128
rect 15841 19119 15899 19125
rect 17402 19116 17408 19128
rect 17460 19116 17466 19168
rect 17770 19156 17776 19168
rect 17731 19128 17776 19156
rect 17770 19116 17776 19128
rect 17828 19156 17834 19168
rect 18385 19156 18413 19184
rect 20990 19156 20996 19168
rect 17828 19128 18413 19156
rect 20951 19128 20996 19156
rect 17828 19116 17834 19128
rect 20990 19116 20996 19128
rect 21048 19116 21054 19168
rect 21450 19156 21456 19168
rect 21411 19128 21456 19156
rect 21450 19116 21456 19128
rect 21508 19116 21514 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 2961 18955 3019 18961
rect 2961 18921 2973 18955
rect 3007 18952 3019 18955
rect 3970 18952 3976 18964
rect 3007 18924 3976 18952
rect 3007 18921 3019 18924
rect 2961 18915 3019 18921
rect 3970 18912 3976 18924
rect 4028 18912 4034 18964
rect 5074 18912 5080 18964
rect 5132 18952 5138 18964
rect 5534 18952 5540 18964
rect 5132 18924 5540 18952
rect 5132 18912 5138 18924
rect 5534 18912 5540 18924
rect 5592 18952 5598 18964
rect 7009 18955 7067 18961
rect 5592 18924 6316 18952
rect 5592 18912 5598 18924
rect 5721 18887 5779 18893
rect 5721 18853 5733 18887
rect 5767 18884 5779 18887
rect 6086 18884 6092 18896
rect 5767 18856 6092 18884
rect 5767 18853 5779 18856
rect 5721 18847 5779 18853
rect 6086 18844 6092 18856
rect 6144 18844 6150 18896
rect 6288 18893 6316 18924
rect 7009 18921 7021 18955
rect 7055 18952 7067 18955
rect 7466 18952 7472 18964
rect 7055 18924 7472 18952
rect 7055 18921 7067 18924
rect 7009 18915 7067 18921
rect 7466 18912 7472 18924
rect 7524 18912 7530 18964
rect 8110 18952 8116 18964
rect 7668 18924 8116 18952
rect 7668 18893 7696 18924
rect 8110 18912 8116 18924
rect 8168 18912 8174 18964
rect 8570 18952 8576 18964
rect 8531 18924 8576 18952
rect 8570 18912 8576 18924
rect 8628 18912 8634 18964
rect 8938 18952 8944 18964
rect 8899 18924 8944 18952
rect 8938 18912 8944 18924
rect 8996 18912 9002 18964
rect 11330 18912 11336 18964
rect 11388 18952 11394 18964
rect 12437 18955 12495 18961
rect 12437 18952 12449 18955
rect 11388 18924 12449 18952
rect 11388 18912 11394 18924
rect 12437 18921 12449 18924
rect 12483 18921 12495 18955
rect 12437 18915 12495 18921
rect 13262 18912 13268 18964
rect 13320 18952 13326 18964
rect 13357 18955 13415 18961
rect 13357 18952 13369 18955
rect 13320 18924 13369 18952
rect 13320 18912 13326 18924
rect 13357 18921 13369 18924
rect 13403 18921 13415 18955
rect 13357 18915 13415 18921
rect 14139 18955 14197 18961
rect 14139 18921 14151 18955
rect 14185 18952 14197 18955
rect 14642 18952 14648 18964
rect 14185 18924 14648 18952
rect 14185 18921 14197 18924
rect 14139 18915 14197 18921
rect 14642 18912 14648 18924
rect 14700 18912 14706 18964
rect 15105 18955 15163 18961
rect 15105 18921 15117 18955
rect 15151 18952 15163 18955
rect 15194 18952 15200 18964
rect 15151 18924 15200 18952
rect 15151 18921 15163 18924
rect 15105 18915 15163 18921
rect 15194 18912 15200 18924
rect 15252 18912 15258 18964
rect 16114 18912 16120 18964
rect 16172 18952 16178 18964
rect 16666 18952 16672 18964
rect 16172 18924 16672 18952
rect 16172 18912 16178 18924
rect 16666 18912 16672 18924
rect 16724 18912 16730 18964
rect 17954 18912 17960 18964
rect 18012 18952 18018 18964
rect 18601 18955 18659 18961
rect 18601 18952 18613 18955
rect 18012 18924 18613 18952
rect 18012 18912 18018 18924
rect 18601 18921 18613 18924
rect 18647 18952 18659 18955
rect 21450 18952 21456 18964
rect 18647 18924 21456 18952
rect 18647 18921 18659 18924
rect 18601 18915 18659 18921
rect 21450 18912 21456 18924
rect 21508 18912 21514 18964
rect 6273 18887 6331 18893
rect 6273 18853 6285 18887
rect 6319 18853 6331 18887
rect 6273 18847 6331 18853
rect 7653 18887 7711 18893
rect 7653 18853 7665 18887
rect 7699 18853 7711 18887
rect 7653 18847 7711 18853
rect 10502 18844 10508 18896
rect 10560 18884 10566 18896
rect 10689 18887 10747 18893
rect 10689 18884 10701 18887
rect 10560 18856 10701 18884
rect 10560 18844 10566 18856
rect 10689 18853 10701 18856
rect 10735 18884 10747 18887
rect 10965 18887 11023 18893
rect 10965 18884 10977 18887
rect 10735 18856 10977 18884
rect 10735 18853 10747 18856
rect 10689 18847 10747 18853
rect 10965 18853 10977 18856
rect 11011 18853 11023 18887
rect 10965 18847 11023 18853
rect 15378 18844 15384 18896
rect 15436 18884 15442 18896
rect 15473 18887 15531 18893
rect 15473 18884 15485 18887
rect 15436 18856 15485 18884
rect 15436 18844 15442 18856
rect 15473 18853 15485 18856
rect 15519 18853 15531 18887
rect 15473 18847 15531 18853
rect 16025 18887 16083 18893
rect 16025 18853 16037 18887
rect 16071 18884 16083 18887
rect 16390 18884 16396 18896
rect 16071 18856 16396 18884
rect 16071 18853 16083 18856
rect 16025 18847 16083 18853
rect 16390 18844 16396 18856
rect 16448 18844 16454 18896
rect 19334 18844 19340 18896
rect 19392 18884 19398 18896
rect 19429 18887 19487 18893
rect 19429 18884 19441 18887
rect 19392 18856 19441 18884
rect 19392 18844 19398 18856
rect 19429 18853 19441 18856
rect 19475 18853 19487 18887
rect 19429 18847 19487 18853
rect 4592 18819 4650 18825
rect 4592 18785 4604 18819
rect 4638 18816 4650 18819
rect 4706 18816 4712 18828
rect 4638 18788 4712 18816
rect 4638 18785 4650 18788
rect 4592 18779 4650 18785
rect 4706 18776 4712 18788
rect 4764 18776 4770 18828
rect 9585 18819 9643 18825
rect 9585 18785 9597 18819
rect 9631 18816 9643 18819
rect 9674 18816 9680 18828
rect 9631 18788 9680 18816
rect 9631 18785 9643 18788
rect 9585 18779 9643 18785
rect 9674 18776 9680 18788
rect 9732 18776 9738 18828
rect 11790 18776 11796 18828
rect 11848 18816 11854 18828
rect 12345 18819 12403 18825
rect 12345 18816 12357 18819
rect 11848 18788 12357 18816
rect 11848 18776 11854 18788
rect 12345 18785 12357 18788
rect 12391 18785 12403 18819
rect 12345 18779 12403 18785
rect 12897 18819 12955 18825
rect 12897 18785 12909 18819
rect 12943 18816 12955 18819
rect 12986 18816 12992 18828
rect 12943 18788 12992 18816
rect 12943 18785 12955 18788
rect 12897 18779 12955 18785
rect 12986 18776 12992 18788
rect 13044 18776 13050 18828
rect 14068 18819 14126 18825
rect 14068 18785 14080 18819
rect 14114 18816 14126 18819
rect 14274 18816 14280 18828
rect 14114 18788 14280 18816
rect 14114 18785 14126 18788
rect 14068 18779 14126 18785
rect 14274 18776 14280 18788
rect 14332 18776 14338 18828
rect 16298 18776 16304 18828
rect 16356 18816 16362 18828
rect 17218 18816 17224 18828
rect 16356 18788 17224 18816
rect 16356 18776 16362 18788
rect 17218 18776 17224 18788
rect 17276 18776 17282 18828
rect 17681 18819 17739 18825
rect 17681 18785 17693 18819
rect 17727 18816 17739 18819
rect 18325 18819 18383 18825
rect 18325 18816 18337 18819
rect 17727 18788 18337 18816
rect 17727 18785 17739 18788
rect 17681 18779 17739 18785
rect 18325 18785 18337 18788
rect 18371 18785 18383 18819
rect 20898 18816 20904 18828
rect 20859 18788 20904 18816
rect 18325 18779 18383 18785
rect 20898 18776 20904 18788
rect 20956 18776 20962 18828
rect 21174 18776 21180 18828
rect 21232 18816 21238 18828
rect 21361 18819 21419 18825
rect 21361 18816 21373 18819
rect 21232 18788 21373 18816
rect 21232 18776 21238 18788
rect 21361 18785 21373 18788
rect 21407 18785 21419 18819
rect 21361 18779 21419 18785
rect 5629 18751 5687 18757
rect 5629 18717 5641 18751
rect 5675 18748 5687 18751
rect 5994 18748 6000 18760
rect 5675 18720 6000 18748
rect 5675 18717 5687 18720
rect 5629 18711 5687 18717
rect 5994 18708 6000 18720
rect 6052 18708 6058 18760
rect 7558 18748 7564 18760
rect 7519 18720 7564 18748
rect 7558 18708 7564 18720
rect 7616 18708 7622 18760
rect 7834 18748 7840 18760
rect 7795 18720 7840 18748
rect 7834 18708 7840 18720
rect 7892 18708 7898 18760
rect 9815 18751 9873 18757
rect 9815 18748 9827 18751
rect 7944 18720 9827 18748
rect 4663 18683 4721 18689
rect 4663 18649 4675 18683
rect 4709 18680 4721 18683
rect 5258 18680 5264 18692
rect 4709 18652 5264 18680
rect 4709 18649 4721 18652
rect 4663 18643 4721 18649
rect 5258 18640 5264 18652
rect 5316 18680 5322 18692
rect 5353 18683 5411 18689
rect 5353 18680 5365 18683
rect 5316 18652 5365 18680
rect 5316 18640 5322 18652
rect 5353 18649 5365 18652
rect 5399 18649 5411 18683
rect 7374 18680 7380 18692
rect 7287 18652 7380 18680
rect 5353 18643 5411 18649
rect 7374 18640 7380 18652
rect 7432 18680 7438 18692
rect 7944 18680 7972 18720
rect 9815 18717 9827 18720
rect 9861 18717 9873 18751
rect 9815 18711 9873 18717
rect 10321 18751 10379 18757
rect 10321 18717 10333 18751
rect 10367 18748 10379 18751
rect 10870 18748 10876 18760
rect 10367 18720 10876 18748
rect 10367 18717 10379 18720
rect 10321 18711 10379 18717
rect 10870 18708 10876 18720
rect 10928 18708 10934 18760
rect 11149 18751 11207 18757
rect 11149 18717 11161 18751
rect 11195 18717 11207 18751
rect 11149 18711 11207 18717
rect 7432 18652 7972 18680
rect 7432 18640 7438 18652
rect 8846 18640 8852 18692
rect 8904 18680 8910 18692
rect 10962 18680 10968 18692
rect 8904 18652 10968 18680
rect 8904 18640 8910 18652
rect 10962 18640 10968 18652
rect 11020 18680 11026 18692
rect 11164 18680 11192 18711
rect 14366 18708 14372 18760
rect 14424 18748 14430 18760
rect 14826 18748 14832 18760
rect 14424 18720 14832 18748
rect 14424 18708 14430 18720
rect 14826 18708 14832 18720
rect 14884 18748 14890 18760
rect 15381 18751 15439 18757
rect 15381 18748 15393 18751
rect 14884 18720 15393 18748
rect 14884 18708 14890 18720
rect 15381 18717 15393 18720
rect 15427 18748 15439 18751
rect 16482 18748 16488 18760
rect 15427 18720 16488 18748
rect 15427 18717 15439 18720
rect 15381 18711 15439 18717
rect 16482 18708 16488 18720
rect 16540 18708 16546 18760
rect 17862 18748 17868 18760
rect 17823 18720 17868 18748
rect 17862 18708 17868 18720
rect 17920 18708 17926 18760
rect 19058 18708 19064 18760
rect 19116 18748 19122 18760
rect 19337 18751 19395 18757
rect 19337 18748 19349 18751
rect 19116 18720 19349 18748
rect 19116 18708 19122 18720
rect 19337 18717 19349 18720
rect 19383 18748 19395 18751
rect 19518 18748 19524 18760
rect 19383 18720 19524 18748
rect 19383 18717 19395 18720
rect 19337 18711 19395 18717
rect 19518 18708 19524 18720
rect 19576 18708 19582 18760
rect 19981 18751 20039 18757
rect 19981 18717 19993 18751
rect 20027 18748 20039 18751
rect 20070 18748 20076 18760
rect 20027 18720 20076 18748
rect 20027 18717 20039 18720
rect 19981 18711 20039 18717
rect 20070 18708 20076 18720
rect 20128 18708 20134 18760
rect 21453 18751 21511 18757
rect 21453 18748 21465 18751
rect 20640 18720 21465 18748
rect 11020 18652 11192 18680
rect 11020 18640 11026 18652
rect 14734 18640 14740 18692
rect 14792 18680 14798 18692
rect 20640 18680 20668 18720
rect 21453 18717 21465 18720
rect 21499 18717 21511 18751
rect 21453 18711 21511 18717
rect 14792 18652 20668 18680
rect 14792 18640 14798 18652
rect 20990 18640 20996 18692
rect 21048 18680 21054 18692
rect 27614 18680 27620 18692
rect 21048 18652 27620 18680
rect 21048 18640 21054 18652
rect 27614 18640 27620 18652
rect 27672 18640 27678 18692
rect 4154 18572 4160 18624
rect 4212 18612 4218 18624
rect 4798 18612 4804 18624
rect 4212 18584 4804 18612
rect 4212 18572 4218 18584
rect 4798 18572 4804 18584
rect 4856 18572 4862 18624
rect 5074 18612 5080 18624
rect 5035 18584 5080 18612
rect 5074 18572 5080 18584
rect 5132 18572 5138 18624
rect 14550 18612 14556 18624
rect 14511 18584 14556 18612
rect 14550 18572 14556 18584
rect 14608 18572 14614 18624
rect 16390 18612 16396 18624
rect 16351 18584 16396 18612
rect 16390 18572 16396 18584
rect 16448 18572 16454 18624
rect 17770 18572 17776 18624
rect 17828 18612 17834 18624
rect 18141 18615 18199 18621
rect 18141 18612 18153 18615
rect 17828 18584 18153 18612
rect 17828 18572 17834 18584
rect 18141 18581 18153 18584
rect 18187 18581 18199 18615
rect 18141 18575 18199 18581
rect 18322 18572 18328 18624
rect 18380 18612 18386 18624
rect 21818 18612 21824 18624
rect 18380 18584 21824 18612
rect 18380 18572 18386 18584
rect 21818 18572 21824 18584
rect 21876 18572 21882 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 6086 18368 6092 18420
rect 6144 18408 6150 18420
rect 6181 18411 6239 18417
rect 6181 18408 6193 18411
rect 6144 18380 6193 18408
rect 6144 18368 6150 18380
rect 6181 18377 6193 18380
rect 6227 18377 6239 18411
rect 6181 18371 6239 18377
rect 8110 18368 8116 18420
rect 8168 18408 8174 18420
rect 8297 18411 8355 18417
rect 8297 18408 8309 18411
rect 8168 18380 8309 18408
rect 8168 18368 8174 18380
rect 8297 18377 8309 18380
rect 8343 18377 8355 18411
rect 8297 18371 8355 18377
rect 9769 18411 9827 18417
rect 9769 18377 9781 18411
rect 9815 18408 9827 18411
rect 9858 18408 9864 18420
rect 9815 18380 9864 18408
rect 9815 18377 9827 18380
rect 9769 18371 9827 18377
rect 9858 18368 9864 18380
rect 9916 18408 9922 18420
rect 10502 18408 10508 18420
rect 9916 18380 10508 18408
rect 9916 18368 9922 18380
rect 10502 18368 10508 18380
rect 10560 18408 10566 18420
rect 10778 18408 10784 18420
rect 10560 18380 10784 18408
rect 10560 18368 10566 18380
rect 10778 18368 10784 18380
rect 10836 18368 10842 18420
rect 14550 18368 14556 18420
rect 14608 18408 14614 18420
rect 16853 18411 16911 18417
rect 16853 18408 16865 18411
rect 14608 18380 16865 18408
rect 14608 18368 14614 18380
rect 7926 18300 7932 18352
rect 7984 18340 7990 18352
rect 9674 18340 9680 18352
rect 7984 18312 9680 18340
rect 7984 18300 7990 18312
rect 9674 18300 9680 18312
rect 9732 18340 9738 18352
rect 10137 18343 10195 18349
rect 10137 18340 10149 18343
rect 9732 18312 10149 18340
rect 9732 18300 9738 18312
rect 10137 18309 10149 18312
rect 10183 18309 10195 18343
rect 10137 18303 10195 18309
rect 4338 18272 4344 18284
rect 4299 18244 4344 18272
rect 4338 18232 4344 18244
rect 4396 18232 4402 18284
rect 5258 18272 5264 18284
rect 5219 18244 5264 18272
rect 5258 18232 5264 18244
rect 5316 18232 5322 18284
rect 5534 18272 5540 18284
rect 5495 18244 5540 18272
rect 5534 18232 5540 18244
rect 5592 18232 5598 18284
rect 7374 18272 7380 18284
rect 7335 18244 7380 18272
rect 7374 18232 7380 18244
rect 7432 18232 7438 18284
rect 7834 18272 7840 18284
rect 7795 18244 7840 18272
rect 7834 18232 7840 18244
rect 7892 18232 7898 18284
rect 8849 18275 8907 18281
rect 8849 18241 8861 18275
rect 8895 18272 8907 18275
rect 8938 18272 8944 18284
rect 8895 18244 8944 18272
rect 8895 18241 8907 18244
rect 8849 18235 8907 18241
rect 8938 18232 8944 18244
rect 8996 18232 9002 18284
rect 10042 18232 10048 18284
rect 10100 18272 10106 18284
rect 10686 18272 10692 18284
rect 10100 18244 10692 18272
rect 10100 18232 10106 18244
rect 10686 18232 10692 18244
rect 10744 18232 10750 18284
rect 11333 18275 11391 18281
rect 11333 18241 11345 18275
rect 11379 18272 11391 18275
rect 12434 18272 12440 18284
rect 11379 18244 12440 18272
rect 11379 18241 11391 18244
rect 11333 18235 11391 18241
rect 12434 18232 12440 18244
rect 12492 18272 12498 18284
rect 12802 18272 12808 18284
rect 12492 18244 12808 18272
rect 12492 18232 12498 18244
rect 12802 18232 12808 18244
rect 12860 18232 12866 18284
rect 3513 18207 3571 18213
rect 3513 18173 3525 18207
rect 3559 18204 3571 18207
rect 4249 18207 4307 18213
rect 4249 18204 4261 18207
rect 3559 18176 4261 18204
rect 3559 18173 3571 18176
rect 3513 18167 3571 18173
rect 4249 18173 4261 18176
rect 4295 18204 4307 18207
rect 4982 18204 4988 18216
rect 4295 18176 4988 18204
rect 4295 18173 4307 18176
rect 4249 18167 4307 18173
rect 4982 18164 4988 18176
rect 5040 18164 5046 18216
rect 12253 18207 12311 18213
rect 12253 18173 12265 18207
rect 12299 18204 12311 18207
rect 12710 18204 12716 18216
rect 12299 18176 12716 18204
rect 12299 18173 12311 18176
rect 12253 18167 12311 18173
rect 12710 18164 12716 18176
rect 12768 18164 12774 18216
rect 12986 18204 12992 18216
rect 12947 18176 12992 18204
rect 12986 18164 12992 18176
rect 13044 18164 13050 18216
rect 14752 18213 14780 18380
rect 16853 18377 16865 18380
rect 16899 18408 16911 18411
rect 18322 18408 18328 18420
rect 16899 18380 18328 18408
rect 16899 18377 16911 18380
rect 16853 18371 16911 18377
rect 18322 18368 18328 18380
rect 18380 18368 18386 18420
rect 18966 18408 18972 18420
rect 18927 18380 18972 18408
rect 18966 18368 18972 18380
rect 19024 18408 19030 18420
rect 19705 18411 19763 18417
rect 19705 18408 19717 18411
rect 19024 18380 19717 18408
rect 19024 18368 19030 18380
rect 19705 18377 19717 18380
rect 19751 18408 19763 18411
rect 20162 18408 20168 18420
rect 19751 18380 20168 18408
rect 19751 18377 19763 18380
rect 19705 18371 19763 18377
rect 20162 18368 20168 18380
rect 20220 18368 20226 18420
rect 20898 18408 20904 18420
rect 20859 18380 20904 18408
rect 20898 18368 20904 18380
rect 20956 18368 20962 18420
rect 24762 18408 24768 18420
rect 24723 18380 24768 18408
rect 24762 18368 24768 18380
rect 24820 18368 24826 18420
rect 17402 18340 17408 18352
rect 15625 18312 17408 18340
rect 14921 18275 14979 18281
rect 14921 18241 14933 18275
rect 14967 18272 14979 18275
rect 15625 18272 15653 18312
rect 17402 18300 17408 18312
rect 17460 18300 17466 18352
rect 20530 18340 20536 18352
rect 20491 18312 20536 18340
rect 20530 18300 20536 18312
rect 20588 18300 20594 18352
rect 14967 18244 15653 18272
rect 15841 18275 15899 18281
rect 14967 18241 14979 18244
rect 14921 18235 14979 18241
rect 15841 18241 15853 18275
rect 15887 18272 15899 18275
rect 16298 18272 16304 18284
rect 15887 18244 16304 18272
rect 15887 18241 15899 18244
rect 15841 18235 15899 18241
rect 16298 18232 16304 18244
rect 16356 18232 16362 18284
rect 16482 18272 16488 18284
rect 16443 18244 16488 18272
rect 16482 18232 16488 18244
rect 16540 18232 16546 18284
rect 17862 18232 17868 18284
rect 17920 18272 17926 18284
rect 18049 18275 18107 18281
rect 18049 18272 18061 18275
rect 17920 18244 18061 18272
rect 17920 18232 17926 18244
rect 18049 18241 18061 18244
rect 18095 18241 18107 18275
rect 18049 18235 18107 18241
rect 14185 18207 14243 18213
rect 14185 18204 14197 18207
rect 13786 18176 14197 18204
rect 5077 18139 5135 18145
rect 5077 18105 5089 18139
rect 5123 18136 5135 18139
rect 5350 18136 5356 18148
rect 5123 18108 5356 18136
rect 5123 18105 5135 18108
rect 5077 18099 5135 18105
rect 5350 18096 5356 18108
rect 5408 18096 5414 18148
rect 7193 18139 7251 18145
rect 7193 18105 7205 18139
rect 7239 18136 7251 18139
rect 7469 18139 7527 18145
rect 7469 18136 7481 18139
rect 7239 18108 7481 18136
rect 7239 18105 7251 18108
rect 7193 18099 7251 18105
rect 7469 18105 7481 18108
rect 7515 18136 7527 18139
rect 8570 18136 8576 18148
rect 7515 18108 8576 18136
rect 7515 18105 7527 18108
rect 7469 18099 7527 18105
rect 8570 18096 8576 18108
rect 8628 18096 8634 18148
rect 8754 18096 8760 18148
rect 8812 18136 8818 18148
rect 9211 18139 9269 18145
rect 9211 18136 9223 18139
rect 8812 18108 9223 18136
rect 8812 18096 8818 18108
rect 9211 18105 9223 18108
rect 9257 18136 9269 18139
rect 10134 18136 10140 18148
rect 9257 18108 10140 18136
rect 9257 18105 9269 18108
rect 9211 18099 9269 18105
rect 10134 18096 10140 18108
rect 10192 18096 10198 18148
rect 10778 18096 10784 18148
rect 10836 18136 10842 18148
rect 10836 18108 10881 18136
rect 10836 18096 10842 18108
rect 4706 18068 4712 18080
rect 4619 18040 4712 18068
rect 4706 18028 4712 18040
rect 4764 18068 4770 18080
rect 7006 18068 7012 18080
rect 4764 18040 7012 18068
rect 4764 18028 4770 18040
rect 7006 18028 7012 18040
rect 7064 18028 7070 18080
rect 11790 18068 11796 18080
rect 11751 18040 11796 18068
rect 11790 18028 11796 18040
rect 11848 18028 11854 18080
rect 12526 18068 12532 18080
rect 12487 18040 12532 18068
rect 12526 18028 12532 18040
rect 12584 18028 12590 18080
rect 13630 18068 13636 18080
rect 13591 18040 13636 18068
rect 13630 18028 13636 18040
rect 13688 18068 13694 18080
rect 13786 18068 13814 18176
rect 14185 18173 14197 18176
rect 14231 18173 14243 18207
rect 14185 18167 14243 18173
rect 14737 18207 14795 18213
rect 14737 18173 14749 18207
rect 14783 18173 14795 18207
rect 14737 18167 14795 18173
rect 24210 18164 24216 18216
rect 24268 18204 24274 18216
rect 24581 18207 24639 18213
rect 24581 18204 24593 18207
rect 24268 18176 24593 18204
rect 24268 18164 24274 18176
rect 24581 18173 24593 18176
rect 24627 18204 24639 18207
rect 25133 18207 25191 18213
rect 25133 18204 25145 18207
rect 24627 18176 25145 18204
rect 24627 18173 24639 18176
rect 24581 18167 24639 18173
rect 25133 18173 25145 18176
rect 25179 18173 25191 18207
rect 25133 18167 25191 18173
rect 15470 18096 15476 18148
rect 15528 18136 15534 18148
rect 15657 18139 15715 18145
rect 15657 18136 15669 18139
rect 15528 18108 15669 18136
rect 15528 18096 15534 18108
rect 15657 18105 15669 18108
rect 15703 18136 15715 18139
rect 15933 18139 15991 18145
rect 15933 18136 15945 18139
rect 15703 18108 15945 18136
rect 15703 18105 15715 18108
rect 15657 18099 15715 18105
rect 15933 18105 15945 18108
rect 15979 18105 15991 18139
rect 15933 18099 15991 18105
rect 18370 18139 18428 18145
rect 18370 18105 18382 18139
rect 18416 18105 18428 18139
rect 19978 18136 19984 18148
rect 19939 18108 19984 18136
rect 18370 18099 18428 18105
rect 13688 18040 13814 18068
rect 14093 18071 14151 18077
rect 13688 18028 13694 18040
rect 14093 18037 14105 18071
rect 14139 18068 14151 18071
rect 14274 18068 14280 18080
rect 14139 18040 14280 18068
rect 14139 18037 14151 18040
rect 14093 18031 14151 18037
rect 14274 18028 14280 18040
rect 14332 18028 14338 18080
rect 15286 18068 15292 18080
rect 15247 18040 15292 18068
rect 15286 18028 15292 18040
rect 15344 18028 15350 18080
rect 17218 18068 17224 18080
rect 17179 18040 17224 18068
rect 17218 18028 17224 18040
rect 17276 18028 17282 18080
rect 17770 18068 17776 18080
rect 17731 18040 17776 18068
rect 17770 18028 17776 18040
rect 17828 18068 17834 18080
rect 18385 18068 18413 18099
rect 19978 18096 19984 18108
rect 20036 18096 20042 18148
rect 20073 18139 20131 18145
rect 20073 18105 20085 18139
rect 20119 18136 20131 18139
rect 20162 18136 20168 18148
rect 20119 18108 20168 18136
rect 20119 18105 20131 18108
rect 20073 18099 20131 18105
rect 20162 18096 20168 18108
rect 20220 18096 20226 18148
rect 19242 18068 19248 18080
rect 17828 18040 18413 18068
rect 19203 18040 19248 18068
rect 17828 18028 17834 18040
rect 19242 18028 19248 18040
rect 19300 18028 19306 18080
rect 21174 18028 21180 18080
rect 21232 18068 21238 18080
rect 21269 18071 21327 18077
rect 21269 18068 21281 18071
rect 21232 18040 21281 18068
rect 21232 18028 21238 18040
rect 21269 18037 21281 18040
rect 21315 18037 21327 18071
rect 21269 18031 21327 18037
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 4798 17864 4804 17876
rect 4759 17836 4804 17864
rect 4798 17824 4804 17836
rect 4856 17824 4862 17876
rect 5721 17867 5779 17873
rect 5721 17833 5733 17867
rect 5767 17864 5779 17867
rect 5994 17864 6000 17876
rect 5767 17836 6000 17864
rect 5767 17833 5779 17836
rect 5721 17827 5779 17833
rect 5994 17824 6000 17836
rect 6052 17824 6058 17876
rect 10686 17864 10692 17876
rect 10647 17836 10692 17864
rect 10686 17824 10692 17836
rect 10744 17824 10750 17876
rect 11333 17867 11391 17873
rect 11333 17833 11345 17867
rect 11379 17864 11391 17867
rect 12526 17864 12532 17876
rect 11379 17836 12532 17864
rect 11379 17833 11391 17836
rect 11333 17827 11391 17833
rect 5350 17756 5356 17808
rect 5408 17796 5414 17808
rect 6181 17799 6239 17805
rect 6181 17796 6193 17799
rect 5408 17768 6193 17796
rect 5408 17756 5414 17768
rect 6181 17765 6193 17768
rect 6227 17765 6239 17799
rect 8202 17796 8208 17808
rect 8163 17768 8208 17796
rect 6181 17759 6239 17765
rect 8202 17756 8208 17768
rect 8260 17756 8266 17808
rect 9858 17796 9864 17808
rect 9819 17768 9864 17796
rect 9858 17756 9864 17768
rect 9916 17756 9922 17808
rect 6086 17688 6092 17740
rect 6144 17728 6150 17740
rect 11440 17737 11468 17836
rect 12526 17824 12532 17836
rect 12584 17824 12590 17876
rect 14826 17824 14832 17876
rect 14884 17864 14890 17876
rect 15013 17867 15071 17873
rect 15013 17864 15025 17867
rect 14884 17836 15025 17864
rect 14884 17824 14890 17836
rect 15013 17833 15025 17836
rect 15059 17833 15071 17867
rect 15013 17827 15071 17833
rect 15286 17824 15292 17876
rect 15344 17864 15350 17876
rect 16209 17867 16267 17873
rect 16209 17864 16221 17867
rect 15344 17836 16221 17864
rect 15344 17824 15350 17836
rect 16209 17833 16221 17836
rect 16255 17833 16267 17867
rect 16209 17827 16267 17833
rect 17862 17824 17868 17876
rect 17920 17864 17926 17876
rect 18049 17867 18107 17873
rect 18049 17864 18061 17867
rect 17920 17836 18061 17864
rect 17920 17824 17926 17836
rect 18049 17833 18061 17836
rect 18095 17833 18107 17867
rect 18049 17827 18107 17833
rect 19245 17867 19303 17873
rect 19245 17833 19257 17867
rect 19291 17864 19303 17867
rect 19291 17836 21128 17864
rect 19291 17833 19303 17836
rect 19245 17827 19303 17833
rect 11606 17756 11612 17808
rect 11664 17796 11670 17808
rect 11746 17799 11804 17805
rect 11746 17796 11758 17799
rect 11664 17768 11758 17796
rect 11664 17756 11670 17768
rect 11746 17765 11758 17768
rect 11792 17765 11804 17799
rect 11746 17759 11804 17765
rect 15470 17756 15476 17808
rect 15528 17796 15534 17808
rect 15610 17799 15668 17805
rect 15610 17796 15622 17799
rect 15528 17768 15622 17796
rect 15528 17756 15534 17768
rect 15610 17765 15622 17768
rect 15656 17765 15668 17799
rect 15610 17759 15668 17765
rect 17770 17756 17776 17808
rect 17828 17796 17834 17808
rect 18646 17799 18704 17805
rect 18646 17796 18658 17799
rect 17828 17768 18658 17796
rect 17828 17756 17834 17768
rect 18646 17765 18658 17768
rect 18692 17765 18704 17799
rect 20530 17796 20536 17808
rect 20491 17768 20536 17796
rect 18646 17759 18704 17765
rect 20530 17756 20536 17768
rect 20588 17756 20594 17808
rect 20806 17756 20812 17808
rect 20864 17796 20870 17808
rect 21100 17805 21128 17836
rect 20993 17799 21051 17805
rect 20993 17796 21005 17799
rect 20864 17768 21005 17796
rect 20864 17756 20870 17768
rect 20993 17765 21005 17768
rect 21039 17765 21051 17799
rect 20993 17759 21051 17765
rect 21085 17799 21143 17805
rect 21085 17765 21097 17799
rect 21131 17796 21143 17799
rect 21450 17796 21456 17808
rect 21131 17768 21456 17796
rect 21131 17765 21143 17768
rect 21085 17759 21143 17765
rect 21450 17756 21456 17768
rect 21508 17756 21514 17808
rect 6273 17731 6331 17737
rect 6273 17728 6285 17731
rect 6144 17700 6285 17728
rect 6144 17688 6150 17700
rect 6273 17697 6285 17700
rect 6319 17697 6331 17731
rect 6273 17691 6331 17697
rect 11425 17731 11483 17737
rect 11425 17697 11437 17731
rect 11471 17697 11483 17731
rect 13630 17728 13636 17740
rect 13591 17700 13636 17728
rect 11425 17691 11483 17697
rect 13630 17688 13636 17700
rect 13688 17688 13694 17740
rect 14182 17728 14188 17740
rect 14143 17700 14188 17728
rect 14182 17688 14188 17700
rect 14240 17688 14246 17740
rect 4246 17620 4252 17672
rect 4304 17660 4310 17672
rect 4433 17663 4491 17669
rect 4433 17660 4445 17663
rect 4304 17632 4445 17660
rect 4304 17620 4310 17632
rect 4433 17629 4445 17632
rect 4479 17629 4491 17663
rect 4433 17623 4491 17629
rect 5534 17620 5540 17672
rect 5592 17660 5598 17672
rect 7469 17663 7527 17669
rect 7469 17660 7481 17663
rect 5592 17632 7481 17660
rect 5592 17620 5598 17632
rect 7469 17629 7481 17632
rect 7515 17660 7527 17663
rect 7558 17660 7564 17672
rect 7515 17632 7564 17660
rect 7515 17629 7527 17632
rect 7469 17623 7527 17629
rect 7558 17620 7564 17632
rect 7616 17620 7622 17672
rect 7834 17620 7840 17672
rect 7892 17660 7898 17672
rect 8113 17663 8171 17669
rect 8113 17660 8125 17663
rect 7892 17632 8125 17660
rect 7892 17620 7898 17632
rect 8113 17629 8125 17632
rect 8159 17629 8171 17663
rect 8113 17623 8171 17629
rect 8389 17663 8447 17669
rect 8389 17629 8401 17663
rect 8435 17629 8447 17663
rect 9766 17660 9772 17672
rect 9727 17632 9772 17660
rect 8389 17623 8447 17629
rect 5074 17552 5080 17604
rect 5132 17592 5138 17604
rect 5353 17595 5411 17601
rect 5353 17592 5365 17595
rect 5132 17564 5365 17592
rect 5132 17552 5138 17564
rect 5353 17561 5365 17564
rect 5399 17561 5411 17595
rect 8404 17592 8432 17623
rect 9766 17620 9772 17632
rect 9824 17620 9830 17672
rect 10042 17660 10048 17672
rect 10003 17632 10048 17660
rect 10042 17620 10048 17632
rect 10100 17620 10106 17672
rect 14369 17663 14427 17669
rect 14369 17629 14381 17663
rect 14415 17660 14427 17663
rect 14826 17660 14832 17672
rect 14415 17632 14832 17660
rect 14415 17629 14427 17632
rect 14369 17623 14427 17629
rect 14826 17620 14832 17632
rect 14884 17620 14890 17672
rect 15286 17660 15292 17672
rect 15247 17632 15292 17660
rect 15286 17620 15292 17632
rect 15344 17620 15350 17672
rect 17678 17620 17684 17672
rect 17736 17660 17742 17672
rect 18325 17663 18383 17669
rect 18325 17660 18337 17663
rect 17736 17632 18337 17660
rect 17736 17620 17742 17632
rect 18325 17629 18337 17632
rect 18371 17629 18383 17663
rect 21266 17660 21272 17672
rect 21227 17632 21272 17660
rect 18325 17623 18383 17629
rect 21266 17620 21272 17632
rect 21324 17620 21330 17672
rect 11146 17592 11152 17604
rect 5353 17555 5411 17561
rect 7392 17564 11152 17592
rect 2038 17484 2044 17536
rect 2096 17524 2102 17536
rect 7392 17524 7420 17564
rect 11146 17552 11152 17564
rect 11204 17552 11210 17604
rect 12342 17524 12348 17536
rect 2096 17496 7420 17524
rect 12303 17496 12348 17524
rect 2096 17484 2102 17496
rect 12342 17484 12348 17496
rect 12400 17484 12406 17536
rect 12713 17527 12771 17533
rect 12713 17493 12725 17527
rect 12759 17524 12771 17527
rect 12986 17524 12992 17536
rect 12759 17496 12992 17524
rect 12759 17493 12771 17496
rect 12713 17487 12771 17493
rect 12986 17484 12992 17496
rect 13044 17524 13050 17536
rect 13081 17527 13139 17533
rect 13081 17524 13093 17527
rect 13044 17496 13093 17524
rect 13044 17484 13050 17496
rect 13081 17493 13093 17496
rect 13127 17524 13139 17527
rect 13354 17524 13360 17536
rect 13127 17496 13360 17524
rect 13127 17493 13139 17496
rect 13081 17487 13139 17493
rect 13354 17484 13360 17496
rect 13412 17484 13418 17536
rect 19518 17524 19524 17536
rect 19479 17496 19524 17524
rect 19518 17484 19524 17496
rect 19576 17484 19582 17536
rect 19978 17524 19984 17536
rect 19891 17496 19984 17524
rect 19978 17484 19984 17496
rect 20036 17524 20042 17536
rect 20254 17524 20260 17536
rect 20036 17496 20260 17524
rect 20036 17484 20042 17496
rect 20254 17484 20260 17496
rect 20312 17484 20318 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 2823 17323 2881 17329
rect 2823 17289 2835 17323
rect 2869 17320 2881 17323
rect 5534 17320 5540 17332
rect 2869 17292 5540 17320
rect 2869 17289 2881 17292
rect 2823 17283 2881 17289
rect 5534 17280 5540 17292
rect 5592 17280 5598 17332
rect 5629 17323 5687 17329
rect 5629 17289 5641 17323
rect 5675 17320 5687 17323
rect 6086 17320 6092 17332
rect 5675 17292 6092 17320
rect 5675 17289 5687 17292
rect 5629 17283 5687 17289
rect 6086 17280 6092 17292
rect 6144 17320 6150 17332
rect 6181 17323 6239 17329
rect 6181 17320 6193 17323
rect 6144 17292 6193 17320
rect 6144 17280 6150 17292
rect 6181 17289 6193 17292
rect 6227 17289 6239 17323
rect 6181 17283 6239 17289
rect 7834 17280 7840 17332
rect 7892 17320 7898 17332
rect 9125 17323 9183 17329
rect 9125 17320 9137 17323
rect 7892 17292 9137 17320
rect 7892 17280 7898 17292
rect 9125 17289 9137 17292
rect 9171 17320 9183 17323
rect 10042 17320 10048 17332
rect 9171 17292 10048 17320
rect 9171 17289 9183 17292
rect 9125 17283 9183 17289
rect 10042 17280 10048 17292
rect 10100 17280 10106 17332
rect 10597 17323 10655 17329
rect 10597 17289 10609 17323
rect 10643 17320 10655 17323
rect 10778 17320 10784 17332
rect 10643 17292 10784 17320
rect 10643 17289 10655 17292
rect 10597 17283 10655 17289
rect 10778 17280 10784 17292
rect 10836 17280 10842 17332
rect 11606 17280 11612 17332
rect 11664 17320 11670 17332
rect 11793 17323 11851 17329
rect 11793 17320 11805 17323
rect 11664 17292 11805 17320
rect 11664 17280 11670 17292
rect 11793 17289 11805 17292
rect 11839 17289 11851 17323
rect 11793 17283 11851 17289
rect 12253 17323 12311 17329
rect 12253 17289 12265 17323
rect 12299 17320 12311 17323
rect 12342 17320 12348 17332
rect 12299 17292 12348 17320
rect 12299 17289 12311 17292
rect 12253 17283 12311 17289
rect 12342 17280 12348 17292
rect 12400 17280 12406 17332
rect 13446 17280 13452 17332
rect 13504 17320 13510 17332
rect 14553 17323 14611 17329
rect 14553 17320 14565 17323
rect 13504 17292 14565 17320
rect 13504 17280 13510 17292
rect 14553 17289 14565 17292
rect 14599 17320 14611 17323
rect 14642 17320 14648 17332
rect 14599 17292 14648 17320
rect 14599 17289 14611 17292
rect 14553 17283 14611 17289
rect 14642 17280 14648 17292
rect 14700 17280 14706 17332
rect 15654 17320 15660 17332
rect 15615 17292 15660 17320
rect 15654 17280 15660 17292
rect 15712 17280 15718 17332
rect 16298 17280 16304 17332
rect 16356 17320 16362 17332
rect 21269 17323 21327 17329
rect 21269 17320 21281 17323
rect 16356 17292 21281 17320
rect 16356 17280 16362 17292
rect 21269 17289 21281 17292
rect 21315 17289 21327 17323
rect 21450 17320 21456 17332
rect 21411 17292 21456 17320
rect 21269 17283 21327 17289
rect 21450 17280 21456 17292
rect 21508 17280 21514 17332
rect 23799 17323 23857 17329
rect 23799 17289 23811 17323
rect 23845 17320 23857 17323
rect 24210 17320 24216 17332
rect 23845 17292 24216 17320
rect 23845 17289 23857 17292
rect 23799 17283 23857 17289
rect 24210 17280 24216 17292
rect 24268 17280 24274 17332
rect 8202 17212 8208 17264
rect 8260 17252 8266 17264
rect 8849 17255 8907 17261
rect 8849 17252 8861 17255
rect 8260 17224 8861 17252
rect 8260 17212 8266 17224
rect 8849 17221 8861 17224
rect 8895 17221 8907 17255
rect 8849 17215 8907 17221
rect 9585 17255 9643 17261
rect 9585 17221 9597 17255
rect 9631 17252 9643 17255
rect 9766 17252 9772 17264
rect 9631 17224 9772 17252
rect 9631 17221 9643 17224
rect 9585 17215 9643 17221
rect 9766 17212 9772 17224
rect 9824 17212 9830 17264
rect 9861 17255 9919 17261
rect 9861 17221 9873 17255
rect 9907 17252 9919 17255
rect 11238 17252 11244 17264
rect 9907 17224 11244 17252
rect 9907 17221 9919 17224
rect 9861 17215 9919 17221
rect 11238 17212 11244 17224
rect 11296 17252 11302 17264
rect 12986 17252 12992 17264
rect 11296 17224 12992 17252
rect 11296 17212 11302 17224
rect 12986 17212 12992 17224
rect 13044 17212 13050 17264
rect 15286 17212 15292 17264
rect 15344 17252 15350 17264
rect 16393 17255 16451 17261
rect 16393 17252 16405 17255
rect 15344 17224 16405 17252
rect 15344 17212 15350 17224
rect 16393 17221 16405 17224
rect 16439 17252 16451 17255
rect 16439 17224 21496 17252
rect 16439 17221 16451 17224
rect 16393 17215 16451 17221
rect 7098 17184 7104 17196
rect 4126 17156 7104 17184
rect 2752 17119 2810 17125
rect 2752 17085 2764 17119
rect 2798 17116 2810 17119
rect 3697 17119 3755 17125
rect 2798 17088 3280 17116
rect 2798 17085 2810 17088
rect 2752 17079 2810 17085
rect 3252 16992 3280 17088
rect 3697 17085 3709 17119
rect 3743 17116 3755 17119
rect 4126 17116 4154 17156
rect 7098 17144 7104 17156
rect 7156 17144 7162 17196
rect 7650 17144 7656 17196
rect 7708 17184 7714 17196
rect 7929 17187 7987 17193
rect 7929 17184 7941 17187
rect 7708 17156 7941 17184
rect 7708 17144 7714 17156
rect 7929 17153 7941 17156
rect 7975 17153 7987 17187
rect 7929 17147 7987 17153
rect 10686 17144 10692 17196
rect 10744 17184 10750 17196
rect 10873 17187 10931 17193
rect 10873 17184 10885 17187
rect 10744 17156 10885 17184
rect 10744 17144 10750 17156
rect 10873 17153 10885 17156
rect 10919 17184 10931 17187
rect 10962 17184 10968 17196
rect 10919 17156 10968 17184
rect 10919 17153 10931 17156
rect 10873 17147 10931 17153
rect 10962 17144 10968 17156
rect 11020 17144 11026 17196
rect 11146 17184 11152 17196
rect 11107 17156 11152 17184
rect 11146 17144 11152 17156
rect 11204 17184 11210 17196
rect 12805 17187 12863 17193
rect 12805 17184 12817 17187
rect 11204 17156 12817 17184
rect 11204 17144 11210 17156
rect 12805 17153 12817 17156
rect 12851 17153 12863 17187
rect 12805 17147 12863 17153
rect 14093 17187 14151 17193
rect 14093 17153 14105 17187
rect 14139 17184 14151 17187
rect 14182 17184 14188 17196
rect 14139 17156 14188 17184
rect 14139 17153 14151 17156
rect 14093 17147 14151 17153
rect 14182 17144 14188 17156
rect 14240 17184 14246 17196
rect 15562 17184 15568 17196
rect 14240 17156 15568 17184
rect 14240 17144 14246 17156
rect 15562 17144 15568 17156
rect 15620 17144 15626 17196
rect 20070 17144 20076 17196
rect 20128 17184 20134 17196
rect 20809 17187 20867 17193
rect 20809 17184 20821 17187
rect 20128 17156 20821 17184
rect 20128 17144 20134 17156
rect 20809 17153 20821 17156
rect 20855 17184 20867 17187
rect 21266 17184 21272 17196
rect 20855 17156 21272 17184
rect 20855 17153 20867 17156
rect 20809 17147 20867 17153
rect 21266 17144 21272 17156
rect 21324 17144 21330 17196
rect 21468 17184 21496 17224
rect 22557 17187 22615 17193
rect 22557 17184 22569 17187
rect 21468 17156 22569 17184
rect 22557 17153 22569 17156
rect 22603 17153 22615 17187
rect 22557 17147 22615 17153
rect 3743 17088 4154 17116
rect 3743 17085 3755 17088
rect 3697 17079 3755 17085
rect 4614 17076 4620 17128
rect 4672 17116 4678 17128
rect 4709 17119 4767 17125
rect 4709 17116 4721 17119
rect 4672 17088 4721 17116
rect 4672 17076 4678 17088
rect 4709 17085 4721 17088
rect 4755 17085 4767 17119
rect 4709 17079 4767 17085
rect 6892 17119 6950 17125
rect 6892 17085 6904 17119
rect 6938 17116 6950 17119
rect 6938 17088 7420 17116
rect 6938 17085 6950 17088
rect 6892 17079 6950 17085
rect 3605 17051 3663 17057
rect 3605 17017 3617 17051
rect 3651 17048 3663 17051
rect 3651 17020 3924 17048
rect 3651 17017 3663 17020
rect 3605 17011 3663 17017
rect 3234 16980 3240 16992
rect 3195 16952 3240 16980
rect 3234 16940 3240 16952
rect 3292 16940 3298 16992
rect 3896 16980 3924 17020
rect 7392 16992 7420 17088
rect 8570 17076 8576 17128
rect 8628 17116 8634 17128
rect 9677 17119 9735 17125
rect 9677 17116 9689 17119
rect 8628 17088 9689 17116
rect 8628 17076 8634 17088
rect 9677 17085 9689 17088
rect 9723 17116 9735 17119
rect 10137 17119 10195 17125
rect 10137 17116 10149 17119
rect 9723 17088 10149 17116
rect 9723 17085 9735 17088
rect 9677 17079 9735 17085
rect 10137 17085 10149 17088
rect 10183 17085 10195 17119
rect 14734 17116 14740 17128
rect 14695 17088 14740 17116
rect 10137 17079 10195 17085
rect 14734 17076 14740 17088
rect 14792 17076 14798 17128
rect 16482 17116 16488 17128
rect 16443 17088 16488 17116
rect 16482 17076 16488 17088
rect 16540 17116 16546 17128
rect 16945 17119 17003 17125
rect 16945 17116 16957 17119
rect 16540 17088 16957 17116
rect 16540 17076 16546 17088
rect 16945 17085 16957 17088
rect 16991 17085 17003 17119
rect 16945 17079 17003 17085
rect 18693 17119 18751 17125
rect 18693 17085 18705 17119
rect 18739 17116 18751 17119
rect 19334 17116 19340 17128
rect 18739 17088 19340 17116
rect 18739 17085 18751 17088
rect 18693 17079 18751 17085
rect 19334 17076 19340 17088
rect 19392 17076 19398 17128
rect 22005 17119 22063 17125
rect 22005 17085 22017 17119
rect 22051 17085 22063 17119
rect 22462 17116 22468 17128
rect 22423 17088 22468 17116
rect 22005 17079 22063 17085
rect 7837 17051 7895 17057
rect 7837 17017 7849 17051
rect 7883 17048 7895 17051
rect 8018 17048 8024 17060
rect 7883 17020 8024 17048
rect 7883 17017 7895 17020
rect 7837 17011 7895 17017
rect 8018 17008 8024 17020
rect 8076 17048 8082 17060
rect 8291 17051 8349 17057
rect 8291 17048 8303 17051
rect 8076 17020 8303 17048
rect 8076 17008 8082 17020
rect 8291 17017 8303 17020
rect 8337 17048 8349 17051
rect 8754 17048 8760 17060
rect 8337 17020 8760 17048
rect 8337 17017 8349 17020
rect 8291 17011 8349 17017
rect 8754 17008 8760 17020
rect 8812 17008 8818 17060
rect 10962 17008 10968 17060
rect 11020 17048 11026 17060
rect 12526 17048 12532 17060
rect 11020 17020 11065 17048
rect 12487 17020 12532 17048
rect 11020 17008 11026 17020
rect 12526 17008 12532 17020
rect 12584 17008 12590 17060
rect 12621 17051 12679 17057
rect 12621 17017 12633 17051
rect 12667 17017 12679 17051
rect 12621 17011 12679 17017
rect 4246 16980 4252 16992
rect 3896 16952 4252 16980
rect 4246 16940 4252 16952
rect 4304 16940 4310 16992
rect 4525 16983 4583 16989
rect 4525 16949 4537 16983
rect 4571 16980 4583 16983
rect 4798 16980 4804 16992
rect 4571 16952 4804 16980
rect 4571 16949 4583 16952
rect 4525 16943 4583 16949
rect 4798 16940 4804 16952
rect 4856 16980 4862 16992
rect 5074 16980 5080 16992
rect 4856 16952 5080 16980
rect 4856 16940 4862 16952
rect 5074 16940 5080 16952
rect 5132 16940 5138 16992
rect 6822 16940 6828 16992
rect 6880 16980 6886 16992
rect 6963 16983 7021 16989
rect 6963 16980 6975 16983
rect 6880 16952 6975 16980
rect 6880 16940 6886 16952
rect 6963 16949 6975 16952
rect 7009 16949 7021 16983
rect 7374 16980 7380 16992
rect 7335 16952 7380 16980
rect 6963 16943 7021 16949
rect 7374 16940 7380 16952
rect 7432 16940 7438 16992
rect 12342 16940 12348 16992
rect 12400 16980 12406 16992
rect 12636 16980 12664 17011
rect 14642 17008 14648 17060
rect 14700 17048 14706 17060
rect 15058 17051 15116 17057
rect 15058 17048 15070 17051
rect 14700 17020 15070 17048
rect 14700 17008 14706 17020
rect 15058 17017 15070 17020
rect 15104 17048 15116 17051
rect 15470 17048 15476 17060
rect 15104 17020 15476 17048
rect 15104 17017 15116 17020
rect 15058 17011 15116 17017
rect 15470 17008 15476 17020
rect 15528 17048 15534 17060
rect 15933 17051 15991 17057
rect 15933 17048 15945 17051
rect 15528 17020 15945 17048
rect 15528 17008 15534 17020
rect 15933 17017 15945 17020
rect 15979 17017 15991 17051
rect 19014 17051 19072 17057
rect 19014 17048 19026 17051
rect 15933 17011 15991 17017
rect 18524 17020 19026 17048
rect 12400 16952 12664 16980
rect 12400 16940 12406 16952
rect 13262 16940 13268 16992
rect 13320 16980 13326 16992
rect 13630 16980 13636 16992
rect 13320 16952 13636 16980
rect 13320 16940 13326 16952
rect 13630 16940 13636 16952
rect 13688 16940 13694 16992
rect 16669 16983 16727 16989
rect 16669 16949 16681 16983
rect 16715 16980 16727 16983
rect 16942 16980 16948 16992
rect 16715 16952 16948 16980
rect 16715 16949 16727 16952
rect 16669 16943 16727 16949
rect 16942 16940 16948 16952
rect 17000 16940 17006 16992
rect 17497 16983 17555 16989
rect 17497 16949 17509 16983
rect 17543 16980 17555 16983
rect 17678 16980 17684 16992
rect 17543 16952 17684 16980
rect 17543 16949 17555 16952
rect 17497 16943 17555 16949
rect 17678 16940 17684 16952
rect 17736 16940 17742 16992
rect 17770 16940 17776 16992
rect 17828 16980 17834 16992
rect 18524 16989 18552 17020
rect 19014 17017 19026 17020
rect 19060 17017 19072 17051
rect 20530 17048 20536 17060
rect 20491 17020 20536 17048
rect 19014 17011 19072 17017
rect 20530 17008 20536 17020
rect 20588 17008 20594 17060
rect 20625 17051 20683 17057
rect 20625 17017 20637 17051
rect 20671 17017 20683 17051
rect 20625 17011 20683 17017
rect 21269 17051 21327 17057
rect 21269 17017 21281 17051
rect 21315 17048 21327 17051
rect 21821 17051 21879 17057
rect 21821 17048 21833 17051
rect 21315 17020 21833 17048
rect 21315 17017 21327 17020
rect 21269 17011 21327 17017
rect 21821 17017 21833 17020
rect 21867 17048 21879 17051
rect 22020 17048 22048 17079
rect 22462 17076 22468 17088
rect 22520 17076 22526 17128
rect 23728 17119 23786 17125
rect 23728 17085 23740 17119
rect 23774 17116 23786 17119
rect 24118 17116 24124 17128
rect 23774 17088 24124 17116
rect 23774 17085 23786 17088
rect 23728 17079 23786 17085
rect 24118 17076 24124 17088
rect 24176 17076 24182 17128
rect 23290 17048 23296 17060
rect 21867 17020 23296 17048
rect 21867 17017 21879 17020
rect 21821 17011 21879 17017
rect 18509 16983 18567 16989
rect 18509 16980 18521 16983
rect 17828 16952 18521 16980
rect 17828 16940 17834 16952
rect 18509 16949 18521 16952
rect 18555 16949 18567 16983
rect 18509 16943 18567 16949
rect 19613 16983 19671 16989
rect 19613 16949 19625 16983
rect 19659 16980 19671 16983
rect 20257 16983 20315 16989
rect 20257 16980 20269 16983
rect 19659 16952 20269 16980
rect 19659 16949 19671 16952
rect 19613 16943 19671 16949
rect 20257 16949 20269 16952
rect 20303 16980 20315 16983
rect 20640 16980 20668 17011
rect 23290 17008 23296 17020
rect 23348 17008 23354 17060
rect 20303 16952 20668 16980
rect 20303 16949 20315 16952
rect 20257 16943 20315 16949
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 4801 16779 4859 16785
rect 4801 16745 4813 16779
rect 4847 16776 4859 16779
rect 5074 16776 5080 16788
rect 4847 16748 5080 16776
rect 4847 16745 4859 16748
rect 4801 16739 4859 16745
rect 5074 16736 5080 16748
rect 5132 16776 5138 16788
rect 8018 16776 8024 16788
rect 5132 16748 8024 16776
rect 5132 16736 5138 16748
rect 8018 16736 8024 16748
rect 8076 16736 8082 16788
rect 8202 16776 8208 16788
rect 8163 16748 8208 16776
rect 8202 16736 8208 16748
rect 8260 16736 8266 16788
rect 10505 16779 10563 16785
rect 10505 16745 10517 16779
rect 10551 16776 10563 16779
rect 10686 16776 10692 16788
rect 10551 16748 10692 16776
rect 10551 16745 10563 16748
rect 10505 16739 10563 16745
rect 10686 16736 10692 16748
rect 10744 16736 10750 16788
rect 12434 16776 12440 16788
rect 12395 16748 12440 16776
rect 12434 16736 12440 16748
rect 12492 16736 12498 16788
rect 14734 16776 14740 16788
rect 14695 16748 14740 16776
rect 14734 16736 14740 16748
rect 14792 16736 14798 16788
rect 15746 16736 15752 16788
rect 15804 16776 15810 16788
rect 16209 16779 16267 16785
rect 16209 16776 16221 16779
rect 15804 16748 16221 16776
rect 15804 16736 15810 16748
rect 16209 16745 16221 16748
rect 16255 16745 16267 16779
rect 16209 16739 16267 16745
rect 16298 16736 16304 16788
rect 16356 16776 16362 16788
rect 16485 16779 16543 16785
rect 16485 16776 16497 16779
rect 16356 16748 16497 16776
rect 16356 16736 16362 16748
rect 16485 16745 16497 16748
rect 16531 16745 16543 16779
rect 16485 16739 16543 16745
rect 18969 16779 19027 16785
rect 18969 16745 18981 16779
rect 19015 16776 19027 16779
rect 19242 16776 19248 16788
rect 19015 16748 19248 16776
rect 19015 16745 19027 16748
rect 18969 16739 19027 16745
rect 19242 16736 19248 16748
rect 19300 16736 19306 16788
rect 19334 16736 19340 16788
rect 19392 16776 19398 16788
rect 20993 16779 21051 16785
rect 20993 16776 21005 16779
rect 19392 16748 21005 16776
rect 19392 16736 19398 16748
rect 20993 16745 21005 16748
rect 21039 16745 21051 16779
rect 20993 16739 21051 16745
rect 21174 16736 21180 16788
rect 21232 16776 21238 16788
rect 22005 16779 22063 16785
rect 22005 16776 22017 16779
rect 21232 16748 22017 16776
rect 21232 16736 21238 16748
rect 22005 16745 22017 16748
rect 22051 16776 22063 16779
rect 22462 16776 22468 16788
rect 22051 16748 22468 16776
rect 22051 16745 22063 16748
rect 22005 16739 22063 16745
rect 22462 16736 22468 16748
rect 22520 16776 22526 16788
rect 22520 16748 22784 16776
rect 22520 16736 22526 16748
rect 5166 16708 5172 16720
rect 5127 16680 5172 16708
rect 5166 16668 5172 16680
rect 5224 16668 5230 16720
rect 7650 16668 7656 16720
rect 7708 16708 7714 16720
rect 8573 16711 8631 16717
rect 8573 16708 8585 16711
rect 7708 16680 8585 16708
rect 7708 16668 7714 16680
rect 8573 16677 8585 16680
rect 8619 16677 8631 16711
rect 8573 16671 8631 16677
rect 11511 16711 11569 16717
rect 11511 16677 11523 16711
rect 11557 16708 11569 16711
rect 11606 16708 11612 16720
rect 11557 16680 11612 16708
rect 11557 16677 11569 16680
rect 11511 16671 11569 16677
rect 11606 16668 11612 16680
rect 11664 16668 11670 16720
rect 15470 16668 15476 16720
rect 15528 16708 15534 16720
rect 15610 16711 15668 16717
rect 15610 16708 15622 16711
rect 15528 16680 15622 16708
rect 15528 16668 15534 16680
rect 15610 16677 15622 16680
rect 15656 16677 15668 16711
rect 15610 16671 15668 16677
rect 17770 16668 17776 16720
rect 17828 16708 17834 16720
rect 18370 16711 18428 16717
rect 18370 16708 18382 16711
rect 17828 16680 18382 16708
rect 17828 16668 17834 16680
rect 18370 16677 18382 16680
rect 18416 16677 18428 16711
rect 18370 16671 18428 16677
rect 20717 16711 20775 16717
rect 20717 16677 20729 16711
rect 20763 16708 20775 16711
rect 20806 16708 20812 16720
rect 20763 16680 20812 16708
rect 20763 16677 20775 16680
rect 20717 16671 20775 16677
rect 20806 16668 20812 16680
rect 20864 16668 20870 16720
rect 21100 16680 22508 16708
rect 21100 16652 21128 16680
rect 1740 16643 1798 16649
rect 1740 16609 1752 16643
rect 1786 16640 1798 16643
rect 2038 16640 2044 16652
rect 1786 16612 2044 16640
rect 1786 16609 1798 16612
rect 1740 16603 1798 16609
rect 2038 16600 2044 16612
rect 2096 16600 2102 16652
rect 7282 16640 7288 16652
rect 7243 16612 7288 16640
rect 7282 16600 7288 16612
rect 7340 16600 7346 16652
rect 9582 16640 9588 16652
rect 9543 16612 9588 16640
rect 9582 16600 9588 16612
rect 9640 16600 9646 16652
rect 10873 16643 10931 16649
rect 10873 16609 10885 16643
rect 10919 16640 10931 16643
rect 10962 16640 10968 16652
rect 10919 16612 10968 16640
rect 10919 16609 10931 16612
rect 10873 16603 10931 16609
rect 10962 16600 10968 16612
rect 11020 16640 11026 16652
rect 12069 16643 12127 16649
rect 12069 16640 12081 16643
rect 11020 16612 12081 16640
rect 11020 16600 11026 16612
rect 12069 16609 12081 16612
rect 12115 16609 12127 16643
rect 12069 16603 12127 16609
rect 12618 16600 12624 16652
rect 12676 16640 12682 16652
rect 12897 16643 12955 16649
rect 12897 16640 12909 16643
rect 12676 16612 12909 16640
rect 12676 16600 12682 16612
rect 12897 16609 12909 16612
rect 12943 16609 12955 16643
rect 13354 16640 13360 16652
rect 13315 16612 13360 16640
rect 12897 16603 12955 16609
rect 13354 16600 13360 16612
rect 13412 16600 13418 16652
rect 15286 16640 15292 16652
rect 15199 16612 15292 16640
rect 15286 16600 15292 16612
rect 15344 16640 15350 16652
rect 19864 16643 19922 16649
rect 15344 16612 18322 16640
rect 15344 16600 15350 16612
rect 2961 16575 3019 16581
rect 2961 16541 2973 16575
rect 3007 16572 3019 16575
rect 4430 16572 4436 16584
rect 3007 16544 4436 16572
rect 3007 16541 3019 16544
rect 2961 16535 3019 16541
rect 4430 16532 4436 16544
rect 4488 16572 4494 16584
rect 5077 16575 5135 16581
rect 5077 16572 5089 16575
rect 4488 16544 5089 16572
rect 4488 16532 4494 16544
rect 5077 16541 5089 16544
rect 5123 16541 5135 16575
rect 5534 16572 5540 16584
rect 5495 16544 5540 16572
rect 5077 16535 5135 16541
rect 5534 16532 5540 16544
rect 5592 16532 5598 16584
rect 11149 16575 11207 16581
rect 11149 16541 11161 16575
rect 11195 16572 11207 16575
rect 11238 16572 11244 16584
rect 11195 16544 11244 16572
rect 11195 16541 11207 16544
rect 11149 16535 11207 16541
rect 11238 16532 11244 16544
rect 11296 16572 11302 16584
rect 13449 16575 13507 16581
rect 13449 16572 13461 16575
rect 11296 16544 13461 16572
rect 11296 16532 11302 16544
rect 13449 16541 13461 16544
rect 13495 16541 13507 16575
rect 13449 16535 13507 16541
rect 17494 16532 17500 16584
rect 17552 16572 17558 16584
rect 18049 16575 18107 16581
rect 18049 16572 18061 16575
rect 17552 16544 18061 16572
rect 17552 16532 17558 16544
rect 18049 16541 18061 16544
rect 18095 16541 18107 16575
rect 18294 16572 18322 16612
rect 19864 16609 19876 16643
rect 19910 16640 19922 16643
rect 20070 16640 20076 16652
rect 19910 16612 20076 16640
rect 19910 16609 19922 16612
rect 19864 16603 19922 16609
rect 20070 16600 20076 16612
rect 20128 16600 20134 16652
rect 21082 16640 21088 16652
rect 21043 16612 21088 16640
rect 21082 16600 21088 16612
rect 21140 16600 21146 16652
rect 21358 16600 21364 16652
rect 21416 16640 21422 16652
rect 21453 16643 21511 16649
rect 21453 16640 21465 16643
rect 21416 16612 21465 16640
rect 21416 16600 21422 16612
rect 21453 16609 21465 16612
rect 21499 16640 21511 16643
rect 21818 16640 21824 16652
rect 21499 16612 21824 16640
rect 21499 16609 21511 16612
rect 21453 16603 21511 16609
rect 21818 16600 21824 16612
rect 21876 16600 21882 16652
rect 22480 16649 22508 16680
rect 22465 16643 22523 16649
rect 22465 16609 22477 16643
rect 22511 16640 22523 16643
rect 22646 16640 22652 16652
rect 22511 16612 22652 16640
rect 22511 16609 22523 16612
rect 22465 16603 22523 16609
rect 22646 16600 22652 16612
rect 22704 16600 22710 16652
rect 22756 16640 22784 16748
rect 22922 16640 22928 16652
rect 22756 16612 22928 16640
rect 22922 16600 22928 16612
rect 22980 16600 22986 16652
rect 23017 16575 23075 16581
rect 23017 16572 23029 16575
rect 18294 16544 23029 16572
rect 18049 16535 18107 16541
rect 23017 16541 23029 16544
rect 23063 16541 23075 16575
rect 23017 16535 23075 16541
rect 1670 16464 1676 16516
rect 1728 16504 1734 16516
rect 9306 16504 9312 16516
rect 1728 16476 9312 16504
rect 1728 16464 1734 16476
rect 9306 16464 9312 16476
rect 9364 16464 9370 16516
rect 12710 16464 12716 16516
rect 12768 16504 12774 16516
rect 15746 16504 15752 16516
rect 12768 16476 15752 16504
rect 12768 16464 12774 16476
rect 15746 16464 15752 16476
rect 15804 16464 15810 16516
rect 1394 16396 1400 16448
rect 1452 16436 1458 16448
rect 1811 16439 1869 16445
rect 1811 16436 1823 16439
rect 1452 16408 1823 16436
rect 1452 16396 1458 16408
rect 1811 16405 1823 16408
rect 1857 16405 1869 16439
rect 1811 16399 1869 16405
rect 4433 16439 4491 16445
rect 4433 16405 4445 16439
rect 4479 16436 4491 16439
rect 4614 16436 4620 16448
rect 4479 16408 4620 16436
rect 4479 16405 4491 16408
rect 4433 16399 4491 16405
rect 4614 16396 4620 16408
rect 4672 16396 4678 16448
rect 7466 16436 7472 16448
rect 7427 16408 7472 16436
rect 7466 16396 7472 16408
rect 7524 16396 7530 16448
rect 9815 16439 9873 16445
rect 9815 16405 9827 16439
rect 9861 16436 9873 16439
rect 10134 16436 10140 16448
rect 9861 16408 10140 16436
rect 9861 16405 9873 16408
rect 9815 16399 9873 16405
rect 10134 16396 10140 16408
rect 10192 16396 10198 16448
rect 13906 16436 13912 16448
rect 13867 16408 13912 16436
rect 13906 16396 13912 16408
rect 13964 16396 13970 16448
rect 16942 16436 16948 16448
rect 16903 16408 16948 16436
rect 16942 16396 16948 16408
rect 17000 16396 17006 16448
rect 19610 16436 19616 16448
rect 19571 16408 19616 16436
rect 19610 16396 19616 16408
rect 19668 16396 19674 16448
rect 19935 16439 19993 16445
rect 19935 16405 19947 16439
rect 19981 16436 19993 16439
rect 20070 16436 20076 16448
rect 19981 16408 20076 16436
rect 19981 16405 19993 16408
rect 19935 16399 19993 16405
rect 20070 16396 20076 16408
rect 20128 16396 20134 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 2038 16232 2044 16244
rect 1999 16204 2044 16232
rect 2038 16192 2044 16204
rect 2096 16192 2102 16244
rect 4430 16232 4436 16244
rect 4391 16204 4436 16232
rect 4430 16192 4436 16204
rect 4488 16192 4494 16244
rect 4801 16235 4859 16241
rect 4801 16201 4813 16235
rect 4847 16232 4859 16235
rect 5166 16232 5172 16244
rect 4847 16204 5172 16232
rect 4847 16201 4859 16204
rect 4801 16195 4859 16201
rect 4617 16167 4675 16173
rect 4617 16164 4629 16167
rect 3988 16136 4629 16164
rect 1394 16028 1400 16040
rect 1355 16000 1400 16028
rect 1394 15988 1400 16000
rect 1452 15988 1458 16040
rect 3988 16037 4016 16136
rect 4617 16133 4629 16136
rect 4663 16133 4675 16167
rect 4617 16127 4675 16133
rect 4065 16099 4123 16105
rect 4065 16065 4077 16099
rect 4111 16096 4123 16099
rect 4816 16096 4844 16195
rect 5166 16192 5172 16204
rect 5224 16192 5230 16244
rect 7098 16232 7104 16244
rect 7059 16204 7104 16232
rect 7098 16192 7104 16204
rect 7156 16192 7162 16244
rect 7466 16232 7472 16244
rect 7427 16204 7472 16232
rect 7466 16192 7472 16204
rect 7524 16192 7530 16244
rect 9582 16192 9588 16244
rect 9640 16232 9646 16244
rect 10229 16235 10287 16241
rect 10229 16232 10241 16235
rect 9640 16204 10241 16232
rect 9640 16192 9646 16204
rect 10229 16201 10241 16204
rect 10275 16201 10287 16235
rect 10229 16195 10287 16201
rect 11606 16192 11612 16244
rect 11664 16232 11670 16244
rect 11793 16235 11851 16241
rect 11793 16232 11805 16235
rect 11664 16204 11805 16232
rect 11664 16192 11670 16204
rect 11793 16201 11805 16204
rect 11839 16201 11851 16235
rect 11793 16195 11851 16201
rect 12621 16235 12679 16241
rect 12621 16201 12633 16235
rect 12667 16232 12679 16235
rect 12894 16232 12900 16244
rect 12667 16204 12900 16232
rect 12667 16201 12679 16204
rect 12621 16195 12679 16201
rect 12894 16192 12900 16204
rect 12952 16192 12958 16244
rect 15013 16235 15071 16241
rect 15013 16201 15025 16235
rect 15059 16232 15071 16235
rect 15286 16232 15292 16244
rect 15059 16204 15292 16232
rect 15059 16201 15071 16204
rect 15013 16195 15071 16201
rect 15286 16192 15292 16204
rect 15344 16192 15350 16244
rect 15470 16192 15476 16244
rect 15528 16232 15534 16244
rect 15930 16232 15936 16244
rect 15528 16204 15936 16232
rect 15528 16192 15534 16204
rect 15930 16192 15936 16204
rect 15988 16192 15994 16244
rect 17494 16232 17500 16244
rect 17455 16204 17500 16232
rect 17494 16192 17500 16204
rect 17552 16192 17558 16244
rect 18966 16232 18972 16244
rect 18927 16204 18972 16232
rect 18966 16192 18972 16204
rect 19024 16192 19030 16244
rect 20162 16232 20168 16244
rect 20123 16204 20168 16232
rect 20162 16192 20168 16204
rect 20220 16192 20226 16244
rect 21358 16232 21364 16244
rect 21319 16204 21364 16232
rect 21358 16192 21364 16204
rect 21416 16192 21422 16244
rect 22646 16232 22652 16244
rect 22607 16204 22652 16232
rect 22646 16192 22652 16204
rect 22704 16192 22710 16244
rect 22922 16192 22928 16244
rect 22980 16232 22986 16244
rect 23017 16235 23075 16241
rect 23017 16232 23029 16235
rect 22980 16204 23029 16232
rect 22980 16192 22986 16204
rect 23017 16201 23029 16204
rect 23063 16201 23075 16235
rect 23017 16195 23075 16201
rect 5534 16164 5540 16176
rect 5495 16136 5540 16164
rect 5534 16124 5540 16136
rect 5592 16124 5598 16176
rect 4982 16096 4988 16108
rect 4111 16068 4844 16096
rect 4895 16068 4988 16096
rect 4111 16065 4123 16068
rect 4065 16059 4123 16065
rect 4982 16056 4988 16068
rect 5040 16096 5046 16108
rect 5905 16099 5963 16105
rect 5905 16096 5917 16099
rect 5040 16068 5917 16096
rect 5040 16056 5046 16068
rect 5905 16065 5917 16068
rect 5951 16065 5963 16099
rect 7116 16096 7144 16192
rect 9861 16167 9919 16173
rect 9861 16133 9873 16167
rect 9907 16164 9919 16167
rect 11425 16167 11483 16173
rect 11425 16164 11437 16167
rect 9907 16136 11437 16164
rect 9907 16133 9919 16136
rect 9861 16127 9919 16133
rect 11425 16133 11437 16136
rect 11471 16164 11483 16167
rect 14182 16164 14188 16176
rect 11471 16136 14188 16164
rect 11471 16133 11483 16136
rect 11425 16127 11483 16133
rect 14182 16124 14188 16136
rect 14240 16124 14246 16176
rect 7745 16099 7803 16105
rect 7745 16096 7757 16099
rect 7116 16068 7757 16096
rect 5905 16059 5963 16065
rect 7745 16065 7757 16068
rect 7791 16065 7803 16099
rect 9306 16096 9312 16108
rect 9267 16068 9312 16096
rect 7745 16059 7803 16065
rect 9306 16056 9312 16068
rect 9364 16056 9370 16108
rect 10873 16099 10931 16105
rect 10873 16065 10885 16099
rect 10919 16096 10931 16099
rect 11054 16096 11060 16108
rect 10919 16068 11060 16096
rect 10919 16065 10931 16068
rect 10873 16059 10931 16065
rect 11054 16056 11060 16068
rect 11112 16056 11118 16108
rect 12253 16099 12311 16105
rect 12253 16065 12265 16099
rect 12299 16096 12311 16099
rect 13354 16096 13360 16108
rect 12299 16068 13360 16096
rect 12299 16065 12311 16068
rect 12253 16059 12311 16065
rect 13354 16056 13360 16068
rect 13412 16056 13418 16108
rect 17129 16099 17187 16105
rect 17129 16065 17141 16099
rect 17175 16096 17187 16099
rect 17512 16096 17540 16192
rect 19518 16124 19524 16176
rect 19576 16164 19582 16176
rect 19797 16167 19855 16173
rect 19797 16164 19809 16167
rect 19576 16136 19809 16164
rect 19576 16124 19582 16136
rect 19797 16133 19809 16136
rect 19843 16133 19855 16167
rect 19797 16127 19855 16133
rect 17175 16068 17540 16096
rect 18279 16099 18337 16105
rect 17175 16065 17187 16068
rect 17129 16059 17187 16065
rect 18279 16065 18291 16099
rect 18325 16096 18337 16099
rect 19245 16099 19303 16105
rect 19245 16096 19257 16099
rect 18325 16068 19257 16096
rect 18325 16065 18337 16068
rect 18279 16059 18337 16065
rect 19245 16065 19257 16068
rect 19291 16096 19303 16099
rect 19610 16096 19616 16108
rect 19291 16068 19616 16096
rect 19291 16065 19303 16068
rect 19245 16059 19303 16065
rect 19610 16056 19616 16068
rect 19668 16056 19674 16108
rect 21729 16099 21787 16105
rect 21729 16065 21741 16099
rect 21775 16096 21787 16099
rect 22186 16096 22192 16108
rect 21775 16068 22192 16096
rect 21775 16065 21787 16068
rect 21729 16059 21787 16065
rect 22186 16056 22192 16068
rect 22244 16056 22250 16108
rect 3237 16031 3295 16037
rect 3237 15997 3249 16031
rect 3283 16028 3295 16031
rect 3973 16031 4031 16037
rect 3973 16028 3985 16031
rect 3283 16000 3985 16028
rect 3283 15997 3295 16000
rect 3237 15991 3295 15997
rect 3973 15997 3985 16000
rect 4019 15997 4031 16031
rect 3973 15991 4031 15997
rect 12342 15988 12348 16040
rect 12400 16028 12406 16040
rect 12437 16031 12495 16037
rect 12437 16028 12449 16031
rect 12400 16000 12449 16028
rect 12400 15988 12406 16000
rect 12437 15997 12449 16000
rect 12483 15997 12495 16031
rect 12437 15991 12495 15997
rect 4617 15963 4675 15969
rect 4617 15929 4629 15963
rect 4663 15960 4675 15963
rect 5077 15963 5135 15969
rect 5077 15960 5089 15963
rect 4663 15932 5089 15960
rect 4663 15929 4675 15932
rect 4617 15923 4675 15929
rect 5077 15929 5089 15932
rect 5123 15960 5135 15963
rect 5258 15960 5264 15972
rect 5123 15932 5264 15960
rect 5123 15929 5135 15932
rect 5077 15923 5135 15929
rect 5258 15920 5264 15932
rect 5316 15920 5322 15972
rect 7837 15963 7895 15969
rect 7837 15929 7849 15963
rect 7883 15929 7895 15963
rect 7837 15923 7895 15929
rect 8389 15963 8447 15969
rect 8389 15929 8401 15963
rect 8435 15960 8447 15963
rect 8478 15960 8484 15972
rect 8435 15932 8484 15960
rect 8435 15929 8447 15932
rect 8389 15923 8447 15929
rect 198 15852 204 15904
rect 256 15892 262 15904
rect 1581 15895 1639 15901
rect 1581 15892 1593 15895
rect 256 15864 1593 15892
rect 256 15852 262 15864
rect 1581 15861 1593 15864
rect 1627 15861 1639 15895
rect 1581 15855 1639 15861
rect 7466 15852 7472 15904
rect 7524 15892 7530 15904
rect 7852 15892 7880 15923
rect 8478 15920 8484 15932
rect 8536 15920 8542 15972
rect 9398 15920 9404 15972
rect 9456 15960 9462 15972
rect 10965 15963 11023 15969
rect 9456 15932 9501 15960
rect 9456 15920 9462 15932
rect 10965 15929 10977 15963
rect 11011 15929 11023 15963
rect 12452 15960 12480 15991
rect 12618 15988 12624 16040
rect 12676 16028 12682 16040
rect 12897 16031 12955 16037
rect 12897 16028 12909 16031
rect 12676 16000 12909 16028
rect 12676 15988 12682 16000
rect 12897 15997 12909 16000
rect 12943 15997 12955 16031
rect 12897 15991 12955 15997
rect 14642 15988 14648 16040
rect 14700 16028 14706 16040
rect 15140 16031 15198 16037
rect 15140 16028 15152 16031
rect 14700 16000 15152 16028
rect 14700 15988 14706 16000
rect 15140 15997 15152 16000
rect 15186 16028 15198 16031
rect 15565 16031 15623 16037
rect 15565 16028 15577 16031
rect 15186 16000 15577 16028
rect 15186 15997 15198 16000
rect 15140 15991 15198 15997
rect 15565 15997 15577 16000
rect 15611 15997 15623 16031
rect 15565 15991 15623 15997
rect 16298 15988 16304 16040
rect 16356 16028 16362 16040
rect 16393 16031 16451 16037
rect 16393 16028 16405 16031
rect 16356 16000 16405 16028
rect 16356 15988 16362 16000
rect 16393 15997 16405 16000
rect 16439 15997 16451 16031
rect 16942 16028 16948 16040
rect 16855 16000 16948 16028
rect 16393 15991 16451 15997
rect 16942 15988 16948 16000
rect 17000 15988 17006 16040
rect 18192 16031 18250 16037
rect 18192 15997 18204 16031
rect 18238 16028 18250 16031
rect 18598 16028 18604 16040
rect 18238 16000 18604 16028
rect 18238 15997 18250 16000
rect 18192 15991 18250 15997
rect 18598 15988 18604 16000
rect 18656 15988 18662 16040
rect 13265 15963 13323 15969
rect 13265 15960 13277 15963
rect 12452 15932 13277 15960
rect 10965 15923 11023 15929
rect 13265 15929 13277 15932
rect 13311 15929 13323 15963
rect 13265 15923 13323 15929
rect 7524 15864 7880 15892
rect 9125 15895 9183 15901
rect 7524 15852 7530 15864
rect 9125 15861 9137 15895
rect 9171 15892 9183 15895
rect 9416 15892 9444 15920
rect 10686 15892 10692 15904
rect 9171 15864 9444 15892
rect 10647 15864 10692 15892
rect 9171 15861 9183 15864
rect 9125 15855 9183 15861
rect 10686 15852 10692 15864
rect 10744 15892 10750 15904
rect 10980 15892 11008 15923
rect 13446 15920 13452 15972
rect 13504 15960 13510 15972
rect 13633 15963 13691 15969
rect 13633 15960 13645 15963
rect 13504 15932 13645 15960
rect 13504 15920 13510 15932
rect 13633 15929 13645 15932
rect 13679 15929 13691 15963
rect 13633 15923 13691 15929
rect 13725 15963 13783 15969
rect 13725 15929 13737 15963
rect 13771 15960 13783 15963
rect 13906 15960 13912 15972
rect 13771 15932 13912 15960
rect 13771 15929 13783 15932
rect 13725 15923 13783 15929
rect 10744 15864 11008 15892
rect 13648 15892 13676 15923
rect 13906 15920 13912 15932
rect 13964 15920 13970 15972
rect 14277 15963 14335 15969
rect 14277 15929 14289 15963
rect 14323 15960 14335 15963
rect 14734 15960 14740 15972
rect 14323 15932 14740 15960
rect 14323 15929 14335 15932
rect 14277 15923 14335 15929
rect 14734 15920 14740 15932
rect 14792 15920 14798 15972
rect 16960 15960 16988 15988
rect 18322 15960 18328 15972
rect 16960 15932 18328 15960
rect 18322 15920 18328 15932
rect 18380 15920 18386 15972
rect 18966 15920 18972 15972
rect 19024 15960 19030 15972
rect 19337 15963 19395 15969
rect 19337 15960 19349 15963
rect 19024 15932 19349 15960
rect 19024 15920 19030 15932
rect 19337 15929 19349 15932
rect 19383 15929 19395 15963
rect 21818 15960 21824 15972
rect 21779 15932 21824 15960
rect 19337 15923 19395 15929
rect 21818 15920 21824 15932
rect 21876 15920 21882 15972
rect 22373 15963 22431 15969
rect 22373 15929 22385 15963
rect 22419 15960 22431 15963
rect 22830 15960 22836 15972
rect 22419 15932 22836 15960
rect 22419 15929 22431 15932
rect 22373 15923 22431 15929
rect 22830 15920 22836 15932
rect 22888 15920 22894 15972
rect 14553 15895 14611 15901
rect 14553 15892 14565 15895
rect 13648 15864 14565 15892
rect 10744 15852 10750 15864
rect 14553 15861 14565 15864
rect 14599 15861 14611 15895
rect 14553 15855 14611 15861
rect 15243 15895 15301 15901
rect 15243 15861 15255 15895
rect 15289 15892 15301 15895
rect 15470 15892 15476 15904
rect 15289 15864 15476 15892
rect 15289 15861 15301 15864
rect 15243 15855 15301 15861
rect 15470 15852 15476 15864
rect 15528 15852 15534 15904
rect 15930 15852 15936 15904
rect 15988 15892 15994 15904
rect 17770 15892 17776 15904
rect 15988 15864 17776 15892
rect 15988 15852 15994 15864
rect 17770 15852 17776 15864
rect 17828 15852 17834 15904
rect 20993 15895 21051 15901
rect 20993 15861 21005 15895
rect 21039 15892 21051 15895
rect 21082 15892 21088 15904
rect 21039 15864 21088 15892
rect 21039 15861 21051 15864
rect 20993 15855 21051 15861
rect 21082 15852 21088 15864
rect 21140 15852 21146 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1394 15648 1400 15700
rect 1452 15688 1458 15700
rect 1581 15691 1639 15697
rect 1581 15688 1593 15691
rect 1452 15660 1593 15688
rect 1452 15648 1458 15660
rect 1581 15657 1593 15660
rect 1627 15657 1639 15691
rect 5258 15688 5264 15700
rect 5219 15660 5264 15688
rect 1581 15651 1639 15657
rect 5258 15648 5264 15660
rect 5316 15648 5322 15700
rect 7282 15688 7288 15700
rect 7243 15660 7288 15688
rect 7282 15648 7288 15660
rect 7340 15688 7346 15700
rect 7834 15688 7840 15700
rect 7340 15660 7840 15688
rect 7340 15648 7346 15660
rect 7834 15648 7840 15660
rect 7892 15688 7898 15700
rect 9214 15688 9220 15700
rect 7892 15660 7972 15688
rect 9175 15660 9220 15688
rect 7892 15648 7898 15660
rect 4430 15620 4436 15632
rect 4391 15592 4436 15620
rect 4430 15580 4436 15592
rect 4488 15580 4494 15632
rect 4982 15620 4988 15632
rect 4943 15592 4988 15620
rect 4982 15580 4988 15592
rect 5040 15580 5046 15632
rect 6270 15580 6276 15632
rect 6328 15620 6334 15632
rect 7944 15629 7972 15660
rect 9214 15648 9220 15660
rect 9272 15648 9278 15700
rect 11238 15688 11244 15700
rect 11199 15660 11244 15688
rect 11238 15648 11244 15660
rect 11296 15648 11302 15700
rect 17678 15688 17684 15700
rect 17639 15660 17684 15688
rect 17678 15648 17684 15660
rect 17736 15648 17742 15700
rect 19518 15688 19524 15700
rect 19431 15660 19524 15688
rect 6365 15623 6423 15629
rect 6365 15620 6377 15623
rect 6328 15592 6377 15620
rect 6328 15580 6334 15592
rect 6365 15589 6377 15592
rect 6411 15589 6423 15623
rect 6365 15583 6423 15589
rect 7929 15623 7987 15629
rect 7929 15589 7941 15623
rect 7975 15589 7987 15623
rect 8478 15620 8484 15632
rect 8439 15592 8484 15620
rect 7929 15583 7987 15589
rect 8478 15580 8484 15592
rect 8536 15580 8542 15632
rect 10134 15620 10140 15632
rect 10095 15592 10140 15620
rect 10134 15580 10140 15592
rect 10192 15580 10198 15632
rect 10229 15623 10287 15629
rect 10229 15589 10241 15623
rect 10275 15620 10287 15623
rect 10594 15620 10600 15632
rect 10275 15592 10600 15620
rect 10275 15589 10287 15592
rect 10229 15583 10287 15589
rect 10594 15580 10600 15592
rect 10652 15580 10658 15632
rect 11054 15580 11060 15632
rect 11112 15620 11118 15632
rect 11517 15623 11575 15629
rect 11517 15620 11529 15623
rect 11112 15592 11529 15620
rect 11112 15580 11118 15592
rect 11517 15589 11529 15592
rect 11563 15589 11575 15623
rect 13170 15620 13176 15632
rect 13131 15592 13176 15620
rect 11517 15583 11575 15589
rect 13170 15580 13176 15592
rect 13228 15580 13234 15632
rect 15930 15580 15936 15632
rect 15988 15620 15994 15632
rect 19444 15629 19472 15660
rect 19518 15648 19524 15660
rect 19576 15688 19582 15700
rect 21818 15688 21824 15700
rect 19576 15660 21824 15688
rect 19576 15648 19582 15660
rect 21818 15648 21824 15660
rect 21876 15688 21882 15700
rect 21913 15691 21971 15697
rect 21913 15688 21925 15691
rect 21876 15660 21925 15688
rect 21876 15648 21882 15660
rect 21913 15657 21925 15660
rect 21959 15657 21971 15691
rect 22278 15688 22284 15700
rect 22239 15660 22284 15688
rect 21913 15651 21971 15657
rect 22278 15648 22284 15660
rect 22336 15648 22342 15700
rect 16162 15623 16220 15629
rect 16162 15620 16174 15623
rect 15988 15592 16174 15620
rect 15988 15580 15994 15592
rect 16162 15589 16174 15592
rect 16208 15589 16220 15623
rect 19429 15623 19487 15629
rect 19429 15620 19441 15623
rect 16162 15583 16220 15589
rect 16776 15592 19441 15620
rect 2958 15552 2964 15564
rect 2919 15524 2964 15552
rect 2958 15512 2964 15524
rect 3016 15512 3022 15564
rect 11882 15512 11888 15564
rect 11940 15552 11946 15564
rect 12012 15555 12070 15561
rect 12012 15552 12024 15555
rect 11940 15524 12024 15552
rect 11940 15512 11946 15524
rect 12012 15521 12024 15524
rect 12058 15521 12070 15555
rect 12012 15515 12070 15521
rect 14826 15512 14832 15564
rect 14884 15552 14890 15564
rect 15841 15555 15899 15561
rect 15841 15552 15853 15555
rect 14884 15524 15853 15552
rect 14884 15512 14890 15524
rect 15841 15521 15853 15524
rect 15887 15521 15899 15555
rect 15841 15515 15899 15521
rect 16298 15512 16304 15564
rect 16356 15552 16362 15564
rect 16776 15561 16804 15592
rect 19429 15589 19441 15592
rect 19475 15589 19487 15623
rect 19429 15583 19487 15589
rect 21085 15623 21143 15629
rect 21085 15589 21097 15623
rect 21131 15620 21143 15623
rect 21450 15620 21456 15632
rect 21131 15592 21456 15620
rect 21131 15589 21143 15592
rect 21085 15583 21143 15589
rect 21450 15580 21456 15592
rect 21508 15580 21514 15632
rect 22554 15620 22560 15632
rect 22515 15592 22560 15620
rect 22554 15580 22560 15592
rect 22612 15580 22618 15632
rect 22646 15580 22652 15632
rect 22704 15620 22710 15632
rect 22704 15592 22749 15620
rect 22704 15580 22710 15592
rect 16761 15555 16819 15561
rect 16761 15552 16773 15555
rect 16356 15524 16773 15552
rect 16356 15512 16362 15524
rect 16761 15521 16773 15524
rect 16807 15521 16819 15555
rect 16761 15515 16819 15521
rect 17678 15512 17684 15564
rect 17736 15552 17742 15564
rect 17865 15555 17923 15561
rect 17865 15552 17877 15555
rect 17736 15524 17877 15552
rect 17736 15512 17742 15524
rect 17865 15521 17877 15524
rect 17911 15521 17923 15555
rect 17865 15515 17923 15521
rect 18141 15555 18199 15561
rect 18141 15521 18153 15555
rect 18187 15552 18199 15555
rect 18322 15552 18328 15564
rect 18187 15524 18328 15552
rect 18187 15521 18199 15524
rect 18141 15515 18199 15521
rect 18322 15512 18328 15524
rect 18380 15512 18386 15564
rect 24581 15555 24639 15561
rect 24581 15521 24593 15555
rect 24627 15552 24639 15555
rect 24670 15552 24676 15564
rect 24627 15524 24676 15552
rect 24627 15521 24639 15524
rect 24581 15515 24639 15521
rect 24670 15512 24676 15524
rect 24728 15512 24734 15564
rect 4341 15487 4399 15493
rect 4341 15484 4353 15487
rect 4126 15456 4353 15484
rect 3142 15348 3148 15360
rect 3103 15320 3148 15348
rect 3142 15308 3148 15320
rect 3200 15308 3206 15360
rect 3418 15308 3424 15360
rect 3476 15348 3482 15360
rect 3789 15351 3847 15357
rect 3789 15348 3801 15351
rect 3476 15320 3801 15348
rect 3476 15308 3482 15320
rect 3789 15317 3801 15320
rect 3835 15348 3847 15351
rect 4126 15348 4154 15456
rect 4341 15453 4353 15456
rect 4387 15453 4399 15487
rect 6273 15487 6331 15493
rect 6273 15484 6285 15487
rect 4341 15447 4399 15453
rect 6012 15456 6285 15484
rect 3835 15320 4154 15348
rect 3835 15317 3847 15320
rect 3789 15311 3847 15317
rect 4338 15308 4344 15360
rect 4396 15348 4402 15360
rect 6012 15357 6040 15456
rect 6273 15453 6285 15456
rect 6319 15453 6331 15487
rect 6273 15447 6331 15453
rect 6917 15487 6975 15493
rect 6917 15453 6929 15487
rect 6963 15484 6975 15487
rect 7466 15484 7472 15496
rect 6963 15456 7472 15484
rect 6963 15453 6975 15456
rect 6917 15447 6975 15453
rect 7466 15444 7472 15456
rect 7524 15484 7530 15496
rect 7837 15487 7895 15493
rect 7837 15484 7849 15487
rect 7524 15456 7849 15484
rect 7524 15444 7530 15456
rect 7837 15453 7849 15456
rect 7883 15453 7895 15487
rect 10410 15484 10416 15496
rect 10371 15456 10416 15484
rect 7837 15447 7895 15453
rect 10410 15444 10416 15456
rect 10468 15444 10474 15496
rect 12115 15487 12173 15493
rect 12115 15453 12127 15487
rect 12161 15484 12173 15487
rect 13078 15484 13084 15496
rect 12161 15456 13084 15484
rect 12161 15453 12173 15456
rect 12115 15447 12173 15453
rect 13078 15444 13084 15456
rect 13136 15444 13142 15496
rect 13357 15487 13415 15493
rect 13357 15453 13369 15487
rect 13403 15484 13415 15487
rect 13446 15484 13452 15496
rect 13403 15456 13452 15484
rect 13403 15453 13415 15456
rect 13357 15447 13415 15453
rect 10428 15416 10456 15444
rect 13372 15416 13400 15447
rect 13446 15444 13452 15456
rect 13504 15444 13510 15496
rect 18782 15484 18788 15496
rect 18695 15456 18788 15484
rect 18782 15444 18788 15456
rect 18840 15484 18846 15496
rect 19337 15487 19395 15493
rect 19337 15484 19349 15487
rect 18840 15456 19349 15484
rect 18840 15444 18846 15456
rect 19337 15453 19349 15456
rect 19383 15453 19395 15487
rect 20990 15484 20996 15496
rect 20951 15456 20996 15484
rect 19337 15447 19395 15453
rect 20990 15444 20996 15456
rect 21048 15444 21054 15496
rect 21269 15487 21327 15493
rect 21269 15484 21281 15487
rect 21100 15456 21281 15484
rect 10428 15388 13400 15416
rect 19889 15419 19947 15425
rect 19889 15385 19901 15419
rect 19935 15416 19947 15419
rect 20530 15416 20536 15428
rect 19935 15388 20536 15416
rect 19935 15385 19947 15388
rect 19889 15379 19947 15385
rect 20530 15376 20536 15388
rect 20588 15416 20594 15428
rect 21100 15416 21128 15456
rect 21269 15453 21281 15456
rect 21315 15453 21327 15487
rect 22830 15484 22836 15496
rect 22791 15456 22836 15484
rect 21269 15447 21327 15453
rect 22830 15444 22836 15456
rect 22888 15444 22894 15496
rect 24762 15416 24768 15428
rect 20588 15388 21128 15416
rect 24723 15388 24768 15416
rect 20588 15376 20594 15388
rect 24762 15376 24768 15388
rect 24820 15376 24826 15428
rect 5997 15351 6055 15357
rect 5997 15348 6009 15351
rect 4396 15320 6009 15348
rect 4396 15308 4402 15320
rect 5997 15317 6009 15320
rect 6043 15317 6055 15351
rect 7558 15348 7564 15360
rect 7519 15320 7564 15348
rect 5997 15311 6055 15317
rect 7558 15308 7564 15320
rect 7616 15308 7622 15360
rect 13998 15348 14004 15360
rect 13959 15320 14004 15348
rect 13998 15308 14004 15320
rect 14056 15308 14062 15360
rect 15654 15348 15660 15360
rect 15615 15320 15660 15348
rect 15654 15308 15660 15320
rect 15712 15308 15718 15360
rect 19058 15348 19064 15360
rect 19019 15320 19064 15348
rect 19058 15308 19064 15320
rect 19116 15308 19122 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 4430 15104 4436 15156
rect 4488 15144 4494 15156
rect 4798 15144 4804 15156
rect 4488 15116 4804 15144
rect 4488 15104 4494 15116
rect 4798 15104 4804 15116
rect 4856 15144 4862 15156
rect 5537 15147 5595 15153
rect 5537 15144 5549 15147
rect 4856 15116 5549 15144
rect 4856 15104 4862 15116
rect 5537 15113 5549 15116
rect 5583 15113 5595 15147
rect 7834 15144 7840 15156
rect 7795 15116 7840 15144
rect 5537 15107 5595 15113
rect 7834 15104 7840 15116
rect 7892 15144 7898 15156
rect 8113 15147 8171 15153
rect 8113 15144 8125 15147
rect 7892 15116 8125 15144
rect 7892 15104 7898 15116
rect 8113 15113 8125 15116
rect 8159 15113 8171 15147
rect 8113 15107 8171 15113
rect 10134 15104 10140 15156
rect 10192 15144 10198 15156
rect 10781 15147 10839 15153
rect 10781 15144 10793 15147
rect 10192 15116 10793 15144
rect 10192 15104 10198 15116
rect 10781 15113 10793 15116
rect 10827 15113 10839 15147
rect 10781 15107 10839 15113
rect 11882 15104 11888 15156
rect 11940 15144 11946 15156
rect 11977 15147 12035 15153
rect 11977 15144 11989 15147
rect 11940 15116 11989 15144
rect 11940 15104 11946 15116
rect 11977 15113 11989 15116
rect 12023 15113 12035 15147
rect 11977 15107 12035 15113
rect 13078 15104 13084 15156
rect 13136 15144 13142 15156
rect 14553 15147 14611 15153
rect 14553 15144 14565 15147
rect 13136 15116 14565 15144
rect 13136 15104 13142 15116
rect 14553 15113 14565 15116
rect 14599 15113 14611 15147
rect 14553 15107 14611 15113
rect 14826 15104 14832 15156
rect 14884 15144 14890 15156
rect 14921 15147 14979 15153
rect 14921 15144 14933 15147
rect 14884 15116 14933 15144
rect 14884 15104 14890 15116
rect 14921 15113 14933 15116
rect 14967 15113 14979 15147
rect 14921 15107 14979 15113
rect 15243 15147 15301 15153
rect 15243 15113 15255 15147
rect 15289 15144 15301 15147
rect 15654 15144 15660 15156
rect 15289 15116 15660 15144
rect 15289 15113 15301 15116
rect 15243 15107 15301 15113
rect 15654 15104 15660 15116
rect 15712 15104 15718 15156
rect 15930 15144 15936 15156
rect 15891 15116 15936 15144
rect 15930 15104 15936 15116
rect 15988 15104 15994 15156
rect 16942 15104 16948 15156
rect 17000 15144 17006 15156
rect 17221 15147 17279 15153
rect 17221 15144 17233 15147
rect 17000 15116 17233 15144
rect 17000 15104 17006 15116
rect 17221 15113 17233 15116
rect 17267 15113 17279 15147
rect 17678 15144 17684 15156
rect 17639 15116 17684 15144
rect 17221 15107 17279 15113
rect 17678 15104 17684 15116
rect 17736 15104 17742 15156
rect 18187 15147 18245 15153
rect 18187 15113 18199 15147
rect 18233 15144 18245 15147
rect 18782 15144 18788 15156
rect 18233 15116 18788 15144
rect 18233 15113 18245 15116
rect 18187 15107 18245 15113
rect 18782 15104 18788 15116
rect 18840 15104 18846 15156
rect 22554 15104 22560 15156
rect 22612 15144 22618 15156
rect 22833 15147 22891 15153
rect 22833 15144 22845 15147
rect 22612 15116 22845 15144
rect 22612 15104 22618 15116
rect 22833 15113 22845 15116
rect 22879 15113 22891 15147
rect 22833 15107 22891 15113
rect 5258 15076 5264 15088
rect 5219 15048 5264 15076
rect 5258 15036 5264 15048
rect 5316 15036 5322 15088
rect 7466 15036 7472 15088
rect 7524 15076 7530 15088
rect 8481 15079 8539 15085
rect 8481 15076 8493 15079
rect 7524 15048 8493 15076
rect 7524 15036 7530 15048
rect 8481 15045 8493 15048
rect 8527 15045 8539 15079
rect 14182 15076 14188 15088
rect 14143 15048 14188 15076
rect 8481 15039 8539 15045
rect 14182 15036 14188 15048
rect 14240 15036 14246 15088
rect 6914 15008 6920 15020
rect 6827 14980 6920 15008
rect 6914 14968 6920 14980
rect 6972 15008 6978 15020
rect 7558 15008 7564 15020
rect 6972 14980 7564 15008
rect 6972 14968 6978 14980
rect 7558 14968 7564 14980
rect 7616 14968 7622 15020
rect 10137 15011 10195 15017
rect 10137 14977 10149 15011
rect 10183 15008 10195 15011
rect 10410 15008 10416 15020
rect 10183 14980 10416 15008
rect 10183 14977 10195 14980
rect 10137 14971 10195 14977
rect 10410 14968 10416 14980
rect 10468 14968 10474 15020
rect 13081 15011 13139 15017
rect 13081 14977 13093 15011
rect 13127 15008 13139 15011
rect 13170 15008 13176 15020
rect 13127 14980 13176 15008
rect 13127 14977 13139 14980
rect 13081 14971 13139 14977
rect 13170 14968 13176 14980
rect 13228 15008 13234 15020
rect 13357 15011 13415 15017
rect 13357 15008 13369 15011
rect 13228 14980 13369 15008
rect 13228 14968 13234 14980
rect 13357 14977 13369 14980
rect 13403 14977 13415 15011
rect 13357 14971 13415 14977
rect 13633 15011 13691 15017
rect 13633 14977 13645 15011
rect 13679 15008 13691 15011
rect 13998 15008 14004 15020
rect 13679 14980 14004 15008
rect 13679 14977 13691 14980
rect 13633 14971 13691 14977
rect 1302 14900 1308 14952
rect 1360 14940 1366 14952
rect 3234 14940 3240 14952
rect 1360 14912 3240 14940
rect 1360 14900 1366 14912
rect 3234 14900 3240 14912
rect 3292 14940 3298 14952
rect 3364 14943 3422 14949
rect 3364 14940 3376 14943
rect 3292 14912 3376 14940
rect 3292 14900 3298 14912
rect 3364 14909 3376 14912
rect 3410 14940 3422 14943
rect 3789 14943 3847 14949
rect 3789 14940 3801 14943
rect 3410 14912 3801 14940
rect 3410 14909 3422 14912
rect 3364 14903 3422 14909
rect 3789 14909 3801 14912
rect 3835 14909 3847 14943
rect 3789 14903 3847 14909
rect 4062 14900 4068 14952
rect 4120 14940 4126 14952
rect 4341 14943 4399 14949
rect 4341 14940 4353 14943
rect 4120 14912 4353 14940
rect 4120 14900 4126 14912
rect 4341 14909 4353 14912
rect 4387 14909 4399 14943
rect 4341 14903 4399 14909
rect 10965 14943 11023 14949
rect 10965 14909 10977 14943
rect 11011 14940 11023 14943
rect 11425 14943 11483 14949
rect 11425 14940 11437 14943
rect 11011 14912 11437 14940
rect 11011 14909 11023 14912
rect 10965 14903 11023 14909
rect 11425 14909 11437 14912
rect 11471 14909 11483 14943
rect 11425 14903 11483 14909
rect 4249 14875 4307 14881
rect 4249 14841 4261 14875
rect 4295 14872 4307 14875
rect 4522 14872 4528 14884
rect 4295 14844 4528 14872
rect 4295 14841 4307 14844
rect 4249 14835 4307 14841
rect 4522 14832 4528 14844
rect 4580 14872 4586 14884
rect 4703 14875 4761 14881
rect 4703 14872 4715 14875
rect 4580 14844 4715 14872
rect 4580 14832 4586 14844
rect 4703 14841 4715 14844
rect 4749 14872 4761 14875
rect 6638 14872 6644 14884
rect 4749 14844 6644 14872
rect 4749 14841 4761 14844
rect 4703 14835 4761 14841
rect 6638 14832 6644 14844
rect 6696 14872 6702 14884
rect 7279 14875 7337 14881
rect 7279 14872 7291 14875
rect 6696 14844 7291 14872
rect 6696 14832 6702 14844
rect 7279 14841 7291 14844
rect 7325 14872 7337 14875
rect 8018 14872 8024 14884
rect 7325 14844 8024 14872
rect 7325 14841 7337 14844
rect 7279 14835 7337 14841
rect 8018 14832 8024 14844
rect 8076 14832 8082 14884
rect 9490 14872 9496 14884
rect 9451 14844 9496 14872
rect 9490 14832 9496 14844
rect 9548 14832 9554 14884
rect 9585 14875 9643 14881
rect 9585 14841 9597 14875
rect 9631 14841 9643 14875
rect 10980 14872 11008 14903
rect 13262 14872 13268 14884
rect 9585 14835 9643 14841
rect 10244 14844 11008 14872
rect 11164 14844 13268 14872
rect 1578 14804 1584 14816
rect 1539 14776 1584 14804
rect 1578 14764 1584 14776
rect 1636 14764 1642 14816
rect 2958 14804 2964 14816
rect 2919 14776 2964 14804
rect 2958 14764 2964 14776
rect 3016 14764 3022 14816
rect 3467 14807 3525 14813
rect 3467 14773 3479 14807
rect 3513 14804 3525 14807
rect 3602 14804 3608 14816
rect 3513 14776 3608 14804
rect 3513 14773 3525 14776
rect 3467 14767 3525 14773
rect 3602 14764 3608 14776
rect 3660 14764 3666 14816
rect 6178 14804 6184 14816
rect 6139 14776 6184 14804
rect 6178 14764 6184 14776
rect 6236 14764 6242 14816
rect 9306 14804 9312 14816
rect 9267 14776 9312 14804
rect 9306 14764 9312 14776
rect 9364 14804 9370 14816
rect 9600 14804 9628 14835
rect 9364 14776 9628 14804
rect 9364 14764 9370 14776
rect 10042 14764 10048 14816
rect 10100 14804 10106 14816
rect 10244 14804 10272 14844
rect 10100 14776 10272 14804
rect 10505 14807 10563 14813
rect 10100 14764 10106 14776
rect 10505 14773 10517 14807
rect 10551 14804 10563 14807
rect 10686 14804 10692 14816
rect 10551 14776 10692 14804
rect 10551 14773 10563 14776
rect 10505 14767 10563 14773
rect 10686 14764 10692 14776
rect 10744 14764 10750 14816
rect 10778 14764 10784 14816
rect 10836 14804 10842 14816
rect 11164 14813 11192 14844
rect 13262 14832 13268 14844
rect 13320 14832 13326 14884
rect 13372 14872 13400 14971
rect 13998 14968 14004 14980
rect 14056 14968 14062 15020
rect 15672 15008 15700 15104
rect 15746 15036 15752 15088
rect 15804 15076 15810 15088
rect 17696 15076 17724 15104
rect 15804 15048 17724 15076
rect 19981 15079 20039 15085
rect 15804 15036 15810 15048
rect 19981 15045 19993 15079
rect 20027 15076 20039 15079
rect 20441 15079 20499 15085
rect 20441 15076 20453 15079
rect 20027 15048 20453 15076
rect 20027 15045 20039 15048
rect 19981 15039 20039 15045
rect 20441 15045 20453 15048
rect 20487 15076 20499 15079
rect 20809 15079 20867 15085
rect 20809 15076 20821 15079
rect 20487 15048 20821 15076
rect 20487 15045 20499 15048
rect 20441 15039 20499 15045
rect 20809 15045 20821 15048
rect 20855 15076 20867 15079
rect 21450 15076 21456 15088
rect 20855 15048 21456 15076
rect 20855 15045 20867 15048
rect 20809 15039 20867 15045
rect 21450 15036 21456 15048
rect 21508 15036 21514 15088
rect 21913 15079 21971 15085
rect 21913 15045 21925 15079
rect 21959 15076 21971 15079
rect 22738 15076 22744 15088
rect 21959 15048 22744 15076
rect 21959 15045 21971 15048
rect 21913 15039 21971 15045
rect 16209 15011 16267 15017
rect 16209 15008 16221 15011
rect 15672 14980 16221 15008
rect 16209 14977 16221 14980
rect 16255 14977 16267 15011
rect 16850 15008 16856 15020
rect 16763 14980 16856 15008
rect 16209 14971 16267 14977
rect 16850 14968 16856 14980
rect 16908 15008 16914 15020
rect 21928 15008 21956 15039
rect 22738 15036 22744 15048
rect 22796 15036 22802 15088
rect 16908 14980 21956 15008
rect 22557 15011 22615 15017
rect 16908 14968 16914 14980
rect 22557 14977 22569 15011
rect 22603 15008 22615 15011
rect 22646 15008 22652 15020
rect 22603 14980 22652 15008
rect 22603 14977 22615 14980
rect 22557 14971 22615 14977
rect 15010 14900 15016 14952
rect 15068 14940 15074 14952
rect 15140 14943 15198 14949
rect 15140 14940 15152 14943
rect 15068 14912 15152 14940
rect 15068 14900 15074 14912
rect 15140 14909 15152 14912
rect 15186 14940 15198 14943
rect 15565 14943 15623 14949
rect 15565 14940 15577 14943
rect 15186 14912 15577 14940
rect 15186 14909 15198 14912
rect 15140 14903 15198 14909
rect 15565 14909 15577 14912
rect 15611 14909 15623 14943
rect 15565 14903 15623 14909
rect 18116 14943 18174 14949
rect 18116 14909 18128 14943
rect 18162 14940 18174 14943
rect 18506 14940 18512 14952
rect 18162 14912 18512 14940
rect 18162 14909 18174 14912
rect 18116 14903 18174 14909
rect 18506 14900 18512 14912
rect 18564 14900 18570 14952
rect 19058 14940 19064 14952
rect 19019 14912 19064 14940
rect 19058 14900 19064 14912
rect 19116 14900 19122 14952
rect 13725 14875 13783 14881
rect 13725 14872 13737 14875
rect 13372 14844 13737 14872
rect 13725 14841 13737 14844
rect 13771 14841 13783 14875
rect 16298 14872 16304 14884
rect 16259 14844 16304 14872
rect 13725 14835 13783 14841
rect 16298 14832 16304 14844
rect 16356 14832 16362 14884
rect 19382 14875 19440 14881
rect 19382 14872 19394 14875
rect 18892 14844 19394 14872
rect 11149 14807 11207 14813
rect 11149 14804 11161 14807
rect 10836 14776 11161 14804
rect 10836 14764 10842 14776
rect 11149 14773 11161 14776
rect 11195 14773 11207 14807
rect 11149 14767 11207 14773
rect 12529 14807 12587 14813
rect 12529 14773 12541 14807
rect 12575 14804 12587 14807
rect 12894 14804 12900 14816
rect 12575 14776 12900 14804
rect 12575 14773 12587 14776
rect 12529 14767 12587 14773
rect 12894 14764 12900 14776
rect 12952 14764 12958 14816
rect 18230 14764 18236 14816
rect 18288 14804 18294 14816
rect 18892 14813 18920 14844
rect 19382 14841 19394 14844
rect 19428 14841 19440 14875
rect 21361 14875 21419 14881
rect 21361 14872 21373 14875
rect 19382 14835 19440 14841
rect 21100 14844 21373 14872
rect 18877 14807 18935 14813
rect 18877 14804 18889 14807
rect 18288 14776 18889 14804
rect 18288 14764 18294 14776
rect 18877 14773 18889 14776
rect 18923 14773 18935 14807
rect 18877 14767 18935 14773
rect 20898 14764 20904 14816
rect 20956 14804 20962 14816
rect 21100 14813 21128 14844
rect 21361 14841 21373 14844
rect 21407 14841 21419 14875
rect 21361 14835 21419 14841
rect 21450 14832 21456 14884
rect 21508 14872 21514 14884
rect 21508 14844 21601 14872
rect 21508 14832 21514 14844
rect 21085 14807 21143 14813
rect 21085 14804 21097 14807
rect 20956 14776 21097 14804
rect 20956 14764 20962 14776
rect 21085 14773 21097 14776
rect 21131 14773 21143 14807
rect 21468 14804 21496 14832
rect 22572 14804 22600 14971
rect 22646 14968 22652 14980
rect 22704 14968 22710 15020
rect 24670 15008 24676 15020
rect 24631 14980 24676 15008
rect 24670 14968 24676 14980
rect 24728 14968 24734 15020
rect 23661 14943 23719 14949
rect 23661 14940 23673 14943
rect 23584 14912 23673 14940
rect 23474 14872 23480 14884
rect 23387 14844 23480 14872
rect 23474 14832 23480 14844
rect 23532 14872 23538 14884
rect 23584 14872 23612 14912
rect 23661 14909 23673 14912
rect 23707 14909 23719 14943
rect 24118 14940 24124 14952
rect 24079 14912 24124 14940
rect 23661 14903 23719 14909
rect 24118 14900 24124 14912
rect 24176 14900 24182 14952
rect 23532 14844 23612 14872
rect 23532 14832 23538 14844
rect 23750 14804 23756 14816
rect 21468 14776 22600 14804
rect 23711 14776 23756 14804
rect 21085 14767 21143 14773
rect 23750 14764 23756 14776
rect 23808 14764 23814 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 934 14560 940 14612
rect 992 14600 998 14612
rect 1581 14603 1639 14609
rect 1581 14600 1593 14603
rect 992 14572 1593 14600
rect 992 14560 998 14572
rect 1581 14569 1593 14572
rect 1627 14569 1639 14603
rect 1581 14563 1639 14569
rect 3099 14603 3157 14609
rect 3099 14569 3111 14603
rect 3145 14600 3157 14603
rect 3418 14600 3424 14612
rect 3145 14572 3424 14600
rect 3145 14569 3157 14572
rect 3099 14563 3157 14569
rect 3418 14560 3424 14572
rect 3476 14560 3482 14612
rect 3513 14603 3571 14609
rect 3513 14569 3525 14603
rect 3559 14600 3571 14603
rect 3602 14600 3608 14612
rect 3559 14572 3608 14600
rect 3559 14569 3571 14572
rect 3513 14563 3571 14569
rect 3602 14560 3608 14572
rect 3660 14600 3666 14612
rect 6641 14603 6699 14609
rect 3660 14572 4384 14600
rect 3660 14560 3666 14572
rect 4356 14541 4384 14572
rect 6641 14569 6653 14603
rect 6687 14600 6699 14603
rect 8435 14603 8493 14609
rect 6687 14572 6960 14600
rect 6687 14569 6699 14572
rect 6641 14563 6699 14569
rect 4341 14535 4399 14541
rect 4341 14501 4353 14535
rect 4387 14501 4399 14535
rect 4341 14495 4399 14501
rect 4430 14492 4436 14544
rect 4488 14532 4494 14544
rect 4982 14532 4988 14544
rect 4488 14504 4533 14532
rect 4943 14504 4988 14532
rect 4488 14492 4494 14504
rect 4982 14492 4988 14504
rect 5040 14492 5046 14544
rect 6822 14532 6828 14544
rect 6783 14504 6828 14532
rect 6822 14492 6828 14504
rect 6880 14492 6886 14544
rect 6932 14541 6960 14572
rect 8435 14569 8447 14603
rect 8481 14600 8493 14603
rect 9490 14600 9496 14612
rect 8481 14572 9496 14600
rect 8481 14569 8493 14572
rect 8435 14563 8493 14569
rect 9490 14560 9496 14572
rect 9548 14560 9554 14612
rect 13078 14560 13084 14612
rect 13136 14600 13142 14612
rect 13173 14603 13231 14609
rect 13173 14600 13185 14603
rect 13136 14572 13185 14600
rect 13136 14560 13142 14572
rect 13173 14569 13185 14572
rect 13219 14569 13231 14603
rect 13173 14563 13231 14569
rect 13725 14603 13783 14609
rect 13725 14569 13737 14603
rect 13771 14600 13783 14603
rect 13906 14600 13912 14612
rect 13771 14572 13912 14600
rect 13771 14569 13783 14572
rect 13725 14563 13783 14569
rect 13906 14560 13912 14572
rect 13964 14560 13970 14612
rect 16209 14603 16267 14609
rect 16209 14569 16221 14603
rect 16255 14600 16267 14603
rect 16298 14600 16304 14612
rect 16255 14572 16304 14600
rect 16255 14569 16267 14572
rect 16209 14563 16267 14569
rect 16298 14560 16304 14572
rect 16356 14560 16362 14612
rect 18230 14560 18236 14612
rect 18288 14600 18294 14612
rect 18325 14603 18383 14609
rect 18325 14600 18337 14603
rect 18288 14572 18337 14600
rect 18288 14560 18294 14572
rect 18325 14569 18337 14572
rect 18371 14569 18383 14603
rect 18325 14563 18383 14569
rect 18877 14603 18935 14609
rect 18877 14569 18889 14603
rect 18923 14600 18935 14603
rect 19935 14603 19993 14609
rect 18923 14572 19886 14600
rect 18923 14569 18935 14572
rect 18877 14563 18935 14569
rect 6917 14535 6975 14541
rect 6917 14501 6929 14535
rect 6963 14532 6975 14535
rect 7006 14532 7012 14544
rect 6963 14504 7012 14532
rect 6963 14501 6975 14504
rect 6917 14495 6975 14501
rect 7006 14492 7012 14504
rect 7064 14492 7070 14544
rect 7466 14532 7472 14544
rect 7427 14504 7472 14532
rect 7466 14492 7472 14504
rect 7524 14492 7530 14544
rect 10502 14532 10508 14544
rect 10463 14504 10508 14532
rect 10502 14492 10508 14504
rect 10560 14492 10566 14544
rect 16574 14532 16580 14544
rect 16535 14504 16580 14532
rect 16574 14492 16580 14504
rect 16632 14492 16638 14544
rect 19518 14532 19524 14544
rect 19479 14504 19524 14532
rect 19518 14492 19524 14504
rect 19576 14492 19582 14544
rect 19858 14532 19886 14572
rect 19935 14569 19947 14603
rect 19981 14600 19993 14603
rect 20717 14603 20775 14609
rect 20717 14600 20729 14603
rect 19981 14572 20729 14600
rect 19981 14569 19993 14572
rect 19935 14563 19993 14569
rect 20717 14569 20729 14572
rect 20763 14600 20775 14603
rect 20990 14600 20996 14612
rect 20763 14572 20996 14600
rect 20763 14569 20775 14572
rect 20717 14563 20775 14569
rect 20990 14560 20996 14572
rect 21048 14560 21054 14612
rect 22554 14600 22560 14612
rect 22515 14572 22560 14600
rect 22554 14560 22560 14572
rect 22612 14560 22618 14612
rect 23753 14603 23811 14609
rect 23753 14600 23765 14603
rect 23446 14572 23765 14600
rect 21085 14535 21143 14541
rect 21085 14532 21097 14535
rect 19858 14504 21097 14532
rect 21085 14501 21097 14504
rect 21131 14532 21143 14535
rect 21450 14532 21456 14544
rect 21131 14504 21456 14532
rect 21131 14501 21143 14504
rect 21085 14495 21143 14501
rect 21450 14492 21456 14504
rect 21508 14492 21514 14544
rect 1397 14467 1455 14473
rect 1397 14433 1409 14467
rect 1443 14464 1455 14467
rect 2130 14464 2136 14476
rect 1443 14436 2136 14464
rect 1443 14433 1455 14436
rect 1397 14427 1455 14433
rect 2130 14424 2136 14436
rect 2188 14424 2194 14476
rect 3028 14467 3086 14473
rect 3028 14433 3040 14467
rect 3074 14464 3086 14467
rect 3418 14464 3424 14476
rect 3074 14436 3424 14464
rect 3074 14433 3086 14436
rect 3028 14427 3086 14433
rect 3418 14424 3424 14436
rect 3476 14424 3482 14476
rect 7926 14424 7932 14476
rect 7984 14464 7990 14476
rect 8294 14464 8300 14476
rect 8352 14473 8358 14476
rect 8352 14467 8390 14473
rect 7984 14436 8300 14464
rect 7984 14424 7990 14436
rect 8294 14424 8300 14436
rect 8378 14433 8390 14467
rect 8352 14427 8390 14433
rect 15289 14467 15347 14473
rect 15289 14433 15301 14467
rect 15335 14464 15347 14467
rect 15378 14464 15384 14476
rect 15335 14436 15384 14464
rect 15335 14433 15347 14436
rect 15289 14427 15347 14433
rect 8352 14424 8358 14427
rect 15378 14424 15384 14436
rect 15436 14424 15442 14476
rect 19864 14467 19922 14473
rect 19864 14433 19876 14467
rect 19910 14433 19922 14467
rect 22462 14464 22468 14476
rect 22423 14436 22468 14464
rect 19864 14427 19922 14433
rect 10410 14396 10416 14408
rect 10371 14368 10416 14396
rect 10410 14356 10416 14368
rect 10468 14356 10474 14408
rect 12802 14396 12808 14408
rect 12763 14368 12808 14396
rect 12802 14356 12808 14368
rect 12860 14356 12866 14408
rect 13998 14356 14004 14408
rect 14056 14396 14062 14408
rect 14182 14396 14188 14408
rect 14056 14368 14188 14396
rect 14056 14356 14062 14368
rect 14182 14356 14188 14368
rect 14240 14356 14246 14408
rect 16485 14399 16543 14405
rect 16485 14365 16497 14399
rect 16531 14396 16543 14399
rect 16850 14396 16856 14408
rect 16531 14368 16856 14396
rect 16531 14365 16543 14368
rect 16485 14359 16543 14365
rect 16850 14356 16856 14368
rect 16908 14356 16914 14408
rect 17494 14356 17500 14408
rect 17552 14396 17558 14408
rect 17957 14399 18015 14405
rect 17957 14396 17969 14399
rect 17552 14368 17969 14396
rect 17552 14356 17558 14368
rect 17957 14365 17969 14368
rect 18003 14365 18015 14399
rect 17957 14359 18015 14365
rect 10962 14328 10968 14340
rect 10875 14300 10968 14328
rect 10962 14288 10968 14300
rect 11020 14328 11026 14340
rect 14458 14328 14464 14340
rect 11020 14300 14464 14328
rect 11020 14288 11026 14300
rect 14458 14288 14464 14300
rect 14516 14288 14522 14340
rect 17034 14328 17040 14340
rect 16995 14300 17040 14328
rect 17034 14288 17040 14300
rect 17092 14288 17098 14340
rect 19879 14328 19907 14427
rect 22462 14424 22468 14436
rect 22520 14424 22526 14476
rect 22925 14467 22983 14473
rect 22925 14433 22937 14467
rect 22971 14464 22983 14467
rect 23446 14464 23474 14572
rect 23753 14569 23765 14572
rect 23799 14600 23811 14603
rect 24118 14600 24124 14612
rect 23799 14572 24124 14600
rect 23799 14569 23811 14572
rect 23753 14563 23811 14569
rect 24118 14560 24124 14572
rect 24176 14560 24182 14612
rect 22971 14436 23474 14464
rect 24096 14467 24154 14473
rect 22971 14433 22983 14436
rect 22925 14427 22983 14433
rect 24096 14433 24108 14467
rect 24142 14464 24154 14467
rect 24670 14464 24676 14476
rect 24142 14436 24676 14464
rect 24142 14433 24154 14436
rect 24096 14427 24154 14433
rect 20714 14356 20720 14408
rect 20772 14396 20778 14408
rect 20993 14399 21051 14405
rect 20993 14396 21005 14399
rect 20772 14368 21005 14396
rect 20772 14356 20778 14368
rect 20993 14365 21005 14368
rect 21039 14365 21051 14399
rect 20993 14359 21051 14365
rect 21174 14356 21180 14408
rect 21232 14396 21238 14408
rect 21269 14399 21327 14405
rect 21269 14396 21281 14399
rect 21232 14368 21281 14396
rect 21232 14356 21238 14368
rect 21269 14365 21281 14368
rect 21315 14365 21327 14399
rect 21269 14359 21327 14365
rect 21818 14356 21824 14408
rect 21876 14396 21882 14408
rect 22940 14396 22968 14427
rect 24670 14424 24676 14436
rect 24728 14424 24734 14476
rect 21876 14368 22968 14396
rect 21876 14356 21882 14368
rect 19978 14328 19984 14340
rect 19879 14300 19984 14328
rect 19978 14288 19984 14300
rect 20036 14328 20042 14340
rect 23658 14328 23664 14340
rect 20036 14300 23664 14328
rect 20036 14288 20042 14300
rect 23658 14288 23664 14300
rect 23716 14288 23722 14340
rect 2038 14260 2044 14272
rect 1999 14232 2044 14260
rect 2038 14220 2044 14232
rect 2096 14220 2102 14272
rect 3881 14263 3939 14269
rect 3881 14229 3893 14263
rect 3927 14260 3939 14263
rect 4062 14260 4068 14272
rect 3927 14232 4068 14260
rect 3927 14229 3939 14232
rect 3881 14223 3939 14229
rect 4062 14220 4068 14232
rect 4120 14220 4126 14272
rect 6270 14260 6276 14272
rect 6231 14232 6276 14260
rect 6270 14220 6276 14232
rect 6328 14220 6334 14272
rect 9766 14220 9772 14272
rect 9824 14260 9830 14272
rect 9861 14263 9919 14269
rect 9861 14260 9873 14263
rect 9824 14232 9873 14260
rect 9824 14220 9830 14232
rect 9861 14229 9873 14232
rect 9907 14229 9919 14263
rect 12526 14260 12532 14272
rect 12487 14232 12532 14260
rect 9861 14223 9919 14229
rect 12526 14220 12532 14232
rect 12584 14220 12590 14272
rect 14277 14263 14335 14269
rect 14277 14229 14289 14263
rect 14323 14260 14335 14263
rect 14366 14260 14372 14272
rect 14323 14232 14372 14260
rect 14323 14229 14335 14232
rect 14277 14223 14335 14229
rect 14366 14220 14372 14232
rect 14424 14220 14430 14272
rect 15473 14263 15531 14269
rect 15473 14229 15485 14263
rect 15519 14260 15531 14263
rect 15562 14260 15568 14272
rect 15519 14232 15568 14260
rect 15519 14229 15531 14232
rect 15473 14223 15531 14229
rect 15562 14220 15568 14232
rect 15620 14220 15626 14272
rect 15838 14260 15844 14272
rect 15799 14232 15844 14260
rect 15838 14220 15844 14232
rect 15896 14220 15902 14272
rect 19150 14260 19156 14272
rect 19111 14232 19156 14260
rect 19150 14220 19156 14232
rect 19208 14220 19214 14272
rect 22097 14263 22155 14269
rect 22097 14229 22109 14263
rect 22143 14260 22155 14263
rect 22278 14260 22284 14272
rect 22143 14232 22284 14260
rect 22143 14229 22155 14232
rect 22097 14223 22155 14229
rect 22278 14220 22284 14232
rect 22336 14220 22342 14272
rect 23750 14220 23756 14272
rect 23808 14260 23814 14272
rect 24167 14263 24225 14269
rect 24167 14260 24179 14263
rect 23808 14232 24179 14260
rect 23808 14220 23814 14232
rect 24167 14229 24179 14232
rect 24213 14229 24225 14263
rect 24167 14223 24225 14229
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 1535 14059 1593 14065
rect 1535 14025 1547 14059
rect 1581 14056 1593 14059
rect 4338 14056 4344 14068
rect 1581 14028 4344 14056
rect 1581 14025 1593 14028
rect 1535 14019 1593 14025
rect 4338 14016 4344 14028
rect 4396 14016 4402 14068
rect 4430 14016 4436 14068
rect 4488 14056 4494 14068
rect 4801 14059 4859 14065
rect 4801 14056 4813 14059
rect 4488 14028 4813 14056
rect 4488 14016 4494 14028
rect 4801 14025 4813 14028
rect 4847 14056 4859 14059
rect 5074 14056 5080 14068
rect 4847 14028 5080 14056
rect 4847 14025 4859 14028
rect 4801 14019 4859 14025
rect 5074 14016 5080 14028
rect 5132 14016 5138 14068
rect 6454 14016 6460 14068
rect 6512 14056 6518 14068
rect 7006 14056 7012 14068
rect 6512 14028 7012 14056
rect 6512 14016 6518 14028
rect 7006 14016 7012 14028
rect 7064 14056 7070 14068
rect 7745 14059 7803 14065
rect 7745 14056 7757 14059
rect 7064 14028 7757 14056
rect 7064 14016 7070 14028
rect 7745 14025 7757 14028
rect 7791 14025 7803 14059
rect 8294 14056 8300 14068
rect 8255 14028 8300 14056
rect 7745 14019 7803 14025
rect 8294 14016 8300 14028
rect 8352 14016 8358 14068
rect 8895 14059 8953 14065
rect 8895 14025 8907 14059
rect 8941 14056 8953 14059
rect 10410 14056 10416 14068
rect 8941 14028 10416 14056
rect 8941 14025 8953 14028
rect 8895 14019 8953 14025
rect 10410 14016 10416 14028
rect 10468 14056 10474 14068
rect 11333 14059 11391 14065
rect 11333 14056 11345 14059
rect 10468 14028 11345 14056
rect 10468 14016 10474 14028
rect 11333 14025 11345 14028
rect 11379 14025 11391 14059
rect 11333 14019 11391 14025
rect 11606 14016 11612 14068
rect 11664 14056 11670 14068
rect 12161 14059 12219 14065
rect 12161 14056 12173 14059
rect 11664 14028 12173 14056
rect 11664 14016 11670 14028
rect 12161 14025 12173 14028
rect 12207 14025 12219 14059
rect 12161 14019 12219 14025
rect 1949 13991 2007 13997
rect 1949 13957 1961 13991
rect 1995 13988 2007 13991
rect 2130 13988 2136 14000
rect 1995 13960 2136 13988
rect 1995 13957 2007 13960
rect 1949 13951 2007 13957
rect 2130 13948 2136 13960
rect 2188 13948 2194 14000
rect 2406 13948 2412 14000
rect 2464 13988 2470 14000
rect 4982 13988 4988 14000
rect 2464 13960 4988 13988
rect 2464 13948 2470 13960
rect 4982 13948 4988 13960
rect 5040 13988 5046 14000
rect 6638 13988 6644 14000
rect 5040 13948 5073 13988
rect 6599 13960 6644 13988
rect 6638 13948 6644 13960
rect 6696 13948 6702 14000
rect 8018 13948 8024 14000
rect 8076 13988 8082 14000
rect 9585 13991 9643 13997
rect 9585 13988 9597 13991
rect 8076 13960 9597 13988
rect 8076 13948 8082 13960
rect 9585 13957 9597 13960
rect 9631 13957 9643 13991
rect 9585 13951 9643 13957
rect 2225 13923 2283 13929
rect 2225 13920 2237 13923
rect 1447 13892 2237 13920
rect 106 13812 112 13864
rect 164 13852 170 13864
rect 1447 13861 1475 13892
rect 2225 13889 2237 13892
rect 2271 13889 2283 13923
rect 5045 13920 5073 13948
rect 5045 13892 5764 13920
rect 2225 13883 2283 13889
rect 1432 13855 1490 13861
rect 1432 13852 1444 13855
rect 164 13824 1444 13852
rect 164 13812 170 13824
rect 1432 13821 1444 13824
rect 1478 13821 1490 13855
rect 1432 13815 1490 13821
rect 2777 13855 2835 13861
rect 2777 13821 2789 13855
rect 2823 13852 2835 13855
rect 2866 13852 2872 13864
rect 2823 13824 2872 13852
rect 2823 13821 2835 13824
rect 2777 13815 2835 13821
rect 2866 13812 2872 13824
rect 2924 13812 2930 13864
rect 5736 13861 5764 13892
rect 6270 13880 6276 13932
rect 6328 13920 6334 13932
rect 6730 13920 6736 13932
rect 6328 13892 6736 13920
rect 6328 13880 6334 13892
rect 6730 13880 6736 13892
rect 6788 13920 6794 13932
rect 6825 13923 6883 13929
rect 6825 13920 6837 13923
rect 6788 13892 6837 13920
rect 6788 13880 6794 13892
rect 6825 13889 6837 13892
rect 6871 13889 6883 13923
rect 6825 13883 6883 13889
rect 3881 13855 3939 13861
rect 3881 13821 3893 13855
rect 3927 13852 3939 13855
rect 5721 13855 5779 13861
rect 3927 13824 5488 13852
rect 3927 13821 3939 13824
rect 3881 13815 3939 13821
rect 4243 13787 4301 13793
rect 4243 13784 4255 13787
rect 4217 13753 4255 13784
rect 4289 13784 4301 13787
rect 4522 13784 4528 13796
rect 4289 13756 4528 13784
rect 4289 13753 4301 13756
rect 4217 13747 4301 13753
rect 3050 13716 3056 13728
rect 3011 13688 3056 13716
rect 3050 13676 3056 13688
rect 3108 13676 3114 13728
rect 3418 13716 3424 13728
rect 3379 13688 3424 13716
rect 3418 13676 3424 13688
rect 3476 13676 3482 13728
rect 3789 13719 3847 13725
rect 3789 13685 3801 13719
rect 3835 13716 3847 13719
rect 4217 13716 4245 13747
rect 4522 13744 4528 13756
rect 4580 13744 4586 13796
rect 5460 13728 5488 13824
rect 5721 13821 5733 13855
rect 5767 13852 5779 13855
rect 6181 13855 6239 13861
rect 6181 13852 6193 13855
rect 5767 13824 6193 13852
rect 5767 13821 5779 13824
rect 5721 13815 5779 13821
rect 6181 13821 6193 13824
rect 6227 13821 6239 13855
rect 6181 13815 6239 13821
rect 8824 13855 8882 13861
rect 8824 13821 8836 13855
rect 8870 13852 8882 13855
rect 8938 13852 8944 13864
rect 8870 13824 8944 13852
rect 8870 13821 8882 13824
rect 8824 13815 8882 13821
rect 8938 13812 8944 13824
rect 8996 13852 9002 13864
rect 9217 13855 9275 13861
rect 9217 13852 9229 13855
rect 8996 13824 9229 13852
rect 8996 13812 9002 13824
rect 9217 13821 9229 13824
rect 9263 13821 9275 13855
rect 9217 13815 9275 13821
rect 6638 13744 6644 13796
rect 6696 13784 6702 13796
rect 7146 13787 7204 13793
rect 7146 13784 7158 13787
rect 6696 13756 7158 13784
rect 6696 13744 6702 13756
rect 7146 13753 7158 13756
rect 7192 13753 7204 13787
rect 7146 13747 7204 13753
rect 5442 13716 5448 13728
rect 3835 13688 4245 13716
rect 5403 13688 5448 13716
rect 3835 13685 3847 13688
rect 3789 13679 3847 13685
rect 5442 13676 5448 13688
rect 5500 13676 5506 13728
rect 5905 13719 5963 13725
rect 5905 13685 5917 13719
rect 5951 13716 5963 13719
rect 6362 13716 6368 13728
rect 5951 13688 6368 13716
rect 5951 13685 5963 13688
rect 5905 13679 5963 13685
rect 6362 13676 6368 13688
rect 6420 13676 6426 13728
rect 9600 13716 9628 13951
rect 10502 13948 10508 14000
rect 10560 13988 10566 14000
rect 10689 13991 10747 13997
rect 10689 13988 10701 13991
rect 10560 13960 10701 13988
rect 10560 13948 10566 13960
rect 10689 13957 10701 13960
rect 10735 13988 10747 13991
rect 10965 13991 11023 13997
rect 10965 13988 10977 13991
rect 10735 13960 10977 13988
rect 10735 13957 10747 13960
rect 10689 13951 10747 13957
rect 10965 13957 10977 13960
rect 11011 13957 11023 13991
rect 10965 13951 11023 13957
rect 9765 13855 9823 13861
rect 9765 13852 9777 13855
rect 9692 13824 9777 13852
rect 9692 13796 9720 13824
rect 9765 13821 9777 13824
rect 9811 13821 9823 13855
rect 9765 13815 9823 13821
rect 9968 13824 10174 13852
rect 9674 13744 9680 13796
rect 9732 13744 9738 13796
rect 9968 13716 9996 13824
rect 10146 13796 10174 13824
rect 10134 13793 10140 13796
rect 10131 13747 10140 13793
rect 10192 13784 10198 13796
rect 12176 13784 12204 14019
rect 12894 14016 12900 14068
rect 12952 14056 12958 14068
rect 14001 14059 14059 14065
rect 14001 14056 14013 14059
rect 12952 14028 14013 14056
rect 12952 14016 12958 14028
rect 14001 14025 14013 14028
rect 14047 14025 14059 14059
rect 14001 14019 14059 14025
rect 15841 14059 15899 14065
rect 15841 14025 15853 14059
rect 15887 14056 15899 14059
rect 15930 14056 15936 14068
rect 15887 14028 15936 14056
rect 15887 14025 15899 14028
rect 15841 14019 15899 14025
rect 13170 13948 13176 14000
rect 13228 13988 13234 14000
rect 13357 13991 13415 13997
rect 13357 13988 13369 13991
rect 13228 13960 13369 13988
rect 13228 13948 13234 13960
rect 13357 13957 13369 13960
rect 13403 13957 13415 13991
rect 13357 13951 13415 13957
rect 12434 13852 12440 13864
rect 12395 13824 12440 13852
rect 12434 13812 12440 13824
rect 12492 13812 12498 13864
rect 12250 13784 12256 13796
rect 10192 13756 12256 13784
rect 10134 13744 10140 13747
rect 10192 13744 10198 13756
rect 12250 13744 12256 13756
rect 12308 13784 12314 13796
rect 12758 13787 12816 13793
rect 12758 13784 12770 13787
rect 12308 13756 12770 13784
rect 12308 13744 12314 13756
rect 12758 13753 12770 13756
rect 12804 13753 12816 13787
rect 13372 13784 13400 13951
rect 14016 13920 14044 14019
rect 15930 14016 15936 14028
rect 15988 14016 15994 14068
rect 16574 14016 16580 14068
rect 16632 14056 16638 14068
rect 16853 14059 16911 14065
rect 16853 14056 16865 14059
rect 16632 14028 16865 14056
rect 16632 14016 16638 14028
rect 16853 14025 16865 14028
rect 16899 14025 16911 14059
rect 19978 14056 19984 14068
rect 19939 14028 19984 14056
rect 16853 14019 16911 14025
rect 19978 14016 19984 14028
rect 20036 14016 20042 14068
rect 21450 14056 21456 14068
rect 21411 14028 21456 14056
rect 21450 14016 21456 14028
rect 21508 14016 21514 14068
rect 23290 14016 23296 14068
rect 23348 14056 23354 14068
rect 23385 14059 23443 14065
rect 23385 14056 23397 14059
rect 23348 14028 23397 14056
rect 23348 14016 23354 14028
rect 23385 14025 23397 14028
rect 23431 14025 23443 14059
rect 25406 14056 25412 14068
rect 25367 14028 25412 14056
rect 23385 14019 23443 14025
rect 25406 14016 25412 14028
rect 25464 14016 25470 14068
rect 19058 13948 19064 14000
rect 19116 13988 19122 14000
rect 22462 13988 22468 14000
rect 19116 13960 22468 13988
rect 19116 13948 19122 13960
rect 22462 13948 22468 13960
rect 22520 13988 22526 14000
rect 23017 13991 23075 13997
rect 23017 13988 23029 13991
rect 22520 13960 23029 13988
rect 22520 13948 22526 13960
rect 23017 13957 23029 13960
rect 23063 13957 23075 13991
rect 23017 13951 23075 13957
rect 14277 13923 14335 13929
rect 14277 13920 14289 13923
rect 14016 13892 14289 13920
rect 14277 13889 14289 13892
rect 14323 13889 14335 13923
rect 14277 13883 14335 13889
rect 14458 13880 14464 13932
rect 14516 13920 14522 13932
rect 14553 13923 14611 13929
rect 14553 13920 14565 13923
rect 14516 13892 14565 13920
rect 14516 13880 14522 13892
rect 14553 13889 14565 13892
rect 14599 13889 14611 13923
rect 14553 13883 14611 13889
rect 15838 13880 15844 13932
rect 15896 13920 15902 13932
rect 15933 13923 15991 13929
rect 15933 13920 15945 13923
rect 15896 13892 15945 13920
rect 15896 13880 15902 13892
rect 15933 13889 15945 13892
rect 15979 13889 15991 13923
rect 15933 13883 15991 13889
rect 19426 13880 19432 13932
rect 19484 13920 19490 13932
rect 24213 13923 24271 13929
rect 24213 13920 24225 13923
rect 19484 13892 24225 13920
rect 19484 13880 19490 13892
rect 24213 13889 24225 13892
rect 24259 13889 24271 13923
rect 24213 13883 24271 13889
rect 18693 13855 18751 13861
rect 18693 13821 18705 13855
rect 18739 13852 18751 13855
rect 19150 13852 19156 13864
rect 18739 13824 19156 13852
rect 18739 13821 18751 13824
rect 18693 13815 18751 13821
rect 19150 13812 19156 13824
rect 19208 13812 19214 13864
rect 22738 13812 22744 13864
rect 22796 13852 22802 13864
rect 22796 13824 22841 13852
rect 22796 13812 22802 13824
rect 23290 13812 23296 13864
rect 23348 13852 23354 13864
rect 23661 13855 23719 13861
rect 23661 13852 23673 13855
rect 23348 13824 23673 13852
rect 23348 13812 23354 13824
rect 23661 13821 23673 13824
rect 23707 13821 23719 13855
rect 24118 13852 24124 13864
rect 24079 13824 24124 13852
rect 23661 13815 23719 13821
rect 24118 13812 24124 13824
rect 24176 13812 24182 13864
rect 25225 13855 25283 13861
rect 25225 13852 25237 13855
rect 24688 13824 25237 13852
rect 24688 13796 24716 13824
rect 25225 13821 25237 13824
rect 25271 13852 25283 13855
rect 25777 13855 25835 13861
rect 25777 13852 25789 13855
rect 25271 13824 25789 13852
rect 25271 13821 25283 13824
rect 25225 13815 25283 13821
rect 25777 13821 25789 13824
rect 25823 13821 25835 13855
rect 25777 13815 25835 13821
rect 14366 13784 14372 13796
rect 13372 13756 14372 13784
rect 12758 13747 12816 13753
rect 9600 13688 9996 13716
rect 12773 13716 12801 13747
rect 14366 13744 14372 13756
rect 14424 13744 14430 13796
rect 16254 13787 16312 13793
rect 16254 13784 16266 13787
rect 14936 13756 16266 13784
rect 13078 13716 13084 13728
rect 12773 13688 13084 13716
rect 13078 13676 13084 13688
rect 13136 13716 13142 13728
rect 13633 13719 13691 13725
rect 13633 13716 13645 13719
rect 13136 13688 13645 13716
rect 13136 13676 13142 13688
rect 13633 13685 13645 13688
rect 13679 13716 13691 13719
rect 14936 13716 14964 13756
rect 16254 13753 16266 13756
rect 16300 13753 16312 13787
rect 17494 13784 17500 13796
rect 17407 13756 17500 13784
rect 16254 13747 16312 13753
rect 15378 13716 15384 13728
rect 13679 13688 14964 13716
rect 15339 13688 15384 13716
rect 13679 13685 13691 13688
rect 13633 13679 13691 13685
rect 15378 13676 15384 13688
rect 15436 13676 15442 13728
rect 16269 13716 16297 13747
rect 17494 13744 17500 13756
rect 17552 13784 17558 13796
rect 17552 13756 18368 13784
rect 17552 13744 17558 13756
rect 17773 13719 17831 13725
rect 17773 13716 17785 13719
rect 16269 13688 17785 13716
rect 17773 13685 17785 13688
rect 17819 13716 17831 13719
rect 18230 13716 18236 13728
rect 17819 13688 18236 13716
rect 17819 13685 17831 13688
rect 17773 13679 17831 13685
rect 18230 13676 18236 13688
rect 18288 13676 18294 13728
rect 18340 13716 18368 13756
rect 18414 13744 18420 13796
rect 18472 13784 18478 13796
rect 19014 13787 19072 13793
rect 19014 13784 19026 13787
rect 18472 13756 19026 13784
rect 18472 13744 18478 13756
rect 19014 13753 19026 13756
rect 19060 13753 19072 13787
rect 20530 13784 20536 13796
rect 20443 13756 20536 13784
rect 19014 13747 19072 13753
rect 20530 13744 20536 13756
rect 20588 13744 20594 13796
rect 20625 13787 20683 13793
rect 20625 13753 20637 13787
rect 20671 13753 20683 13787
rect 21174 13784 21180 13796
rect 21135 13756 21180 13784
rect 20625 13747 20683 13753
rect 19426 13716 19432 13728
rect 18340 13688 19432 13716
rect 19426 13676 19432 13688
rect 19484 13676 19490 13728
rect 19518 13676 19524 13728
rect 19576 13716 19582 13728
rect 19613 13719 19671 13725
rect 19613 13716 19625 13719
rect 19576 13688 19625 13716
rect 19576 13676 19582 13688
rect 19613 13685 19625 13688
rect 19659 13685 19671 13719
rect 19613 13679 19671 13685
rect 20162 13676 20168 13728
rect 20220 13716 20226 13728
rect 20257 13719 20315 13725
rect 20257 13716 20269 13719
rect 20220 13688 20269 13716
rect 20220 13676 20226 13688
rect 20257 13685 20269 13688
rect 20303 13716 20315 13719
rect 20640 13716 20668 13747
rect 21174 13744 21180 13756
rect 21232 13744 21238 13796
rect 22094 13784 22100 13796
rect 22055 13756 22100 13784
rect 22094 13744 22100 13756
rect 22152 13744 22158 13796
rect 22189 13787 22247 13793
rect 22189 13753 22201 13787
rect 22235 13784 22247 13787
rect 22278 13784 22284 13796
rect 22235 13756 22284 13784
rect 22235 13753 22247 13756
rect 22189 13747 22247 13753
rect 22278 13744 22284 13756
rect 22336 13744 22342 13796
rect 24670 13784 24676 13796
rect 24583 13756 24676 13784
rect 24670 13744 24676 13756
rect 24728 13744 24734 13796
rect 21818 13716 21824 13728
rect 20303 13688 20668 13716
rect 21779 13688 21824 13716
rect 20303 13685 20315 13688
rect 20257 13679 20315 13685
rect 21818 13676 21824 13688
rect 21876 13676 21882 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 3050 13472 3056 13524
rect 3108 13512 3114 13524
rect 3421 13515 3479 13521
rect 3421 13512 3433 13515
rect 3108 13484 3433 13512
rect 3108 13472 3114 13484
rect 3421 13481 3433 13484
rect 3467 13512 3479 13515
rect 4522 13512 4528 13524
rect 3467 13484 4528 13512
rect 3467 13481 3479 13484
rect 3421 13475 3479 13481
rect 4522 13472 4528 13484
rect 4580 13472 4586 13524
rect 5074 13512 5080 13524
rect 5035 13484 5080 13512
rect 5074 13472 5080 13484
rect 5132 13472 5138 13524
rect 6089 13515 6147 13521
rect 6089 13481 6101 13515
rect 6135 13512 6147 13515
rect 6822 13512 6828 13524
rect 6135 13484 6828 13512
rect 6135 13481 6147 13484
rect 6089 13475 6147 13481
rect 6822 13472 6828 13484
rect 6880 13472 6886 13524
rect 10962 13512 10968 13524
rect 10428 13484 10968 13512
rect 4798 13444 4804 13456
rect 4759 13416 4804 13444
rect 4798 13404 4804 13416
rect 4856 13404 4862 13456
rect 1464 13379 1522 13385
rect 1464 13345 1476 13379
rect 1510 13376 1522 13379
rect 2222 13376 2228 13388
rect 1510 13348 2228 13376
rect 1510 13345 1522 13348
rect 1464 13339 1522 13345
rect 2222 13336 2228 13348
rect 2280 13336 2286 13388
rect 2406 13336 2412 13388
rect 2464 13376 2470 13388
rect 2501 13379 2559 13385
rect 2501 13376 2513 13379
rect 2464 13348 2513 13376
rect 2464 13336 2470 13348
rect 2501 13345 2513 13348
rect 2547 13345 2559 13379
rect 2501 13339 2559 13345
rect 4709 13379 4767 13385
rect 4709 13345 4721 13379
rect 4755 13376 4767 13379
rect 5092 13376 5120 13472
rect 10428 13456 10456 13484
rect 10962 13472 10968 13484
rect 11020 13472 11026 13524
rect 12802 13512 12808 13524
rect 12763 13484 12808 13512
rect 12802 13472 12808 13484
rect 12860 13512 12866 13524
rect 12860 13484 13814 13512
rect 12860 13472 12866 13484
rect 6178 13444 6184 13456
rect 6139 13416 6184 13444
rect 6178 13404 6184 13416
rect 6236 13404 6242 13456
rect 10039 13447 10097 13453
rect 10039 13413 10051 13447
rect 10085 13444 10097 13447
rect 10134 13444 10140 13456
rect 10085 13416 10140 13444
rect 10085 13413 10097 13416
rect 10039 13407 10097 13413
rect 10134 13404 10140 13416
rect 10192 13404 10198 13456
rect 10410 13404 10416 13456
rect 10468 13404 10474 13456
rect 12161 13447 12219 13453
rect 11440 13416 12020 13444
rect 11440 13388 11468 13416
rect 6454 13376 6460 13388
rect 4755 13348 5120 13376
rect 6415 13348 6460 13376
rect 4755 13345 4767 13348
rect 4709 13339 4767 13345
rect 6454 13336 6460 13348
rect 6512 13336 6518 13388
rect 8294 13376 8300 13388
rect 8255 13348 8300 13376
rect 8294 13336 8300 13348
rect 8352 13336 8358 13388
rect 8573 13379 8631 13385
rect 8573 13345 8585 13379
rect 8619 13376 8631 13379
rect 8846 13376 8852 13388
rect 8619 13348 8852 13376
rect 8619 13345 8631 13348
rect 8573 13339 8631 13345
rect 8846 13336 8852 13348
rect 8904 13336 8910 13388
rect 11422 13376 11428 13388
rect 11383 13348 11428 13376
rect 11422 13336 11428 13348
rect 11480 13336 11486 13388
rect 11882 13376 11888 13388
rect 11843 13348 11888 13376
rect 11882 13336 11888 13348
rect 11940 13336 11946 13388
rect 11992 13376 12020 13416
rect 12161 13413 12173 13447
rect 12207 13444 12219 13447
rect 12434 13444 12440 13456
rect 12207 13416 12440 13444
rect 12207 13413 12219 13416
rect 12161 13407 12219 13413
rect 12434 13404 12440 13416
rect 12492 13404 12498 13456
rect 13078 13404 13084 13456
rect 13136 13444 13142 13456
rect 13402 13447 13460 13453
rect 13402 13444 13414 13447
rect 13136 13416 13414 13444
rect 13136 13404 13142 13416
rect 13402 13413 13414 13416
rect 13448 13413 13460 13447
rect 13786 13444 13814 13484
rect 13998 13472 14004 13524
rect 14056 13512 14062 13524
rect 14274 13512 14280 13524
rect 14056 13484 14280 13512
rect 14056 13472 14062 13484
rect 14274 13472 14280 13484
rect 14332 13472 14338 13524
rect 15381 13515 15439 13521
rect 15381 13481 15393 13515
rect 15427 13481 15439 13515
rect 15381 13475 15439 13481
rect 15396 13444 15424 13475
rect 16574 13472 16580 13524
rect 16632 13512 16638 13524
rect 16669 13515 16727 13521
rect 16669 13512 16681 13515
rect 16632 13484 16681 13512
rect 16632 13472 16638 13484
rect 16669 13481 16681 13484
rect 16715 13481 16727 13515
rect 16669 13475 16727 13481
rect 16850 13472 16856 13524
rect 16908 13512 16914 13524
rect 17313 13515 17371 13521
rect 17313 13512 17325 13515
rect 16908 13484 17325 13512
rect 16908 13472 16914 13484
rect 17313 13481 17325 13484
rect 17359 13481 17371 13515
rect 17313 13475 17371 13481
rect 19153 13515 19211 13521
rect 19153 13481 19165 13515
rect 19199 13512 19211 13515
rect 20162 13512 20168 13524
rect 19199 13484 20168 13512
rect 19199 13481 19211 13484
rect 19153 13475 19211 13481
rect 20162 13472 20168 13484
rect 20220 13472 20226 13524
rect 20349 13515 20407 13521
rect 20349 13481 20361 13515
rect 20395 13512 20407 13515
rect 20530 13512 20536 13524
rect 20395 13484 20536 13512
rect 20395 13481 20407 13484
rect 20349 13475 20407 13481
rect 20530 13472 20536 13484
rect 20588 13472 20594 13524
rect 20898 13512 20904 13524
rect 20859 13484 20904 13512
rect 20898 13472 20904 13484
rect 20956 13472 20962 13524
rect 22186 13472 22192 13524
rect 22244 13512 22250 13524
rect 22925 13515 22983 13521
rect 22925 13512 22937 13515
rect 22244 13484 22937 13512
rect 22244 13472 22250 13484
rect 22925 13481 22937 13484
rect 22971 13512 22983 13515
rect 23750 13512 23756 13524
rect 22971 13484 23756 13512
rect 22971 13481 22983 13484
rect 22925 13475 22983 13481
rect 23750 13472 23756 13484
rect 23808 13472 23814 13524
rect 13786 13416 15424 13444
rect 13402 13407 13460 13413
rect 18322 13404 18328 13456
rect 18380 13444 18386 13456
rect 18554 13447 18612 13453
rect 18554 13444 18566 13447
rect 18380 13416 18566 13444
rect 18380 13404 18386 13416
rect 18554 13413 18566 13416
rect 18600 13413 18612 13447
rect 18554 13407 18612 13413
rect 19518 13404 19524 13456
rect 19576 13444 19582 13456
rect 22097 13447 22155 13453
rect 22097 13444 22109 13447
rect 19576 13416 22109 13444
rect 19576 13404 19582 13416
rect 22097 13413 22109 13416
rect 22143 13444 22155 13447
rect 22278 13444 22284 13456
rect 22143 13416 22284 13444
rect 22143 13413 22155 13416
rect 22097 13407 22155 13413
rect 22278 13404 22284 13416
rect 22336 13404 22342 13456
rect 22649 13447 22707 13453
rect 22649 13413 22661 13447
rect 22695 13444 22707 13447
rect 22830 13444 22836 13456
rect 22695 13416 22836 13444
rect 22695 13413 22707 13416
rect 22649 13407 22707 13413
rect 15286 13376 15292 13388
rect 11992 13348 15292 13376
rect 15286 13336 15292 13348
rect 15344 13336 15350 13388
rect 15838 13376 15844 13388
rect 15751 13348 15844 13376
rect 15838 13336 15844 13348
rect 15896 13336 15902 13388
rect 16920 13379 16978 13385
rect 16920 13345 16932 13379
rect 16966 13376 16978 13379
rect 17034 13376 17040 13388
rect 16966 13348 17040 13376
rect 16966 13345 16978 13348
rect 16920 13339 16978 13345
rect 17034 13336 17040 13348
rect 17092 13376 17098 13388
rect 21174 13376 21180 13388
rect 17092 13348 21180 13376
rect 17092 13336 17098 13348
rect 21174 13336 21180 13348
rect 21232 13336 21238 13388
rect 8757 13311 8815 13317
rect 8757 13277 8769 13311
rect 8803 13308 8815 13311
rect 9677 13311 9735 13317
rect 9677 13308 9689 13311
rect 8803 13280 9689 13308
rect 8803 13277 8815 13280
rect 8757 13271 8815 13277
rect 9677 13277 9689 13280
rect 9723 13308 9735 13311
rect 10778 13308 10784 13320
rect 9723 13280 10784 13308
rect 9723 13277 9735 13280
rect 9677 13271 9735 13277
rect 10778 13268 10784 13280
rect 10836 13268 10842 13320
rect 13078 13308 13084 13320
rect 13039 13280 13084 13308
rect 13078 13268 13084 13280
rect 13136 13268 13142 13320
rect 15856 13308 15884 13336
rect 16022 13308 16028 13320
rect 15856 13280 16028 13308
rect 16022 13268 16028 13280
rect 16080 13308 16086 13320
rect 18230 13308 18236 13320
rect 16080 13280 17172 13308
rect 18191 13280 18236 13308
rect 16080 13268 16086 13280
rect 17144 13252 17172 13280
rect 18230 13268 18236 13280
rect 18288 13268 18294 13320
rect 18414 13268 18420 13320
rect 18472 13308 18478 13320
rect 21082 13308 21088 13320
rect 18472 13280 21088 13308
rect 18472 13268 18478 13280
rect 21082 13268 21088 13280
rect 21140 13308 21146 13320
rect 21450 13308 21456 13320
rect 21140 13280 21456 13308
rect 21140 13268 21146 13280
rect 21450 13268 21456 13280
rect 21508 13268 21514 13320
rect 22002 13308 22008 13320
rect 21963 13280 22008 13308
rect 22002 13268 22008 13280
rect 22060 13268 22066 13320
rect 1535 13243 1593 13249
rect 1535 13209 1547 13243
rect 1581 13240 1593 13243
rect 1581 13212 2176 13240
rect 1581 13209 1593 13212
rect 1535 13203 1593 13209
rect 2148 13184 2176 13212
rect 8018 13200 8024 13252
rect 8076 13240 8082 13252
rect 12342 13240 12348 13252
rect 8076 13212 12348 13240
rect 8076 13200 8082 13212
rect 12342 13200 12348 13212
rect 12400 13200 12406 13252
rect 14734 13200 14740 13252
rect 14792 13240 14798 13252
rect 16991 13243 17049 13249
rect 16991 13240 17003 13243
rect 14792 13212 17003 13240
rect 14792 13200 14798 13212
rect 16991 13209 17003 13212
rect 17037 13209 17049 13243
rect 16991 13203 17049 13209
rect 17126 13200 17132 13252
rect 17184 13240 17190 13252
rect 20438 13240 20444 13252
rect 17184 13212 20444 13240
rect 17184 13200 17190 13212
rect 20438 13200 20444 13212
rect 20496 13200 20502 13252
rect 20714 13240 20720 13252
rect 20627 13212 20720 13240
rect 20714 13200 20720 13212
rect 20772 13240 20778 13252
rect 22664 13240 22692 13407
rect 22830 13404 22836 13416
rect 22888 13404 22894 13456
rect 23474 13336 23480 13388
rect 23532 13376 23538 13388
rect 23934 13376 23940 13388
rect 23532 13348 23577 13376
rect 23895 13348 23940 13376
rect 23532 13336 23538 13348
rect 23934 13336 23940 13348
rect 23992 13376 23998 13388
rect 24489 13379 24547 13385
rect 24489 13376 24501 13379
rect 23992 13348 24501 13376
rect 23992 13336 23998 13348
rect 24489 13345 24501 13348
rect 24535 13345 24547 13379
rect 24489 13339 24547 13345
rect 25041 13379 25099 13385
rect 25041 13345 25053 13379
rect 25087 13376 25099 13379
rect 25130 13376 25136 13388
rect 25087 13348 25136 13376
rect 25087 13345 25099 13348
rect 25041 13339 25099 13345
rect 25130 13336 25136 13348
rect 25188 13336 25194 13388
rect 24026 13308 24032 13320
rect 23987 13280 24032 13308
rect 24026 13268 24032 13280
rect 24084 13268 24090 13320
rect 20772 13212 22692 13240
rect 20772 13200 20778 13212
rect 1854 13172 1860 13184
rect 1815 13144 1860 13172
rect 1854 13132 1860 13144
rect 1912 13132 1918 13184
rect 2130 13132 2136 13184
rect 2188 13172 2194 13184
rect 2225 13175 2283 13181
rect 2225 13172 2237 13175
rect 2188 13144 2237 13172
rect 2188 13132 2194 13144
rect 2225 13141 2237 13144
rect 2271 13141 2283 13175
rect 2225 13135 2283 13141
rect 2498 13132 2504 13184
rect 2556 13172 2562 13184
rect 2685 13175 2743 13181
rect 2685 13172 2697 13175
rect 2556 13144 2697 13172
rect 2556 13132 2562 13144
rect 2685 13141 2697 13144
rect 2731 13172 2743 13175
rect 2866 13172 2872 13184
rect 2731 13144 2872 13172
rect 2731 13141 2743 13144
rect 2685 13135 2743 13141
rect 2866 13132 2872 13144
rect 2924 13132 2930 13184
rect 3881 13175 3939 13181
rect 3881 13141 3893 13175
rect 3927 13172 3939 13175
rect 5350 13172 5356 13184
rect 3927 13144 5356 13172
rect 3927 13141 3939 13144
rect 3881 13135 3939 13141
rect 5350 13132 5356 13144
rect 5408 13132 5414 13184
rect 7469 13175 7527 13181
rect 7469 13141 7481 13175
rect 7515 13172 7527 13175
rect 7650 13172 7656 13184
rect 7515 13144 7656 13172
rect 7515 13141 7527 13144
rect 7469 13135 7527 13141
rect 7650 13132 7656 13144
rect 7708 13132 7714 13184
rect 9306 13132 9312 13184
rect 9364 13172 9370 13184
rect 10597 13175 10655 13181
rect 10597 13172 10609 13175
rect 9364 13144 10609 13172
rect 9364 13132 9370 13144
rect 10597 13141 10609 13144
rect 10643 13141 10655 13175
rect 13998 13172 14004 13184
rect 13959 13144 14004 13172
rect 10597 13135 10655 13141
rect 13998 13132 14004 13144
rect 14056 13132 14062 13184
rect 15746 13132 15752 13184
rect 15804 13172 15810 13184
rect 16114 13172 16120 13184
rect 15804 13144 16120 13172
rect 15804 13132 15810 13144
rect 16114 13132 16120 13144
rect 16172 13172 16178 13184
rect 16301 13175 16359 13181
rect 16301 13172 16313 13175
rect 16172 13144 16313 13172
rect 16172 13132 16178 13144
rect 16301 13141 16313 13144
rect 16347 13141 16359 13175
rect 16301 13135 16359 13141
rect 18141 13175 18199 13181
rect 18141 13141 18153 13175
rect 18187 13172 18199 13175
rect 18782 13172 18788 13184
rect 18187 13144 18788 13172
rect 18187 13141 18199 13144
rect 18141 13135 18199 13141
rect 18782 13132 18788 13144
rect 18840 13132 18846 13184
rect 19978 13172 19984 13184
rect 19939 13144 19984 13172
rect 19978 13132 19984 13144
rect 20036 13132 20042 13184
rect 21542 13172 21548 13184
rect 21503 13144 21548 13172
rect 21542 13132 21548 13144
rect 21600 13132 21606 13184
rect 24670 13132 24676 13184
rect 24728 13172 24734 13184
rect 25179 13175 25237 13181
rect 25179 13172 25191 13175
rect 24728 13144 25191 13172
rect 24728 13132 24734 13144
rect 25179 13141 25191 13144
rect 25225 13141 25237 13175
rect 25179 13135 25237 13141
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1627 12971 1685 12977
rect 1627 12937 1639 12971
rect 1673 12968 1685 12971
rect 1946 12968 1952 12980
rect 1673 12940 1952 12968
rect 1673 12937 1685 12940
rect 1627 12931 1685 12937
rect 1946 12928 1952 12940
rect 2004 12928 2010 12980
rect 2133 12971 2191 12977
rect 2133 12937 2145 12971
rect 2179 12968 2191 12971
rect 2406 12968 2412 12980
rect 2179 12940 2412 12968
rect 2179 12937 2191 12940
rect 2133 12931 2191 12937
rect 2406 12928 2412 12940
rect 2464 12968 2470 12980
rect 8846 12968 8852 12980
rect 2464 12940 2728 12968
rect 8807 12940 8852 12968
rect 2464 12928 2470 12940
rect 2700 12909 2728 12940
rect 8846 12928 8852 12940
rect 8904 12928 8910 12980
rect 9306 12968 9312 12980
rect 9267 12940 9312 12968
rect 9306 12928 9312 12940
rect 9364 12928 9370 12980
rect 9677 12971 9735 12977
rect 9677 12937 9689 12971
rect 9723 12968 9735 12971
rect 10134 12968 10140 12980
rect 9723 12940 10140 12968
rect 9723 12937 9735 12940
rect 9677 12931 9735 12937
rect 10134 12928 10140 12940
rect 10192 12928 10198 12980
rect 10778 12968 10784 12980
rect 10739 12940 10784 12968
rect 10778 12928 10784 12940
rect 10836 12928 10842 12980
rect 12250 12968 12256 12980
rect 12211 12940 12256 12968
rect 12250 12928 12256 12940
rect 12308 12968 12314 12980
rect 13633 12971 13691 12977
rect 13633 12968 13645 12971
rect 12308 12940 13645 12968
rect 12308 12928 12314 12940
rect 2685 12903 2743 12909
rect 2685 12869 2697 12903
rect 2731 12869 2743 12903
rect 2685 12863 2743 12869
rect 2866 12860 2872 12912
rect 2924 12900 2930 12912
rect 6549 12903 6607 12909
rect 6549 12900 6561 12903
rect 2924 12872 6561 12900
rect 2924 12860 2930 12872
rect 6549 12869 6561 12872
rect 6595 12900 6607 12903
rect 6822 12900 6828 12912
rect 6595 12872 6828 12900
rect 6595 12869 6607 12872
rect 6549 12863 6607 12869
rect 6822 12860 6828 12872
rect 6880 12900 6886 12912
rect 7469 12903 7527 12909
rect 7469 12900 7481 12903
rect 6880 12872 7481 12900
rect 6880 12860 6886 12872
rect 7469 12869 7481 12872
rect 7515 12869 7527 12903
rect 10410 12900 10416 12912
rect 10371 12872 10416 12900
rect 7469 12863 7527 12869
rect 10410 12860 10416 12872
rect 10468 12860 10474 12912
rect 3329 12835 3387 12841
rect 3329 12801 3341 12835
rect 3375 12832 3387 12835
rect 7926 12832 7932 12844
rect 3375 12804 7932 12832
rect 3375 12801 3387 12804
rect 3329 12795 3387 12801
rect 7926 12792 7932 12804
rect 7984 12792 7990 12844
rect 8110 12832 8116 12844
rect 8071 12804 8116 12832
rect 8110 12792 8116 12804
rect 8168 12792 8174 12844
rect 9490 12792 9496 12844
rect 9548 12832 9554 12844
rect 9861 12835 9919 12841
rect 9861 12832 9873 12835
rect 9548 12804 9873 12832
rect 9548 12792 9554 12804
rect 9861 12801 9873 12804
rect 9907 12832 9919 12835
rect 11471 12835 11529 12841
rect 11471 12832 11483 12835
rect 9907 12804 11483 12832
rect 9907 12801 9919 12804
rect 9861 12795 9919 12801
rect 11471 12801 11483 12804
rect 11517 12801 11529 12835
rect 12544 12832 12572 12940
rect 13633 12937 13645 12940
rect 13679 12937 13691 12971
rect 13998 12968 14004 12980
rect 13959 12940 14004 12968
rect 13633 12931 13691 12937
rect 13998 12928 14004 12940
rect 14056 12928 14062 12980
rect 15286 12968 15292 12980
rect 15247 12940 15292 12968
rect 15286 12928 15292 12940
rect 15344 12928 15350 12980
rect 16853 12971 16911 12977
rect 16853 12937 16865 12971
rect 16899 12968 16911 12971
rect 17126 12968 17132 12980
rect 16899 12940 17132 12968
rect 16899 12937 16911 12940
rect 16853 12931 16911 12937
rect 17126 12928 17132 12940
rect 17184 12928 17190 12980
rect 20070 12928 20076 12980
rect 20128 12968 20134 12980
rect 22186 12968 22192 12980
rect 20128 12940 22192 12968
rect 20128 12928 20134 12940
rect 22186 12928 22192 12940
rect 22244 12928 22250 12980
rect 22278 12928 22284 12980
rect 22336 12968 22342 12980
rect 22465 12971 22523 12977
rect 22465 12968 22477 12971
rect 22336 12940 22477 12968
rect 22336 12928 22342 12940
rect 22465 12937 22477 12940
rect 22511 12937 22523 12971
rect 22465 12931 22523 12937
rect 23474 12928 23480 12980
rect 23532 12968 23538 12980
rect 23845 12971 23903 12977
rect 23845 12968 23857 12971
rect 23532 12940 23857 12968
rect 23532 12928 23538 12940
rect 23845 12937 23857 12940
rect 23891 12937 23903 12971
rect 23845 12931 23903 12937
rect 23934 12928 23940 12980
rect 23992 12968 23998 12980
rect 24213 12971 24271 12977
rect 24213 12968 24225 12971
rect 23992 12940 24225 12968
rect 23992 12928 23998 12940
rect 24213 12937 24225 12940
rect 24259 12937 24271 12971
rect 25130 12968 25136 12980
rect 25091 12940 25136 12968
rect 24213 12931 24271 12937
rect 25130 12928 25136 12940
rect 25188 12928 25194 12980
rect 12618 12860 12624 12912
rect 12676 12900 12682 12912
rect 17773 12903 17831 12909
rect 17773 12900 17785 12903
rect 12676 12872 17785 12900
rect 12676 12860 12682 12872
rect 17773 12869 17785 12872
rect 17819 12869 17831 12903
rect 17773 12863 17831 12869
rect 14274 12832 14280 12844
rect 12544 12804 12801 12832
rect 14235 12804 14280 12832
rect 11471 12795 11529 12801
rect 1397 12767 1455 12773
rect 1397 12733 1409 12767
rect 1443 12764 1455 12767
rect 1578 12764 1584 12776
rect 1443 12736 1584 12764
rect 1443 12733 1455 12736
rect 1397 12727 1455 12733
rect 1578 12724 1584 12736
rect 1636 12724 1642 12776
rect 2590 12764 2596 12776
rect 2551 12736 2596 12764
rect 2590 12724 2596 12736
rect 2648 12724 2654 12776
rect 2869 12767 2927 12773
rect 2869 12733 2881 12767
rect 2915 12764 2927 12767
rect 3421 12767 3479 12773
rect 3421 12764 3433 12767
rect 2915 12736 3433 12764
rect 2915 12733 2927 12736
rect 2869 12727 2927 12733
rect 3421 12733 3433 12736
rect 3467 12733 3479 12767
rect 3421 12727 3479 12733
rect 4157 12767 4215 12773
rect 4157 12733 4169 12767
rect 4203 12733 4215 12767
rect 4157 12727 4215 12733
rect 1762 12656 1768 12708
rect 1820 12696 1826 12708
rect 2958 12696 2964 12708
rect 1820 12668 2964 12696
rect 1820 12656 1826 12668
rect 2958 12656 2964 12668
rect 3016 12696 3022 12708
rect 3973 12699 4031 12705
rect 3973 12696 3985 12699
rect 3016 12668 3985 12696
rect 3016 12656 3022 12668
rect 3973 12665 3985 12668
rect 4019 12696 4031 12699
rect 4172 12696 4200 12727
rect 4522 12724 4528 12776
rect 4580 12764 4586 12776
rect 4617 12767 4675 12773
rect 4617 12764 4629 12767
rect 4580 12736 4629 12764
rect 4580 12724 4586 12736
rect 4617 12733 4629 12736
rect 4663 12733 4675 12767
rect 4617 12727 4675 12733
rect 5169 12767 5227 12773
rect 5169 12733 5181 12767
rect 5215 12733 5227 12767
rect 5350 12764 5356 12776
rect 5311 12736 5356 12764
rect 5169 12727 5227 12733
rect 4338 12696 4344 12708
rect 4019 12668 4344 12696
rect 4019 12665 4031 12668
rect 3973 12659 4031 12665
rect 4338 12656 4344 12668
rect 4396 12656 4402 12708
rect 5184 12696 5212 12727
rect 5350 12724 5356 12736
rect 5408 12724 5414 12776
rect 7377 12767 7435 12773
rect 7377 12764 7389 12767
rect 7208 12736 7389 12764
rect 5184 12668 6040 12696
rect 6012 12640 6040 12668
rect 7208 12640 7236 12736
rect 7377 12733 7389 12736
rect 7423 12733 7435 12767
rect 7650 12764 7656 12776
rect 7611 12736 7656 12764
rect 7377 12727 7435 12733
rect 7650 12724 7656 12736
rect 7708 12724 7714 12776
rect 11368 12767 11426 12773
rect 11368 12733 11380 12767
rect 11414 12733 11426 12767
rect 11368 12727 11426 12733
rect 12437 12767 12495 12773
rect 12437 12733 12449 12767
rect 12483 12764 12495 12767
rect 12526 12764 12532 12776
rect 12483 12736 12532 12764
rect 12483 12733 12495 12736
rect 12437 12727 12495 12733
rect 9306 12656 9312 12708
rect 9364 12696 9370 12708
rect 9953 12699 10011 12705
rect 9953 12696 9965 12699
rect 9364 12668 9965 12696
rect 9364 12656 9370 12668
rect 9953 12665 9965 12668
rect 9999 12665 10011 12699
rect 11383 12696 11411 12727
rect 12526 12724 12532 12736
rect 12584 12724 12590 12776
rect 12773 12708 12801 12804
rect 14274 12792 14280 12804
rect 14332 12792 14338 12844
rect 15746 12764 15752 12776
rect 15707 12736 15752 12764
rect 15746 12724 15752 12736
rect 15804 12724 15810 12776
rect 16298 12764 16304 12776
rect 16259 12736 16304 12764
rect 16298 12724 16304 12736
rect 16356 12724 16362 12776
rect 17788 12764 17816 12863
rect 18322 12860 18328 12912
rect 18380 12900 18386 12912
rect 19061 12903 19119 12909
rect 19061 12900 19073 12903
rect 18380 12872 19073 12900
rect 18380 12860 18386 12872
rect 19061 12869 19073 12872
rect 19107 12869 19119 12903
rect 20530 12900 20536 12912
rect 20491 12872 20536 12900
rect 19061 12863 19119 12869
rect 20530 12860 20536 12872
rect 20588 12860 20594 12912
rect 24762 12900 24768 12912
rect 24723 12872 24768 12900
rect 24762 12860 24768 12872
rect 24820 12860 24826 12912
rect 18598 12832 18604 12844
rect 18559 12804 18604 12832
rect 18598 12792 18604 12804
rect 18656 12792 18662 12844
rect 20070 12792 20076 12844
rect 20128 12832 20134 12844
rect 21821 12835 21879 12841
rect 21821 12832 21833 12835
rect 20128 12804 21833 12832
rect 20128 12792 20134 12804
rect 21821 12801 21833 12804
rect 21867 12801 21879 12835
rect 21821 12795 21879 12801
rect 18049 12767 18107 12773
rect 18049 12764 18061 12767
rect 17788 12736 18061 12764
rect 18049 12733 18061 12736
rect 18095 12764 18107 12767
rect 18414 12764 18420 12776
rect 18095 12736 18420 12764
rect 18095 12733 18107 12736
rect 18049 12727 18107 12733
rect 18414 12724 18420 12736
rect 18472 12724 18478 12776
rect 18509 12767 18567 12773
rect 18509 12733 18521 12767
rect 18555 12764 18567 12767
rect 18782 12764 18788 12776
rect 18555 12736 18788 12764
rect 18555 12733 18567 12736
rect 18509 12727 18567 12733
rect 18782 12724 18788 12736
rect 18840 12724 18846 12776
rect 24581 12767 24639 12773
rect 24581 12733 24593 12767
rect 24627 12764 24639 12767
rect 24670 12764 24676 12776
rect 24627 12736 24676 12764
rect 24627 12733 24639 12736
rect 24581 12727 24639 12733
rect 24670 12724 24676 12736
rect 24728 12724 24734 12776
rect 11793 12699 11851 12705
rect 11793 12696 11805 12699
rect 9953 12659 10011 12665
rect 10146 12668 11805 12696
rect 3421 12631 3479 12637
rect 3421 12597 3433 12631
rect 3467 12628 3479 12631
rect 3697 12631 3755 12637
rect 3697 12628 3709 12631
rect 3467 12600 3709 12628
rect 3467 12597 3479 12600
rect 3421 12591 3479 12597
rect 3697 12597 3709 12600
rect 3743 12628 3755 12631
rect 3878 12628 3884 12640
rect 3743 12600 3884 12628
rect 3743 12597 3755 12600
rect 3697 12591 3755 12597
rect 3878 12588 3884 12600
rect 3936 12588 3942 12640
rect 4246 12628 4252 12640
rect 4207 12600 4252 12628
rect 4246 12588 4252 12600
rect 4304 12588 4310 12640
rect 5994 12628 6000 12640
rect 5955 12600 6000 12628
rect 5994 12588 6000 12600
rect 6052 12588 6058 12640
rect 7190 12628 7196 12640
rect 7151 12600 7196 12628
rect 7190 12588 7196 12600
rect 7248 12588 7254 12640
rect 8294 12588 8300 12640
rect 8352 12628 8358 12640
rect 8481 12631 8539 12637
rect 8481 12628 8493 12631
rect 8352 12600 8493 12628
rect 8352 12588 8358 12600
rect 8481 12597 8493 12600
rect 8527 12628 8539 12631
rect 9030 12628 9036 12640
rect 8527 12600 9036 12628
rect 8527 12597 8539 12600
rect 8481 12591 8539 12597
rect 9030 12588 9036 12600
rect 9088 12588 9094 12640
rect 9674 12588 9680 12640
rect 9732 12628 9738 12640
rect 10146 12628 10174 12668
rect 11793 12665 11805 12668
rect 11839 12665 11851 12699
rect 12710 12696 12716 12708
rect 12668 12668 12716 12696
rect 11793 12659 11851 12665
rect 12710 12656 12716 12668
rect 12768 12705 12801 12708
rect 12768 12699 12816 12705
rect 12768 12665 12770 12699
rect 12804 12665 12816 12699
rect 12768 12659 12816 12665
rect 12768 12656 12774 12659
rect 13170 12656 13176 12708
rect 13228 12696 13234 12708
rect 13722 12696 13728 12708
rect 13228 12668 13728 12696
rect 13228 12656 13234 12668
rect 13722 12656 13728 12668
rect 13780 12656 13786 12708
rect 14369 12699 14427 12705
rect 14369 12665 14381 12699
rect 14415 12665 14427 12699
rect 14918 12696 14924 12708
rect 14879 12668 14924 12696
rect 14369 12659 14427 12665
rect 9732 12600 10174 12628
rect 11241 12631 11299 12637
rect 9732 12588 9738 12600
rect 11241 12597 11253 12631
rect 11287 12628 11299 12631
rect 11422 12628 11428 12640
rect 11287 12600 11428 12628
rect 11287 12597 11299 12600
rect 11241 12591 11299 12597
rect 11422 12588 11428 12600
rect 11480 12588 11486 12640
rect 13357 12631 13415 12637
rect 13357 12597 13369 12631
rect 13403 12628 13415 12631
rect 13538 12628 13544 12640
rect 13403 12600 13544 12628
rect 13403 12597 13415 12600
rect 13357 12591 13415 12597
rect 13538 12588 13544 12600
rect 13596 12588 13602 12640
rect 13998 12588 14004 12640
rect 14056 12628 14062 12640
rect 14384 12628 14412 12659
rect 14918 12656 14924 12668
rect 14976 12656 14982 12708
rect 17497 12699 17555 12705
rect 17497 12665 17509 12699
rect 17543 12696 17555 12699
rect 18230 12696 18236 12708
rect 17543 12668 18236 12696
rect 17543 12665 17555 12668
rect 17497 12659 17555 12665
rect 18230 12656 18236 12668
rect 18288 12656 18294 12708
rect 19978 12696 19984 12708
rect 19939 12668 19984 12696
rect 19978 12656 19984 12668
rect 20036 12656 20042 12708
rect 20073 12699 20131 12705
rect 20073 12665 20085 12699
rect 20119 12665 20131 12699
rect 21542 12696 21548 12708
rect 21503 12668 21548 12696
rect 20073 12659 20131 12665
rect 15838 12628 15844 12640
rect 14056 12600 14412 12628
rect 15799 12600 15844 12628
rect 14056 12588 14062 12600
rect 15838 12588 15844 12600
rect 15896 12588 15902 12640
rect 19518 12588 19524 12640
rect 19576 12628 19582 12640
rect 19797 12631 19855 12637
rect 19797 12628 19809 12631
rect 19576 12600 19809 12628
rect 19576 12588 19582 12600
rect 19797 12597 19809 12600
rect 19843 12628 19855 12631
rect 20088 12628 20116 12659
rect 21542 12656 21548 12668
rect 21600 12656 21606 12708
rect 21637 12699 21695 12705
rect 21637 12665 21649 12699
rect 21683 12665 21695 12699
rect 21637 12659 21695 12665
rect 19843 12600 20116 12628
rect 19843 12597 19855 12600
rect 19797 12591 19855 12597
rect 21082 12588 21088 12640
rect 21140 12628 21146 12640
rect 21269 12631 21327 12637
rect 21269 12628 21281 12631
rect 21140 12600 21281 12628
rect 21140 12588 21146 12600
rect 21269 12597 21281 12600
rect 21315 12628 21327 12631
rect 21652 12628 21680 12659
rect 21315 12600 21680 12628
rect 21315 12597 21327 12600
rect 21269 12591 21327 12597
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1581 12427 1639 12433
rect 1581 12393 1593 12427
rect 1627 12424 1639 12427
rect 1762 12424 1768 12436
rect 1627 12396 1768 12424
rect 1627 12393 1639 12396
rect 1581 12387 1639 12393
rect 1762 12384 1768 12396
rect 1820 12384 1826 12436
rect 1949 12427 2007 12433
rect 1949 12393 1961 12427
rect 1995 12424 2007 12427
rect 2222 12424 2228 12436
rect 1995 12396 2228 12424
rect 1995 12393 2007 12396
rect 1949 12387 2007 12393
rect 2222 12384 2228 12396
rect 2280 12384 2286 12436
rect 3142 12384 3148 12436
rect 3200 12424 3206 12436
rect 3789 12427 3847 12433
rect 3789 12424 3801 12427
rect 3200 12396 3801 12424
rect 3200 12384 3206 12396
rect 3789 12393 3801 12396
rect 3835 12424 3847 12427
rect 3970 12424 3976 12436
rect 3835 12396 3976 12424
rect 3835 12393 3847 12396
rect 3789 12387 3847 12393
rect 3970 12384 3976 12396
rect 4028 12384 4034 12436
rect 4614 12424 4620 12436
rect 4575 12396 4620 12424
rect 4614 12384 4620 12396
rect 4672 12384 4678 12436
rect 6454 12424 6460 12436
rect 6415 12396 6460 12424
rect 6454 12384 6460 12396
rect 6512 12384 6518 12436
rect 6822 12424 6828 12436
rect 6783 12396 6828 12424
rect 6822 12384 6828 12396
rect 6880 12424 6886 12436
rect 9490 12424 9496 12436
rect 6880 12396 7512 12424
rect 9451 12396 9496 12424
rect 6880 12384 6886 12396
rect 2590 12316 2596 12368
rect 2648 12356 2654 12368
rect 3513 12359 3571 12365
rect 3513 12356 3525 12359
rect 2648 12328 3525 12356
rect 2648 12316 2654 12328
rect 3513 12325 3525 12328
rect 3559 12356 3571 12359
rect 5994 12356 6000 12368
rect 3559 12328 6000 12356
rect 3559 12325 3571 12328
rect 3513 12319 3571 12325
rect 1394 12288 1400 12300
rect 1355 12260 1400 12288
rect 1394 12248 1400 12260
rect 1452 12248 1458 12300
rect 2406 12288 2412 12300
rect 2367 12260 2412 12288
rect 2406 12248 2412 12260
rect 2464 12248 2470 12300
rect 2685 12291 2743 12297
rect 2685 12257 2697 12291
rect 2731 12288 2743 12291
rect 3050 12288 3056 12300
rect 2731 12260 3056 12288
rect 2731 12257 2743 12260
rect 2685 12251 2743 12257
rect 3050 12248 3056 12260
rect 3108 12248 3114 12300
rect 4338 12288 4344 12300
rect 4299 12260 4344 12288
rect 4338 12248 4344 12260
rect 4396 12248 4402 12300
rect 4522 12248 4528 12300
rect 4580 12288 4586 12300
rect 5368 12297 5396 12328
rect 5994 12316 6000 12328
rect 6052 12316 6058 12368
rect 6362 12316 6368 12368
rect 6420 12356 6426 12368
rect 7193 12359 7251 12365
rect 7193 12356 7205 12359
rect 6420 12328 7205 12356
rect 6420 12316 6426 12328
rect 7193 12325 7205 12328
rect 7239 12356 7251 12359
rect 7282 12356 7288 12368
rect 7239 12328 7288 12356
rect 7239 12325 7251 12328
rect 7193 12319 7251 12325
rect 7282 12316 7288 12328
rect 7340 12316 7346 12368
rect 4801 12291 4859 12297
rect 4801 12288 4813 12291
rect 4580 12260 4813 12288
rect 4580 12248 4586 12260
rect 4801 12257 4813 12260
rect 4847 12257 4859 12291
rect 4801 12251 4859 12257
rect 5353 12291 5411 12297
rect 5353 12257 5365 12291
rect 5399 12257 5411 12291
rect 5353 12251 5411 12257
rect 5721 12291 5779 12297
rect 5721 12257 5733 12291
rect 5767 12288 5779 12291
rect 6178 12288 6184 12300
rect 5767 12260 6184 12288
rect 5767 12257 5779 12260
rect 5721 12251 5779 12257
rect 2317 12223 2375 12229
rect 2317 12189 2329 12223
rect 2363 12220 2375 12223
rect 2498 12220 2504 12232
rect 2363 12192 2504 12220
rect 2363 12189 2375 12192
rect 2317 12183 2375 12189
rect 2498 12180 2504 12192
rect 2556 12180 2562 12232
rect 3142 12220 3148 12232
rect 3103 12192 3148 12220
rect 3142 12180 3148 12192
rect 3200 12180 3206 12232
rect 4816 12220 4844 12251
rect 6178 12248 6184 12260
rect 6236 12248 6242 12300
rect 7374 12288 7380 12300
rect 7335 12260 7380 12288
rect 7374 12248 7380 12260
rect 7432 12248 7438 12300
rect 7484 12297 7512 12396
rect 9490 12384 9496 12396
rect 9548 12384 9554 12436
rect 9766 12424 9772 12436
rect 9727 12396 9772 12424
rect 9766 12384 9772 12396
rect 9824 12384 9830 12436
rect 11517 12427 11575 12433
rect 11517 12393 11529 12427
rect 11563 12424 11575 12427
rect 11882 12424 11888 12436
rect 11563 12396 11888 12424
rect 11563 12393 11575 12396
rect 11517 12387 11575 12393
rect 11882 12384 11888 12396
rect 11940 12424 11946 12436
rect 14826 12424 14832 12436
rect 11940 12396 14832 12424
rect 11940 12384 11946 12396
rect 14826 12384 14832 12396
rect 14884 12384 14890 12436
rect 17034 12424 17040 12436
rect 16995 12396 17040 12424
rect 17034 12384 17040 12396
rect 17092 12384 17098 12436
rect 18322 12424 18328 12436
rect 18283 12396 18328 12424
rect 18322 12384 18328 12396
rect 18380 12384 18386 12436
rect 20346 12384 20352 12436
rect 20404 12424 20410 12436
rect 20625 12427 20683 12433
rect 20625 12424 20637 12427
rect 20404 12396 20637 12424
rect 20404 12384 20410 12396
rect 20625 12393 20637 12396
rect 20671 12393 20683 12427
rect 20625 12387 20683 12393
rect 8113 12359 8171 12365
rect 8113 12325 8125 12359
rect 8159 12356 8171 12359
rect 8478 12356 8484 12368
rect 8159 12328 8484 12356
rect 8159 12325 8171 12328
rect 8113 12319 8171 12325
rect 8478 12316 8484 12328
rect 8536 12316 8542 12368
rect 12529 12359 12587 12365
rect 12529 12325 12541 12359
rect 12575 12356 12587 12359
rect 13078 12356 13084 12368
rect 12575 12328 13084 12356
rect 12575 12325 12587 12328
rect 12529 12319 12587 12325
rect 13078 12316 13084 12328
rect 13136 12316 13142 12368
rect 13538 12356 13544 12368
rect 13499 12328 13544 12356
rect 13538 12316 13544 12328
rect 13596 12316 13602 12368
rect 14093 12359 14151 12365
rect 14093 12325 14105 12359
rect 14139 12356 14151 12359
rect 14918 12356 14924 12368
rect 14139 12328 14924 12356
rect 14139 12325 14151 12328
rect 14093 12319 14151 12325
rect 14918 12316 14924 12328
rect 14976 12316 14982 12368
rect 19426 12356 19432 12368
rect 19387 12328 19432 12356
rect 19426 12316 19432 12328
rect 19484 12316 19490 12368
rect 19981 12359 20039 12365
rect 19981 12325 19993 12359
rect 20027 12356 20039 12359
rect 20070 12356 20076 12368
rect 20027 12328 20076 12356
rect 20027 12325 20039 12328
rect 19981 12319 20039 12325
rect 20070 12316 20076 12328
rect 20128 12316 20134 12368
rect 20640 12356 20668 12387
rect 21542 12384 21548 12436
rect 21600 12424 21606 12436
rect 23615 12427 23673 12433
rect 23615 12424 23627 12427
rect 21600 12396 23627 12424
rect 21600 12384 21606 12396
rect 23615 12393 23627 12396
rect 23661 12393 23673 12427
rect 24670 12424 24676 12436
rect 24631 12396 24676 12424
rect 23615 12387 23673 12393
rect 24670 12384 24676 12396
rect 24728 12384 24734 12436
rect 20993 12359 21051 12365
rect 20993 12356 21005 12359
rect 20640 12328 21005 12356
rect 20993 12325 21005 12328
rect 21039 12325 21051 12359
rect 20993 12319 21051 12325
rect 21082 12316 21088 12368
rect 21140 12356 21146 12368
rect 21140 12328 21185 12356
rect 21140 12316 21146 12328
rect 7469 12291 7527 12297
rect 7469 12257 7481 12291
rect 7515 12257 7527 12291
rect 7650 12288 7656 12300
rect 7563 12260 7656 12288
rect 7469 12251 7527 12257
rect 7650 12248 7656 12260
rect 7708 12248 7714 12300
rect 9953 12291 10011 12297
rect 9953 12257 9965 12291
rect 9999 12257 10011 12291
rect 9953 12251 10011 12257
rect 10229 12291 10287 12297
rect 10229 12257 10241 12291
rect 10275 12288 10287 12291
rect 10686 12288 10692 12300
rect 10275 12260 10692 12288
rect 10275 12257 10287 12260
rect 10229 12251 10287 12257
rect 6089 12223 6147 12229
rect 6089 12220 6101 12223
rect 4816 12192 6101 12220
rect 6089 12189 6101 12192
rect 6135 12189 6147 12223
rect 6089 12183 6147 12189
rect 3050 12112 3056 12164
rect 3108 12152 3114 12164
rect 7668 12152 7696 12248
rect 9030 12180 9036 12232
rect 9088 12220 9094 12232
rect 9968 12220 9996 12251
rect 10686 12248 10692 12260
rect 10744 12288 10750 12300
rect 11330 12288 11336 12300
rect 10744 12260 11336 12288
rect 10744 12248 10750 12260
rect 11330 12248 11336 12260
rect 11388 12248 11394 12300
rect 11422 12248 11428 12300
rect 11480 12288 11486 12300
rect 11882 12288 11888 12300
rect 11480 12260 11888 12288
rect 11480 12248 11486 12260
rect 11882 12248 11888 12260
rect 11940 12248 11946 12300
rect 12345 12291 12403 12297
rect 12345 12257 12357 12291
rect 12391 12257 12403 12291
rect 15562 12288 15568 12300
rect 15523 12260 15568 12288
rect 12345 12251 12403 12257
rect 11440 12220 11468 12248
rect 9088 12192 11468 12220
rect 9088 12180 9094 12192
rect 8570 12152 8576 12164
rect 3108 12124 8576 12152
rect 3108 12112 3114 12124
rect 6104 12096 6132 12124
rect 8570 12112 8576 12124
rect 8628 12112 8634 12164
rect 12250 12112 12256 12164
rect 12308 12152 12314 12164
rect 12360 12152 12388 12251
rect 15562 12248 15568 12260
rect 15620 12248 15626 12300
rect 15654 12248 15660 12300
rect 15712 12288 15718 12300
rect 16025 12291 16083 12297
rect 16025 12288 16037 12291
rect 15712 12260 16037 12288
rect 15712 12248 15718 12260
rect 16025 12257 16037 12260
rect 16071 12288 16083 12291
rect 16298 12288 16304 12300
rect 16071 12260 16304 12288
rect 16071 12257 16083 12260
rect 16025 12251 16083 12257
rect 16298 12248 16304 12260
rect 16356 12288 16362 12300
rect 17218 12288 17224 12300
rect 16356 12260 16712 12288
rect 17179 12260 17224 12288
rect 16356 12248 16362 12260
rect 13446 12220 13452 12232
rect 13407 12192 13452 12220
rect 13446 12180 13452 12192
rect 13504 12180 13510 12232
rect 15746 12220 15752 12232
rect 13786 12192 15752 12220
rect 13786 12152 13814 12192
rect 15746 12180 15752 12192
rect 15804 12180 15810 12232
rect 16114 12220 16120 12232
rect 16075 12192 16120 12220
rect 16114 12180 16120 12192
rect 16172 12180 16178 12232
rect 16684 12229 16712 12260
rect 17218 12248 17224 12260
rect 17276 12248 17282 12300
rect 17678 12288 17684 12300
rect 17639 12260 17684 12288
rect 17678 12248 17684 12260
rect 17736 12248 17742 12300
rect 22462 12288 22468 12300
rect 22423 12260 22468 12288
rect 22462 12248 22468 12260
rect 22520 12248 22526 12300
rect 23544 12291 23602 12297
rect 23544 12257 23556 12291
rect 23590 12288 23602 12291
rect 23658 12288 23664 12300
rect 23590 12260 23664 12288
rect 23590 12257 23602 12260
rect 23544 12251 23602 12257
rect 23658 12248 23664 12260
rect 23716 12248 23722 12300
rect 16669 12223 16727 12229
rect 16669 12189 16681 12223
rect 16715 12220 16727 12223
rect 17696 12220 17724 12248
rect 16715 12192 17724 12220
rect 17957 12223 18015 12229
rect 16715 12189 16727 12192
rect 16669 12183 16727 12189
rect 17957 12189 17969 12223
rect 18003 12220 18015 12223
rect 18322 12220 18328 12232
rect 18003 12192 18328 12220
rect 18003 12189 18015 12192
rect 17957 12183 18015 12189
rect 18322 12180 18328 12192
rect 18380 12220 18386 12232
rect 18693 12223 18751 12229
rect 18693 12220 18705 12223
rect 18380 12192 18705 12220
rect 18380 12180 18386 12192
rect 18693 12189 18705 12192
rect 18739 12189 18751 12223
rect 18693 12183 18751 12189
rect 19150 12180 19156 12232
rect 19208 12220 19214 12232
rect 19337 12223 19395 12229
rect 19337 12220 19349 12223
rect 19208 12192 19349 12220
rect 19208 12180 19214 12192
rect 19337 12189 19349 12192
rect 19383 12220 19395 12223
rect 21266 12220 21272 12232
rect 19383 12192 20116 12220
rect 21227 12192 21272 12220
rect 19383 12189 19395 12192
rect 19337 12183 19395 12189
rect 12308 12124 13814 12152
rect 20088 12152 20116 12192
rect 21266 12180 21272 12192
rect 21324 12180 21330 12232
rect 22603 12155 22661 12161
rect 22603 12152 22615 12155
rect 20088 12124 22615 12152
rect 12308 12112 12314 12124
rect 22603 12121 22615 12124
rect 22649 12121 22661 12155
rect 22603 12115 22661 12121
rect 6086 12044 6092 12096
rect 6144 12044 6150 12096
rect 9950 12044 9956 12096
rect 10008 12084 10014 12096
rect 10689 12087 10747 12093
rect 10689 12084 10701 12087
rect 10008 12056 10701 12084
rect 10008 12044 10014 12056
rect 10689 12053 10701 12056
rect 10735 12053 10747 12087
rect 10689 12047 10747 12053
rect 11238 12044 11244 12096
rect 11296 12084 11302 12096
rect 14090 12084 14096 12096
rect 11296 12056 14096 12084
rect 11296 12044 11302 12056
rect 14090 12044 14096 12056
rect 14148 12084 14154 12096
rect 14642 12084 14648 12096
rect 14148 12056 14648 12084
rect 14148 12044 14154 12056
rect 14642 12044 14648 12056
rect 14700 12044 14706 12096
rect 21358 12044 21364 12096
rect 21416 12084 21422 12096
rect 21913 12087 21971 12093
rect 21913 12084 21925 12087
rect 21416 12056 21925 12084
rect 21416 12044 21422 12056
rect 21913 12053 21925 12056
rect 21959 12084 21971 12087
rect 22002 12084 22008 12096
rect 21959 12056 22008 12084
rect 21959 12053 21971 12056
rect 21913 12047 21971 12053
rect 22002 12044 22008 12056
rect 22060 12044 22066 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 2406 11840 2412 11892
rect 2464 11880 2470 11892
rect 2869 11883 2927 11889
rect 2869 11880 2881 11883
rect 2464 11852 2881 11880
rect 2464 11840 2470 11852
rect 2869 11849 2881 11852
rect 2915 11880 2927 11883
rect 4154 11880 4160 11892
rect 2915 11852 4160 11880
rect 2915 11849 2927 11852
rect 2869 11843 2927 11849
rect 4154 11840 4160 11852
rect 4212 11840 4218 11892
rect 5813 11883 5871 11889
rect 5813 11849 5825 11883
rect 5859 11880 5871 11883
rect 5994 11880 6000 11892
rect 5859 11852 6000 11880
rect 5859 11849 5871 11852
rect 5813 11843 5871 11849
rect 5994 11840 6000 11852
rect 6052 11880 6058 11892
rect 7374 11880 7380 11892
rect 6052 11852 7380 11880
rect 6052 11840 6058 11852
rect 7374 11840 7380 11852
rect 7432 11880 7438 11892
rect 8570 11880 8576 11892
rect 7432 11852 8340 11880
rect 8531 11852 8576 11880
rect 7432 11840 7438 11852
rect 3881 11815 3939 11821
rect 3881 11781 3893 11815
rect 3927 11812 3939 11815
rect 4338 11812 4344 11824
rect 3927 11784 4344 11812
rect 3927 11781 3939 11784
rect 3881 11775 3939 11781
rect 4338 11772 4344 11784
rect 4396 11812 4402 11824
rect 7009 11815 7067 11821
rect 7009 11812 7021 11815
rect 4396 11784 7021 11812
rect 4396 11772 4402 11784
rect 7009 11781 7021 11784
rect 7055 11812 7067 11815
rect 7055 11784 7512 11812
rect 7055 11781 7067 11784
rect 7009 11775 7067 11781
rect 1394 11704 1400 11756
rect 1452 11744 1458 11756
rect 1673 11747 1731 11753
rect 1673 11744 1685 11747
rect 1452 11716 1685 11744
rect 1452 11704 1458 11716
rect 1673 11713 1685 11716
rect 1719 11744 1731 11747
rect 3786 11744 3792 11756
rect 1719 11716 3792 11744
rect 1719 11713 1731 11716
rect 1673 11707 1731 11713
rect 3786 11704 3792 11716
rect 3844 11704 3850 11756
rect 7282 11744 7288 11756
rect 7243 11716 7288 11744
rect 7282 11704 7288 11716
rect 7340 11704 7346 11756
rect 1854 11676 1860 11688
rect 1815 11648 1860 11676
rect 1854 11636 1860 11648
rect 1912 11636 1918 11688
rect 3970 11676 3976 11688
rect 3931 11648 3976 11676
rect 3970 11636 3976 11648
rect 4028 11636 4034 11688
rect 4522 11676 4528 11688
rect 4483 11648 4528 11676
rect 4522 11636 4528 11648
rect 4580 11636 4586 11688
rect 4801 11679 4859 11685
rect 4801 11645 4813 11679
rect 4847 11645 4859 11679
rect 5350 11676 5356 11688
rect 5311 11648 5356 11676
rect 4801 11639 4859 11645
rect 3513 11611 3571 11617
rect 3513 11577 3525 11611
rect 3559 11608 3571 11611
rect 4430 11608 4436 11620
rect 3559 11580 4436 11608
rect 3559 11577 3571 11580
rect 3513 11571 3571 11577
rect 4430 11568 4436 11580
rect 4488 11608 4494 11620
rect 4816 11608 4844 11639
rect 5350 11636 5356 11648
rect 5408 11636 5414 11688
rect 6917 11679 6975 11685
rect 6917 11645 6929 11679
rect 6963 11676 6975 11679
rect 7190 11676 7196 11688
rect 6963 11648 7196 11676
rect 6963 11645 6975 11648
rect 6917 11639 6975 11645
rect 7190 11636 7196 11648
rect 7248 11636 7254 11688
rect 7374 11636 7380 11688
rect 7432 11676 7438 11688
rect 7484 11685 7512 11784
rect 7929 11747 7987 11753
rect 7929 11713 7941 11747
rect 7975 11744 7987 11747
rect 8018 11744 8024 11756
rect 7975 11716 8024 11744
rect 7975 11713 7987 11716
rect 7929 11707 7987 11713
rect 8018 11704 8024 11716
rect 8076 11704 8082 11756
rect 8312 11753 8340 11852
rect 8570 11840 8576 11852
rect 8628 11840 8634 11892
rect 9030 11880 9036 11892
rect 8991 11852 9036 11880
rect 9030 11840 9036 11852
rect 9088 11840 9094 11892
rect 9309 11883 9367 11889
rect 9309 11849 9321 11883
rect 9355 11880 9367 11883
rect 9858 11880 9864 11892
rect 9355 11852 9864 11880
rect 9355 11849 9367 11852
rect 9309 11843 9367 11849
rect 9858 11840 9864 11852
rect 9916 11840 9922 11892
rect 12250 11880 12256 11892
rect 12211 11852 12256 11880
rect 12250 11840 12256 11852
rect 12308 11840 12314 11892
rect 13446 11840 13452 11892
rect 13504 11880 13510 11892
rect 14458 11880 14464 11892
rect 13504 11852 14464 11880
rect 13504 11840 13510 11852
rect 14458 11840 14464 11852
rect 14516 11840 14522 11892
rect 14826 11840 14832 11892
rect 14884 11880 14890 11892
rect 15197 11883 15255 11889
rect 15197 11880 15209 11883
rect 14884 11852 15209 11880
rect 14884 11840 14890 11852
rect 15197 11849 15209 11852
rect 15243 11880 15255 11883
rect 17310 11880 17316 11892
rect 15243 11852 17316 11880
rect 15243 11849 15255 11852
rect 15197 11843 15255 11849
rect 17310 11840 17316 11852
rect 17368 11840 17374 11892
rect 18690 11840 18696 11892
rect 18748 11880 18754 11892
rect 22462 11880 22468 11892
rect 18748 11852 22468 11880
rect 18748 11840 18754 11852
rect 22462 11840 22468 11852
rect 22520 11880 22526 11892
rect 22741 11883 22799 11889
rect 22741 11880 22753 11883
rect 22520 11852 22753 11880
rect 22520 11840 22526 11852
rect 22741 11849 22753 11852
rect 22787 11849 22799 11883
rect 22741 11843 22799 11849
rect 23658 11840 23664 11892
rect 23716 11880 23722 11892
rect 23845 11883 23903 11889
rect 23845 11880 23857 11883
rect 23716 11852 23857 11880
rect 23716 11840 23722 11852
rect 23845 11849 23857 11852
rect 23891 11849 23903 11883
rect 23845 11843 23903 11849
rect 11238 11812 11244 11824
rect 9692 11784 11244 11812
rect 8297 11747 8355 11753
rect 8297 11713 8309 11747
rect 8343 11744 8355 11747
rect 8570 11744 8576 11756
rect 8343 11716 8576 11744
rect 8343 11713 8355 11716
rect 8297 11707 8355 11713
rect 8570 11704 8576 11716
rect 8628 11704 8634 11756
rect 7469 11679 7527 11685
rect 7469 11676 7481 11679
rect 7432 11648 7481 11676
rect 7432 11636 7438 11648
rect 7469 11645 7481 11648
rect 7515 11645 7527 11679
rect 7469 11639 7527 11645
rect 7650 11636 7656 11688
rect 7708 11676 7714 11688
rect 9692 11685 9720 11784
rect 11238 11772 11244 11784
rect 11296 11772 11302 11824
rect 11330 11772 11336 11824
rect 11388 11812 11394 11824
rect 15562 11812 15568 11824
rect 11388 11784 15568 11812
rect 11388 11772 11394 11784
rect 15562 11772 15568 11784
rect 15620 11772 15626 11824
rect 17218 11812 17224 11824
rect 15948 11784 17224 11812
rect 10042 11704 10048 11756
rect 10100 11744 10106 11756
rect 10689 11747 10747 11753
rect 10689 11744 10701 11747
rect 10100 11716 10701 11744
rect 10100 11704 10106 11716
rect 10689 11713 10701 11716
rect 10735 11713 10747 11747
rect 10689 11707 10747 11713
rect 13354 11704 13360 11756
rect 13412 11744 13418 11756
rect 13541 11747 13599 11753
rect 13541 11744 13553 11747
rect 13412 11716 13553 11744
rect 13412 11704 13418 11716
rect 13541 11713 13553 11716
rect 13587 11713 13599 11747
rect 13541 11707 13599 11713
rect 14182 11704 14188 11756
rect 14240 11744 14246 11756
rect 15948 11744 15976 11784
rect 17218 11772 17224 11784
rect 17276 11772 17282 11824
rect 18046 11772 18052 11824
rect 18104 11812 18110 11824
rect 21174 11812 21180 11824
rect 18104 11784 20300 11812
rect 21135 11784 21180 11812
rect 18104 11772 18110 11784
rect 14240 11716 15976 11744
rect 16025 11747 16083 11753
rect 14240 11704 14246 11716
rect 16025 11713 16037 11747
rect 16071 11744 16083 11747
rect 16114 11744 16120 11756
rect 16071 11716 16120 11744
rect 16071 11713 16083 11716
rect 16025 11707 16083 11713
rect 16114 11704 16120 11716
rect 16172 11704 16178 11756
rect 18322 11744 18328 11756
rect 18283 11716 18328 11744
rect 18322 11704 18328 11716
rect 18380 11704 18386 11756
rect 20272 11753 20300 11784
rect 21174 11772 21180 11784
rect 21232 11812 21238 11824
rect 21232 11784 21864 11812
rect 21232 11772 21238 11784
rect 20257 11747 20315 11753
rect 20257 11713 20269 11747
rect 20303 11744 20315 11747
rect 20346 11744 20352 11756
rect 20303 11716 20352 11744
rect 20303 11713 20315 11716
rect 20257 11707 20315 11713
rect 20346 11704 20352 11716
rect 20404 11704 20410 11756
rect 20901 11747 20959 11753
rect 20901 11713 20913 11747
rect 20947 11744 20959 11747
rect 21266 11744 21272 11756
rect 20947 11716 21272 11744
rect 20947 11713 20959 11716
rect 20901 11707 20959 11713
rect 21266 11704 21272 11716
rect 21324 11704 21330 11756
rect 21450 11704 21456 11756
rect 21508 11744 21514 11756
rect 21545 11747 21603 11753
rect 21545 11744 21557 11747
rect 21508 11716 21557 11744
rect 21508 11704 21514 11716
rect 21545 11713 21557 11716
rect 21591 11744 21603 11747
rect 21591 11716 21772 11744
rect 21591 11713 21603 11716
rect 21545 11707 21603 11713
rect 9125 11679 9183 11685
rect 9125 11676 9137 11679
rect 7708 11648 9137 11676
rect 7708 11636 7714 11648
rect 9125 11645 9137 11648
rect 9171 11676 9183 11679
rect 9677 11679 9735 11685
rect 9677 11676 9689 11679
rect 9171 11648 9689 11676
rect 9171 11645 9183 11648
rect 9125 11639 9183 11645
rect 9677 11645 9689 11648
rect 9723 11645 9735 11679
rect 9677 11639 9735 11645
rect 9950 11636 9956 11688
rect 10008 11676 10014 11688
rect 10229 11679 10287 11685
rect 10229 11676 10241 11679
rect 10008 11648 10241 11676
rect 10008 11636 10014 11648
rect 10229 11645 10241 11648
rect 10275 11645 10287 11679
rect 10229 11639 10287 11645
rect 10318 11636 10324 11688
rect 10376 11676 10382 11688
rect 10505 11679 10563 11685
rect 10376 11648 10421 11676
rect 10376 11636 10382 11648
rect 10505 11645 10517 11679
rect 10551 11676 10563 11679
rect 10778 11676 10784 11688
rect 10551 11648 10784 11676
rect 10551 11645 10563 11648
rect 10505 11639 10563 11645
rect 10778 11636 10784 11648
rect 10836 11636 10842 11688
rect 12437 11679 12495 11685
rect 12437 11645 12449 11679
rect 12483 11645 12495 11679
rect 15013 11679 15071 11685
rect 15013 11676 15025 11679
rect 12437 11639 12495 11645
rect 14384 11648 15025 11676
rect 4890 11608 4896 11620
rect 4488 11580 4896 11608
rect 4488 11568 4494 11580
rect 4890 11568 4896 11580
rect 4948 11608 4954 11620
rect 6178 11608 6184 11620
rect 4948 11580 6040 11608
rect 6091 11580 6184 11608
rect 4948 11568 4954 11580
rect 2222 11540 2228 11552
rect 2183 11512 2228 11540
rect 2222 11500 2228 11512
rect 2280 11500 2286 11552
rect 4062 11540 4068 11552
rect 4023 11512 4068 11540
rect 4062 11500 4068 11512
rect 4120 11500 4126 11552
rect 6012 11540 6040 11580
rect 6178 11568 6184 11580
rect 6236 11608 6242 11620
rect 8294 11608 8300 11620
rect 6236 11580 8300 11608
rect 6236 11568 6242 11580
rect 8294 11568 8300 11580
rect 8352 11568 8358 11620
rect 8478 11568 8484 11620
rect 8536 11608 8542 11620
rect 12452 11608 12480 11639
rect 12897 11611 12955 11617
rect 12897 11608 12909 11611
rect 8536 11580 12909 11608
rect 8536 11568 8542 11580
rect 12897 11577 12909 11580
rect 12943 11577 12955 11611
rect 12897 11571 12955 11577
rect 13630 11568 13636 11620
rect 13688 11608 13694 11620
rect 14185 11611 14243 11617
rect 13688 11580 13733 11608
rect 13688 11568 13694 11580
rect 14185 11577 14197 11611
rect 14231 11608 14243 11611
rect 14274 11608 14280 11620
rect 14231 11580 14280 11608
rect 14231 11577 14243 11580
rect 14185 11571 14243 11577
rect 14274 11568 14280 11580
rect 14332 11568 14338 11620
rect 6549 11543 6607 11549
rect 6549 11540 6561 11543
rect 6012 11512 6561 11540
rect 6549 11509 6561 11512
rect 6595 11540 6607 11543
rect 6917 11543 6975 11549
rect 6917 11540 6929 11543
rect 6595 11512 6929 11540
rect 6595 11509 6607 11512
rect 6549 11503 6607 11509
rect 6917 11509 6929 11512
rect 6963 11509 6975 11543
rect 6917 11503 6975 11509
rect 10137 11543 10195 11549
rect 10137 11509 10149 11543
rect 10183 11540 10195 11543
rect 10778 11540 10784 11552
rect 10183 11512 10784 11540
rect 10183 11509 10195 11512
rect 10137 11503 10195 11509
rect 10778 11500 10784 11512
rect 10836 11500 10842 11552
rect 11882 11540 11888 11552
rect 11795 11512 11888 11540
rect 11882 11500 11888 11512
rect 11940 11540 11946 11552
rect 12621 11543 12679 11549
rect 12621 11540 12633 11543
rect 11940 11512 12633 11540
rect 11940 11500 11946 11512
rect 12621 11509 12633 11512
rect 12667 11540 12679 11543
rect 12802 11540 12808 11552
rect 12667 11512 12808 11540
rect 12667 11509 12679 11512
rect 12621 11503 12679 11509
rect 12802 11500 12808 11512
rect 12860 11500 12866 11552
rect 13262 11540 13268 11552
rect 13223 11512 13268 11540
rect 13262 11500 13268 11512
rect 13320 11500 13326 11552
rect 13354 11500 13360 11552
rect 13412 11540 13418 11552
rect 14384 11540 14412 11648
rect 15013 11645 15025 11648
rect 15059 11676 15071 11679
rect 15473 11679 15531 11685
rect 15473 11676 15485 11679
rect 15059 11648 15485 11676
rect 15059 11645 15071 11648
rect 15013 11639 15071 11645
rect 15473 11645 15485 11648
rect 15519 11645 15531 11679
rect 17678 11676 17684 11688
rect 17591 11648 17684 11676
rect 15473 11639 15531 11645
rect 17678 11636 17684 11648
rect 17736 11676 17742 11688
rect 18782 11676 18788 11688
rect 17736 11648 18788 11676
rect 17736 11636 17742 11648
rect 18782 11636 18788 11648
rect 18840 11676 18846 11688
rect 20070 11676 20076 11688
rect 18840 11648 20076 11676
rect 18840 11636 18846 11648
rect 20070 11636 20076 11648
rect 20128 11636 20134 11688
rect 21744 11685 21772 11716
rect 21729 11679 21787 11685
rect 21729 11645 21741 11679
rect 21775 11645 21787 11679
rect 21836 11676 21864 11784
rect 22189 11679 22247 11685
rect 22189 11676 22201 11679
rect 21836 11648 22201 11676
rect 21729 11639 21787 11645
rect 22189 11645 22201 11648
rect 22235 11645 22247 11679
rect 22189 11639 22247 11645
rect 14921 11611 14979 11617
rect 14921 11577 14933 11611
rect 14967 11608 14979 11611
rect 15654 11608 15660 11620
rect 14967 11580 15660 11608
rect 14967 11577 14979 11580
rect 14921 11571 14979 11577
rect 15654 11568 15660 11580
rect 15712 11568 15718 11620
rect 16346 11611 16404 11617
rect 16346 11577 16358 11611
rect 16392 11577 16404 11611
rect 16346 11571 16404 11577
rect 20349 11611 20407 11617
rect 20349 11577 20361 11611
rect 20395 11608 20407 11611
rect 21082 11608 21088 11620
rect 20395 11580 21088 11608
rect 20395 11577 20407 11580
rect 20349 11571 20407 11577
rect 15930 11540 15936 11552
rect 13412 11512 14412 11540
rect 15891 11512 15936 11540
rect 13412 11500 13418 11512
rect 15930 11500 15936 11512
rect 15988 11540 15994 11552
rect 16361 11540 16389 11571
rect 15988 11512 16389 11540
rect 15988 11500 15994 11512
rect 16482 11500 16488 11552
rect 16540 11540 16546 11552
rect 16945 11543 17003 11549
rect 16945 11540 16957 11543
rect 16540 11512 16957 11540
rect 16540 11500 16546 11512
rect 16945 11509 16957 11512
rect 16991 11509 17003 11543
rect 18690 11540 18696 11552
rect 18651 11512 18696 11540
rect 16945 11503 17003 11509
rect 18690 11500 18696 11512
rect 18748 11500 18754 11552
rect 19245 11543 19303 11549
rect 19245 11509 19257 11543
rect 19291 11540 19303 11543
rect 19426 11540 19432 11552
rect 19291 11512 19432 11540
rect 19291 11509 19303 11512
rect 19245 11503 19303 11509
rect 19426 11500 19432 11512
rect 19484 11540 19490 11552
rect 19613 11543 19671 11549
rect 19613 11540 19625 11543
rect 19484 11512 19625 11540
rect 19484 11500 19490 11512
rect 19613 11509 19625 11512
rect 19659 11540 19671 11543
rect 20073 11543 20131 11549
rect 20073 11540 20085 11543
rect 19659 11512 20085 11540
rect 19659 11509 19671 11512
rect 19613 11503 19671 11509
rect 20073 11509 20085 11512
rect 20119 11540 20131 11543
rect 20364 11540 20392 11571
rect 21082 11568 21088 11580
rect 21140 11568 21146 11620
rect 21818 11540 21824 11552
rect 20119 11512 20392 11540
rect 21779 11512 21824 11540
rect 20119 11509 20131 11512
rect 20073 11503 20131 11509
rect 21818 11500 21824 11512
rect 21876 11500 21882 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1854 11336 1860 11348
rect 1815 11308 1860 11336
rect 1854 11296 1860 11308
rect 1912 11336 1918 11348
rect 3050 11336 3056 11348
rect 1912 11308 2268 11336
rect 3011 11308 3056 11336
rect 1912 11296 1918 11308
rect 1946 11228 1952 11280
rect 2004 11268 2010 11280
rect 2240 11277 2268 11308
rect 3050 11296 3056 11308
rect 3108 11296 3114 11348
rect 3881 11339 3939 11345
rect 3881 11305 3893 11339
rect 3927 11336 3939 11339
rect 3970 11336 3976 11348
rect 3927 11308 3976 11336
rect 3927 11305 3939 11308
rect 3881 11299 3939 11305
rect 3970 11296 3976 11308
rect 4028 11296 4034 11348
rect 5442 11336 5448 11348
rect 5403 11308 5448 11336
rect 5442 11296 5448 11308
rect 5500 11296 5506 11348
rect 6641 11339 6699 11345
rect 6641 11305 6653 11339
rect 6687 11336 6699 11339
rect 6822 11336 6828 11348
rect 6687 11308 6828 11336
rect 6687 11305 6699 11308
rect 6641 11299 6699 11305
rect 6822 11296 6828 11308
rect 6880 11336 6886 11348
rect 6917 11339 6975 11345
rect 6917 11336 6929 11339
rect 6880 11308 6929 11336
rect 6880 11296 6886 11308
rect 6917 11305 6929 11308
rect 6963 11305 6975 11339
rect 6917 11299 6975 11305
rect 2133 11271 2191 11277
rect 2133 11268 2145 11271
rect 2004 11240 2145 11268
rect 2004 11228 2010 11240
rect 2133 11237 2145 11240
rect 2179 11237 2191 11271
rect 2133 11231 2191 11237
rect 2225 11271 2283 11277
rect 2225 11237 2237 11271
rect 2271 11268 2283 11271
rect 2774 11268 2780 11280
rect 2271 11240 2780 11268
rect 2271 11237 2283 11240
rect 2225 11231 2283 11237
rect 2774 11228 2780 11240
rect 2832 11228 2838 11280
rect 3988 11268 4016 11296
rect 5813 11271 5871 11277
rect 5813 11268 5825 11271
rect 3988 11240 4200 11268
rect 4172 11209 4200 11240
rect 4540 11240 5825 11268
rect 4540 11212 4568 11240
rect 5813 11237 5825 11240
rect 5859 11237 5871 11271
rect 6932 11268 6960 11299
rect 10134 11296 10140 11348
rect 10192 11336 10198 11348
rect 10229 11339 10287 11345
rect 10229 11336 10241 11339
rect 10192 11308 10241 11336
rect 10192 11296 10198 11308
rect 10229 11305 10241 11308
rect 10275 11305 10287 11339
rect 13538 11336 13544 11348
rect 13499 11308 13544 11336
rect 10229 11299 10287 11305
rect 13538 11296 13544 11308
rect 13596 11296 13602 11348
rect 14182 11336 14188 11348
rect 14143 11308 14188 11336
rect 14182 11296 14188 11308
rect 14240 11296 14246 11348
rect 15562 11336 15568 11348
rect 15523 11308 15568 11336
rect 15562 11296 15568 11308
rect 15620 11296 15626 11348
rect 16114 11336 16120 11348
rect 16075 11308 16120 11336
rect 16114 11296 16120 11308
rect 16172 11296 16178 11348
rect 18371 11339 18429 11345
rect 18371 11305 18383 11339
rect 18417 11336 18429 11339
rect 19978 11336 19984 11348
rect 18417 11308 19984 11336
rect 18417 11305 18429 11308
rect 18371 11299 18429 11305
rect 19978 11296 19984 11308
rect 20036 11296 20042 11348
rect 20346 11336 20352 11348
rect 20307 11308 20352 11336
rect 20346 11296 20352 11308
rect 20404 11296 20410 11348
rect 22649 11339 22707 11345
rect 22649 11336 22661 11339
rect 20548 11308 22661 11336
rect 12615 11271 12673 11277
rect 6932 11240 7604 11268
rect 5813 11231 5871 11237
rect 4157 11203 4215 11209
rect 4157 11169 4169 11203
rect 4203 11169 4215 11203
rect 4522 11200 4528 11212
rect 4483 11172 4528 11200
rect 4157 11163 4215 11169
rect 4522 11160 4528 11172
rect 4580 11160 4586 11212
rect 4890 11200 4896 11212
rect 4851 11172 4896 11200
rect 4890 11160 4896 11172
rect 4948 11160 4954 11212
rect 5445 11203 5503 11209
rect 5445 11169 5457 11203
rect 5491 11200 5503 11203
rect 6178 11200 6184 11212
rect 5491 11172 6184 11200
rect 5491 11169 5503 11172
rect 5445 11163 5503 11169
rect 6178 11160 6184 11172
rect 6236 11160 6242 11212
rect 7374 11200 7380 11212
rect 7335 11172 7380 11200
rect 7374 11160 7380 11172
rect 7432 11160 7438 11212
rect 7576 11209 7604 11240
rect 12615 11237 12627 11271
rect 12661 11268 12673 11271
rect 12710 11268 12716 11280
rect 12661 11240 12716 11268
rect 12661 11237 12673 11240
rect 12615 11231 12673 11237
rect 12710 11228 12716 11240
rect 12768 11228 12774 11280
rect 15470 11228 15476 11280
rect 15528 11268 15534 11280
rect 16298 11268 16304 11280
rect 15528 11240 16304 11268
rect 15528 11228 15534 11240
rect 16298 11228 16304 11240
rect 16356 11228 16362 11280
rect 16393 11271 16451 11277
rect 16393 11237 16405 11271
rect 16439 11268 16451 11271
rect 16482 11268 16488 11280
rect 16439 11240 16488 11268
rect 16439 11237 16451 11240
rect 16393 11231 16451 11237
rect 16482 11228 16488 11240
rect 16540 11268 16546 11280
rect 18969 11271 19027 11277
rect 18969 11268 18981 11271
rect 16540 11240 18981 11268
rect 16540 11228 16546 11240
rect 18969 11237 18981 11240
rect 19015 11237 19027 11271
rect 19150 11268 19156 11280
rect 19111 11240 19156 11268
rect 18969 11231 19027 11237
rect 19150 11228 19156 11240
rect 19208 11228 19214 11280
rect 19429 11271 19487 11277
rect 19429 11237 19441 11271
rect 19475 11268 19487 11271
rect 19794 11268 19800 11280
rect 19475 11240 19800 11268
rect 19475 11237 19487 11240
rect 19429 11231 19487 11237
rect 19794 11228 19800 11240
rect 19852 11228 19858 11280
rect 20070 11228 20076 11280
rect 20128 11268 20134 11280
rect 20548 11268 20576 11308
rect 22649 11305 22661 11308
rect 22695 11305 22707 11339
rect 22649 11299 22707 11305
rect 21082 11268 21088 11280
rect 20128 11240 20576 11268
rect 21043 11240 21088 11268
rect 20128 11228 20134 11240
rect 21082 11228 21088 11240
rect 21140 11228 21146 11280
rect 7561 11203 7619 11209
rect 7561 11169 7573 11203
rect 7607 11200 7619 11203
rect 7650 11200 7656 11212
rect 7607 11172 7656 11200
rect 7607 11169 7619 11172
rect 7561 11163 7619 11169
rect 7650 11160 7656 11172
rect 7708 11160 7714 11212
rect 7929 11203 7987 11209
rect 7929 11169 7941 11203
rect 7975 11169 7987 11203
rect 7929 11163 7987 11169
rect 1578 11092 1584 11144
rect 1636 11132 1642 11144
rect 2314 11132 2320 11144
rect 1636 11104 2320 11132
rect 1636 11092 1642 11104
rect 2314 11092 2320 11104
rect 2372 11132 2378 11144
rect 2409 11135 2467 11141
rect 2409 11132 2421 11135
rect 2372 11104 2421 11132
rect 2372 11092 2378 11104
rect 2409 11101 2421 11104
rect 2455 11101 2467 11135
rect 2409 11095 2467 11101
rect 3418 11092 3424 11144
rect 3476 11132 3482 11144
rect 3513 11135 3571 11141
rect 3513 11132 3525 11135
rect 3476 11104 3525 11132
rect 3476 11092 3482 11104
rect 3513 11101 3525 11104
rect 3559 11101 3571 11135
rect 3513 11095 3571 11101
rect 6273 10999 6331 11005
rect 6273 10965 6285 10999
rect 6319 10996 6331 10999
rect 7944 10996 7972 11163
rect 8294 11160 8300 11212
rect 8352 11200 8358 11212
rect 8481 11203 8539 11209
rect 8481 11200 8493 11203
rect 8352 11172 8493 11200
rect 8352 11160 8358 11172
rect 8481 11169 8493 11172
rect 8527 11200 8539 11203
rect 8849 11203 8907 11209
rect 8849 11200 8861 11203
rect 8527 11172 8861 11200
rect 8527 11169 8539 11172
rect 8481 11163 8539 11169
rect 8849 11169 8861 11172
rect 8895 11169 8907 11203
rect 8849 11163 8907 11169
rect 9582 11160 9588 11212
rect 9640 11200 9646 11212
rect 9677 11203 9735 11209
rect 9677 11200 9689 11203
rect 9640 11172 9689 11200
rect 9640 11160 9646 11172
rect 9677 11169 9689 11172
rect 9723 11169 9735 11203
rect 11330 11200 11336 11212
rect 11291 11172 11336 11200
rect 9677 11163 9735 11169
rect 11330 11160 11336 11172
rect 11388 11200 11394 11212
rect 13173 11203 13231 11209
rect 13173 11200 13185 11203
rect 11388 11172 13185 11200
rect 11388 11160 11394 11172
rect 13173 11169 13185 11172
rect 13219 11200 13231 11203
rect 13262 11200 13268 11212
rect 13219 11172 13268 11200
rect 13219 11169 13231 11172
rect 13173 11163 13231 11169
rect 13262 11160 13268 11172
rect 13320 11200 13326 11212
rect 13630 11200 13636 11212
rect 13320 11172 13636 11200
rect 13320 11160 13326 11172
rect 13630 11160 13636 11172
rect 13688 11160 13694 11212
rect 13998 11200 14004 11212
rect 13959 11172 14004 11200
rect 13998 11160 14004 11172
rect 14056 11160 14062 11212
rect 17954 11160 17960 11212
rect 18012 11200 18018 11212
rect 18690 11200 18696 11212
rect 18012 11172 18696 11200
rect 18012 11160 18018 11172
rect 18690 11160 18696 11172
rect 18748 11160 18754 11212
rect 22465 11203 22523 11209
rect 22465 11169 22477 11203
rect 22511 11200 22523 11203
rect 22738 11200 22744 11212
rect 22511 11172 22744 11200
rect 22511 11169 22523 11172
rect 22465 11163 22523 11169
rect 22738 11160 22744 11172
rect 22796 11160 22802 11212
rect 8573 11135 8631 11141
rect 8573 11101 8585 11135
rect 8619 11132 8631 11135
rect 11790 11132 11796 11144
rect 8619 11104 11796 11132
rect 8619 11101 8631 11104
rect 8573 11095 8631 11101
rect 11790 11092 11796 11104
rect 11848 11132 11854 11144
rect 12253 11135 12311 11141
rect 12253 11132 12265 11135
rect 11848 11104 12265 11132
rect 11848 11092 11854 11104
rect 12253 11101 12265 11104
rect 12299 11101 12311 11135
rect 12253 11095 12311 11101
rect 19337 11135 19395 11141
rect 19337 11101 19349 11135
rect 19383 11132 19395 11135
rect 19426 11132 19432 11144
rect 19383 11104 19432 11132
rect 19383 11101 19395 11104
rect 19337 11095 19395 11101
rect 19426 11092 19432 11104
rect 19484 11092 19490 11144
rect 20993 11135 21051 11141
rect 20993 11101 21005 11135
rect 21039 11132 21051 11135
rect 21726 11132 21732 11144
rect 21039 11104 21732 11132
rect 21039 11101 21051 11104
rect 20993 11095 21051 11101
rect 21726 11092 21732 11104
rect 21784 11092 21790 11144
rect 9861 11067 9919 11073
rect 9861 11033 9873 11067
rect 9907 11064 9919 11067
rect 11149 11067 11207 11073
rect 9907 11036 10542 11064
rect 9907 11033 9919 11036
rect 9861 11027 9919 11033
rect 8202 10996 8208 11008
rect 6319 10968 8208 10996
rect 6319 10965 6331 10968
rect 6273 10959 6331 10965
rect 8202 10956 8208 10968
rect 8260 10956 8266 11008
rect 10514 10996 10542 11036
rect 11149 11033 11161 11067
rect 11195 11064 11207 11067
rect 13722 11064 13728 11076
rect 11195 11036 13728 11064
rect 11195 11033 11207 11036
rect 11149 11027 11207 11033
rect 13722 11024 13728 11036
rect 13780 11024 13786 11076
rect 16666 11024 16672 11076
rect 16724 11064 16730 11076
rect 16853 11067 16911 11073
rect 16853 11064 16865 11067
rect 16724 11036 16865 11064
rect 16724 11024 16730 11036
rect 16853 11033 16865 11036
rect 16899 11064 16911 11067
rect 19889 11067 19947 11073
rect 19889 11064 19901 11067
rect 16899 11036 19901 11064
rect 16899 11033 16911 11036
rect 16853 11027 16911 11033
rect 19889 11033 19901 11036
rect 19935 11064 19947 11067
rect 21545 11067 21603 11073
rect 21545 11064 21557 11067
rect 19935 11036 21557 11064
rect 19935 11033 19947 11036
rect 19889 11027 19947 11033
rect 21545 11033 21557 11036
rect 21591 11033 21603 11067
rect 21545 11027 21603 11033
rect 12618 10996 12624 11008
rect 10514 10968 12624 10996
rect 12618 10956 12624 10968
rect 12676 10956 12682 11008
rect 13446 10956 13452 11008
rect 13504 10996 13510 11008
rect 13817 10999 13875 11005
rect 13817 10996 13829 10999
rect 13504 10968 13829 10996
rect 13504 10956 13510 10968
rect 13817 10965 13829 10968
rect 13863 10965 13875 10999
rect 18138 10996 18144 11008
rect 18099 10968 18144 10996
rect 13817 10959 13875 10965
rect 18138 10956 18144 10968
rect 18196 10956 18202 11008
rect 18969 10999 19027 11005
rect 18969 10965 18981 10999
rect 19015 10996 19027 10999
rect 20625 10999 20683 11005
rect 20625 10996 20637 10999
rect 19015 10968 20637 10996
rect 19015 10965 19027 10968
rect 18969 10959 19027 10965
rect 20625 10965 20637 10968
rect 20671 10996 20683 10999
rect 20990 10996 20996 11008
rect 20671 10968 20996 10996
rect 20671 10965 20683 10968
rect 20625 10959 20683 10965
rect 20990 10956 20996 10968
rect 21048 10956 21054 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 14 10752 20 10804
rect 72 10792 78 10804
rect 3145 10795 3203 10801
rect 72 10764 3096 10792
rect 72 10752 78 10764
rect 2038 10684 2044 10736
rect 2096 10724 2102 10736
rect 3068 10724 3096 10764
rect 3145 10761 3157 10795
rect 3191 10792 3203 10795
rect 3234 10792 3240 10804
rect 3191 10764 3240 10792
rect 3191 10761 3203 10764
rect 3145 10755 3203 10761
rect 3234 10752 3240 10764
rect 3292 10752 3298 10804
rect 4982 10792 4988 10804
rect 4943 10764 4988 10792
rect 4982 10752 4988 10764
rect 5040 10752 5046 10804
rect 6641 10795 6699 10801
rect 6641 10761 6653 10795
rect 6687 10792 6699 10795
rect 7009 10795 7067 10801
rect 7009 10792 7021 10795
rect 6687 10764 7021 10792
rect 6687 10761 6699 10764
rect 6641 10755 6699 10761
rect 7009 10761 7021 10764
rect 7055 10792 7067 10795
rect 7374 10792 7380 10804
rect 7055 10764 7380 10792
rect 7055 10761 7067 10764
rect 7009 10755 7067 10761
rect 7374 10752 7380 10764
rect 7432 10752 7438 10804
rect 11330 10792 11336 10804
rect 11291 10764 11336 10792
rect 11330 10752 11336 10764
rect 11388 10752 11394 10804
rect 11790 10792 11796 10804
rect 11751 10764 11796 10792
rect 11790 10752 11796 10764
rect 11848 10752 11854 10804
rect 12253 10795 12311 10801
rect 12253 10761 12265 10795
rect 12299 10792 12311 10795
rect 12710 10792 12716 10804
rect 12299 10764 12716 10792
rect 12299 10761 12311 10764
rect 12253 10755 12311 10761
rect 12710 10752 12716 10764
rect 12768 10752 12774 10804
rect 13998 10792 14004 10804
rect 13786 10764 14004 10792
rect 3421 10727 3479 10733
rect 3421 10724 3433 10727
rect 2096 10696 2452 10724
rect 3068 10696 3433 10724
rect 2096 10684 2102 10696
rect 2130 10656 2136 10668
rect 2091 10628 2136 10656
rect 2130 10616 2136 10628
rect 2188 10616 2194 10668
rect 2424 10665 2452 10696
rect 3421 10693 3433 10696
rect 3467 10693 3479 10727
rect 5000 10724 5028 10752
rect 5261 10727 5319 10733
rect 5261 10724 5273 10727
rect 5000 10696 5273 10724
rect 3421 10687 3479 10693
rect 5261 10693 5273 10696
rect 5307 10693 5319 10727
rect 5261 10687 5319 10693
rect 2409 10659 2467 10665
rect 2409 10625 2421 10659
rect 2455 10625 2467 10659
rect 2409 10619 2467 10625
rect 3436 10588 3464 10687
rect 5350 10684 5356 10736
rect 5408 10724 5414 10736
rect 9125 10727 9183 10733
rect 5408 10696 8616 10724
rect 5408 10684 5414 10696
rect 3878 10616 3884 10668
rect 3936 10656 3942 10668
rect 4617 10659 4675 10665
rect 4617 10656 4629 10659
rect 3936 10628 4629 10656
rect 3936 10616 3942 10628
rect 4617 10625 4629 10628
rect 4663 10656 4675 10659
rect 5905 10659 5963 10665
rect 4663 10628 5488 10656
rect 4663 10625 4675 10628
rect 4617 10619 4675 10625
rect 3697 10591 3755 10597
rect 3697 10588 3709 10591
rect 3436 10560 3709 10588
rect 3697 10557 3709 10560
rect 3743 10588 3755 10591
rect 5166 10588 5172 10600
rect 3743 10560 4154 10588
rect 5127 10560 5172 10588
rect 3743 10557 3755 10560
rect 3697 10551 3755 10557
rect 2225 10523 2283 10529
rect 2225 10489 2237 10523
rect 2271 10489 2283 10523
rect 4126 10520 4154 10560
rect 5166 10548 5172 10560
rect 5224 10548 5230 10600
rect 5460 10597 5488 10628
rect 5905 10625 5917 10659
rect 5951 10656 5963 10659
rect 8478 10656 8484 10668
rect 5951 10628 8484 10656
rect 5951 10625 5963 10628
rect 5905 10619 5963 10625
rect 8478 10616 8484 10628
rect 8536 10616 8542 10668
rect 5445 10591 5503 10597
rect 5445 10557 5457 10591
rect 5491 10557 5503 10591
rect 7374 10588 7380 10600
rect 7335 10560 7380 10588
rect 5445 10551 5503 10557
rect 7374 10548 7380 10560
rect 7432 10548 7438 10600
rect 7650 10588 7656 10600
rect 7611 10560 7656 10588
rect 7650 10548 7656 10560
rect 7708 10548 7714 10600
rect 8202 10588 8208 10600
rect 8163 10560 8208 10588
rect 8202 10548 8208 10560
rect 8260 10548 8266 10600
rect 8588 10597 8616 10696
rect 9125 10693 9137 10727
rect 9171 10724 9183 10727
rect 9582 10724 9588 10736
rect 9171 10696 9588 10724
rect 9171 10693 9183 10696
rect 9125 10687 9183 10693
rect 9582 10684 9588 10696
rect 9640 10724 9646 10736
rect 13078 10724 13084 10736
rect 9640 10696 13084 10724
rect 9640 10684 9646 10696
rect 13078 10684 13084 10696
rect 13136 10684 13142 10736
rect 8665 10659 8723 10665
rect 8665 10625 8677 10659
rect 8711 10656 8723 10659
rect 12805 10659 12863 10665
rect 12805 10656 12817 10659
rect 8711 10628 12817 10656
rect 8711 10625 8723 10628
rect 8665 10619 8723 10625
rect 12805 10625 12817 10628
rect 12851 10656 12863 10659
rect 12894 10656 12900 10668
rect 12851 10628 12900 10656
rect 12851 10625 12863 10628
rect 12805 10619 12863 10625
rect 12894 10616 12900 10628
rect 12952 10616 12958 10668
rect 12986 10616 12992 10668
rect 13044 10656 13050 10668
rect 13786 10656 13814 10764
rect 13998 10752 14004 10764
rect 14056 10752 14062 10804
rect 14737 10795 14795 10801
rect 14737 10761 14749 10795
rect 14783 10792 14795 10795
rect 16022 10792 16028 10804
rect 14783 10764 16028 10792
rect 14783 10761 14795 10764
rect 14737 10755 14795 10761
rect 16022 10752 16028 10764
rect 16080 10752 16086 10804
rect 16298 10752 16304 10804
rect 16356 10792 16362 10804
rect 17129 10795 17187 10801
rect 17129 10792 17141 10795
rect 16356 10764 17141 10792
rect 16356 10752 16362 10764
rect 17129 10761 17141 10764
rect 17175 10761 17187 10795
rect 17129 10755 17187 10761
rect 19334 10752 19340 10804
rect 19392 10792 19398 10804
rect 19794 10792 19800 10804
rect 19392 10764 19800 10792
rect 19392 10752 19398 10764
rect 19794 10752 19800 10764
rect 19852 10752 19858 10804
rect 21082 10752 21088 10804
rect 21140 10792 21146 10804
rect 21361 10795 21419 10801
rect 21361 10792 21373 10795
rect 21140 10764 21373 10792
rect 21140 10752 21146 10764
rect 21361 10761 21373 10764
rect 21407 10761 21419 10795
rect 21726 10792 21732 10804
rect 21687 10764 21732 10792
rect 21361 10755 21419 10761
rect 21726 10752 21732 10764
rect 21784 10792 21790 10804
rect 22051 10795 22109 10801
rect 22051 10792 22063 10795
rect 21784 10764 22063 10792
rect 21784 10752 21790 10764
rect 22051 10761 22063 10764
rect 22097 10761 22109 10795
rect 22051 10755 22109 10761
rect 13044 10628 13814 10656
rect 15473 10659 15531 10665
rect 13044 10616 13050 10628
rect 15473 10625 15485 10659
rect 15519 10656 15531 10659
rect 15838 10656 15844 10668
rect 15519 10628 15844 10656
rect 15519 10625 15531 10628
rect 15473 10619 15531 10625
rect 15838 10616 15844 10628
rect 15896 10656 15902 10668
rect 15933 10659 15991 10665
rect 15933 10656 15945 10659
rect 15896 10628 15945 10656
rect 15896 10616 15902 10628
rect 15933 10625 15945 10628
rect 15979 10625 15991 10659
rect 15933 10619 15991 10625
rect 17865 10659 17923 10665
rect 17865 10625 17877 10659
rect 17911 10656 17923 10659
rect 18598 10656 18604 10668
rect 17911 10628 18604 10656
rect 17911 10625 17923 10628
rect 17865 10619 17923 10625
rect 18598 10616 18604 10628
rect 18656 10616 18662 10668
rect 20438 10656 20444 10668
rect 20351 10628 20444 10656
rect 20438 10616 20444 10628
rect 20496 10656 20502 10668
rect 21266 10656 21272 10668
rect 20496 10628 21272 10656
rect 20496 10616 20502 10628
rect 21266 10616 21272 10628
rect 21324 10616 21330 10668
rect 22465 10659 22523 10665
rect 22465 10625 22477 10659
rect 22511 10656 22523 10659
rect 27614 10656 27620 10668
rect 22511 10628 27620 10656
rect 22511 10625 22523 10628
rect 22465 10619 22523 10625
rect 8573 10591 8631 10597
rect 8573 10557 8585 10591
rect 8619 10588 8631 10591
rect 8754 10588 8760 10600
rect 8619 10560 8760 10588
rect 8619 10557 8631 10560
rect 8573 10551 8631 10557
rect 8754 10548 8760 10560
rect 8812 10548 8818 10600
rect 9306 10548 9312 10600
rect 9364 10588 9370 10600
rect 9953 10591 10011 10597
rect 9953 10588 9965 10591
rect 9364 10560 9965 10588
rect 9364 10548 9370 10560
rect 9953 10557 9965 10560
rect 9999 10557 10011 10591
rect 9953 10551 10011 10557
rect 10045 10591 10103 10597
rect 10045 10557 10057 10591
rect 10091 10588 10103 10591
rect 10134 10588 10140 10600
rect 10091 10560 10140 10588
rect 10091 10557 10103 10560
rect 10045 10551 10103 10557
rect 9861 10523 9919 10529
rect 9861 10520 9873 10523
rect 4126 10492 9873 10520
rect 2225 10483 2283 10489
rect 9861 10489 9873 10492
rect 9907 10520 9919 10523
rect 10060 10520 10088 10551
rect 10134 10548 10140 10560
rect 10192 10548 10198 10600
rect 10229 10591 10287 10597
rect 10229 10557 10241 10591
rect 10275 10588 10287 10591
rect 14550 10588 14556 10600
rect 10275 10560 11100 10588
rect 14511 10560 14556 10588
rect 10275 10557 10287 10560
rect 10229 10551 10287 10557
rect 10686 10520 10692 10532
rect 9907 10492 10088 10520
rect 10647 10492 10692 10520
rect 9907 10489 9919 10492
rect 9861 10483 9919 10489
rect 1946 10452 1952 10464
rect 1907 10424 1952 10452
rect 1946 10412 1952 10424
rect 2004 10452 2010 10464
rect 2240 10452 2268 10483
rect 10686 10480 10692 10492
rect 10744 10480 10750 10532
rect 4062 10452 4068 10464
rect 2004 10424 2268 10452
rect 4023 10424 4068 10452
rect 2004 10412 2010 10424
rect 4062 10412 4068 10424
rect 4120 10412 4126 10464
rect 5166 10412 5172 10464
rect 5224 10452 5230 10464
rect 6181 10455 6239 10461
rect 6181 10452 6193 10455
rect 5224 10424 6193 10452
rect 5224 10412 5230 10424
rect 6181 10421 6193 10424
rect 6227 10452 6239 10455
rect 6546 10452 6552 10464
rect 6227 10424 6552 10452
rect 6227 10421 6239 10424
rect 6181 10415 6239 10421
rect 6546 10412 6552 10424
rect 6604 10412 6610 10464
rect 9306 10412 9312 10464
rect 9364 10452 9370 10464
rect 11072 10461 11100 10560
rect 14550 10548 14556 10560
rect 14608 10588 14614 10600
rect 15013 10591 15071 10597
rect 15013 10588 15025 10591
rect 14608 10560 15025 10588
rect 14608 10548 14614 10560
rect 15013 10557 15025 10560
rect 15059 10557 15071 10591
rect 15013 10551 15071 10557
rect 19521 10591 19579 10597
rect 19521 10557 19533 10591
rect 19567 10588 19579 10591
rect 20165 10591 20223 10597
rect 20165 10588 20177 10591
rect 19567 10560 20177 10588
rect 19567 10557 19579 10560
rect 19521 10551 19579 10557
rect 20165 10557 20177 10560
rect 20211 10557 20223 10591
rect 20165 10551 20223 10557
rect 12710 10480 12716 10532
rect 12768 10520 12774 10532
rect 13126 10523 13184 10529
rect 13126 10520 13138 10523
rect 12768 10492 13138 10520
rect 12768 10480 12774 10492
rect 13126 10489 13138 10492
rect 13172 10520 13184 10523
rect 13998 10520 14004 10532
rect 13172 10492 14004 10520
rect 13172 10489 13184 10492
rect 13126 10483 13184 10489
rect 13998 10480 14004 10492
rect 14056 10520 14062 10532
rect 15749 10523 15807 10529
rect 15749 10520 15761 10523
rect 14056 10492 15761 10520
rect 14056 10480 14062 10492
rect 15749 10489 15761 10492
rect 15795 10520 15807 10523
rect 15930 10520 15936 10532
rect 15795 10492 15936 10520
rect 15795 10489 15807 10492
rect 15749 10483 15807 10489
rect 15930 10480 15936 10492
rect 15988 10520 15994 10532
rect 16254 10523 16312 10529
rect 16254 10520 16266 10523
rect 15988 10492 16266 10520
rect 15988 10480 15994 10492
rect 16254 10489 16266 10492
rect 16300 10520 16312 10523
rect 17954 10520 17960 10532
rect 16300 10492 17960 10520
rect 16300 10489 16312 10492
rect 16254 10483 16312 10489
rect 17954 10480 17960 10492
rect 18012 10520 18018 10532
rect 18922 10523 18980 10529
rect 18922 10520 18934 10523
rect 18012 10492 18934 10520
rect 18012 10480 18018 10492
rect 18922 10489 18934 10492
rect 18968 10489 18980 10523
rect 18922 10483 18980 10489
rect 9401 10455 9459 10461
rect 9401 10452 9413 10455
rect 9364 10424 9413 10452
rect 9364 10412 9370 10424
rect 9401 10421 9413 10424
rect 9447 10421 9459 10455
rect 9401 10415 9459 10421
rect 11057 10455 11115 10461
rect 11057 10421 11069 10455
rect 11103 10452 11115 10455
rect 11330 10452 11336 10464
rect 11103 10424 11336 10452
rect 11103 10421 11115 10424
rect 11057 10415 11115 10421
rect 11330 10412 11336 10424
rect 11388 10412 11394 10464
rect 13630 10412 13636 10464
rect 13688 10452 13694 10464
rect 13725 10455 13783 10461
rect 13725 10452 13737 10455
rect 13688 10424 13737 10452
rect 13688 10412 13694 10424
rect 13725 10421 13737 10424
rect 13771 10421 13783 10455
rect 16850 10452 16856 10464
rect 16811 10424 16856 10452
rect 13725 10415 13783 10421
rect 16850 10412 16856 10424
rect 16908 10412 16914 10464
rect 17402 10412 17408 10464
rect 17460 10452 17466 10464
rect 18138 10452 18144 10464
rect 17460 10424 18144 10452
rect 17460 10412 17466 10424
rect 18138 10412 18144 10424
rect 18196 10452 18202 10464
rect 18233 10455 18291 10461
rect 18233 10452 18245 10455
rect 18196 10424 18245 10452
rect 18196 10412 18202 10424
rect 18233 10421 18245 10424
rect 18279 10421 18291 10455
rect 20180 10452 20208 10551
rect 21634 10548 21640 10600
rect 21692 10588 21698 10600
rect 21980 10591 22038 10597
rect 21980 10588 21992 10591
rect 21692 10560 21992 10588
rect 21692 10548 21698 10560
rect 21980 10557 21992 10560
rect 22026 10588 22038 10591
rect 22480 10588 22508 10619
rect 27614 10616 27620 10628
rect 27672 10616 27678 10668
rect 22026 10560 22508 10588
rect 22026 10557 22038 10560
rect 21980 10551 22038 10557
rect 20533 10523 20591 10529
rect 20533 10489 20545 10523
rect 20579 10489 20591 10523
rect 20533 10483 20591 10489
rect 20548 10452 20576 10483
rect 20898 10480 20904 10532
rect 20956 10520 20962 10532
rect 21085 10523 21143 10529
rect 21085 10520 21097 10523
rect 20956 10492 21097 10520
rect 20956 10480 20962 10492
rect 21085 10489 21097 10492
rect 21131 10489 21143 10523
rect 21085 10483 21143 10489
rect 22738 10452 22744 10464
rect 20180 10424 20576 10452
rect 22699 10424 22744 10452
rect 18233 10415 18291 10421
rect 22738 10412 22744 10424
rect 22796 10412 22802 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 2774 10248 2780 10260
rect 2735 10220 2780 10248
rect 2774 10208 2780 10220
rect 2832 10208 2838 10260
rect 4157 10251 4215 10257
rect 4157 10248 4169 10251
rect 2884 10220 4169 10248
rect 2038 10140 2044 10192
rect 2096 10180 2102 10192
rect 2178 10183 2236 10189
rect 2178 10180 2190 10183
rect 2096 10152 2190 10180
rect 2096 10140 2102 10152
rect 2178 10149 2190 10152
rect 2224 10149 2236 10183
rect 2178 10143 2236 10149
rect 1854 10112 1860 10124
rect 1767 10084 1860 10112
rect 1854 10072 1860 10084
rect 1912 10112 1918 10124
rect 2884 10112 2912 10220
rect 4157 10217 4169 10220
rect 4203 10217 4215 10251
rect 4522 10248 4528 10260
rect 4157 10211 4215 10217
rect 4356 10220 4528 10248
rect 3145 10183 3203 10189
rect 3145 10149 3157 10183
rect 3191 10180 3203 10183
rect 4356 10180 4384 10220
rect 4522 10208 4528 10220
rect 4580 10248 4586 10260
rect 6825 10251 6883 10257
rect 4580 10220 4660 10248
rect 4580 10208 4586 10220
rect 3191 10152 4384 10180
rect 3191 10149 3203 10152
rect 3145 10143 3203 10149
rect 4632 10124 4660 10220
rect 6825 10217 6837 10251
rect 6871 10248 6883 10251
rect 6914 10248 6920 10260
rect 6871 10220 6920 10248
rect 6871 10217 6883 10220
rect 6825 10211 6883 10217
rect 6914 10208 6920 10220
rect 6972 10208 6978 10260
rect 8754 10248 8760 10260
rect 8715 10220 8760 10248
rect 8754 10208 8760 10220
rect 8812 10208 8818 10260
rect 12618 10248 12624 10260
rect 12579 10220 12624 10248
rect 12618 10208 12624 10220
rect 12676 10208 12682 10260
rect 12894 10248 12900 10260
rect 12855 10220 12900 10248
rect 12894 10208 12900 10220
rect 12952 10208 12958 10260
rect 15473 10251 15531 10257
rect 15473 10217 15485 10251
rect 15519 10248 15531 10251
rect 15746 10248 15752 10260
rect 15519 10220 15752 10248
rect 15519 10217 15531 10220
rect 15473 10211 15531 10217
rect 15746 10208 15752 10220
rect 15804 10208 15810 10260
rect 16301 10251 16359 10257
rect 16301 10217 16313 10251
rect 16347 10248 16359 10251
rect 16482 10248 16488 10260
rect 16347 10220 16488 10248
rect 16347 10217 16359 10220
rect 16301 10211 16359 10217
rect 16482 10208 16488 10220
rect 16540 10208 16546 10260
rect 19334 10248 19340 10260
rect 19295 10220 19340 10248
rect 19334 10208 19340 10220
rect 19392 10208 19398 10260
rect 20438 10248 20444 10260
rect 20399 10220 20444 10248
rect 20438 10208 20444 10220
rect 20496 10208 20502 10260
rect 7190 10140 7196 10192
rect 7248 10180 7254 10192
rect 9950 10180 9956 10192
rect 7248 10152 7420 10180
rect 9911 10152 9956 10180
rect 7248 10140 7254 10152
rect 1912 10084 2912 10112
rect 1912 10072 1918 10084
rect 3234 10072 3240 10124
rect 3292 10112 3298 10124
rect 3421 10115 3479 10121
rect 3421 10112 3433 10115
rect 3292 10084 3433 10112
rect 3292 10072 3298 10084
rect 3421 10081 3433 10084
rect 3467 10081 3479 10115
rect 3421 10075 3479 10081
rect 3970 10072 3976 10124
rect 4028 10112 4034 10124
rect 4065 10115 4123 10121
rect 4065 10112 4077 10115
rect 4028 10084 4077 10112
rect 4028 10072 4034 10084
rect 4065 10081 4077 10084
rect 4111 10112 4123 10115
rect 4338 10112 4344 10124
rect 4111 10084 4344 10112
rect 4111 10081 4123 10084
rect 4065 10075 4123 10081
rect 4338 10072 4344 10084
rect 4396 10072 4402 10124
rect 4614 10072 4620 10124
rect 4672 10112 4678 10124
rect 4893 10115 4951 10121
rect 4672 10084 4765 10112
rect 4672 10072 4678 10084
rect 4893 10081 4905 10115
rect 4939 10112 4951 10115
rect 5166 10112 5172 10124
rect 4939 10084 5172 10112
rect 4939 10081 4951 10084
rect 4893 10075 4951 10081
rect 4154 10004 4160 10056
rect 4212 10044 4218 10056
rect 4908 10044 4936 10075
rect 5166 10072 5172 10084
rect 5224 10072 5230 10124
rect 5350 10112 5356 10124
rect 5311 10084 5356 10112
rect 5350 10072 5356 10084
rect 5408 10072 5414 10124
rect 7392 10121 7420 10152
rect 9950 10140 9956 10152
rect 10008 10140 10014 10192
rect 11330 10140 11336 10192
rect 11388 10180 11394 10192
rect 12253 10183 12311 10189
rect 11388 10152 11836 10180
rect 11388 10140 11394 10152
rect 6825 10115 6883 10121
rect 6825 10081 6837 10115
rect 6871 10081 6883 10115
rect 6825 10075 6883 10081
rect 7285 10115 7343 10121
rect 7285 10081 7297 10115
rect 7331 10081 7343 10115
rect 7285 10075 7343 10081
rect 7377 10115 7435 10121
rect 7377 10081 7389 10115
rect 7423 10112 7435 10115
rect 7650 10112 7656 10124
rect 7423 10084 7656 10112
rect 7423 10081 7435 10084
rect 7377 10075 7435 10081
rect 4212 10016 4936 10044
rect 6840 10044 6868 10075
rect 7190 10044 7196 10056
rect 6840 10016 7196 10044
rect 4212 10004 4218 10016
rect 7190 10004 7196 10016
rect 7248 10004 7254 10056
rect 3881 9979 3939 9985
rect 3881 9945 3893 9979
rect 3927 9976 3939 9979
rect 4430 9976 4436 9988
rect 3927 9948 4436 9976
rect 3927 9945 3939 9948
rect 3881 9939 3939 9945
rect 4430 9936 4436 9948
rect 4488 9936 4494 9988
rect 1762 9908 1768 9920
rect 1723 9880 1768 9908
rect 1762 9868 1768 9880
rect 1820 9868 1826 9920
rect 6089 9911 6147 9917
rect 6089 9877 6101 9911
rect 6135 9908 6147 9911
rect 6365 9911 6423 9917
rect 6365 9908 6377 9911
rect 6135 9880 6377 9908
rect 6135 9877 6147 9880
rect 6089 9871 6147 9877
rect 6365 9877 6377 9880
rect 6411 9908 6423 9911
rect 7300 9908 7328 10075
rect 7650 10072 7656 10084
rect 7708 10072 7714 10124
rect 7926 10112 7932 10124
rect 7887 10084 7932 10112
rect 7926 10072 7932 10084
rect 7984 10072 7990 10124
rect 10502 10112 10508 10124
rect 10463 10084 10508 10112
rect 10502 10072 10508 10084
rect 10560 10072 10566 10124
rect 11517 10115 11575 10121
rect 11517 10081 11529 10115
rect 11563 10112 11575 10115
rect 11698 10112 11704 10124
rect 11563 10084 11704 10112
rect 11563 10081 11575 10084
rect 11517 10075 11575 10081
rect 11698 10072 11704 10084
rect 11756 10072 11762 10124
rect 11808 10121 11836 10152
rect 12253 10149 12265 10183
rect 12299 10180 12311 10183
rect 13354 10180 13360 10192
rect 12299 10152 13360 10180
rect 12299 10149 12311 10152
rect 12253 10143 12311 10149
rect 13354 10140 13360 10152
rect 13412 10140 13418 10192
rect 13722 10180 13728 10192
rect 13464 10152 13728 10180
rect 11793 10115 11851 10121
rect 11793 10081 11805 10115
rect 11839 10081 11851 10115
rect 11793 10075 11851 10081
rect 13262 10072 13268 10124
rect 13320 10112 13326 10124
rect 13464 10112 13492 10152
rect 13722 10140 13728 10152
rect 13780 10140 13786 10192
rect 13814 10140 13820 10192
rect 13872 10180 13878 10192
rect 14274 10180 14280 10192
rect 13872 10152 14280 10180
rect 13872 10140 13878 10152
rect 14274 10140 14280 10152
rect 14332 10180 14338 10192
rect 14553 10183 14611 10189
rect 14553 10180 14565 10183
rect 14332 10152 14565 10180
rect 14332 10140 14338 10152
rect 14553 10149 14565 10152
rect 14599 10149 14611 10183
rect 16666 10180 16672 10192
rect 16627 10152 16672 10180
rect 14553 10143 14611 10149
rect 16666 10140 16672 10152
rect 16724 10140 16730 10192
rect 16761 10183 16819 10189
rect 16761 10149 16773 10183
rect 16807 10180 16819 10183
rect 16850 10180 16856 10192
rect 16807 10152 16856 10180
rect 16807 10149 16819 10152
rect 16761 10143 16819 10149
rect 16850 10140 16856 10152
rect 16908 10140 16914 10192
rect 17954 10140 17960 10192
rect 18012 10180 18018 10192
rect 18738 10183 18796 10189
rect 18738 10180 18750 10183
rect 18012 10152 18750 10180
rect 18012 10140 18018 10152
rect 18738 10149 18750 10152
rect 18784 10149 18796 10183
rect 19352 10180 19380 10208
rect 20070 10180 20076 10192
rect 19352 10152 20076 10180
rect 18738 10143 18796 10149
rect 20070 10140 20076 10152
rect 20128 10180 20134 10192
rect 21085 10183 21143 10189
rect 21085 10180 21097 10183
rect 20128 10152 21097 10180
rect 20128 10140 20134 10152
rect 21085 10149 21097 10152
rect 21131 10180 21143 10183
rect 21450 10180 21456 10192
rect 21131 10152 21456 10180
rect 21131 10149 21143 10152
rect 21085 10143 21143 10149
rect 21450 10140 21456 10152
rect 21508 10140 21514 10192
rect 13320 10084 13492 10112
rect 13320 10072 13326 10084
rect 14734 10072 14740 10124
rect 14792 10112 14798 10124
rect 15289 10115 15347 10121
rect 15289 10112 15301 10115
rect 14792 10084 15301 10112
rect 14792 10072 14798 10084
rect 15289 10081 15301 10084
rect 15335 10081 15347 10115
rect 15289 10075 15347 10081
rect 17313 10115 17371 10121
rect 17313 10081 17325 10115
rect 17359 10112 17371 10115
rect 18598 10112 18604 10124
rect 17359 10084 18604 10112
rect 17359 10081 17371 10084
rect 17313 10075 17371 10081
rect 18598 10072 18604 10084
rect 18656 10112 18662 10124
rect 20806 10112 20812 10124
rect 18656 10084 20812 10112
rect 18656 10072 18662 10084
rect 20806 10072 20812 10084
rect 20864 10072 20870 10124
rect 22462 10112 22468 10124
rect 22423 10084 22468 10112
rect 22462 10072 22468 10084
rect 22520 10072 22526 10124
rect 24581 10115 24639 10121
rect 24581 10081 24593 10115
rect 24627 10112 24639 10115
rect 24670 10112 24676 10124
rect 24627 10084 24676 10112
rect 24627 10081 24639 10084
rect 24581 10075 24639 10081
rect 24670 10072 24676 10084
rect 24728 10072 24734 10124
rect 13354 10004 13360 10056
rect 13412 10044 13418 10056
rect 13633 10047 13691 10053
rect 13633 10044 13645 10047
rect 13412 10016 13645 10044
rect 13412 10004 13418 10016
rect 13633 10013 13645 10016
rect 13679 10013 13691 10047
rect 18414 10044 18420 10056
rect 18375 10016 18420 10044
rect 13633 10007 13691 10013
rect 18414 10004 18420 10016
rect 18472 10004 18478 10056
rect 20990 10044 20996 10056
rect 20951 10016 20996 10044
rect 20990 10004 20996 10016
rect 21048 10004 21054 10056
rect 21266 10044 21272 10056
rect 21227 10016 21272 10044
rect 21266 10004 21272 10016
rect 21324 10004 21330 10056
rect 11606 9976 11612 9988
rect 11567 9948 11612 9976
rect 11606 9936 11612 9948
rect 11664 9936 11670 9988
rect 13538 9936 13544 9988
rect 13596 9976 13602 9988
rect 14090 9976 14096 9988
rect 13596 9948 14096 9976
rect 13596 9936 13602 9948
rect 14090 9936 14096 9948
rect 14148 9936 14154 9988
rect 19426 9936 19432 9988
rect 19484 9976 19490 9988
rect 19705 9979 19763 9985
rect 19705 9976 19717 9979
rect 19484 9948 19717 9976
rect 19484 9936 19490 9948
rect 19705 9945 19717 9948
rect 19751 9976 19763 9979
rect 22603 9979 22661 9985
rect 22603 9976 22615 9979
rect 19751 9948 22615 9976
rect 19751 9945 19763 9948
rect 19705 9939 19763 9945
rect 22603 9945 22615 9948
rect 22649 9945 22661 9979
rect 22603 9939 22661 9945
rect 7374 9908 7380 9920
rect 6411 9880 7380 9908
rect 6411 9877 6423 9880
rect 6365 9871 6423 9877
rect 7374 9868 7380 9880
rect 7432 9868 7438 9920
rect 8202 9868 8208 9920
rect 8260 9908 8266 9920
rect 8297 9911 8355 9917
rect 8297 9908 8309 9911
rect 8260 9880 8309 9908
rect 8260 9868 8266 9880
rect 8297 9877 8309 9880
rect 8343 9877 8355 9911
rect 8297 9871 8355 9877
rect 9125 9911 9183 9917
rect 9125 9877 9137 9911
rect 9171 9908 9183 9911
rect 9214 9908 9220 9920
rect 9171 9880 9220 9908
rect 9171 9877 9183 9880
rect 9125 9871 9183 9877
rect 9214 9868 9220 9880
rect 9272 9868 9278 9920
rect 10778 9868 10784 9920
rect 10836 9908 10842 9920
rect 10965 9911 11023 9917
rect 10965 9908 10977 9911
rect 10836 9880 10977 9908
rect 10836 9868 10842 9880
rect 10965 9877 10977 9880
rect 11011 9877 11023 9911
rect 11330 9908 11336 9920
rect 11291 9880 11336 9908
rect 10965 9871 11023 9877
rect 11330 9868 11336 9880
rect 11388 9868 11394 9920
rect 15838 9908 15844 9920
rect 15799 9880 15844 9908
rect 15838 9868 15844 9880
rect 15896 9868 15902 9920
rect 16482 9868 16488 9920
rect 16540 9908 16546 9920
rect 24719 9911 24777 9917
rect 24719 9908 24731 9911
rect 16540 9880 24731 9908
rect 16540 9868 16546 9880
rect 24719 9877 24731 9880
rect 24765 9877 24777 9911
rect 24719 9871 24777 9877
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 9401 9707 9459 9713
rect 9401 9673 9413 9707
rect 9447 9704 9459 9707
rect 9950 9704 9956 9716
rect 9447 9676 9956 9704
rect 9447 9673 9459 9676
rect 9401 9667 9459 9673
rect 2958 9636 2964 9648
rect 2193 9608 2964 9636
rect 2041 9571 2099 9577
rect 2041 9537 2053 9571
rect 2087 9568 2099 9571
rect 2193 9568 2221 9608
rect 2958 9596 2964 9608
rect 3016 9596 3022 9648
rect 4154 9596 4160 9648
rect 4212 9636 4218 9648
rect 6641 9639 6699 9645
rect 4212 9608 4660 9636
rect 4212 9596 4218 9608
rect 2314 9568 2320 9580
rect 2087 9540 2221 9568
rect 2275 9540 2320 9568
rect 2087 9537 2099 9540
rect 2041 9531 2099 9537
rect 2314 9528 2320 9540
rect 2372 9528 2378 9580
rect 3878 9528 3884 9580
rect 3936 9568 3942 9580
rect 4522 9568 4528 9580
rect 3936 9540 4528 9568
rect 3936 9528 3942 9540
rect 4522 9528 4528 9540
rect 4580 9528 4586 9580
rect 4632 9568 4660 9608
rect 6641 9605 6653 9639
rect 6687 9636 6699 9639
rect 7926 9636 7932 9648
rect 6687 9608 7932 9636
rect 6687 9605 6699 9608
rect 6641 9599 6699 9605
rect 7926 9596 7932 9608
rect 7984 9596 7990 9648
rect 8573 9571 8631 9577
rect 8573 9568 8585 9571
rect 4632 9540 4844 9568
rect 3786 9460 3792 9512
rect 3844 9500 3850 9512
rect 4249 9503 4307 9509
rect 4249 9500 4261 9503
rect 3844 9472 4261 9500
rect 3844 9460 3850 9472
rect 4249 9469 4261 9472
rect 4295 9469 4307 9503
rect 4614 9500 4620 9512
rect 4575 9472 4620 9500
rect 4249 9463 4307 9469
rect 2133 9435 2191 9441
rect 2133 9401 2145 9435
rect 2179 9432 2191 9435
rect 2222 9432 2228 9444
rect 2179 9404 2228 9432
rect 2179 9401 2191 9404
rect 2133 9395 2191 9401
rect 2222 9392 2228 9404
rect 2280 9392 2286 9444
rect 4154 9432 4160 9444
rect 3804 9404 4160 9432
rect 1857 9367 1915 9373
rect 1857 9333 1869 9367
rect 1903 9364 1915 9367
rect 2038 9364 2044 9376
rect 1903 9336 2044 9364
rect 1903 9333 1915 9336
rect 1857 9327 1915 9333
rect 2038 9324 2044 9336
rect 2096 9324 2102 9376
rect 2240 9364 2268 9392
rect 3804 9373 3832 9404
rect 4154 9392 4160 9404
rect 4212 9392 4218 9444
rect 4264 9432 4292 9463
rect 4614 9460 4620 9472
rect 4672 9460 4678 9512
rect 4816 9509 4844 9540
rect 7668 9540 8585 9568
rect 7668 9512 7696 9540
rect 8573 9537 8585 9540
rect 8619 9537 8631 9571
rect 8573 9531 8631 9537
rect 4801 9503 4859 9509
rect 4801 9469 4813 9503
rect 4847 9469 4859 9503
rect 5350 9500 5356 9512
rect 5311 9472 5356 9500
rect 4801 9463 4859 9469
rect 5350 9460 5356 9472
rect 5408 9460 5414 9512
rect 7101 9503 7159 9509
rect 7101 9469 7113 9503
rect 7147 9500 7159 9503
rect 7190 9500 7196 9512
rect 7147 9472 7196 9500
rect 7147 9469 7159 9472
rect 7101 9463 7159 9469
rect 7190 9460 7196 9472
rect 7248 9460 7254 9512
rect 7374 9500 7380 9512
rect 7335 9472 7380 9500
rect 7374 9460 7380 9472
rect 7432 9460 7438 9512
rect 7650 9500 7656 9512
rect 7611 9472 7656 9500
rect 7650 9460 7656 9472
rect 7708 9460 7714 9512
rect 9508 9509 9536 9676
rect 9950 9664 9956 9676
rect 10008 9664 10014 9716
rect 13262 9664 13268 9716
rect 13320 9704 13326 9716
rect 13541 9707 13599 9713
rect 13541 9704 13553 9707
rect 13320 9676 13553 9704
rect 13320 9664 13326 9676
rect 13541 9673 13553 9676
rect 13587 9673 13599 9707
rect 16850 9704 16856 9716
rect 16811 9676 16856 9704
rect 13541 9667 13599 9673
rect 16850 9664 16856 9676
rect 16908 9664 16914 9716
rect 17865 9707 17923 9713
rect 17865 9673 17877 9707
rect 17911 9704 17923 9707
rect 18046 9704 18052 9716
rect 17911 9676 18052 9704
rect 17911 9673 17923 9676
rect 17865 9667 17923 9673
rect 18046 9664 18052 9676
rect 18104 9704 18110 9716
rect 18414 9704 18420 9716
rect 18104 9676 18420 9704
rect 18104 9664 18110 9676
rect 18414 9664 18420 9676
rect 18472 9664 18478 9716
rect 19029 9676 20392 9704
rect 10042 9596 10048 9648
rect 10100 9636 10106 9648
rect 10597 9639 10655 9645
rect 10597 9636 10609 9639
rect 10100 9608 10609 9636
rect 10100 9596 10106 9608
rect 10597 9605 10609 9608
rect 10643 9636 10655 9639
rect 11517 9639 11575 9645
rect 11517 9636 11529 9639
rect 10643 9608 11529 9636
rect 10643 9605 10655 9608
rect 10597 9599 10655 9605
rect 11517 9605 11529 9608
rect 11563 9636 11575 9639
rect 11606 9636 11612 9648
rect 11563 9608 11612 9636
rect 11563 9605 11575 9608
rect 11517 9599 11575 9605
rect 11606 9596 11612 9608
rect 11664 9636 11670 9648
rect 11885 9639 11943 9645
rect 11885 9636 11897 9639
rect 11664 9608 11897 9636
rect 11664 9596 11670 9608
rect 11885 9605 11897 9608
rect 11931 9605 11943 9639
rect 11885 9599 11943 9605
rect 13630 9596 13636 9648
rect 13688 9636 13694 9648
rect 13814 9636 13820 9648
rect 13688 9608 13820 9636
rect 13688 9596 13694 9608
rect 13814 9596 13820 9608
rect 13872 9596 13878 9648
rect 14734 9596 14740 9648
rect 14792 9636 14798 9648
rect 15197 9639 15255 9645
rect 15197 9636 15209 9639
rect 14792 9608 15209 9636
rect 14792 9596 14798 9608
rect 15197 9605 15209 9608
rect 15243 9605 15255 9639
rect 15197 9599 15255 9605
rect 16666 9596 16672 9648
rect 16724 9636 16730 9648
rect 17129 9639 17187 9645
rect 17129 9636 17141 9639
rect 16724 9608 17141 9636
rect 16724 9596 16730 9608
rect 17129 9605 17141 9608
rect 17175 9605 17187 9639
rect 17129 9599 17187 9605
rect 17402 9596 17408 9648
rect 17460 9636 17466 9648
rect 19029 9636 19057 9676
rect 17460 9608 19057 9636
rect 17460 9596 17466 9608
rect 20162 9596 20168 9648
rect 20220 9636 20226 9648
rect 20364 9636 20392 9676
rect 20990 9664 20996 9716
rect 21048 9704 21054 9716
rect 21177 9707 21235 9713
rect 21177 9704 21189 9707
rect 21048 9676 21189 9704
rect 21048 9664 21054 9676
rect 21177 9673 21189 9676
rect 21223 9673 21235 9707
rect 21177 9667 21235 9673
rect 21450 9664 21456 9716
rect 21508 9704 21514 9716
rect 21545 9707 21603 9713
rect 21545 9704 21557 9707
rect 21508 9676 21557 9704
rect 21508 9664 21514 9676
rect 21545 9673 21557 9676
rect 21591 9673 21603 9707
rect 24670 9704 24676 9716
rect 24631 9676 24676 9704
rect 21545 9667 21603 9673
rect 24670 9664 24676 9676
rect 24728 9664 24734 9716
rect 22462 9636 22468 9648
rect 20220 9608 20300 9636
rect 20364 9608 22468 9636
rect 20220 9596 20226 9608
rect 11241 9571 11299 9577
rect 11241 9537 11253 9571
rect 11287 9568 11299 9571
rect 12986 9568 12992 9580
rect 11287 9540 12992 9568
rect 11287 9537 11299 9540
rect 11241 9531 11299 9537
rect 12986 9528 12992 9540
rect 13044 9528 13050 9580
rect 13722 9528 13728 9580
rect 13780 9568 13786 9580
rect 14277 9571 14335 9577
rect 14277 9568 14289 9571
rect 13780 9540 14289 9568
rect 13780 9528 13786 9540
rect 14277 9537 14289 9540
rect 14323 9537 14335 9571
rect 14277 9531 14335 9537
rect 14921 9571 14979 9577
rect 14921 9537 14933 9571
rect 14967 9568 14979 9571
rect 16114 9568 16120 9580
rect 14967 9540 16120 9568
rect 14967 9537 14979 9540
rect 14921 9531 14979 9537
rect 16114 9528 16120 9540
rect 16172 9528 16178 9580
rect 17954 9528 17960 9580
rect 18012 9568 18018 9580
rect 18233 9571 18291 9577
rect 18233 9568 18245 9571
rect 18012 9540 18245 9568
rect 18012 9528 18018 9540
rect 18233 9537 18245 9540
rect 18279 9537 18291 9571
rect 18233 9531 18291 9537
rect 18417 9571 18475 9577
rect 18417 9537 18429 9571
rect 18463 9568 18475 9571
rect 18782 9568 18788 9580
rect 18463 9540 18788 9568
rect 18463 9537 18475 9540
rect 18417 9531 18475 9537
rect 8205 9503 8263 9509
rect 8205 9469 8217 9503
rect 8251 9469 8263 9503
rect 8205 9463 8263 9469
rect 9493 9503 9551 9509
rect 9493 9469 9505 9503
rect 9539 9469 9551 9503
rect 10502 9500 10508 9512
rect 10415 9472 10508 9500
rect 9493 9463 9551 9469
rect 4338 9432 4344 9444
rect 4264 9404 4344 9432
rect 4338 9392 4344 9404
rect 4396 9432 4402 9444
rect 6273 9435 6331 9441
rect 4396 9404 5304 9432
rect 4396 9392 4402 9404
rect 5276 9376 5304 9404
rect 6273 9401 6285 9435
rect 6319 9432 6331 9435
rect 8220 9432 8248 9463
rect 10502 9460 10508 9472
rect 10560 9460 10566 9512
rect 10778 9500 10784 9512
rect 10739 9472 10784 9500
rect 10778 9460 10784 9472
rect 10836 9460 10842 9512
rect 12618 9500 12624 9512
rect 12579 9472 12624 9500
rect 12618 9460 12624 9472
rect 12676 9460 12682 9512
rect 12802 9460 12808 9512
rect 12860 9500 12866 9512
rect 12897 9503 12955 9509
rect 12897 9500 12909 9503
rect 12860 9472 12909 9500
rect 12860 9460 12866 9472
rect 12897 9469 12909 9472
rect 12943 9469 12955 9503
rect 12897 9463 12955 9469
rect 9122 9432 9128 9444
rect 6319 9404 7144 9432
rect 6319 9401 6331 9404
rect 6273 9395 6331 9401
rect 7116 9376 7144 9404
rect 8220 9404 9128 9432
rect 2961 9367 3019 9373
rect 2961 9364 2973 9367
rect 2240 9336 2973 9364
rect 2961 9333 2973 9336
rect 3007 9333 3019 9367
rect 2961 9327 3019 9333
rect 3513 9367 3571 9373
rect 3513 9333 3525 9367
rect 3559 9364 3571 9367
rect 3789 9367 3847 9373
rect 3789 9364 3801 9367
rect 3559 9336 3801 9364
rect 3559 9333 3571 9336
rect 3513 9327 3571 9333
rect 3789 9333 3801 9336
rect 3835 9333 3847 9367
rect 3789 9327 3847 9333
rect 3970 9324 3976 9376
rect 4028 9364 4034 9376
rect 4065 9367 4123 9373
rect 4065 9364 4077 9367
rect 4028 9336 4077 9364
rect 4028 9324 4034 9336
rect 4065 9333 4077 9336
rect 4111 9333 4123 9367
rect 4065 9327 4123 9333
rect 5258 9324 5264 9376
rect 5316 9364 5322 9376
rect 5721 9367 5779 9373
rect 5721 9364 5733 9367
rect 5316 9336 5733 9364
rect 5316 9324 5322 9336
rect 5721 9333 5733 9336
rect 5767 9333 5779 9367
rect 5721 9327 5779 9333
rect 6730 9324 6736 9376
rect 6788 9364 6794 9376
rect 6917 9367 6975 9373
rect 6917 9364 6929 9367
rect 6788 9336 6929 9364
rect 6788 9324 6794 9336
rect 6917 9333 6929 9336
rect 6963 9333 6975 9367
rect 6917 9327 6975 9333
rect 7098 9324 7104 9376
rect 7156 9364 7162 9376
rect 8220 9364 8248 9404
rect 9122 9392 9128 9404
rect 9180 9432 9186 9444
rect 10134 9432 10140 9444
rect 9180 9404 10140 9432
rect 9180 9392 9186 9404
rect 10134 9392 10140 9404
rect 10192 9392 10198 9444
rect 7156 9336 8248 9364
rect 9033 9367 9091 9373
rect 7156 9324 7162 9336
rect 9033 9333 9045 9367
rect 9079 9364 9091 9367
rect 9214 9364 9220 9376
rect 9079 9336 9220 9364
rect 9079 9333 9091 9336
rect 9033 9327 9091 9333
rect 9214 9324 9220 9336
rect 9272 9324 9278 9376
rect 9306 9324 9312 9376
rect 9364 9364 9370 9376
rect 9677 9367 9735 9373
rect 9677 9364 9689 9367
rect 9364 9336 9689 9364
rect 9364 9324 9370 9336
rect 9677 9333 9689 9336
rect 9723 9333 9735 9367
rect 10042 9364 10048 9376
rect 9955 9336 10048 9364
rect 9677 9327 9735 9333
rect 10042 9324 10048 9336
rect 10100 9364 10106 9376
rect 10413 9367 10471 9373
rect 10413 9364 10425 9367
rect 10100 9336 10425 9364
rect 10100 9324 10106 9336
rect 10413 9333 10425 9336
rect 10459 9364 10471 9367
rect 10520 9364 10548 9460
rect 14369 9435 14427 9441
rect 14369 9432 14381 9435
rect 14016 9404 14381 9432
rect 11238 9364 11244 9376
rect 10459 9336 11244 9364
rect 10459 9333 10471 9336
rect 10413 9327 10471 9333
rect 11238 9324 11244 9336
rect 11296 9324 11302 9376
rect 12526 9364 12532 9376
rect 12487 9336 12532 9364
rect 12526 9324 12532 9336
rect 12584 9324 12590 9376
rect 13814 9324 13820 9376
rect 13872 9364 13878 9376
rect 14016 9373 14044 9404
rect 14369 9401 14381 9404
rect 14415 9401 14427 9435
rect 15838 9432 15844 9444
rect 15799 9404 15844 9432
rect 14369 9395 14427 9401
rect 15838 9392 15844 9404
rect 15896 9392 15902 9444
rect 15933 9435 15991 9441
rect 15933 9401 15945 9435
rect 15979 9401 15991 9435
rect 18248 9432 18276 9531
rect 18782 9528 18788 9540
rect 18840 9528 18846 9580
rect 20272 9577 20300 9608
rect 22462 9596 22468 9608
rect 22520 9596 22526 9648
rect 20257 9571 20315 9577
rect 20257 9537 20269 9571
rect 20303 9537 20315 9571
rect 20898 9568 20904 9580
rect 20859 9540 20904 9568
rect 20257 9531 20315 9537
rect 20898 9528 20904 9540
rect 20956 9528 20962 9580
rect 18738 9435 18796 9441
rect 18738 9432 18750 9435
rect 18248 9404 18750 9432
rect 15933 9395 15991 9401
rect 18738 9401 18750 9404
rect 18784 9401 18796 9435
rect 18738 9395 18796 9401
rect 20349 9435 20407 9441
rect 20349 9401 20361 9435
rect 20395 9401 20407 9435
rect 20349 9395 20407 9401
rect 14001 9367 14059 9373
rect 14001 9364 14013 9367
rect 13872 9336 14013 9364
rect 13872 9324 13878 9336
rect 14001 9333 14013 9336
rect 14047 9333 14059 9367
rect 15562 9364 15568 9376
rect 15523 9336 15568 9364
rect 14001 9327 14059 9333
rect 15562 9324 15568 9336
rect 15620 9364 15626 9376
rect 15948 9364 15976 9395
rect 15620 9336 15976 9364
rect 19337 9367 19395 9373
rect 15620 9324 15626 9336
rect 19337 9333 19349 9367
rect 19383 9364 19395 9367
rect 19981 9367 20039 9373
rect 19981 9364 19993 9367
rect 19383 9336 19993 9364
rect 19383 9333 19395 9336
rect 19337 9327 19395 9333
rect 19981 9333 19993 9336
rect 20027 9364 20039 9367
rect 20364 9364 20392 9395
rect 20027 9336 20392 9364
rect 20027 9333 20039 9336
rect 19981 9327 20039 9333
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 1765 9163 1823 9169
rect 1765 9129 1777 9163
rect 1811 9160 1823 9163
rect 1854 9160 1860 9172
rect 1811 9132 1860 9160
rect 1811 9129 1823 9132
rect 1765 9123 1823 9129
rect 1854 9120 1860 9132
rect 1912 9120 1918 9172
rect 2038 9120 2044 9172
rect 2096 9120 2102 9172
rect 3786 9160 3792 9172
rect 3747 9132 3792 9160
rect 3786 9120 3792 9132
rect 3844 9120 3850 9172
rect 7282 9120 7288 9172
rect 7340 9160 7346 9172
rect 8386 9160 8392 9172
rect 7340 9132 8392 9160
rect 7340 9120 7346 9132
rect 8386 9120 8392 9132
rect 8444 9160 8450 9172
rect 8665 9163 8723 9169
rect 8665 9160 8677 9163
rect 8444 9132 8677 9160
rect 8444 9120 8450 9132
rect 8665 9129 8677 9132
rect 8711 9129 8723 9163
rect 8665 9123 8723 9129
rect 10134 9120 10140 9172
rect 10192 9160 10198 9172
rect 11517 9163 11575 9169
rect 11517 9160 11529 9163
rect 10192 9132 11529 9160
rect 10192 9120 10198 9132
rect 11517 9129 11529 9132
rect 11563 9160 11575 9163
rect 11698 9160 11704 9172
rect 11563 9132 11704 9160
rect 11563 9129 11575 9132
rect 11517 9123 11575 9129
rect 11698 9120 11704 9132
rect 11756 9120 11762 9172
rect 12802 9160 12808 9172
rect 12763 9132 12808 9160
rect 12802 9120 12808 9132
rect 12860 9120 12866 9172
rect 17954 9120 17960 9172
rect 18012 9160 18018 9172
rect 18417 9163 18475 9169
rect 18417 9160 18429 9163
rect 18012 9132 18429 9160
rect 18012 9120 18018 9132
rect 18417 9129 18429 9132
rect 18463 9129 18475 9163
rect 20162 9160 20168 9172
rect 20123 9132 20168 9160
rect 18417 9123 18475 9129
rect 20162 9120 20168 9132
rect 20220 9120 20226 9172
rect 20901 9163 20959 9169
rect 20901 9129 20913 9163
rect 20947 9160 20959 9163
rect 20990 9160 20996 9172
rect 20947 9132 20996 9160
rect 20947 9129 20959 9132
rect 20901 9123 20959 9129
rect 20990 9120 20996 9132
rect 21048 9120 21054 9172
rect 22465 9163 22523 9169
rect 22465 9129 22477 9163
rect 22511 9160 22523 9163
rect 27614 9160 27620 9172
rect 22511 9132 27620 9160
rect 22511 9129 22523 9132
rect 22465 9123 22523 9129
rect 27614 9120 27620 9132
rect 27672 9120 27678 9172
rect 2056 9092 2084 9120
rect 2219 9095 2277 9101
rect 2219 9092 2231 9095
rect 2056 9064 2231 9092
rect 2219 9061 2231 9064
rect 2265 9092 2277 9095
rect 2866 9092 2872 9104
rect 2265 9064 2872 9092
rect 2265 9061 2277 9064
rect 2219 9055 2277 9061
rect 2866 9052 2872 9064
rect 2924 9052 2930 9104
rect 3418 9092 3424 9104
rect 3379 9064 3424 9092
rect 3418 9052 3424 9064
rect 3476 9052 3482 9104
rect 4246 9092 4252 9104
rect 4207 9064 4252 9092
rect 4246 9052 4252 9064
rect 4304 9052 4310 9104
rect 5350 9052 5356 9104
rect 5408 9092 5414 9104
rect 5813 9095 5871 9101
rect 5813 9092 5825 9095
rect 5408 9064 5825 9092
rect 5408 9052 5414 9064
rect 5813 9061 5825 9064
rect 5859 9092 5871 9095
rect 10873 9095 10931 9101
rect 5859 9064 8340 9092
rect 5859 9061 5871 9064
rect 5813 9055 5871 9061
rect 8312 9036 8340 9064
rect 10873 9061 10885 9095
rect 10919 9092 10931 9095
rect 11330 9092 11336 9104
rect 10919 9064 11336 9092
rect 10919 9061 10931 9064
rect 10873 9055 10931 9061
rect 11330 9052 11336 9064
rect 11388 9052 11394 9104
rect 14369 9095 14427 9101
rect 11532 9064 11928 9092
rect 1857 9027 1915 9033
rect 1857 8993 1869 9027
rect 1903 9024 1915 9027
rect 2038 9024 2044 9036
rect 1903 8996 2044 9024
rect 1903 8993 1915 8996
rect 1857 8987 1915 8993
rect 2038 8984 2044 8996
rect 2096 9024 2102 9036
rect 3970 9024 3976 9036
rect 2096 8996 3976 9024
rect 2096 8984 2102 8996
rect 3970 8984 3976 8996
rect 4028 8984 4034 9036
rect 5905 9027 5963 9033
rect 5905 8993 5917 9027
rect 5951 9024 5963 9027
rect 5994 9024 6000 9036
rect 5951 8996 6000 9024
rect 5951 8993 5963 8996
rect 5905 8987 5963 8993
rect 5994 8984 6000 8996
rect 6052 8984 6058 9036
rect 7190 9024 7196 9036
rect 7151 8996 7196 9024
rect 7190 8984 7196 8996
rect 7248 8984 7254 9036
rect 7374 9024 7380 9036
rect 7335 8996 7380 9024
rect 7374 8984 7380 8996
rect 7432 8984 7438 9036
rect 7745 9027 7803 9033
rect 7745 8993 7757 9027
rect 7791 8993 7803 9027
rect 8294 9024 8300 9036
rect 8255 8996 8300 9024
rect 7745 8987 7803 8993
rect 4154 8916 4160 8968
rect 4212 8956 4218 8968
rect 4430 8956 4436 8968
rect 4212 8928 4257 8956
rect 4391 8928 4436 8956
rect 4212 8916 4218 8928
rect 4430 8916 4436 8928
rect 4488 8916 4494 8968
rect 6086 8916 6092 8968
rect 6144 8956 6150 8968
rect 7006 8956 7012 8968
rect 6144 8928 7012 8956
rect 6144 8916 6150 8928
rect 7006 8916 7012 8928
rect 7064 8916 7070 8968
rect 7760 8956 7788 8987
rect 8294 8984 8300 8996
rect 8352 8984 8358 9036
rect 10778 9024 10784 9036
rect 10691 8996 10784 9024
rect 10778 8984 10784 8996
rect 10836 9024 10842 9036
rect 11532 9024 11560 9064
rect 11900 9036 11928 9064
rect 14369 9061 14381 9095
rect 14415 9092 14427 9095
rect 15562 9092 15568 9104
rect 14415 9064 15568 9092
rect 14415 9061 14427 9064
rect 14369 9055 14427 9061
rect 15562 9052 15568 9064
rect 15620 9052 15626 9104
rect 18046 9092 18052 9104
rect 18007 9064 18052 9092
rect 18046 9052 18052 9064
rect 18104 9052 18110 9104
rect 11698 9024 11704 9036
rect 10836 8996 11560 9024
rect 11659 8996 11704 9024
rect 10836 8984 10842 8996
rect 11698 8984 11704 8996
rect 11756 8984 11762 9036
rect 11882 8984 11888 9036
rect 11940 9024 11946 9036
rect 11977 9027 12035 9033
rect 11977 9024 11989 9027
rect 11940 8996 11989 9024
rect 11940 8984 11946 8996
rect 11977 8993 11989 8996
rect 12023 8993 12035 9027
rect 11977 8987 12035 8993
rect 13814 8984 13820 9036
rect 13872 9024 13878 9036
rect 15378 9024 15384 9036
rect 13872 8996 13917 9024
rect 15339 8996 15384 9024
rect 13872 8984 13878 8996
rect 15378 8984 15384 8996
rect 15436 8984 15442 9036
rect 17310 9024 17316 9036
rect 17271 8996 17316 9024
rect 17310 8984 17316 8996
rect 17368 8984 17374 9036
rect 17678 8984 17684 9036
rect 17736 9024 17742 9036
rect 17773 9027 17831 9033
rect 17773 9024 17785 9027
rect 17736 8996 17785 9024
rect 17736 8984 17742 8996
rect 17773 8993 17785 8996
rect 17819 8993 17831 9027
rect 17773 8987 17831 8993
rect 19705 9027 19763 9033
rect 19705 8993 19717 9027
rect 19751 9024 19763 9027
rect 19794 9024 19800 9036
rect 19751 8996 19800 9024
rect 19751 8993 19763 8996
rect 19705 8987 19763 8993
rect 19794 8984 19800 8996
rect 19852 8984 19858 9036
rect 22186 8984 22192 9036
rect 22244 9024 22250 9036
rect 22281 9027 22339 9033
rect 22281 9024 22293 9027
rect 22244 8996 22293 9024
rect 22244 8984 22250 8996
rect 22281 8993 22293 8996
rect 22327 8993 22339 9027
rect 22281 8987 22339 8993
rect 7161 8928 7788 8956
rect 8389 8959 8447 8965
rect 3145 8891 3203 8897
rect 3145 8857 3157 8891
rect 3191 8888 3203 8891
rect 3510 8888 3516 8900
rect 3191 8860 3516 8888
rect 3191 8857 3203 8860
rect 3145 8851 3203 8857
rect 3510 8848 3516 8860
rect 3568 8888 3574 8900
rect 3568 8860 4292 8888
rect 3568 8848 3574 8860
rect 2774 8820 2780 8832
rect 2735 8792 2780 8820
rect 2774 8780 2780 8792
rect 2832 8780 2838 8832
rect 4264 8820 4292 8860
rect 4338 8848 4344 8900
rect 4396 8888 4402 8900
rect 6549 8891 6607 8897
rect 6549 8888 6561 8891
rect 4396 8860 6561 8888
rect 4396 8848 4402 8860
rect 6549 8857 6561 8860
rect 6595 8857 6607 8891
rect 6549 8851 6607 8857
rect 6638 8848 6644 8900
rect 6696 8888 6702 8900
rect 7161 8888 7189 8928
rect 8389 8925 8401 8959
rect 8435 8956 8447 8959
rect 12342 8956 12348 8968
rect 8435 8928 12348 8956
rect 8435 8925 8447 8928
rect 8389 8919 8447 8925
rect 12342 8916 12348 8928
rect 12400 8916 12406 8968
rect 12437 8959 12495 8965
rect 12437 8925 12449 8959
rect 12483 8956 12495 8959
rect 14550 8956 14556 8968
rect 12483 8928 14556 8956
rect 12483 8925 12495 8928
rect 12437 8919 12495 8925
rect 14550 8916 14556 8928
rect 14608 8916 14614 8968
rect 6696 8860 7189 8888
rect 6696 8848 6702 8860
rect 11698 8848 11704 8900
rect 11756 8888 11762 8900
rect 11793 8891 11851 8897
rect 11793 8888 11805 8891
rect 11756 8860 11805 8888
rect 11756 8848 11762 8860
rect 11793 8857 11805 8860
rect 11839 8857 11851 8891
rect 11793 8851 11851 8857
rect 4614 8820 4620 8832
rect 4264 8792 4620 8820
rect 4614 8780 4620 8792
rect 4672 8780 4678 8832
rect 5074 8820 5080 8832
rect 5035 8792 5080 8820
rect 5074 8780 5080 8792
rect 5132 8780 5138 8832
rect 6089 8823 6147 8829
rect 6089 8789 6101 8823
rect 6135 8820 6147 8823
rect 7190 8820 7196 8832
rect 6135 8792 7196 8820
rect 6135 8789 6147 8792
rect 6089 8783 6147 8789
rect 7190 8780 7196 8792
rect 7248 8820 7254 8832
rect 7558 8820 7564 8832
rect 7248 8792 7564 8820
rect 7248 8780 7254 8792
rect 7558 8780 7564 8792
rect 7616 8780 7622 8832
rect 9125 8823 9183 8829
rect 9125 8789 9137 8823
rect 9171 8820 9183 8823
rect 9214 8820 9220 8832
rect 9171 8792 9220 8820
rect 9171 8789 9183 8792
rect 9125 8783 9183 8789
rect 9214 8780 9220 8792
rect 9272 8780 9278 8832
rect 13354 8780 13360 8832
rect 13412 8820 13418 8832
rect 13541 8823 13599 8829
rect 13541 8820 13553 8823
rect 13412 8792 13553 8820
rect 13412 8780 13418 8792
rect 13541 8789 13553 8792
rect 13587 8820 13599 8823
rect 13722 8820 13728 8832
rect 13587 8792 13728 8820
rect 13587 8789 13599 8792
rect 13541 8783 13599 8789
rect 13722 8780 13728 8792
rect 13780 8780 13786 8832
rect 15746 8820 15752 8832
rect 15707 8792 15752 8820
rect 15746 8780 15752 8792
rect 15804 8780 15810 8832
rect 18782 8820 18788 8832
rect 18743 8792 18788 8820
rect 18782 8780 18788 8792
rect 18840 8780 18846 8832
rect 19843 8823 19901 8829
rect 19843 8789 19855 8823
rect 19889 8820 19901 8823
rect 19978 8820 19984 8832
rect 19889 8792 19984 8820
rect 19889 8789 19901 8792
rect 19843 8783 19901 8789
rect 19978 8780 19984 8792
rect 20036 8780 20042 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 3234 8576 3240 8628
rect 3292 8616 3298 8628
rect 3605 8619 3663 8625
rect 3605 8616 3617 8619
rect 3292 8588 3617 8616
rect 3292 8576 3298 8588
rect 3605 8585 3617 8588
rect 3651 8616 3663 8619
rect 3786 8616 3792 8628
rect 3651 8588 3792 8616
rect 3651 8585 3663 8588
rect 3605 8579 3663 8585
rect 3786 8576 3792 8588
rect 3844 8616 3850 8628
rect 5350 8616 5356 8628
rect 3844 8588 5356 8616
rect 3844 8576 3850 8588
rect 5350 8576 5356 8588
rect 5408 8576 5414 8628
rect 5534 8576 5540 8628
rect 5592 8616 5598 8628
rect 5994 8616 6000 8628
rect 5592 8588 6000 8616
rect 5592 8576 5598 8588
rect 5994 8576 6000 8588
rect 6052 8616 6058 8628
rect 6181 8619 6239 8625
rect 6181 8616 6193 8619
rect 6052 8588 6193 8616
rect 6052 8576 6058 8588
rect 6181 8585 6193 8588
rect 6227 8585 6239 8619
rect 6546 8616 6552 8628
rect 6507 8588 6552 8616
rect 6181 8579 6239 8585
rect 6546 8576 6552 8588
rect 6604 8576 6610 8628
rect 7098 8616 7104 8628
rect 6656 8588 7104 8616
rect 3329 8551 3387 8557
rect 3329 8517 3341 8551
rect 3375 8548 3387 8551
rect 6656 8548 6684 8588
rect 7098 8576 7104 8588
rect 7156 8576 7162 8628
rect 7469 8619 7527 8625
rect 7469 8585 7481 8619
rect 7515 8616 7527 8619
rect 10042 8616 10048 8628
rect 7515 8588 10048 8616
rect 7515 8585 7527 8588
rect 7469 8579 7527 8585
rect 3375 8520 6684 8548
rect 3375 8517 3387 8520
rect 3329 8511 3387 8517
rect 2130 8480 2136 8492
rect 2091 8452 2136 8480
rect 2130 8440 2136 8452
rect 2188 8440 2194 8492
rect 3436 8421 3464 8520
rect 3421 8415 3479 8421
rect 3421 8381 3433 8415
rect 3467 8381 3479 8415
rect 4706 8412 4712 8424
rect 4667 8384 4712 8412
rect 3421 8375 3479 8381
rect 4706 8372 4712 8384
rect 4764 8372 4770 8424
rect 5166 8412 5172 8424
rect 5127 8384 5172 8412
rect 5166 8372 5172 8384
rect 5224 8372 5230 8424
rect 5261 8415 5319 8421
rect 5261 8381 5273 8415
rect 5307 8381 5319 8415
rect 5261 8375 5319 8381
rect 1762 8344 1768 8356
rect 1723 8316 1768 8344
rect 1762 8304 1768 8316
rect 1820 8304 1826 8356
rect 1854 8304 1860 8356
rect 1912 8344 1918 8356
rect 1912 8316 1957 8344
rect 1912 8304 1918 8316
rect 5074 8304 5080 8356
rect 5132 8344 5138 8356
rect 5276 8344 5304 8375
rect 5350 8372 5356 8424
rect 5408 8412 5414 8424
rect 5629 8415 5687 8421
rect 5629 8412 5641 8415
rect 5408 8384 5641 8412
rect 5408 8372 5414 8384
rect 5629 8381 5641 8384
rect 5675 8381 5687 8415
rect 5629 8375 5687 8381
rect 6917 8415 6975 8421
rect 6917 8381 6929 8415
rect 6963 8412 6975 8415
rect 7484 8412 7512 8579
rect 10042 8576 10048 8588
rect 10100 8576 10106 8628
rect 10229 8619 10287 8625
rect 10229 8585 10241 8619
rect 10275 8616 10287 8619
rect 10778 8616 10784 8628
rect 10275 8588 10784 8616
rect 10275 8585 10287 8588
rect 10229 8579 10287 8585
rect 10778 8576 10784 8588
rect 10836 8576 10842 8628
rect 13449 8619 13507 8625
rect 13449 8585 13461 8619
rect 13495 8616 13507 8619
rect 14185 8619 14243 8625
rect 14185 8616 14197 8619
rect 13495 8588 14197 8616
rect 13495 8585 13507 8588
rect 13449 8579 13507 8585
rect 14185 8585 14197 8588
rect 14231 8616 14243 8619
rect 14458 8616 14464 8628
rect 14231 8588 14464 8616
rect 14231 8585 14243 8588
rect 14185 8579 14243 8585
rect 14458 8576 14464 8588
rect 14516 8616 14522 8628
rect 15378 8616 15384 8628
rect 14516 8588 15384 8616
rect 14516 8576 14522 8588
rect 15378 8576 15384 8588
rect 15436 8576 15442 8628
rect 15746 8616 15752 8628
rect 15707 8588 15752 8616
rect 15746 8576 15752 8588
rect 15804 8576 15810 8628
rect 17310 8616 17316 8628
rect 17271 8588 17316 8616
rect 17310 8576 17316 8588
rect 17368 8576 17374 8628
rect 22186 8576 22192 8628
rect 22244 8616 22250 8628
rect 22281 8619 22339 8625
rect 22281 8616 22293 8619
rect 22244 8588 22293 8616
rect 22244 8576 22250 8588
rect 22281 8585 22293 8588
rect 22327 8585 22339 8619
rect 22281 8579 22339 8585
rect 23382 8576 23388 8628
rect 23440 8616 23446 8628
rect 23799 8619 23857 8625
rect 23799 8616 23811 8619
rect 23440 8588 23811 8616
rect 23440 8576 23446 8588
rect 23799 8585 23811 8588
rect 23845 8585 23857 8619
rect 23799 8579 23857 8585
rect 13814 8508 13820 8560
rect 13872 8548 13878 8560
rect 13872 8520 13917 8548
rect 13872 8508 13878 8520
rect 16022 8508 16028 8560
rect 16080 8548 16086 8560
rect 17037 8551 17095 8557
rect 16080 8520 16942 8548
rect 16080 8508 16086 8520
rect 8570 8440 8576 8492
rect 8628 8480 8634 8492
rect 9582 8480 9588 8492
rect 8628 8452 9588 8480
rect 8628 8440 8634 8452
rect 6963 8384 7512 8412
rect 6963 8381 6975 8384
rect 6917 8375 6975 8381
rect 7558 8372 7564 8424
rect 7616 8412 7622 8424
rect 7929 8415 7987 8421
rect 7929 8412 7941 8415
rect 7616 8384 7941 8412
rect 7616 8372 7622 8384
rect 7929 8381 7941 8384
rect 7975 8381 7987 8415
rect 8386 8412 8392 8424
rect 8347 8384 8392 8412
rect 7929 8375 7987 8381
rect 8386 8372 8392 8384
rect 8444 8372 8450 8424
rect 8956 8421 8984 8452
rect 9582 8440 9588 8452
rect 9640 8440 9646 8492
rect 12342 8440 12348 8492
rect 12400 8480 12406 8492
rect 12529 8483 12587 8489
rect 12529 8480 12541 8483
rect 12400 8452 12541 8480
rect 12400 8440 12406 8452
rect 12529 8449 12541 8452
rect 12575 8449 12587 8483
rect 12529 8443 12587 8449
rect 15013 8483 15071 8489
rect 15013 8449 15025 8483
rect 15059 8480 15071 8483
rect 15378 8480 15384 8492
rect 15059 8452 15384 8480
rect 15059 8449 15071 8452
rect 15013 8443 15071 8449
rect 15378 8440 15384 8452
rect 15436 8480 15442 8492
rect 16209 8483 16267 8489
rect 16209 8480 16221 8483
rect 15436 8452 16221 8480
rect 15436 8440 15442 8452
rect 16209 8449 16221 8452
rect 16255 8449 16267 8483
rect 16209 8443 16267 8449
rect 8941 8415 8999 8421
rect 8941 8381 8953 8415
rect 8987 8381 8999 8415
rect 8941 8375 8999 8381
rect 9125 8415 9183 8421
rect 9125 8381 9137 8415
rect 9171 8412 9183 8415
rect 9306 8412 9312 8424
rect 9171 8384 9312 8412
rect 9171 8381 9183 8384
rect 9125 8375 9183 8381
rect 5132 8316 5304 8344
rect 5132 8304 5138 8316
rect 2777 8279 2835 8285
rect 2777 8245 2789 8279
rect 2823 8276 2835 8279
rect 2866 8276 2872 8288
rect 2823 8248 2872 8276
rect 2823 8245 2835 8248
rect 2777 8239 2835 8245
rect 2866 8236 2872 8248
rect 2924 8236 2930 8288
rect 3970 8236 3976 8288
rect 4028 8276 4034 8288
rect 4065 8279 4123 8285
rect 4065 8276 4077 8279
rect 4028 8248 4077 8276
rect 4028 8236 4034 8248
rect 4065 8245 4077 8248
rect 4111 8276 4123 8279
rect 4246 8276 4252 8288
rect 4111 8248 4252 8276
rect 4111 8245 4123 8248
rect 4065 8239 4123 8245
rect 4246 8236 4252 8248
rect 4304 8236 4310 8288
rect 5276 8276 5304 8316
rect 5905 8347 5963 8353
rect 5905 8313 5917 8347
rect 5951 8344 5963 8347
rect 9030 8344 9036 8356
rect 5951 8316 9036 8344
rect 5951 8313 5963 8316
rect 5905 8307 5963 8313
rect 9030 8304 9036 8316
rect 9088 8304 9094 8356
rect 5994 8276 6000 8288
rect 5276 8248 6000 8276
rect 5994 8236 6000 8248
rect 6052 8236 6058 8288
rect 7837 8279 7895 8285
rect 7837 8245 7849 8279
rect 7883 8276 7895 8279
rect 7926 8276 7932 8288
rect 7883 8248 7932 8276
rect 7883 8245 7895 8248
rect 7837 8239 7895 8245
rect 7926 8236 7932 8248
rect 7984 8276 7990 8288
rect 9140 8276 9168 8375
rect 9306 8372 9312 8384
rect 9364 8372 9370 8424
rect 11793 8415 11851 8421
rect 11793 8381 11805 8415
rect 11839 8412 11851 8415
rect 11882 8412 11888 8424
rect 11839 8384 11888 8412
rect 11839 8381 11851 8384
rect 11793 8375 11851 8381
rect 11882 8372 11888 8384
rect 11940 8412 11946 8424
rect 13354 8412 13360 8424
rect 11940 8384 13360 8412
rect 11940 8372 11946 8384
rect 13354 8372 13360 8384
rect 13412 8372 13418 8424
rect 16914 8412 16942 8520
rect 17037 8517 17049 8551
rect 17083 8548 17095 8551
rect 17678 8548 17684 8560
rect 17083 8520 17684 8548
rect 17083 8517 17095 8520
rect 17037 8511 17095 8517
rect 17678 8508 17684 8520
rect 17736 8508 17742 8560
rect 19794 8548 19800 8560
rect 19707 8520 19800 8548
rect 19794 8508 19800 8520
rect 19852 8548 19858 8560
rect 20622 8548 20628 8560
rect 19852 8520 20628 8548
rect 19852 8508 19858 8520
rect 20622 8508 20628 8520
rect 20680 8508 20686 8560
rect 17696 8480 17724 8508
rect 18782 8480 18788 8492
rect 17696 8452 18552 8480
rect 18743 8452 18788 8480
rect 18524 8424 18552 8452
rect 18782 8440 18788 8452
rect 18840 8440 18846 8492
rect 19429 8483 19487 8489
rect 19429 8449 19441 8483
rect 19475 8480 19487 8483
rect 19978 8480 19984 8492
rect 19475 8452 19984 8480
rect 19475 8449 19487 8452
rect 19429 8443 19487 8449
rect 19978 8440 19984 8452
rect 20036 8440 20042 8492
rect 20162 8440 20168 8492
rect 20220 8480 20226 8492
rect 20257 8483 20315 8489
rect 20257 8480 20269 8483
rect 20220 8452 20269 8480
rect 20220 8440 20226 8452
rect 20257 8449 20269 8452
rect 20303 8449 20315 8483
rect 20257 8443 20315 8449
rect 17773 8415 17831 8421
rect 17773 8412 17785 8415
rect 16914 8384 17785 8412
rect 17773 8381 17785 8384
rect 17819 8412 17831 8415
rect 18049 8415 18107 8421
rect 18049 8412 18061 8415
rect 17819 8384 18061 8412
rect 17819 8381 17831 8384
rect 17773 8375 17831 8381
rect 18049 8381 18061 8384
rect 18095 8381 18107 8415
rect 18506 8412 18512 8424
rect 18419 8384 18512 8412
rect 18049 8375 18107 8381
rect 18506 8372 18512 8384
rect 18564 8372 18570 8424
rect 23728 8415 23786 8421
rect 23728 8381 23740 8415
rect 23774 8412 23786 8415
rect 24118 8412 24124 8424
rect 23774 8384 24124 8412
rect 23774 8381 23786 8384
rect 23728 8375 23786 8381
rect 24118 8372 24124 8384
rect 24176 8372 24182 8424
rect 9398 8344 9404 8356
rect 9359 8316 9404 8344
rect 9398 8304 9404 8316
rect 9456 8304 9462 8356
rect 9950 8304 9956 8356
rect 10008 8344 10014 8356
rect 10505 8347 10563 8353
rect 10505 8344 10517 8347
rect 10008 8316 10517 8344
rect 10008 8304 10014 8316
rect 10505 8313 10517 8316
rect 10551 8313 10563 8347
rect 10505 8307 10563 8313
rect 10597 8347 10655 8353
rect 10597 8313 10609 8347
rect 10643 8344 10655 8347
rect 10962 8344 10968 8356
rect 10643 8316 10968 8344
rect 10643 8313 10655 8316
rect 10597 8307 10655 8313
rect 10962 8304 10968 8316
rect 11020 8304 11026 8356
rect 11146 8344 11152 8356
rect 11107 8316 11152 8344
rect 11146 8304 11152 8316
rect 11204 8304 11210 8356
rect 12891 8347 12949 8353
rect 12891 8313 12903 8347
rect 12937 8313 12949 8347
rect 14366 8344 14372 8356
rect 14327 8316 14372 8344
rect 12891 8307 12949 8313
rect 7984 8248 9168 8276
rect 7984 8236 7990 8248
rect 9582 8236 9588 8288
rect 9640 8276 9646 8288
rect 9677 8279 9735 8285
rect 9677 8276 9689 8279
rect 9640 8248 9689 8276
rect 9640 8236 9646 8248
rect 9677 8245 9689 8248
rect 9723 8245 9735 8279
rect 9677 8239 9735 8245
rect 12253 8279 12311 8285
rect 12253 8245 12265 8279
rect 12299 8276 12311 8279
rect 12906 8276 12934 8307
rect 14366 8304 14372 8316
rect 14424 8304 14430 8356
rect 14458 8304 14464 8356
rect 14516 8344 14522 8356
rect 15930 8344 15936 8356
rect 14516 8316 14561 8344
rect 15891 8316 15936 8344
rect 14516 8304 14522 8316
rect 15930 8304 15936 8316
rect 15988 8304 15994 8356
rect 16025 8347 16083 8353
rect 16025 8313 16037 8347
rect 16071 8313 16083 8347
rect 20070 8344 20076 8356
rect 20031 8316 20076 8344
rect 16025 8307 16083 8313
rect 13630 8276 13636 8288
rect 12299 8248 13636 8276
rect 12299 8245 12311 8248
rect 12253 8239 12311 8245
rect 13630 8236 13636 8248
rect 13688 8236 13694 8288
rect 15746 8236 15752 8288
rect 15804 8276 15810 8288
rect 16040 8276 16068 8307
rect 20070 8304 20076 8316
rect 20128 8304 20134 8356
rect 15804 8248 16068 8276
rect 15804 8236 15810 8248
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 2038 8072 2044 8084
rect 1999 8044 2044 8072
rect 2038 8032 2044 8044
rect 2096 8032 2102 8084
rect 3510 8072 3516 8084
rect 3471 8044 3516 8072
rect 3510 8032 3516 8044
rect 3568 8032 3574 8084
rect 3786 8072 3792 8084
rect 3747 8044 3792 8072
rect 3786 8032 3792 8044
rect 3844 8032 3850 8084
rect 6196 8044 8248 8072
rect 1765 8007 1823 8013
rect 1765 7973 1777 8007
rect 1811 8004 1823 8007
rect 1854 8004 1860 8016
rect 1811 7976 1860 8004
rect 1811 7973 1823 7976
rect 1765 7967 1823 7973
rect 1854 7964 1860 7976
rect 1912 8004 1918 8016
rect 2409 8007 2467 8013
rect 2409 8004 2421 8007
rect 1912 7976 2421 8004
rect 1912 7964 1918 7976
rect 2409 7973 2421 7976
rect 2455 8004 2467 8007
rect 2774 8004 2780 8016
rect 2455 7976 2780 8004
rect 2455 7973 2467 7976
rect 2409 7967 2467 7973
rect 2774 7964 2780 7976
rect 2832 7964 2838 8016
rect 2958 8004 2964 8016
rect 2919 7976 2964 8004
rect 2958 7964 2964 7976
rect 3016 8004 3022 8016
rect 4430 8004 4436 8016
rect 3016 7976 4436 8004
rect 3016 7964 3022 7976
rect 4430 7964 4436 7976
rect 4488 7964 4494 8016
rect 5442 7964 5448 8016
rect 5500 8004 5506 8016
rect 6196 8004 6224 8044
rect 5500 7976 6224 8004
rect 5500 7964 5506 7976
rect 4525 7939 4583 7945
rect 4525 7905 4537 7939
rect 4571 7936 4583 7939
rect 4706 7936 4712 7948
rect 4571 7908 4712 7936
rect 4571 7905 4583 7908
rect 4525 7899 4583 7905
rect 4706 7896 4712 7908
rect 4764 7936 4770 7948
rect 5258 7936 5264 7948
rect 4764 7908 5264 7936
rect 4764 7896 4770 7908
rect 5258 7896 5264 7908
rect 5316 7896 5322 7948
rect 5721 7939 5779 7945
rect 5721 7905 5733 7939
rect 5767 7905 5779 7939
rect 5994 7936 6000 7948
rect 5955 7908 6000 7936
rect 5721 7899 5779 7905
rect 2317 7871 2375 7877
rect 2317 7837 2329 7871
rect 2363 7868 2375 7871
rect 3142 7868 3148 7880
rect 2363 7840 3148 7868
rect 2363 7837 2375 7840
rect 2317 7831 2375 7837
rect 3142 7828 3148 7840
rect 3200 7828 3206 7880
rect 4614 7828 4620 7880
rect 4672 7868 4678 7880
rect 4893 7871 4951 7877
rect 4893 7868 4905 7871
rect 4672 7840 4905 7868
rect 4672 7828 4678 7840
rect 4893 7837 4905 7840
rect 4939 7868 4951 7871
rect 5166 7868 5172 7880
rect 4939 7840 5172 7868
rect 4939 7837 4951 7840
rect 4893 7831 4951 7837
rect 5166 7828 5172 7840
rect 5224 7868 5230 7880
rect 5736 7868 5764 7899
rect 5994 7896 6000 7908
rect 6052 7896 6058 7948
rect 6196 7945 6224 7976
rect 6181 7939 6239 7945
rect 6181 7905 6193 7939
rect 6227 7905 6239 7939
rect 7558 7936 7564 7948
rect 7519 7908 7564 7936
rect 6181 7899 6239 7905
rect 7558 7896 7564 7908
rect 7616 7896 7622 7948
rect 7745 7939 7803 7945
rect 7745 7905 7757 7939
rect 7791 7905 7803 7939
rect 7745 7899 7803 7905
rect 6454 7868 6460 7880
rect 5224 7840 5799 7868
rect 6415 7840 6460 7868
rect 5224 7828 5230 7840
rect 3418 7760 3424 7812
rect 3476 7800 3482 7812
rect 4062 7800 4068 7812
rect 3476 7772 4068 7800
rect 3476 7760 3482 7772
rect 4062 7760 4068 7772
rect 4120 7800 4126 7812
rect 5442 7800 5448 7812
rect 4120 7772 5448 7800
rect 4120 7760 4126 7772
rect 5442 7760 5448 7772
rect 5500 7760 5506 7812
rect 5771 7800 5799 7840
rect 6454 7828 6460 7840
rect 6512 7828 6518 7880
rect 7374 7868 7380 7880
rect 6932 7840 7380 7868
rect 5771 7772 6408 7800
rect 6380 7744 6408 7772
rect 6362 7692 6368 7744
rect 6420 7732 6426 7744
rect 6932 7741 6960 7840
rect 7374 7828 7380 7840
rect 7432 7868 7438 7880
rect 7760 7868 7788 7899
rect 7834 7896 7840 7948
rect 7892 7936 7898 7948
rect 8113 7939 8171 7945
rect 8113 7936 8125 7939
rect 7892 7908 8125 7936
rect 7892 7896 7898 7908
rect 8113 7905 8125 7908
rect 8159 7905 8171 7939
rect 8220 7936 8248 8044
rect 12342 8032 12348 8084
rect 12400 8072 12406 8084
rect 12713 8075 12771 8081
rect 12713 8072 12725 8075
rect 12400 8044 12725 8072
rect 12400 8032 12406 8044
rect 12713 8041 12725 8044
rect 12759 8041 12771 8075
rect 12713 8035 12771 8041
rect 14185 8075 14243 8081
rect 14185 8041 14197 8075
rect 14231 8072 14243 8075
rect 14231 8044 15516 8072
rect 14231 8041 14243 8044
rect 14185 8035 14243 8041
rect 15488 8016 15516 8044
rect 15930 8032 15936 8084
rect 15988 8072 15994 8084
rect 16393 8075 16451 8081
rect 16393 8072 16405 8075
rect 15988 8044 16405 8072
rect 15988 8032 15994 8044
rect 16393 8041 16405 8044
rect 16439 8072 16451 8075
rect 16482 8072 16488 8084
rect 16439 8044 16488 8072
rect 16439 8041 16451 8044
rect 16393 8035 16451 8041
rect 16482 8032 16488 8044
rect 16540 8032 16546 8084
rect 18506 8072 18512 8084
rect 18467 8044 18512 8072
rect 18506 8032 18512 8044
rect 18564 8032 18570 8084
rect 19981 8075 20039 8081
rect 19981 8041 19993 8075
rect 20027 8072 20039 8075
rect 20070 8072 20076 8084
rect 20027 8044 20076 8072
rect 20027 8041 20039 8044
rect 19981 8035 20039 8041
rect 20070 8032 20076 8044
rect 20128 8032 20134 8084
rect 9950 7964 9956 8016
rect 10008 8004 10014 8016
rect 11149 8007 11207 8013
rect 11149 8004 11161 8007
rect 10008 7976 11161 8004
rect 10008 7964 10014 7976
rect 11149 7973 11161 7976
rect 11195 7973 11207 8007
rect 11149 7967 11207 7973
rect 11422 7964 11428 8016
rect 11480 8004 11486 8016
rect 11517 8007 11575 8013
rect 11517 8004 11529 8007
rect 11480 7976 11529 8004
rect 11480 7964 11486 7976
rect 11517 7973 11529 7976
rect 11563 7973 11575 8007
rect 11517 7967 11575 7973
rect 11790 7964 11796 8016
rect 11848 8004 11854 8016
rect 13630 8013 13636 8016
rect 12437 8007 12495 8013
rect 12437 8004 12449 8007
rect 11848 7976 12449 8004
rect 11848 7964 11854 7976
rect 12437 7973 12449 7976
rect 12483 7973 12495 8007
rect 13627 8004 13636 8013
rect 13543 7976 13636 8004
rect 12437 7967 12495 7973
rect 13627 7967 13636 7976
rect 13688 8004 13694 8016
rect 13998 8004 14004 8016
rect 13688 7976 14004 8004
rect 13630 7964 13636 7967
rect 13688 7964 13694 7976
rect 13998 7964 14004 7976
rect 14056 7964 14062 8016
rect 15378 8004 15384 8016
rect 15339 7976 15384 8004
rect 15378 7964 15384 7976
rect 15436 7964 15442 8016
rect 15470 7964 15476 8016
rect 15528 8004 15534 8016
rect 15528 7976 15621 8004
rect 15528 7964 15534 7976
rect 8481 7939 8539 7945
rect 8481 7936 8493 7939
rect 8220 7908 8493 7936
rect 8113 7899 8171 7905
rect 8481 7905 8493 7908
rect 8527 7936 8539 7939
rect 8846 7936 8852 7948
rect 8527 7908 8852 7936
rect 8527 7905 8539 7908
rect 8481 7899 8539 7905
rect 8846 7896 8852 7908
rect 8904 7896 8910 7948
rect 10413 7939 10471 7945
rect 10413 7905 10425 7939
rect 10459 7936 10471 7939
rect 10962 7936 10968 7948
rect 10459 7908 10968 7936
rect 10459 7905 10471 7908
rect 10413 7899 10471 7905
rect 10962 7896 10968 7908
rect 11020 7896 11026 7948
rect 13265 7939 13323 7945
rect 13265 7936 13277 7939
rect 12906 7908 13277 7936
rect 7432 7840 7788 7868
rect 7432 7828 7438 7840
rect 11146 7828 11152 7880
rect 11204 7868 11210 7880
rect 11425 7871 11483 7877
rect 11425 7868 11437 7871
rect 11204 7840 11437 7868
rect 11204 7828 11210 7840
rect 11425 7837 11437 7840
rect 11471 7837 11483 7871
rect 11425 7831 11483 7837
rect 12069 7871 12127 7877
rect 12069 7837 12081 7871
rect 12115 7868 12127 7871
rect 12802 7868 12808 7880
rect 12115 7840 12808 7868
rect 12115 7837 12127 7840
rect 12069 7831 12127 7837
rect 12802 7828 12808 7840
rect 12860 7828 12866 7880
rect 8665 7803 8723 7809
rect 8665 7769 8677 7803
rect 8711 7800 8723 7803
rect 12906 7800 12934 7908
rect 13265 7905 13277 7908
rect 13311 7936 13323 7939
rect 13814 7936 13820 7948
rect 13311 7908 13820 7936
rect 13311 7905 13323 7908
rect 13265 7899 13323 7905
rect 13814 7896 13820 7908
rect 13872 7896 13878 7948
rect 16850 7936 16856 7948
rect 16811 7908 16856 7936
rect 16850 7896 16856 7908
rect 16908 7896 16914 7948
rect 16298 7828 16304 7880
rect 16356 7868 16362 7880
rect 17957 7871 18015 7877
rect 17957 7868 17969 7871
rect 16356 7840 17969 7868
rect 16356 7828 16362 7840
rect 17957 7837 17969 7840
rect 18003 7837 18015 7871
rect 17957 7831 18015 7837
rect 14366 7800 14372 7812
rect 8711 7772 12934 7800
rect 13786 7772 14372 7800
rect 8711 7769 8723 7772
rect 8665 7763 8723 7769
rect 6917 7735 6975 7741
rect 6917 7732 6929 7735
rect 6420 7704 6929 7732
rect 6420 7692 6426 7704
rect 6917 7701 6929 7704
rect 6963 7701 6975 7735
rect 6917 7695 6975 7701
rect 9125 7735 9183 7741
rect 9125 7701 9137 7735
rect 9171 7732 9183 7735
rect 9214 7732 9220 7744
rect 9171 7704 9220 7732
rect 9171 7701 9183 7704
rect 9125 7695 9183 7701
rect 9214 7692 9220 7704
rect 9272 7732 9278 7744
rect 9401 7735 9459 7741
rect 9401 7732 9413 7735
rect 9272 7704 9413 7732
rect 9272 7692 9278 7704
rect 9401 7701 9413 7704
rect 9447 7701 9459 7735
rect 10042 7732 10048 7744
rect 10003 7704 10048 7732
rect 9401 7695 9459 7701
rect 10042 7692 10048 7704
rect 10100 7692 10106 7744
rect 10873 7735 10931 7741
rect 10873 7701 10885 7735
rect 10919 7732 10931 7735
rect 10962 7732 10968 7744
rect 10919 7704 10968 7732
rect 10919 7701 10931 7704
rect 10873 7695 10931 7701
rect 10962 7692 10968 7704
rect 11020 7692 11026 7744
rect 12526 7692 12532 7744
rect 12584 7732 12590 7744
rect 13786 7732 13814 7772
rect 14366 7760 14372 7772
rect 14424 7800 14430 7812
rect 14461 7803 14519 7809
rect 14461 7800 14473 7803
rect 14424 7772 14473 7800
rect 14424 7760 14430 7772
rect 14461 7769 14473 7772
rect 14507 7769 14519 7803
rect 15930 7800 15936 7812
rect 15891 7772 15936 7800
rect 14461 7763 14519 7769
rect 15930 7760 15936 7772
rect 15988 7760 15994 7812
rect 12584 7704 13814 7732
rect 17037 7735 17095 7741
rect 12584 7692 12590 7704
rect 17037 7701 17049 7735
rect 17083 7732 17095 7735
rect 18138 7732 18144 7744
rect 17083 7704 18144 7732
rect 17083 7701 17095 7704
rect 17037 7695 17095 7701
rect 18138 7692 18144 7704
rect 18196 7692 18202 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 2774 7528 2780 7540
rect 2735 7500 2780 7528
rect 2774 7488 2780 7500
rect 2832 7488 2838 7540
rect 3510 7488 3516 7540
rect 3568 7528 3574 7540
rect 4154 7528 4160 7540
rect 3568 7500 4160 7528
rect 3568 7488 3574 7500
rect 4154 7488 4160 7500
rect 4212 7488 4218 7540
rect 4614 7528 4620 7540
rect 4575 7500 4620 7528
rect 4614 7488 4620 7500
rect 4672 7488 4678 7540
rect 5258 7488 5264 7540
rect 5316 7528 5322 7540
rect 5537 7531 5595 7537
rect 5537 7528 5549 7531
rect 5316 7500 5549 7528
rect 5316 7488 5322 7500
rect 5537 7497 5549 7500
rect 5583 7497 5595 7531
rect 5537 7491 5595 7497
rect 5905 7531 5963 7537
rect 5905 7497 5917 7531
rect 5951 7528 5963 7531
rect 6546 7528 6552 7540
rect 5951 7500 6552 7528
rect 5951 7497 5963 7500
rect 5905 7491 5963 7497
rect 6546 7488 6552 7500
rect 6604 7488 6610 7540
rect 6963 7531 7021 7537
rect 6963 7497 6975 7531
rect 7009 7528 7021 7531
rect 9950 7528 9956 7540
rect 7009 7500 9956 7528
rect 7009 7497 7021 7500
rect 6963 7491 7021 7497
rect 9950 7488 9956 7500
rect 10008 7488 10014 7540
rect 10962 7488 10968 7540
rect 11020 7528 11026 7540
rect 11333 7531 11391 7537
rect 11333 7528 11345 7531
rect 11020 7500 11345 7528
rect 11020 7488 11026 7500
rect 11333 7497 11345 7500
rect 11379 7497 11391 7531
rect 11698 7528 11704 7540
rect 11659 7500 11704 7528
rect 11333 7491 11391 7497
rect 11698 7488 11704 7500
rect 11756 7488 11762 7540
rect 13446 7488 13452 7540
rect 13504 7528 13510 7540
rect 14139 7531 14197 7537
rect 14139 7528 14151 7531
rect 13504 7500 14151 7528
rect 13504 7488 13510 7500
rect 14139 7497 14151 7500
rect 14185 7497 14197 7531
rect 16298 7528 16304 7540
rect 16259 7500 16304 7528
rect 14139 7491 14197 7497
rect 16298 7488 16304 7500
rect 16356 7488 16362 7540
rect 18598 7528 18604 7540
rect 18559 7500 18604 7528
rect 18598 7488 18604 7500
rect 18656 7488 18662 7540
rect 3881 7463 3939 7469
rect 3881 7429 3893 7463
rect 3927 7460 3939 7463
rect 4338 7460 4344 7472
rect 3927 7432 4344 7460
rect 3927 7429 3939 7432
rect 3881 7423 3939 7429
rect 4338 7420 4344 7432
rect 4396 7420 4402 7472
rect 6564 7460 6592 7488
rect 7653 7463 7711 7469
rect 7653 7460 7665 7463
rect 6564 7432 7665 7460
rect 7653 7429 7665 7432
rect 7699 7460 7711 7463
rect 7834 7460 7840 7472
rect 7699 7432 7840 7460
rect 7699 7429 7711 7432
rect 7653 7423 7711 7429
rect 7834 7420 7840 7432
rect 7892 7420 7898 7472
rect 9214 7460 9220 7472
rect 8036 7432 9220 7460
rect 1946 7352 1952 7404
rect 2004 7392 2010 7404
rect 2409 7395 2467 7401
rect 2409 7392 2421 7395
rect 2004 7364 2421 7392
rect 2004 7352 2010 7364
rect 2409 7361 2421 7364
rect 2455 7392 2467 7395
rect 3970 7392 3976 7404
rect 2455 7364 3976 7392
rect 2455 7361 2467 7364
rect 2409 7355 2467 7361
rect 3970 7352 3976 7364
rect 4028 7352 4034 7404
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7392 7435 7395
rect 7742 7392 7748 7404
rect 7423 7364 7748 7392
rect 7423 7361 7435 7364
rect 7377 7355 7435 7361
rect 2317 7327 2375 7333
rect 2317 7293 2329 7327
rect 2363 7324 2375 7327
rect 2774 7324 2780 7336
rect 2363 7296 2780 7324
rect 2363 7293 2375 7296
rect 2317 7287 2375 7293
rect 2774 7284 2780 7296
rect 2832 7284 2838 7336
rect 3697 7327 3755 7333
rect 3697 7293 3709 7327
rect 3743 7324 3755 7327
rect 4706 7324 4712 7336
rect 3743 7296 4154 7324
rect 4619 7296 4712 7324
rect 3743 7293 3755 7296
rect 3697 7287 3755 7293
rect 4126 7256 4154 7296
rect 4706 7284 4712 7296
rect 4764 7324 4770 7336
rect 5169 7327 5227 7333
rect 5169 7324 5181 7327
rect 4764 7296 5181 7324
rect 4764 7284 4770 7296
rect 5169 7293 5181 7296
rect 5215 7293 5227 7327
rect 5169 7287 5227 7293
rect 5350 7284 5356 7336
rect 5408 7324 5414 7336
rect 5721 7327 5779 7333
rect 5721 7324 5733 7327
rect 5408 7296 5733 7324
rect 5408 7284 5414 7296
rect 5721 7293 5733 7296
rect 5767 7324 5779 7327
rect 6181 7327 6239 7333
rect 6181 7324 6193 7327
rect 5767 7296 6193 7324
rect 5767 7293 5779 7296
rect 5721 7287 5779 7293
rect 6181 7293 6193 7296
rect 6227 7293 6239 7327
rect 6181 7287 6239 7293
rect 6892 7327 6950 7333
rect 6892 7293 6904 7327
rect 6938 7324 6950 7327
rect 7392 7324 7420 7355
rect 7742 7352 7748 7364
rect 7800 7352 7806 7404
rect 6938 7296 7420 7324
rect 6938 7293 6950 7296
rect 6892 7287 6950 7293
rect 7558 7284 7564 7336
rect 7616 7324 7622 7336
rect 8036 7333 8064 7432
rect 9214 7420 9220 7432
rect 9272 7420 9278 7472
rect 13814 7460 13820 7472
rect 13775 7432 13820 7460
rect 13814 7420 13820 7432
rect 13872 7420 13878 7472
rect 16316 7460 16344 7488
rect 16850 7460 16856 7472
rect 15304 7432 16344 7460
rect 16809 7432 16856 7460
rect 9398 7352 9404 7404
rect 9456 7392 9462 7404
rect 10137 7395 10195 7401
rect 10137 7392 10149 7395
rect 9456 7364 10149 7392
rect 9456 7352 9462 7364
rect 10137 7361 10149 7364
rect 10183 7392 10195 7395
rect 10778 7392 10784 7404
rect 10183 7364 10784 7392
rect 10183 7361 10195 7364
rect 10137 7355 10195 7361
rect 10778 7352 10784 7364
rect 10836 7352 10842 7404
rect 12802 7392 12808 7404
rect 12763 7364 12808 7392
rect 12802 7352 12808 7364
rect 12860 7352 12866 7404
rect 15304 7401 15332 7432
rect 16850 7420 16856 7432
rect 16908 7469 16914 7472
rect 16908 7463 16957 7469
rect 16908 7429 16911 7463
rect 16945 7460 16957 7463
rect 17589 7463 17647 7469
rect 17589 7460 17601 7463
rect 16945 7432 17601 7460
rect 16945 7429 16957 7432
rect 16908 7423 16957 7429
rect 17589 7429 17601 7432
rect 17635 7429 17647 7463
rect 17589 7423 17647 7429
rect 16908 7420 16914 7423
rect 15289 7395 15347 7401
rect 15289 7361 15301 7395
rect 15335 7361 15347 7395
rect 15930 7392 15936 7404
rect 15891 7364 15936 7392
rect 15289 7355 15347 7361
rect 15930 7352 15936 7364
rect 15988 7352 15994 7404
rect 8021 7327 8079 7333
rect 8021 7324 8033 7327
rect 7616 7296 8033 7324
rect 7616 7284 7622 7296
rect 8021 7293 8033 7296
rect 8067 7293 8079 7327
rect 8386 7324 8392 7336
rect 8347 7296 8392 7324
rect 8021 7287 8079 7293
rect 8386 7284 8392 7296
rect 8444 7284 8450 7336
rect 8849 7327 8907 7333
rect 8849 7293 8861 7327
rect 8895 7293 8907 7327
rect 9122 7324 9128 7336
rect 9083 7296 9128 7324
rect 8849 7287 8907 7293
rect 4249 7259 4307 7265
rect 4249 7256 4261 7259
rect 4126 7228 4261 7256
rect 4249 7225 4261 7228
rect 4295 7256 4307 7259
rect 5074 7256 5080 7268
rect 4295 7228 5080 7256
rect 4295 7225 4307 7228
rect 4249 7219 4307 7225
rect 5074 7216 5080 7228
rect 5132 7216 5138 7268
rect 8864 7256 8892 7287
rect 9122 7284 9128 7296
rect 9180 7284 9186 7336
rect 11057 7327 11115 7333
rect 11057 7293 11069 7327
rect 11103 7324 11115 7327
rect 11422 7324 11428 7336
rect 11103 7296 11428 7324
rect 11103 7293 11115 7296
rect 11057 7287 11115 7293
rect 11422 7284 11428 7296
rect 11480 7284 11486 7336
rect 13538 7284 13544 7336
rect 13596 7324 13602 7336
rect 14068 7327 14126 7333
rect 14068 7324 14080 7327
rect 13596 7296 14080 7324
rect 13596 7284 13602 7296
rect 14068 7293 14080 7296
rect 14114 7324 14126 7327
rect 14461 7327 14519 7333
rect 14461 7324 14473 7327
rect 14114 7296 14473 7324
rect 14114 7293 14126 7296
rect 14068 7287 14126 7293
rect 14461 7293 14473 7296
rect 14507 7293 14519 7327
rect 14461 7287 14519 7293
rect 16114 7284 16120 7336
rect 16172 7324 16178 7336
rect 16796 7327 16854 7333
rect 16796 7324 16808 7327
rect 16172 7296 16808 7324
rect 16172 7284 16178 7296
rect 16796 7293 16808 7296
rect 16842 7324 16854 7327
rect 17221 7327 17279 7333
rect 17221 7324 17233 7327
rect 16842 7296 17233 7324
rect 16842 7293 16854 7296
rect 16796 7287 16854 7293
rect 17221 7293 17233 7296
rect 17267 7293 17279 7327
rect 17221 7287 17279 7293
rect 18100 7327 18158 7333
rect 18100 7293 18112 7327
rect 18146 7324 18158 7327
rect 18598 7324 18604 7336
rect 18146 7296 18604 7324
rect 18146 7293 18158 7296
rect 18100 7287 18158 7293
rect 18598 7284 18604 7296
rect 18656 7284 18662 7336
rect 24648 7327 24706 7333
rect 24648 7293 24660 7327
rect 24694 7324 24706 7327
rect 24694 7296 25176 7324
rect 24694 7293 24706 7296
rect 24648 7287 24706 7293
rect 9306 7256 9312 7268
rect 5368 7228 8892 7256
rect 9267 7228 9312 7256
rect 3142 7188 3148 7200
rect 3103 7160 3148 7188
rect 3142 7148 3148 7160
rect 3200 7148 3206 7200
rect 3510 7188 3516 7200
rect 3471 7160 3516 7188
rect 3510 7148 3516 7160
rect 3568 7148 3574 7200
rect 4893 7191 4951 7197
rect 4893 7157 4905 7191
rect 4939 7188 4951 7191
rect 5368 7188 5396 7228
rect 4939 7160 5396 7188
rect 4939 7157 4951 7160
rect 4893 7151 4951 7157
rect 6362 7148 6368 7200
rect 6420 7188 6426 7200
rect 6549 7191 6607 7197
rect 6549 7188 6561 7191
rect 6420 7160 6561 7188
rect 6420 7148 6426 7160
rect 6549 7157 6561 7160
rect 6595 7157 6607 7191
rect 8864 7188 8892 7228
rect 9306 7216 9312 7228
rect 9364 7216 9370 7268
rect 10458 7259 10516 7265
rect 10458 7256 10470 7259
rect 9968 7228 10470 7256
rect 9968 7200 9996 7228
rect 10458 7225 10470 7228
rect 10504 7225 10516 7259
rect 10458 7219 10516 7225
rect 12529 7259 12587 7265
rect 12529 7225 12541 7259
rect 12575 7225 12587 7259
rect 12529 7219 12587 7225
rect 9582 7188 9588 7200
rect 8864 7160 9588 7188
rect 6549 7151 6607 7157
rect 9582 7148 9588 7160
rect 9640 7148 9646 7200
rect 9950 7188 9956 7200
rect 9911 7160 9956 7188
rect 9950 7148 9956 7160
rect 10008 7148 10014 7200
rect 12158 7188 12164 7200
rect 12119 7160 12164 7188
rect 12158 7148 12164 7160
rect 12216 7148 12222 7200
rect 12434 7148 12440 7200
rect 12492 7188 12498 7200
rect 12544 7188 12572 7219
rect 12618 7216 12624 7268
rect 12676 7256 12682 7268
rect 12676 7228 12721 7256
rect 12676 7216 12682 7228
rect 15378 7216 15384 7268
rect 15436 7256 15442 7268
rect 15436 7228 15481 7256
rect 15436 7216 15442 7228
rect 16942 7216 16948 7268
rect 17000 7256 17006 7268
rect 18187 7259 18245 7265
rect 18187 7256 18199 7259
rect 17000 7228 18199 7256
rect 17000 7216 17006 7228
rect 18187 7225 18199 7228
rect 18233 7225 18245 7259
rect 18187 7219 18245 7225
rect 13446 7188 13452 7200
rect 12492 7160 12572 7188
rect 13407 7160 13452 7188
rect 12492 7148 12498 7160
rect 13446 7148 13452 7160
rect 13504 7148 13510 7200
rect 15105 7191 15163 7197
rect 15105 7157 15117 7191
rect 15151 7188 15163 7191
rect 15396 7188 15424 7216
rect 25148 7200 25176 7296
rect 15151 7160 15424 7188
rect 15151 7157 15163 7160
rect 15105 7151 15163 7157
rect 15470 7148 15476 7200
rect 15528 7188 15534 7200
rect 16577 7191 16635 7197
rect 16577 7188 16589 7191
rect 15528 7160 16589 7188
rect 15528 7148 15534 7160
rect 16577 7157 16589 7160
rect 16623 7157 16635 7191
rect 16577 7151 16635 7157
rect 18598 7148 18604 7200
rect 18656 7188 18662 7200
rect 24719 7191 24777 7197
rect 24719 7188 24731 7191
rect 18656 7160 24731 7188
rect 18656 7148 18662 7160
rect 24719 7157 24731 7160
rect 24765 7157 24777 7191
rect 25130 7188 25136 7200
rect 25091 7160 25136 7188
rect 24719 7151 24777 7157
rect 25130 7148 25136 7160
rect 25188 7148 25194 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 1397 6987 1455 6993
rect 1397 6953 1409 6987
rect 1443 6984 1455 6987
rect 3510 6984 3516 6996
rect 1443 6956 3516 6984
rect 1443 6953 1455 6956
rect 1397 6947 1455 6953
rect 3510 6944 3516 6956
rect 3568 6944 3574 6996
rect 4062 6944 4068 6996
rect 4120 6984 4126 6996
rect 4249 6987 4307 6993
rect 4249 6984 4261 6987
rect 4120 6956 4261 6984
rect 4120 6944 4126 6956
rect 4249 6953 4261 6956
rect 4295 6953 4307 6987
rect 6638 6984 6644 6996
rect 6599 6956 6644 6984
rect 4249 6947 4307 6953
rect 6638 6944 6644 6956
rect 6696 6944 6702 6996
rect 8386 6944 8392 6996
rect 8444 6984 8450 6996
rect 8481 6987 8539 6993
rect 8481 6984 8493 6987
rect 8444 6956 8493 6984
rect 8444 6944 8450 6956
rect 8481 6953 8493 6956
rect 8527 6953 8539 6987
rect 8846 6984 8852 6996
rect 8807 6956 8852 6984
rect 8481 6947 8539 6953
rect 8846 6944 8852 6956
rect 8904 6944 8910 6996
rect 9214 6984 9220 6996
rect 9175 6956 9220 6984
rect 9214 6944 9220 6956
rect 9272 6944 9278 6996
rect 9950 6944 9956 6996
rect 10008 6984 10014 6996
rect 10045 6987 10103 6993
rect 10045 6984 10057 6987
rect 10008 6956 10057 6984
rect 10008 6944 10014 6956
rect 10045 6953 10057 6956
rect 10091 6953 10103 6987
rect 10045 6947 10103 6953
rect 10597 6987 10655 6993
rect 10597 6953 10609 6987
rect 10643 6984 10655 6987
rect 10962 6984 10968 6996
rect 10643 6956 10968 6984
rect 10643 6953 10655 6956
rect 10597 6947 10655 6953
rect 10962 6944 10968 6956
rect 11020 6944 11026 6996
rect 11146 6944 11152 6996
rect 11204 6984 11210 6996
rect 12805 6987 12863 6993
rect 12805 6984 12817 6987
rect 11204 6956 12817 6984
rect 11204 6944 11210 6956
rect 12805 6953 12817 6956
rect 12851 6953 12863 6987
rect 12805 6947 12863 6953
rect 13078 6944 13084 6996
rect 13136 6984 13142 6996
rect 13449 6987 13507 6993
rect 13449 6984 13461 6987
rect 13136 6956 13461 6984
rect 13136 6944 13142 6956
rect 13449 6953 13461 6956
rect 13495 6953 13507 6987
rect 13449 6947 13507 6953
rect 15105 6987 15163 6993
rect 15105 6953 15117 6987
rect 15151 6984 15163 6987
rect 15286 6984 15292 6996
rect 15151 6956 15292 6984
rect 15151 6953 15163 6956
rect 15105 6947 15163 6953
rect 15286 6944 15292 6956
rect 15344 6944 15350 6996
rect 15378 6944 15384 6996
rect 15436 6984 15442 6996
rect 15565 6987 15623 6993
rect 15565 6984 15577 6987
rect 15436 6956 15577 6984
rect 15436 6944 15442 6956
rect 15565 6953 15577 6956
rect 15611 6953 15623 6987
rect 24762 6984 24768 6996
rect 24723 6956 24768 6984
rect 15565 6947 15623 6953
rect 24762 6944 24768 6956
rect 24820 6944 24826 6996
rect 1854 6916 1860 6928
rect 1815 6888 1860 6916
rect 1854 6876 1860 6888
rect 1912 6876 1918 6928
rect 2317 6919 2375 6925
rect 2317 6885 2329 6919
rect 2363 6916 2375 6919
rect 2958 6916 2964 6928
rect 2363 6888 2964 6916
rect 2363 6885 2375 6888
rect 2317 6879 2375 6885
rect 2958 6876 2964 6888
rect 3016 6876 3022 6928
rect 3145 6919 3203 6925
rect 3145 6885 3157 6919
rect 3191 6916 3203 6919
rect 4706 6916 4712 6928
rect 3191 6888 4712 6916
rect 3191 6885 3203 6888
rect 3145 6879 3203 6885
rect 4706 6876 4712 6888
rect 4764 6876 4770 6928
rect 5534 6916 5540 6928
rect 5495 6888 5540 6916
rect 5534 6876 5540 6888
rect 5592 6916 5598 6928
rect 6730 6916 6736 6928
rect 5592 6888 6736 6916
rect 5592 6876 5598 6888
rect 2409 6851 2467 6857
rect 2409 6817 2421 6851
rect 2455 6848 2467 6851
rect 2590 6848 2596 6860
rect 2455 6820 2596 6848
rect 2455 6817 2467 6820
rect 2409 6811 2467 6817
rect 2590 6808 2596 6820
rect 2648 6808 2654 6860
rect 2685 6851 2743 6857
rect 2685 6817 2697 6851
rect 2731 6848 2743 6851
rect 2774 6848 2780 6860
rect 2731 6820 2780 6848
rect 2731 6817 2743 6820
rect 2685 6811 2743 6817
rect 2774 6808 2780 6820
rect 2832 6808 2838 6860
rect 4522 6808 4528 6860
rect 4580 6848 4586 6860
rect 6380 6857 6408 6888
rect 6730 6876 6736 6888
rect 6788 6876 6794 6928
rect 7742 6916 7748 6928
rect 7116 6888 7748 6916
rect 4893 6851 4951 6857
rect 4893 6848 4905 6851
rect 4580 6820 4905 6848
rect 4580 6808 4586 6820
rect 4893 6817 4905 6820
rect 4939 6817 4951 6851
rect 4893 6811 4951 6817
rect 6365 6851 6423 6857
rect 6365 6817 6377 6851
rect 6411 6817 6423 6851
rect 6365 6811 6423 6817
rect 6546 6808 6552 6860
rect 6604 6848 6610 6860
rect 7116 6857 7144 6888
rect 7742 6876 7748 6888
rect 7800 6916 7806 6928
rect 8404 6916 8432 6944
rect 7800 6888 8432 6916
rect 7800 6876 7806 6888
rect 10778 6876 10784 6928
rect 10836 6916 10842 6928
rect 10873 6919 10931 6925
rect 10873 6916 10885 6919
rect 10836 6888 10885 6916
rect 10836 6876 10842 6888
rect 10873 6885 10885 6888
rect 10919 6885 10931 6919
rect 12158 6916 12164 6928
rect 12119 6888 12164 6916
rect 10873 6879 10931 6885
rect 12158 6876 12164 6888
rect 12216 6916 12222 6928
rect 12618 6916 12624 6928
rect 12216 6888 12624 6916
rect 12216 6876 12222 6888
rect 12618 6876 12624 6888
rect 12676 6876 12682 6928
rect 7101 6851 7159 6857
rect 7101 6848 7113 6851
rect 6604 6820 7113 6848
rect 6604 6808 6610 6820
rect 7101 6817 7113 6820
rect 7147 6817 7159 6851
rect 7101 6811 7159 6817
rect 7193 6851 7251 6857
rect 7193 6817 7205 6851
rect 7239 6817 7251 6851
rect 7193 6811 7251 6817
rect 7208 6780 7236 6811
rect 7282 6808 7288 6860
rect 7340 6848 7346 6860
rect 7653 6851 7711 6857
rect 7653 6848 7665 6851
rect 7340 6820 7665 6848
rect 7340 6808 7346 6820
rect 7653 6817 7665 6820
rect 7699 6848 7711 6851
rect 8205 6851 8263 6857
rect 8205 6848 8217 6851
rect 7699 6820 8217 6848
rect 7699 6817 7711 6820
rect 7653 6811 7711 6817
rect 8205 6817 8217 6820
rect 8251 6848 8263 6851
rect 9122 6848 9128 6860
rect 8251 6820 9128 6848
rect 8251 6817 8263 6820
rect 8205 6811 8263 6817
rect 9122 6808 9128 6820
rect 9180 6808 9186 6860
rect 11422 6808 11428 6860
rect 11480 6848 11486 6860
rect 11517 6851 11575 6857
rect 11517 6848 11529 6851
rect 11480 6820 11529 6848
rect 11480 6808 11486 6820
rect 11517 6817 11529 6820
rect 11563 6817 11575 6851
rect 12986 6848 12992 6860
rect 12947 6820 12992 6848
rect 11517 6811 11575 6817
rect 12986 6808 12992 6820
rect 13044 6808 13050 6860
rect 13262 6848 13268 6860
rect 13223 6820 13268 6848
rect 13262 6808 13268 6820
rect 13320 6808 13326 6860
rect 15470 6848 15476 6860
rect 15431 6820 15476 6848
rect 15470 6808 15476 6820
rect 15528 6808 15534 6860
rect 15930 6808 15936 6860
rect 15988 6848 15994 6860
rect 16850 6848 16856 6860
rect 16908 6857 16914 6860
rect 16908 6851 16946 6857
rect 15988 6820 16856 6848
rect 15988 6808 15994 6820
rect 16850 6808 16856 6820
rect 16934 6817 16946 6851
rect 16908 6811 16946 6817
rect 24581 6851 24639 6857
rect 24581 6817 24593 6851
rect 24627 6848 24639 6851
rect 24670 6848 24676 6860
rect 24627 6820 24676 6848
rect 24627 6817 24639 6820
rect 24581 6811 24639 6817
rect 16908 6808 16914 6811
rect 24670 6808 24676 6820
rect 24728 6808 24734 6860
rect 8110 6780 8116 6792
rect 6196 6752 8116 6780
rect 2501 6715 2559 6721
rect 2501 6681 2513 6715
rect 2547 6681 2559 6715
rect 2501 6675 2559 6681
rect 2516 6644 2544 6675
rect 3234 6644 3240 6656
rect 2516 6616 3240 6644
rect 3234 6604 3240 6616
rect 3292 6644 3298 6656
rect 3421 6647 3479 6653
rect 3421 6644 3433 6647
rect 3292 6616 3433 6644
rect 3292 6604 3298 6616
rect 3421 6613 3433 6616
rect 3467 6613 3479 6647
rect 4614 6644 4620 6656
rect 4575 6616 4620 6644
rect 3421 6607 3479 6613
rect 4614 6604 4620 6616
rect 4672 6604 4678 6656
rect 5534 6604 5540 6656
rect 5592 6644 5598 6656
rect 5813 6647 5871 6653
rect 5813 6644 5825 6647
rect 5592 6616 5825 6644
rect 5592 6604 5598 6616
rect 5813 6613 5825 6616
rect 5859 6644 5871 6647
rect 5994 6644 6000 6656
rect 5859 6616 6000 6644
rect 5859 6613 5871 6616
rect 5813 6607 5871 6613
rect 5994 6604 6000 6616
rect 6052 6644 6058 6656
rect 6196 6653 6224 6752
rect 8110 6740 8116 6752
rect 8168 6740 8174 6792
rect 9306 6740 9312 6792
rect 9364 6780 9370 6792
rect 9677 6783 9735 6789
rect 9677 6780 9689 6783
rect 9364 6752 9689 6780
rect 9364 6740 9370 6752
rect 9677 6749 9689 6752
rect 9723 6780 9735 6783
rect 11238 6780 11244 6792
rect 9723 6752 11244 6780
rect 9723 6749 9735 6752
rect 9677 6743 9735 6749
rect 11238 6740 11244 6752
rect 11296 6740 11302 6792
rect 11698 6740 11704 6792
rect 11756 6780 11762 6792
rect 13081 6783 13139 6789
rect 13081 6780 13093 6783
rect 11756 6752 13093 6780
rect 11756 6740 11762 6752
rect 13081 6749 13093 6752
rect 13127 6749 13139 6783
rect 13081 6743 13139 6749
rect 13096 6712 13124 6743
rect 13998 6712 14004 6724
rect 13096 6684 14004 6712
rect 13998 6672 14004 6684
rect 14056 6672 14062 6724
rect 6181 6647 6239 6653
rect 6181 6644 6193 6647
rect 6052 6616 6193 6644
rect 6052 6604 6058 6616
rect 6181 6613 6193 6616
rect 6227 6613 6239 6647
rect 6181 6607 6239 6613
rect 11333 6647 11391 6653
rect 11333 6613 11345 6647
rect 11379 6644 11391 6647
rect 11422 6644 11428 6656
rect 11379 6616 11428 6644
rect 11379 6613 11391 6616
rect 11333 6607 11391 6613
rect 11422 6604 11428 6616
rect 11480 6604 11486 6656
rect 12434 6644 12440 6656
rect 12395 6616 12440 6644
rect 12434 6604 12440 6616
rect 12492 6604 12498 6656
rect 14277 6647 14335 6653
rect 14277 6613 14289 6647
rect 14323 6644 14335 6647
rect 14458 6644 14464 6656
rect 14323 6616 14464 6644
rect 14323 6613 14335 6616
rect 14277 6607 14335 6613
rect 14458 6604 14464 6616
rect 14516 6604 14522 6656
rect 16991 6647 17049 6653
rect 16991 6613 17003 6647
rect 17037 6644 17049 6647
rect 18046 6644 18052 6656
rect 17037 6616 18052 6644
rect 17037 6613 17049 6616
rect 16991 6607 17049 6613
rect 18046 6604 18052 6616
rect 18104 6604 18110 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 1578 6440 1584 6452
rect 1539 6412 1584 6440
rect 1578 6400 1584 6412
rect 1636 6400 1642 6452
rect 5994 6400 6000 6452
rect 6052 6440 6058 6452
rect 6089 6443 6147 6449
rect 6089 6440 6101 6443
rect 6052 6412 6101 6440
rect 6052 6400 6058 6412
rect 6089 6409 6101 6412
rect 6135 6440 6147 6443
rect 6546 6440 6552 6452
rect 6135 6412 6552 6440
rect 6135 6409 6147 6412
rect 6089 6403 6147 6409
rect 6546 6400 6552 6412
rect 6604 6400 6610 6452
rect 10042 6440 10048 6452
rect 10003 6412 10048 6440
rect 10042 6400 10048 6412
rect 10100 6400 10106 6452
rect 11238 6440 11244 6452
rect 11199 6412 11244 6440
rect 11238 6400 11244 6412
rect 11296 6400 11302 6452
rect 13998 6440 14004 6452
rect 13959 6412 14004 6440
rect 13998 6400 14004 6412
rect 14056 6400 14062 6452
rect 15381 6443 15439 6449
rect 15381 6409 15393 6443
rect 15427 6440 15439 6443
rect 15470 6440 15476 6452
rect 15427 6412 15476 6440
rect 15427 6409 15439 6412
rect 15381 6403 15439 6409
rect 15470 6400 15476 6412
rect 15528 6400 15534 6452
rect 16850 6440 16856 6452
rect 16811 6412 16856 6440
rect 16850 6400 16856 6412
rect 16908 6400 16914 6452
rect 23842 6400 23848 6452
rect 23900 6440 23906 6452
rect 23937 6443 23995 6449
rect 23937 6440 23949 6443
rect 23900 6412 23949 6440
rect 23900 6400 23906 6412
rect 23937 6409 23949 6412
rect 23983 6409 23995 6443
rect 23937 6403 23995 6409
rect 3326 6332 3332 6384
rect 3384 6372 3390 6384
rect 4522 6372 4528 6384
rect 3384 6344 4528 6372
rect 3384 6332 3390 6344
rect 4522 6332 4528 6344
rect 4580 6372 4586 6384
rect 5629 6375 5687 6381
rect 5629 6372 5641 6375
rect 4580 6344 5641 6372
rect 4580 6332 4586 6344
rect 5629 6341 5641 6344
rect 5675 6341 5687 6375
rect 5629 6335 5687 6341
rect 6454 6332 6460 6384
rect 6512 6372 6518 6384
rect 11793 6375 11851 6381
rect 11793 6372 11805 6375
rect 6512 6344 11805 6372
rect 6512 6332 6518 6344
rect 11793 6341 11805 6344
rect 11839 6341 11851 6375
rect 11793 6335 11851 6341
rect 3418 6304 3424 6316
rect 3331 6276 3424 6304
rect 1302 6196 1308 6248
rect 1360 6236 1366 6248
rect 1397 6239 1455 6245
rect 1397 6236 1409 6239
rect 1360 6208 1409 6236
rect 1360 6196 1366 6208
rect 1397 6205 1409 6208
rect 1443 6236 1455 6239
rect 1949 6239 2007 6245
rect 1949 6236 1961 6239
rect 1443 6208 1961 6236
rect 1443 6205 1455 6208
rect 1397 6199 1455 6205
rect 1949 6205 1961 6208
rect 1995 6205 2007 6239
rect 3053 6239 3111 6245
rect 3053 6236 3065 6239
rect 1949 6199 2007 6205
rect 2884 6208 3065 6236
rect 2682 6128 2688 6180
rect 2740 6168 2746 6180
rect 2884 6177 2912 6208
rect 3053 6205 3065 6208
rect 3099 6205 3111 6239
rect 3053 6199 3111 6205
rect 3145 6239 3203 6245
rect 3145 6205 3157 6239
rect 3191 6236 3203 6239
rect 3234 6236 3240 6248
rect 3191 6208 3240 6236
rect 3191 6205 3203 6208
rect 3145 6199 3203 6205
rect 3234 6196 3240 6208
rect 3292 6196 3298 6248
rect 3344 6245 3372 6276
rect 3418 6264 3424 6276
rect 3476 6304 3482 6316
rect 5074 6304 5080 6316
rect 3476 6276 4936 6304
rect 5035 6276 5080 6304
rect 3476 6264 3482 6276
rect 4908 6248 4936 6276
rect 5074 6264 5080 6276
rect 5132 6264 5138 6316
rect 6730 6264 6736 6316
rect 6788 6304 6794 6316
rect 9033 6307 9091 6313
rect 9033 6304 9045 6307
rect 6788 6276 7328 6304
rect 6788 6264 6794 6276
rect 3329 6239 3387 6245
rect 3329 6205 3341 6239
rect 3375 6205 3387 6239
rect 4614 6236 4620 6248
rect 3329 6199 3387 6205
rect 4080 6208 4620 6236
rect 2869 6171 2927 6177
rect 2869 6168 2881 6171
rect 2740 6140 2881 6168
rect 2740 6128 2746 6140
rect 2869 6137 2881 6140
rect 2915 6137 2927 6171
rect 3786 6168 3792 6180
rect 3747 6140 3792 6168
rect 2869 6131 2927 6137
rect 2501 6103 2559 6109
rect 2501 6069 2513 6103
rect 2547 6100 2559 6103
rect 2774 6100 2780 6112
rect 2547 6072 2780 6100
rect 2547 6069 2559 6072
rect 2501 6063 2559 6069
rect 2774 6060 2780 6072
rect 2832 6060 2838 6112
rect 2884 6100 2912 6131
rect 3786 6128 3792 6140
rect 3844 6128 3850 6180
rect 4080 6109 4108 6208
rect 4614 6196 4620 6208
rect 4672 6196 4678 6248
rect 4709 6239 4767 6245
rect 4709 6205 4721 6239
rect 4755 6205 4767 6239
rect 4890 6236 4896 6248
rect 4851 6208 4896 6236
rect 4709 6199 4767 6205
rect 4724 6168 4752 6199
rect 4890 6196 4896 6208
rect 4948 6196 4954 6248
rect 7300 6245 7328 6276
rect 8128 6276 9045 6304
rect 8128 6248 8156 6276
rect 9033 6273 9045 6276
rect 9079 6273 9091 6307
rect 9033 6267 9091 6273
rect 10321 6307 10379 6313
rect 10321 6273 10333 6307
rect 10367 6304 10379 6307
rect 10686 6304 10692 6316
rect 10367 6276 10692 6304
rect 10367 6273 10379 6276
rect 10321 6267 10379 6273
rect 10686 6264 10692 6276
rect 10744 6264 10750 6316
rect 10965 6307 11023 6313
rect 10965 6273 10977 6307
rect 11011 6304 11023 6307
rect 11146 6304 11152 6316
rect 11011 6276 11152 6304
rect 11011 6273 11023 6276
rect 10965 6267 11023 6273
rect 11146 6264 11152 6276
rect 11204 6264 11210 6316
rect 11808 6304 11836 6335
rect 12437 6307 12495 6313
rect 12437 6304 12449 6307
rect 11808 6276 12449 6304
rect 12437 6273 12449 6276
rect 12483 6273 12495 6307
rect 12437 6267 12495 6273
rect 15749 6307 15807 6313
rect 15749 6273 15761 6307
rect 15795 6304 15807 6307
rect 15838 6304 15844 6316
rect 15795 6276 15844 6304
rect 15795 6273 15807 6276
rect 15749 6267 15807 6273
rect 15838 6264 15844 6276
rect 15896 6264 15902 6316
rect 7285 6239 7343 6245
rect 7285 6205 7297 6239
rect 7331 6205 7343 6239
rect 7742 6236 7748 6248
rect 7703 6208 7748 6236
rect 7285 6199 7343 6205
rect 7742 6196 7748 6208
rect 7800 6196 7806 6248
rect 8110 6236 8116 6248
rect 8071 6208 8116 6236
rect 8110 6196 8116 6208
rect 8168 6196 8174 6248
rect 8662 6236 8668 6248
rect 8623 6208 8668 6236
rect 8662 6196 8668 6208
rect 8720 6196 8726 6248
rect 13357 6239 13415 6245
rect 13357 6205 13369 6239
rect 13403 6236 13415 6239
rect 14458 6236 14464 6248
rect 13403 6208 14320 6236
rect 14419 6208 14464 6236
rect 13403 6205 13415 6208
rect 13357 6199 13415 6205
rect 4448 6140 4752 6168
rect 4065 6103 4123 6109
rect 4065 6100 4077 6103
rect 2884 6072 4077 6100
rect 4065 6069 4077 6072
rect 4111 6069 4123 6103
rect 4065 6063 4123 6069
rect 4154 6060 4160 6112
rect 4212 6100 4218 6112
rect 4448 6109 4476 6140
rect 6270 6128 6276 6180
rect 6328 6168 6334 6180
rect 7193 6171 7251 6177
rect 7193 6168 7205 6171
rect 6328 6140 7205 6168
rect 6328 6128 6334 6140
rect 7193 6137 7205 6140
rect 7239 6168 7251 6171
rect 7926 6168 7932 6180
rect 7239 6140 7932 6168
rect 7239 6137 7251 6140
rect 7193 6131 7251 6137
rect 7926 6128 7932 6140
rect 7984 6168 7990 6180
rect 8680 6168 8708 6196
rect 7984 6140 8708 6168
rect 10413 6171 10471 6177
rect 7984 6128 7990 6140
rect 10413 6137 10425 6171
rect 10459 6137 10471 6171
rect 10413 6131 10471 6137
rect 12758 6171 12816 6177
rect 12758 6137 12770 6171
rect 12804 6168 12816 6171
rect 13446 6168 13452 6180
rect 12804 6140 13452 6168
rect 12804 6137 12816 6140
rect 12758 6131 12816 6137
rect 4433 6103 4491 6109
rect 4433 6100 4445 6103
rect 4212 6072 4445 6100
rect 4212 6060 4218 6072
rect 4433 6069 4445 6072
rect 4479 6069 4491 6103
rect 4433 6063 4491 6069
rect 6457 6103 6515 6109
rect 6457 6069 6469 6103
rect 6503 6100 6515 6103
rect 7282 6100 7288 6112
rect 6503 6072 7288 6100
rect 6503 6069 6515 6072
rect 6457 6063 6515 6069
rect 7282 6060 7288 6072
rect 7340 6060 7346 6112
rect 7558 6100 7564 6112
rect 7519 6072 7564 6100
rect 7558 6060 7564 6072
rect 7616 6060 7622 6112
rect 8018 6060 8024 6112
rect 8076 6100 8082 6112
rect 9677 6103 9735 6109
rect 9677 6100 9689 6103
rect 8076 6072 9689 6100
rect 8076 6060 8082 6072
rect 9677 6069 9689 6072
rect 9723 6100 9735 6103
rect 9950 6100 9956 6112
rect 9723 6072 9956 6100
rect 9723 6069 9735 6072
rect 9677 6063 9735 6069
rect 9950 6060 9956 6072
rect 10008 6060 10014 6112
rect 10042 6060 10048 6112
rect 10100 6100 10106 6112
rect 10428 6100 10456 6131
rect 12250 6100 12256 6112
rect 10100 6072 10456 6100
rect 12211 6072 12256 6100
rect 10100 6060 10106 6072
rect 12250 6060 12256 6072
rect 12308 6100 12314 6112
rect 12773 6100 12801 6131
rect 13446 6128 13452 6140
rect 13504 6128 13510 6180
rect 14182 6168 14188 6180
rect 14143 6140 14188 6168
rect 14182 6128 14188 6140
rect 14240 6128 14246 6180
rect 14292 6168 14320 6208
rect 14458 6196 14464 6208
rect 14516 6196 14522 6248
rect 18046 6236 18052 6248
rect 18007 6208 18052 6236
rect 18046 6196 18052 6208
rect 18104 6236 18110 6248
rect 18601 6239 18659 6245
rect 18601 6236 18613 6239
rect 18104 6208 18613 6236
rect 18104 6196 18110 6208
rect 18601 6205 18613 6208
rect 18647 6205 18659 6239
rect 18601 6199 18659 6205
rect 23728 6239 23786 6245
rect 23728 6205 23740 6239
rect 23774 6236 23786 6239
rect 24118 6236 24124 6248
rect 23774 6208 24124 6236
rect 23774 6205 23786 6208
rect 23728 6199 23786 6205
rect 24118 6196 24124 6208
rect 24176 6196 24182 6248
rect 15654 6168 15660 6180
rect 14292 6140 15660 6168
rect 15654 6128 15660 6140
rect 15712 6128 15718 6180
rect 16850 6128 16856 6180
rect 16908 6168 16914 6180
rect 18966 6168 18972 6180
rect 16908 6140 18972 6168
rect 16908 6128 16914 6140
rect 18966 6128 18972 6140
rect 19024 6168 19030 6180
rect 24581 6171 24639 6177
rect 24581 6168 24593 6171
rect 19024 6140 24593 6168
rect 19024 6128 19030 6140
rect 24581 6137 24593 6140
rect 24627 6168 24639 6171
rect 24670 6168 24676 6180
rect 24627 6140 24676 6168
rect 24627 6137 24639 6140
rect 24581 6131 24639 6137
rect 24670 6128 24676 6140
rect 24728 6128 24734 6180
rect 12308 6072 12801 6100
rect 12308 6060 12314 6072
rect 13262 6060 13268 6112
rect 13320 6100 13326 6112
rect 13725 6103 13783 6109
rect 13725 6100 13737 6103
rect 13320 6072 13737 6100
rect 13320 6060 13326 6072
rect 13725 6069 13737 6072
rect 13771 6100 13783 6103
rect 13998 6100 14004 6112
rect 13771 6072 14004 6100
rect 13771 6069 13783 6072
rect 13725 6063 13783 6069
rect 13998 6060 14004 6072
rect 14056 6060 14062 6112
rect 18230 6100 18236 6112
rect 18191 6072 18236 6100
rect 18230 6060 18236 6072
rect 18288 6060 18294 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 3418 5896 3424 5908
rect 3160 5868 3424 5896
rect 3160 5837 3188 5868
rect 3418 5856 3424 5868
rect 3476 5856 3482 5908
rect 4890 5856 4896 5908
rect 4948 5896 4954 5908
rect 5077 5899 5135 5905
rect 5077 5896 5089 5899
rect 4948 5868 5089 5896
rect 4948 5856 4954 5868
rect 5077 5865 5089 5868
rect 5123 5865 5135 5899
rect 5077 5859 5135 5865
rect 5442 5856 5448 5908
rect 5500 5896 5506 5908
rect 5997 5899 6055 5905
rect 5997 5896 6009 5899
rect 5500 5868 6009 5896
rect 5500 5856 5506 5868
rect 5997 5865 6009 5868
rect 6043 5865 6055 5899
rect 5997 5859 6055 5865
rect 6457 5899 6515 5905
rect 6457 5865 6469 5899
rect 6503 5896 6515 5899
rect 6730 5896 6736 5908
rect 6503 5868 6736 5896
rect 6503 5865 6515 5868
rect 6457 5859 6515 5865
rect 6730 5856 6736 5868
rect 6788 5856 6794 5908
rect 7377 5899 7435 5905
rect 7377 5865 7389 5899
rect 7423 5896 7435 5899
rect 7742 5896 7748 5908
rect 7423 5868 7748 5896
rect 7423 5865 7435 5868
rect 7377 5859 7435 5865
rect 7742 5856 7748 5868
rect 7800 5856 7806 5908
rect 8757 5899 8815 5905
rect 8757 5865 8769 5899
rect 8803 5896 8815 5899
rect 11422 5896 11428 5908
rect 8803 5868 9674 5896
rect 11383 5868 11428 5896
rect 8803 5865 8815 5868
rect 8757 5859 8815 5865
rect 3145 5831 3203 5837
rect 3145 5797 3157 5831
rect 3191 5797 3203 5831
rect 3145 5791 3203 5797
rect 3234 5788 3240 5840
rect 3292 5828 3298 5840
rect 4065 5831 4123 5837
rect 4065 5828 4077 5831
rect 3292 5800 4077 5828
rect 3292 5788 3298 5800
rect 4065 5797 4077 5800
rect 4111 5797 4123 5831
rect 6748 5828 6776 5856
rect 7653 5831 7711 5837
rect 7653 5828 7665 5831
rect 6748 5800 7665 5828
rect 4065 5791 4123 5797
rect 7653 5797 7665 5800
rect 7699 5797 7711 5831
rect 7653 5791 7711 5797
rect 8018 5788 8024 5840
rect 8076 5828 8082 5840
rect 8158 5831 8216 5837
rect 8158 5828 8170 5831
rect 8076 5800 8170 5828
rect 8076 5788 8082 5800
rect 8158 5797 8170 5800
rect 8204 5797 8216 5831
rect 9646 5828 9674 5868
rect 11422 5856 11428 5868
rect 11480 5856 11486 5908
rect 13081 5899 13139 5905
rect 13081 5865 13093 5899
rect 13127 5896 13139 5899
rect 13127 5868 13670 5896
rect 13127 5865 13139 5868
rect 13081 5859 13139 5865
rect 9858 5828 9864 5840
rect 9646 5800 9864 5828
rect 8158 5791 8216 5797
rect 9858 5788 9864 5800
rect 9916 5788 9922 5840
rect 12250 5788 12256 5840
rect 12308 5828 12314 5840
rect 12482 5831 12540 5837
rect 12482 5828 12494 5831
rect 12308 5800 12494 5828
rect 12308 5788 12314 5800
rect 12482 5797 12494 5800
rect 12528 5797 12540 5831
rect 12482 5791 12540 5797
rect 12986 5788 12992 5840
rect 13044 5828 13050 5840
rect 13357 5831 13415 5837
rect 13357 5828 13369 5831
rect 13044 5800 13369 5828
rect 13044 5788 13050 5800
rect 13357 5797 13369 5800
rect 13403 5797 13415 5831
rect 13642 5828 13670 5868
rect 13722 5856 13728 5908
rect 13780 5896 13786 5908
rect 14047 5899 14105 5905
rect 14047 5896 14059 5899
rect 13780 5868 14059 5896
rect 13780 5856 13786 5868
rect 14047 5865 14059 5868
rect 14093 5865 14105 5899
rect 14047 5859 14105 5865
rect 14458 5828 14464 5840
rect 13642 5800 14464 5828
rect 13357 5791 13415 5797
rect 14458 5788 14464 5800
rect 14516 5788 14522 5840
rect 15470 5828 15476 5840
rect 15431 5800 15476 5828
rect 15470 5788 15476 5800
rect 15528 5788 15534 5840
rect 2774 5760 2780 5772
rect 2735 5732 2780 5760
rect 2774 5720 2780 5732
rect 2832 5720 2838 5772
rect 2317 5695 2375 5701
rect 2317 5661 2329 5695
rect 2363 5692 2375 5695
rect 3252 5692 3280 5788
rect 4154 5720 4160 5772
rect 4212 5760 4218 5772
rect 5813 5763 5871 5769
rect 4212 5732 4257 5760
rect 4212 5720 4218 5732
rect 5813 5729 5825 5763
rect 5859 5760 5871 5763
rect 6270 5760 6276 5772
rect 5859 5732 6276 5760
rect 5859 5729 5871 5732
rect 5813 5723 5871 5729
rect 6270 5720 6276 5732
rect 6328 5720 6334 5772
rect 6546 5720 6552 5772
rect 6604 5760 6610 5772
rect 6860 5763 6918 5769
rect 6860 5760 6872 5763
rect 6604 5732 6872 5760
rect 6604 5720 6610 5732
rect 6860 5729 6872 5732
rect 6906 5729 6918 5763
rect 6860 5723 6918 5729
rect 7558 5720 7564 5772
rect 7616 5760 7622 5772
rect 7837 5763 7895 5769
rect 7837 5760 7849 5763
rect 7616 5732 7849 5760
rect 7616 5720 7622 5732
rect 7837 5729 7849 5732
rect 7883 5760 7895 5763
rect 8386 5760 8392 5772
rect 7883 5732 8392 5760
rect 7883 5729 7895 5732
rect 7837 5723 7895 5729
rect 8386 5720 8392 5732
rect 8444 5720 8450 5772
rect 12158 5760 12164 5772
rect 11348 5732 12164 5760
rect 2363 5664 3280 5692
rect 2363 5661 2375 5664
rect 2317 5655 2375 5661
rect 9306 5652 9312 5704
rect 9364 5692 9370 5704
rect 9769 5695 9827 5701
rect 9769 5692 9781 5695
rect 9364 5664 9781 5692
rect 9364 5652 9370 5664
rect 9769 5661 9781 5664
rect 9815 5661 9827 5695
rect 9769 5655 9827 5661
rect 10413 5695 10471 5701
rect 10413 5661 10425 5695
rect 10459 5692 10471 5695
rect 10962 5692 10968 5704
rect 10459 5664 10968 5692
rect 10459 5661 10471 5664
rect 10413 5655 10471 5661
rect 10962 5652 10968 5664
rect 11020 5652 11026 5704
rect 9030 5584 9036 5636
rect 9088 5624 9094 5636
rect 11348 5624 11376 5732
rect 12158 5720 12164 5732
rect 12216 5720 12222 5772
rect 13170 5720 13176 5772
rect 13228 5760 13234 5772
rect 13722 5760 13728 5772
rect 13228 5732 13728 5760
rect 13228 5720 13234 5732
rect 13722 5720 13728 5732
rect 13780 5760 13786 5772
rect 13944 5763 14002 5769
rect 13944 5760 13956 5763
rect 13780 5732 13956 5760
rect 13780 5720 13786 5732
rect 13944 5729 13956 5732
rect 13990 5729 14002 5763
rect 13944 5723 14002 5729
rect 15378 5692 15384 5704
rect 15339 5664 15384 5692
rect 15378 5652 15384 5664
rect 15436 5652 15442 5704
rect 16022 5692 16028 5704
rect 15983 5664 16028 5692
rect 16022 5652 16028 5664
rect 16080 5652 16086 5704
rect 9088 5596 11376 5624
rect 9088 5584 9094 5596
rect 6963 5559 7021 5565
rect 6963 5525 6975 5559
rect 7009 5556 7021 5559
rect 7190 5556 7196 5568
rect 7009 5528 7196 5556
rect 7009 5525 7021 5528
rect 6963 5519 7021 5525
rect 7190 5516 7196 5528
rect 7248 5516 7254 5568
rect 10686 5556 10692 5568
rect 10647 5528 10692 5556
rect 10686 5516 10692 5528
rect 10744 5516 10750 5568
rect 14458 5556 14464 5568
rect 14419 5528 14464 5556
rect 14458 5516 14464 5528
rect 14516 5516 14522 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 4525 5355 4583 5361
rect 4525 5321 4537 5355
rect 4571 5352 4583 5355
rect 5534 5352 5540 5364
rect 4571 5324 5540 5352
rect 4571 5321 4583 5324
rect 4525 5315 4583 5321
rect 5534 5312 5540 5324
rect 5592 5312 5598 5364
rect 5905 5355 5963 5361
rect 5905 5321 5917 5355
rect 5951 5352 5963 5355
rect 6362 5352 6368 5364
rect 5951 5324 6368 5352
rect 5951 5321 5963 5324
rect 5905 5315 5963 5321
rect 6362 5312 6368 5324
rect 6420 5312 6426 5364
rect 9950 5312 9956 5364
rect 10008 5352 10014 5364
rect 12161 5355 12219 5361
rect 12161 5352 12173 5355
rect 10008 5324 12173 5352
rect 10008 5312 10014 5324
rect 12161 5321 12173 5324
rect 12207 5352 12219 5355
rect 12250 5352 12256 5364
rect 12207 5324 12256 5352
rect 12207 5321 12219 5324
rect 12161 5315 12219 5321
rect 12250 5312 12256 5324
rect 12308 5312 12314 5364
rect 13722 5312 13728 5364
rect 13780 5352 13786 5364
rect 13909 5355 13967 5361
rect 13909 5352 13921 5355
rect 13780 5324 13921 5352
rect 13780 5312 13786 5324
rect 13909 5321 13921 5324
rect 13955 5321 13967 5355
rect 13909 5315 13967 5321
rect 15378 5312 15384 5364
rect 15436 5352 15442 5364
rect 16853 5355 16911 5361
rect 16853 5352 16865 5355
rect 15436 5324 16865 5352
rect 15436 5312 15442 5324
rect 16853 5321 16865 5324
rect 16899 5321 16911 5355
rect 16853 5315 16911 5321
rect 5629 5287 5687 5293
rect 5629 5253 5641 5287
rect 5675 5284 5687 5287
rect 5994 5284 6000 5296
rect 5675 5256 6000 5284
rect 5675 5253 5687 5256
rect 5629 5247 5687 5253
rect 2038 5176 2044 5228
rect 2096 5216 2102 5228
rect 2869 5219 2927 5225
rect 2869 5216 2881 5219
rect 2096 5188 2881 5216
rect 2096 5176 2102 5188
rect 2869 5185 2881 5188
rect 2915 5216 2927 5219
rect 4065 5219 4123 5225
rect 4065 5216 4077 5219
rect 2915 5188 4077 5216
rect 2915 5185 2927 5188
rect 2869 5179 2927 5185
rect 4065 5185 4077 5188
rect 4111 5216 4123 5219
rect 4154 5216 4160 5228
rect 4111 5188 4160 5216
rect 4111 5185 4123 5188
rect 4065 5179 4123 5185
rect 4154 5176 4160 5188
rect 4212 5176 4218 5228
rect 2682 5108 2688 5160
rect 2740 5148 2746 5160
rect 2777 5151 2835 5157
rect 2777 5148 2789 5151
rect 2740 5120 2789 5148
rect 2740 5108 2746 5120
rect 2777 5117 2789 5120
rect 2823 5117 2835 5151
rect 2777 5111 2835 5117
rect 3053 5151 3111 5157
rect 3053 5117 3065 5151
rect 3099 5117 3111 5151
rect 3053 5111 3111 5117
rect 3068 5080 3096 5111
rect 3786 5108 3792 5160
rect 3844 5148 3850 5160
rect 5736 5157 5764 5256
rect 5994 5244 6000 5256
rect 6052 5244 6058 5296
rect 6270 5284 6276 5296
rect 6231 5256 6276 5284
rect 6270 5244 6276 5256
rect 6328 5244 6334 5296
rect 14921 5287 14979 5293
rect 14921 5284 14933 5287
rect 13786 5256 14933 5284
rect 6638 5176 6644 5228
rect 6696 5216 6702 5228
rect 6825 5219 6883 5225
rect 6825 5216 6837 5219
rect 6696 5188 6837 5216
rect 6696 5176 6702 5188
rect 6825 5185 6837 5188
rect 6871 5185 6883 5219
rect 6825 5179 6883 5185
rect 10873 5219 10931 5225
rect 10873 5185 10885 5219
rect 10919 5216 10931 5219
rect 10962 5216 10968 5228
rect 10919 5188 10968 5216
rect 10919 5185 10931 5188
rect 10873 5179 10931 5185
rect 10962 5176 10968 5188
rect 11020 5176 11026 5228
rect 13449 5219 13507 5225
rect 13449 5185 13461 5219
rect 13495 5216 13507 5219
rect 13786 5216 13814 5256
rect 14921 5253 14933 5256
rect 14967 5284 14979 5287
rect 15396 5284 15424 5312
rect 15654 5284 15660 5296
rect 14967 5256 15424 5284
rect 15615 5256 15660 5284
rect 14967 5253 14979 5256
rect 14921 5247 14979 5253
rect 15654 5244 15660 5256
rect 15712 5284 15718 5296
rect 15712 5256 15976 5284
rect 15712 5244 15718 5256
rect 13495 5188 13814 5216
rect 15381 5219 15439 5225
rect 13495 5185 13507 5188
rect 13449 5179 13507 5185
rect 15381 5185 15393 5219
rect 15427 5216 15439 5219
rect 15470 5216 15476 5228
rect 15427 5188 15476 5216
rect 15427 5185 15439 5188
rect 15381 5179 15439 5185
rect 15470 5176 15476 5188
rect 15528 5216 15534 5228
rect 15841 5219 15899 5225
rect 15841 5216 15853 5219
rect 15528 5188 15853 5216
rect 15528 5176 15534 5188
rect 15841 5185 15853 5188
rect 15887 5185 15899 5219
rect 15841 5179 15899 5185
rect 15948 5157 15976 5256
rect 4341 5151 4399 5157
rect 4341 5148 4353 5151
rect 3844 5120 4353 5148
rect 3844 5108 3850 5120
rect 4341 5117 4353 5120
rect 4387 5148 4399 5151
rect 4801 5151 4859 5157
rect 4801 5148 4813 5151
rect 4387 5120 4813 5148
rect 4387 5117 4399 5120
rect 4341 5111 4399 5117
rect 4801 5117 4813 5120
rect 4847 5117 4859 5151
rect 4801 5111 4859 5117
rect 5721 5151 5779 5157
rect 5721 5117 5733 5151
rect 5767 5117 5779 5151
rect 5721 5111 5779 5117
rect 15933 5151 15991 5157
rect 15933 5117 15945 5151
rect 15979 5117 15991 5151
rect 15933 5111 15991 5117
rect 2792 5052 3096 5080
rect 3513 5083 3571 5089
rect 2792 5024 2820 5052
rect 3513 5049 3525 5083
rect 3559 5080 3571 5083
rect 5350 5080 5356 5092
rect 3559 5052 5356 5080
rect 3559 5049 3571 5052
rect 3513 5043 3571 5049
rect 5350 5040 5356 5052
rect 5408 5040 5414 5092
rect 6546 5080 6552 5092
rect 6507 5052 6552 5080
rect 6546 5040 6552 5052
rect 6604 5040 6610 5092
rect 6822 5040 6828 5092
rect 6880 5080 6886 5092
rect 7146 5083 7204 5089
rect 7146 5080 7158 5083
rect 6880 5052 7158 5080
rect 6880 5040 6886 5052
rect 7146 5049 7158 5052
rect 7192 5080 7204 5083
rect 8018 5080 8024 5092
rect 7192 5052 8024 5080
rect 7192 5049 7204 5052
rect 7146 5043 7204 5049
rect 8018 5040 8024 5052
rect 8076 5040 8082 5092
rect 8662 5080 8668 5092
rect 8623 5052 8668 5080
rect 8662 5040 8668 5052
rect 8720 5040 8726 5092
rect 8757 5083 8815 5089
rect 8757 5049 8769 5083
rect 8803 5049 8815 5083
rect 9306 5080 9312 5092
rect 9267 5052 9312 5080
rect 8757 5043 8815 5049
rect 2038 5012 2044 5024
rect 1999 4984 2044 5012
rect 2038 4972 2044 4984
rect 2096 4972 2102 5024
rect 2501 5015 2559 5021
rect 2501 4981 2513 5015
rect 2547 5012 2559 5015
rect 2774 5012 2780 5024
rect 2547 4984 2780 5012
rect 2547 4981 2559 4984
rect 2501 4975 2559 4981
rect 2774 4972 2780 4984
rect 2832 4972 2838 5024
rect 7742 5012 7748 5024
rect 7703 4984 7748 5012
rect 7742 4972 7748 4984
rect 7800 4972 7806 5024
rect 8294 4972 8300 5024
rect 8352 5012 8358 5024
rect 8389 5015 8447 5021
rect 8389 5012 8401 5015
rect 8352 4984 8401 5012
rect 8352 4972 8358 4984
rect 8389 4981 8401 4984
rect 8435 5012 8447 5015
rect 8772 5012 8800 5043
rect 9306 5040 9312 5052
rect 9364 5040 9370 5092
rect 9677 5083 9735 5089
rect 9677 5049 9689 5083
rect 9723 5080 9735 5083
rect 10042 5080 10048 5092
rect 9723 5052 10048 5080
rect 9723 5049 9735 5052
rect 9677 5043 9735 5049
rect 10042 5040 10048 5052
rect 10100 5080 10106 5092
rect 10229 5083 10287 5089
rect 10229 5080 10241 5083
rect 10100 5052 10241 5080
rect 10100 5040 10106 5052
rect 10229 5049 10241 5052
rect 10275 5049 10287 5083
rect 10229 5043 10287 5049
rect 10321 5083 10379 5089
rect 10321 5049 10333 5083
rect 10367 5049 10379 5083
rect 10321 5043 10379 5049
rect 11885 5083 11943 5089
rect 11885 5049 11897 5083
rect 11931 5080 11943 5083
rect 12802 5080 12808 5092
rect 11931 5052 12808 5080
rect 11931 5049 11943 5052
rect 11885 5043 11943 5049
rect 9950 5012 9956 5024
rect 8435 4984 8800 5012
rect 9911 4984 9956 5012
rect 8435 4981 8447 4984
rect 8389 4975 8447 4981
rect 9950 4972 9956 4984
rect 10008 5012 10014 5024
rect 10336 5012 10364 5043
rect 12802 5040 12808 5052
rect 12860 5040 12866 5092
rect 12894 5040 12900 5092
rect 12952 5080 12958 5092
rect 14366 5080 14372 5092
rect 12952 5052 12997 5080
rect 14327 5052 14372 5080
rect 12952 5040 12958 5052
rect 14366 5040 14372 5052
rect 14424 5040 14430 5092
rect 14458 5040 14464 5092
rect 14516 5080 14522 5092
rect 14516 5052 14561 5080
rect 14516 5040 14522 5052
rect 11146 5012 11152 5024
rect 10008 4984 10364 5012
rect 11107 4984 11152 5012
rect 10008 4972 10014 4984
rect 11146 4972 11152 4984
rect 11204 4972 11210 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 6638 4768 6644 4820
rect 6696 4808 6702 4820
rect 7285 4811 7343 4817
rect 7285 4808 7297 4811
rect 6696 4780 7297 4808
rect 6696 4768 6702 4780
rect 7285 4777 7297 4780
rect 7331 4777 7343 4811
rect 8386 4808 8392 4820
rect 8347 4780 8392 4808
rect 7285 4771 7343 4777
rect 8386 4768 8392 4780
rect 8444 4768 8450 4820
rect 9950 4808 9956 4820
rect 9911 4780 9956 4808
rect 9950 4768 9956 4780
rect 10008 4768 10014 4820
rect 11747 4811 11805 4817
rect 11747 4777 11759 4811
rect 11793 4808 11805 4811
rect 12526 4808 12532 4820
rect 11793 4780 12532 4808
rect 11793 4777 11805 4780
rect 11747 4771 11805 4777
rect 12526 4768 12532 4780
rect 12584 4768 12590 4820
rect 14366 4768 14372 4820
rect 14424 4808 14430 4820
rect 14645 4811 14703 4817
rect 14645 4808 14657 4811
rect 14424 4780 14657 4808
rect 14424 4768 14430 4780
rect 14645 4777 14657 4780
rect 14691 4808 14703 4811
rect 14734 4808 14740 4820
rect 14691 4780 14740 4808
rect 14691 4777 14703 4780
rect 14645 4771 14703 4777
rect 14734 4768 14740 4780
rect 14792 4768 14798 4820
rect 2133 4743 2191 4749
rect 2133 4709 2145 4743
rect 2179 4740 2191 4743
rect 2682 4740 2688 4752
rect 2179 4712 2688 4740
rect 2179 4709 2191 4712
rect 2133 4703 2191 4709
rect 2682 4700 2688 4712
rect 2740 4740 2746 4752
rect 3145 4743 3203 4749
rect 3145 4740 3157 4743
rect 2740 4712 3157 4740
rect 2740 4700 2746 4712
rect 3145 4709 3157 4712
rect 3191 4709 3203 4743
rect 3145 4703 3203 4709
rect 7190 4700 7196 4752
rect 7248 4740 7254 4752
rect 7469 4743 7527 4749
rect 7469 4740 7481 4743
rect 7248 4712 7481 4740
rect 7248 4700 7254 4712
rect 7469 4709 7481 4712
rect 7515 4709 7527 4743
rect 7469 4703 7527 4709
rect 7561 4743 7619 4749
rect 7561 4709 7573 4743
rect 7607 4740 7619 4743
rect 7742 4740 7748 4752
rect 7607 4712 7748 4740
rect 7607 4709 7619 4712
rect 7561 4703 7619 4709
rect 7742 4700 7748 4712
rect 7800 4700 7806 4752
rect 8113 4743 8171 4749
rect 8113 4709 8125 4743
rect 8159 4740 8171 4743
rect 9306 4740 9312 4752
rect 8159 4712 9312 4740
rect 8159 4709 8171 4712
rect 8113 4703 8171 4709
rect 9306 4700 9312 4712
rect 9364 4740 9370 4752
rect 9401 4743 9459 4749
rect 9401 4740 9413 4743
rect 9364 4712 9413 4740
rect 9364 4700 9370 4712
rect 9401 4709 9413 4712
rect 9447 4709 9459 4743
rect 12158 4740 12164 4752
rect 12119 4712 12164 4740
rect 9401 4703 9459 4709
rect 12158 4700 12164 4712
rect 12216 4700 12222 4752
rect 13826 4743 13884 4749
rect 13826 4709 13838 4743
rect 13872 4740 13884 4743
rect 14182 4740 14188 4752
rect 13872 4712 14188 4740
rect 13872 4709 13884 4712
rect 13826 4703 13884 4709
rect 14182 4700 14188 4712
rect 14240 4700 14246 4752
rect 15473 4743 15531 4749
rect 15473 4709 15485 4743
rect 15519 4740 15531 4743
rect 15654 4740 15660 4752
rect 15519 4712 15660 4740
rect 15519 4709 15531 4712
rect 15473 4703 15531 4709
rect 15654 4700 15660 4712
rect 15712 4700 15718 4752
rect 16022 4740 16028 4752
rect 15983 4712 16028 4740
rect 16022 4700 16028 4712
rect 16080 4700 16086 4752
rect 27614 4740 27620 4752
rect 24663 4712 27620 4740
rect 24663 4684 24691 4712
rect 27614 4700 27620 4712
rect 27672 4700 27678 4752
rect 1486 4672 1492 4684
rect 1447 4644 1492 4672
rect 1486 4632 1492 4644
rect 1544 4632 1550 4684
rect 5442 4632 5448 4684
rect 5500 4672 5506 4684
rect 5756 4675 5814 4681
rect 5756 4672 5768 4675
rect 5500 4644 5768 4672
rect 5500 4632 5506 4644
rect 5756 4641 5768 4644
rect 5802 4641 5814 4675
rect 5756 4635 5814 4641
rect 9858 4632 9864 4684
rect 9916 4672 9922 4684
rect 10318 4672 10324 4684
rect 9916 4644 10324 4672
rect 9916 4632 9922 4644
rect 10318 4632 10324 4644
rect 10376 4672 10382 4684
rect 11146 4672 11152 4684
rect 10376 4644 11152 4672
rect 10376 4632 10382 4644
rect 11146 4632 11152 4644
rect 11204 4632 11210 4684
rect 11514 4632 11520 4684
rect 11572 4672 11578 4684
rect 11644 4675 11702 4681
rect 11644 4672 11656 4675
rect 11572 4644 11656 4672
rect 11572 4632 11578 4644
rect 11644 4641 11656 4644
rect 11690 4641 11702 4675
rect 11644 4635 11702 4641
rect 11974 4632 11980 4684
rect 12032 4672 12038 4684
rect 24663 4681 24676 4684
rect 12656 4675 12714 4681
rect 12656 4672 12668 4675
rect 12032 4644 12668 4672
rect 12032 4632 12038 4644
rect 12656 4641 12668 4644
rect 12702 4641 12714 4675
rect 24648 4675 24676 4681
rect 24648 4672 24660 4675
rect 24583 4644 24660 4672
rect 12656 4635 12714 4641
rect 24648 4641 24660 4644
rect 24648 4635 24676 4641
rect 24670 4632 24676 4635
rect 24728 4632 24734 4684
rect 5859 4607 5917 4613
rect 5859 4573 5871 4607
rect 5905 4604 5917 4607
rect 8662 4604 8668 4616
rect 5905 4576 8668 4604
rect 5905 4573 5917 4576
rect 5859 4567 5917 4573
rect 8662 4564 8668 4576
rect 8720 4604 8726 4616
rect 8757 4607 8815 4613
rect 8757 4604 8769 4607
rect 8720 4576 8769 4604
rect 8720 4564 8726 4576
rect 8757 4573 8769 4576
rect 8803 4573 8815 4607
rect 8757 4567 8815 4573
rect 12759 4607 12817 4613
rect 12759 4573 12771 4607
rect 12805 4604 12817 4607
rect 13722 4604 13728 4616
rect 12805 4576 13728 4604
rect 12805 4573 12817 4576
rect 12759 4567 12817 4573
rect 13722 4564 13728 4576
rect 13780 4564 13786 4616
rect 14369 4607 14427 4613
rect 14369 4573 14381 4607
rect 14415 4604 14427 4607
rect 14550 4604 14556 4616
rect 14415 4576 14556 4604
rect 14415 4573 14427 4576
rect 14369 4567 14427 4573
rect 14550 4564 14556 4576
rect 14608 4604 14614 4616
rect 15381 4607 15439 4613
rect 15381 4604 15393 4607
rect 14608 4576 15393 4604
rect 14608 4564 14614 4576
rect 15381 4573 15393 4576
rect 15427 4573 15439 4607
rect 15381 4567 15439 4573
rect 1670 4496 1676 4548
rect 1728 4536 1734 4548
rect 2866 4536 2872 4548
rect 1728 4508 2872 4536
rect 1728 4496 1734 4508
rect 2866 4496 2872 4508
rect 2924 4536 2930 4548
rect 6822 4536 6828 4548
rect 2924 4508 6828 4536
rect 2924 4496 2930 4508
rect 6822 4496 6828 4508
rect 6880 4496 6886 4548
rect 12894 4496 12900 4548
rect 12952 4536 12958 4548
rect 13173 4539 13231 4545
rect 13173 4536 13185 4539
rect 12952 4508 13185 4536
rect 12952 4496 12958 4508
rect 13173 4505 13185 4508
rect 13219 4536 13231 4539
rect 14182 4536 14188 4548
rect 13219 4508 14188 4536
rect 13219 4505 13231 4508
rect 13173 4499 13231 4505
rect 14182 4496 14188 4508
rect 14240 4496 14246 4548
rect 2774 4468 2780 4480
rect 2735 4440 2780 4468
rect 2774 4428 2780 4440
rect 2832 4428 2838 4480
rect 21542 4428 21548 4480
rect 21600 4468 21606 4480
rect 24719 4471 24777 4477
rect 24719 4468 24731 4471
rect 21600 4440 24731 4468
rect 21600 4428 21606 4440
rect 24719 4437 24731 4440
rect 24765 4437 24777 4471
rect 24719 4431 24777 4437
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 5442 4224 5448 4276
rect 5500 4264 5506 4276
rect 5721 4267 5779 4273
rect 5721 4264 5733 4267
rect 5500 4236 5733 4264
rect 5500 4224 5506 4236
rect 5721 4233 5733 4236
rect 5767 4233 5779 4267
rect 5721 4227 5779 4233
rect 7742 4224 7748 4276
rect 7800 4264 7806 4276
rect 7929 4267 7987 4273
rect 7929 4264 7941 4267
rect 7800 4236 7941 4264
rect 7800 4224 7806 4236
rect 7929 4233 7941 4236
rect 7975 4233 7987 4267
rect 7929 4227 7987 4233
rect 9263 4267 9321 4273
rect 9263 4233 9275 4267
rect 9309 4264 9321 4267
rect 10686 4264 10692 4276
rect 9309 4236 10692 4264
rect 9309 4233 9321 4236
rect 9263 4227 9321 4233
rect 10686 4224 10692 4236
rect 10744 4224 10750 4276
rect 11514 4224 11520 4276
rect 11572 4264 11578 4276
rect 11793 4267 11851 4273
rect 11793 4264 11805 4267
rect 11572 4236 11805 4264
rect 11572 4224 11578 4236
rect 11793 4233 11805 4236
rect 11839 4233 11851 4267
rect 11793 4227 11851 4233
rect 11974 4224 11980 4276
rect 12032 4264 12038 4276
rect 12621 4267 12679 4273
rect 12621 4264 12633 4267
rect 12032 4236 12633 4264
rect 12032 4224 12038 4236
rect 12621 4233 12633 4236
rect 12667 4233 12679 4267
rect 12621 4227 12679 4233
rect 13725 4267 13783 4273
rect 13725 4233 13737 4267
rect 13771 4264 13783 4267
rect 14182 4264 14188 4276
rect 13771 4236 14188 4264
rect 13771 4233 13783 4236
rect 13725 4227 13783 4233
rect 14182 4224 14188 4236
rect 14240 4224 14246 4276
rect 15381 4267 15439 4273
rect 15381 4233 15393 4267
rect 15427 4264 15439 4267
rect 15654 4264 15660 4276
rect 15427 4236 15660 4264
rect 15427 4233 15439 4236
rect 15381 4227 15439 4233
rect 15654 4224 15660 4236
rect 15712 4224 15718 4276
rect 24670 4264 24676 4276
rect 24631 4236 24676 4264
rect 24670 4224 24676 4236
rect 24728 4224 24734 4276
rect 9953 4199 10011 4205
rect 9953 4165 9965 4199
rect 9999 4196 10011 4199
rect 10318 4196 10324 4208
rect 9999 4168 10324 4196
rect 9999 4165 10011 4168
rect 9953 4159 10011 4165
rect 10318 4156 10324 4168
rect 10376 4156 10382 4208
rect 14093 4199 14151 4205
rect 14093 4165 14105 4199
rect 14139 4196 14151 4199
rect 14458 4196 14464 4208
rect 14139 4168 14464 4196
rect 14139 4165 14151 4168
rect 14093 4159 14151 4165
rect 14458 4156 14464 4168
rect 14516 4156 14522 4208
rect 7653 4131 7711 4137
rect 7653 4097 7665 4131
rect 7699 4128 7711 4131
rect 8294 4128 8300 4140
rect 7699 4100 8300 4128
rect 7699 4097 7711 4100
rect 7653 4091 7711 4097
rect 8294 4088 8300 4100
rect 8352 4088 8358 4140
rect 9858 4128 9864 4140
rect 9048 4100 9864 4128
rect 6641 4063 6699 4069
rect 6641 4029 6653 4063
rect 6687 4060 6699 4063
rect 7561 4063 7619 4069
rect 7561 4060 7573 4063
rect 6687 4032 7573 4060
rect 6687 4029 6699 4032
rect 6641 4023 6699 4029
rect 7561 4029 7573 4032
rect 7607 4060 7619 4063
rect 7742 4060 7748 4072
rect 7607 4032 7748 4060
rect 7607 4029 7619 4032
rect 7561 4023 7619 4029
rect 7742 4020 7748 4032
rect 7800 4020 7806 4072
rect 6546 3952 6552 4004
rect 6604 3992 6610 4004
rect 9048 3992 9076 4100
rect 9858 4088 9864 4100
rect 9916 4088 9922 4140
rect 10042 4088 10048 4140
rect 10100 4128 10106 4140
rect 10137 4131 10195 4137
rect 10137 4128 10149 4131
rect 10100 4100 10149 4128
rect 10100 4088 10106 4100
rect 10137 4097 10149 4100
rect 10183 4097 10195 4131
rect 10137 4091 10195 4097
rect 11333 4131 11391 4137
rect 11333 4097 11345 4131
rect 11379 4128 11391 4131
rect 12434 4128 12440 4140
rect 11379 4100 12440 4128
rect 11379 4097 11391 4100
rect 11333 4091 11391 4097
rect 12434 4088 12440 4100
rect 12492 4088 12498 4140
rect 12802 4088 12808 4140
rect 12860 4128 12866 4140
rect 13173 4131 13231 4137
rect 13173 4128 13185 4131
rect 12860 4100 13185 4128
rect 12860 4088 12866 4100
rect 13173 4097 13185 4100
rect 13219 4097 13231 4131
rect 14550 4128 14556 4140
rect 14511 4100 14556 4128
rect 13173 4091 13231 4097
rect 14550 4088 14556 4100
rect 14608 4128 14614 4140
rect 15657 4131 15715 4137
rect 15657 4128 15669 4131
rect 14608 4100 15669 4128
rect 14608 4088 14614 4100
rect 15657 4097 15669 4100
rect 15703 4097 15715 4131
rect 15657 4091 15715 4097
rect 9192 4063 9250 4069
rect 9192 4029 9204 4063
rect 9238 4060 9250 4063
rect 9238 4032 9628 4060
rect 9238 4029 9250 4032
rect 9192 4023 9250 4029
rect 6604 3964 9076 3992
rect 6604 3952 6610 3964
rect 9600 3936 9628 4032
rect 14274 3992 14280 4004
rect 14235 3964 14280 3992
rect 14274 3952 14280 3964
rect 14332 3952 14338 4004
rect 14369 3995 14427 4001
rect 14369 3961 14381 3995
rect 14415 3992 14427 3995
rect 14458 3992 14464 4004
rect 14415 3964 14464 3992
rect 14415 3961 14427 3964
rect 14369 3955 14427 3961
rect 14458 3952 14464 3964
rect 14516 3952 14522 4004
rect 14734 3952 14740 4004
rect 14792 3992 14798 4004
rect 21542 3992 21548 4004
rect 14792 3964 21548 3992
rect 14792 3952 14798 3964
rect 21542 3952 21548 3964
rect 21600 3952 21606 4004
rect 1486 3884 1492 3936
rect 1544 3924 1550 3936
rect 1581 3927 1639 3933
rect 1581 3924 1593 3927
rect 1544 3896 1593 3924
rect 1544 3884 1550 3896
rect 1581 3893 1593 3896
rect 1627 3893 1639 3927
rect 9582 3924 9588 3936
rect 9543 3896 9588 3924
rect 1581 3887 1639 3893
rect 9582 3884 9588 3896
rect 9640 3884 9646 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1535 3723 1593 3729
rect 1535 3689 1547 3723
rect 1581 3720 1593 3723
rect 1762 3720 1768 3732
rect 1581 3692 1768 3720
rect 1581 3689 1593 3692
rect 1535 3683 1593 3689
rect 1762 3680 1768 3692
rect 1820 3680 1826 3732
rect 7190 3680 7196 3732
rect 7248 3720 7254 3732
rect 7377 3723 7435 3729
rect 7377 3720 7389 3723
rect 7248 3692 7389 3720
rect 7248 3680 7254 3692
rect 7377 3689 7389 3692
rect 7423 3689 7435 3723
rect 13722 3720 13728 3732
rect 13683 3692 13728 3720
rect 7377 3683 7435 3689
rect 13722 3680 13728 3692
rect 13780 3680 13786 3732
rect 1394 3584 1400 3596
rect 1355 3556 1400 3584
rect 1394 3544 1400 3556
rect 1452 3544 1458 3596
rect 15378 3593 15384 3596
rect 15356 3587 15384 3593
rect 15356 3584 15368 3587
rect 15291 3556 15368 3584
rect 15356 3553 15368 3556
rect 15436 3584 15442 3596
rect 16022 3584 16028 3596
rect 15436 3556 16028 3584
rect 15356 3547 15384 3553
rect 15378 3544 15384 3547
rect 15436 3544 15442 3556
rect 16022 3544 16028 3556
rect 16080 3544 16086 3596
rect 24670 3593 24676 3596
rect 24648 3587 24676 3593
rect 24648 3584 24660 3587
rect 24583 3556 24660 3584
rect 24648 3553 24660 3556
rect 24728 3584 24734 3596
rect 27614 3584 27620 3596
rect 24728 3556 27620 3584
rect 24648 3547 24676 3553
rect 24670 3544 24676 3547
rect 24728 3544 24734 3556
rect 27614 3544 27620 3556
rect 27672 3544 27678 3596
rect 14274 3448 14280 3460
rect 14187 3420 14280 3448
rect 14274 3408 14280 3420
rect 14332 3448 14338 3460
rect 24719 3451 24777 3457
rect 24719 3448 24731 3451
rect 14332 3420 24731 3448
rect 14332 3408 14338 3420
rect 24719 3417 24731 3420
rect 24765 3417 24777 3451
rect 24719 3411 24777 3417
rect 15427 3383 15485 3389
rect 15427 3349 15439 3383
rect 15473 3380 15485 3383
rect 15654 3380 15660 3392
rect 15473 3352 15660 3380
rect 15473 3349 15485 3352
rect 15427 3343 15485 3349
rect 15654 3340 15660 3352
rect 15712 3340 15718 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 9769 3179 9827 3185
rect 9769 3176 9781 3179
rect 9140 3148 9781 3176
rect 106 3068 112 3120
rect 164 3108 170 3120
rect 1394 3108 1400 3120
rect 164 3080 1400 3108
rect 164 3068 170 3080
rect 1394 3068 1400 3080
rect 1452 3108 1458 3120
rect 1581 3111 1639 3117
rect 1581 3108 1593 3111
rect 1452 3080 1593 3108
rect 1452 3068 1458 3080
rect 1581 3077 1593 3080
rect 1627 3077 1639 3111
rect 1581 3071 1639 3077
rect 9140 2981 9168 3148
rect 9769 3145 9781 3148
rect 9815 3176 9827 3179
rect 9858 3176 9864 3188
rect 9815 3148 9864 3176
rect 9815 3145 9827 3148
rect 9769 3139 9827 3145
rect 9858 3136 9864 3148
rect 9916 3136 9922 3188
rect 11425 3179 11483 3185
rect 11425 3176 11437 3179
rect 10888 3148 11437 3176
rect 9309 3111 9367 3117
rect 9309 3077 9321 3111
rect 9355 3108 9367 3111
rect 10778 3108 10784 3120
rect 9355 3080 10784 3108
rect 9355 3077 9367 3080
rect 9309 3071 9367 3077
rect 10778 3068 10784 3080
rect 10836 3068 10842 3120
rect 9125 2975 9183 2981
rect 9125 2941 9137 2975
rect 9171 2941 9183 2975
rect 9125 2935 9183 2941
rect 10781 2975 10839 2981
rect 10781 2941 10793 2975
rect 10827 2972 10839 2975
rect 10888 2972 10916 3148
rect 11425 3145 11437 3148
rect 11471 3176 11483 3179
rect 11974 3176 11980 3188
rect 11471 3148 11980 3176
rect 11471 3145 11483 3148
rect 11425 3139 11483 3145
rect 11974 3136 11980 3148
rect 12032 3136 12038 3188
rect 15378 3176 15384 3188
rect 15339 3148 15384 3176
rect 15378 3136 15384 3148
rect 15436 3136 15442 3188
rect 24670 3176 24676 3188
rect 24631 3148 24676 3176
rect 24670 3136 24676 3148
rect 24728 3136 24734 3188
rect 10965 3111 11023 3117
rect 10965 3077 10977 3111
rect 11011 3108 11023 3111
rect 12066 3108 12072 3120
rect 11011 3080 12072 3108
rect 11011 3077 11023 3080
rect 10965 3071 11023 3077
rect 12066 3068 12072 3080
rect 12124 3068 12130 3120
rect 13906 3068 13912 3120
rect 13964 3108 13970 3120
rect 23106 3108 23112 3120
rect 13964 3080 23112 3108
rect 13964 3068 13970 3080
rect 23106 3068 23112 3080
rect 23164 3068 23170 3120
rect 15654 2972 15660 2984
rect 10827 2944 10916 2972
rect 15615 2944 15660 2972
rect 10827 2941 10839 2944
rect 10781 2935 10839 2941
rect 15654 2932 15660 2944
rect 15712 2972 15718 2984
rect 16209 2975 16267 2981
rect 16209 2972 16221 2975
rect 15712 2944 16221 2972
rect 15712 2932 15718 2944
rect 16209 2941 16221 2944
rect 16255 2941 16267 2975
rect 16209 2935 16267 2941
rect 15841 2839 15899 2845
rect 15841 2805 15853 2839
rect 15887 2836 15899 2839
rect 16758 2836 16764 2848
rect 15887 2808 16764 2836
rect 15887 2805 15899 2808
rect 15841 2799 15899 2805
rect 16758 2796 16764 2808
rect 16816 2796 16822 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 842 2592 848 2644
rect 900 2632 906 2644
rect 1486 2632 1492 2644
rect 900 2604 1492 2632
rect 900 2592 906 2604
rect 1486 2592 1492 2604
rect 1544 2592 1550 2644
rect 14826 2632 14832 2644
rect 14787 2604 14832 2632
rect 14826 2592 14832 2604
rect 14884 2592 14890 2644
rect 16255 2635 16313 2641
rect 16255 2601 16267 2635
rect 16301 2632 16313 2635
rect 16390 2632 16396 2644
rect 16301 2604 16396 2632
rect 16301 2601 16313 2604
rect 16255 2595 16313 2601
rect 16390 2592 16396 2604
rect 16448 2592 16454 2644
rect 20254 2592 20260 2644
rect 20312 2632 20318 2644
rect 20349 2635 20407 2641
rect 20349 2632 20361 2635
rect 20312 2604 20361 2632
rect 20312 2592 20318 2604
rect 20349 2601 20361 2604
rect 20395 2601 20407 2635
rect 20349 2595 20407 2601
rect 21358 2592 21364 2644
rect 21416 2632 21422 2644
rect 22787 2635 22845 2641
rect 22787 2632 22799 2635
rect 21416 2604 22799 2632
rect 21416 2592 21422 2604
rect 22787 2601 22799 2604
rect 22833 2601 22845 2635
rect 22787 2595 22845 2601
rect 6917 2499 6975 2505
rect 6917 2465 6929 2499
rect 6963 2496 6975 2499
rect 7558 2496 7564 2508
rect 6963 2468 7564 2496
rect 6963 2465 6975 2468
rect 6917 2459 6975 2465
rect 7558 2456 7564 2468
rect 7616 2456 7622 2508
rect 8938 2456 8944 2508
rect 8996 2496 9002 2508
rect 11149 2499 11207 2505
rect 11149 2496 11161 2499
rect 8996 2468 11161 2496
rect 8996 2456 9002 2468
rect 11149 2465 11161 2468
rect 11195 2496 11207 2499
rect 11701 2499 11759 2505
rect 11701 2496 11713 2499
rect 11195 2468 11713 2496
rect 11195 2465 11207 2468
rect 11149 2459 11207 2465
rect 11701 2465 11713 2468
rect 11747 2465 11759 2499
rect 11701 2459 11759 2465
rect 14277 2499 14335 2505
rect 14277 2465 14289 2499
rect 14323 2496 14335 2499
rect 14844 2496 14872 2592
rect 23201 2567 23259 2573
rect 23201 2533 23213 2567
rect 23247 2564 23259 2567
rect 24762 2564 24768 2576
rect 23247 2536 24768 2564
rect 23247 2533 23259 2536
rect 23201 2527 23259 2533
rect 14323 2468 14872 2496
rect 16184 2499 16242 2505
rect 14323 2465 14335 2468
rect 14277 2459 14335 2465
rect 16184 2465 16196 2499
rect 16230 2496 16242 2499
rect 16666 2496 16672 2508
rect 16230 2468 16672 2496
rect 16230 2465 16242 2468
rect 16184 2459 16242 2465
rect 16666 2456 16672 2468
rect 16724 2456 16730 2508
rect 20140 2499 20198 2505
rect 20140 2465 20152 2499
rect 20186 2496 20198 2499
rect 21612 2499 21670 2505
rect 20186 2468 20668 2496
rect 20186 2465 20198 2468
rect 20140 2459 20198 2465
rect 4706 2320 4712 2372
rect 4764 2360 4770 2372
rect 8938 2360 8944 2372
rect 4764 2332 8944 2360
rect 4764 2320 4770 2332
rect 8938 2320 8944 2332
rect 8996 2320 9002 2372
rect 11333 2363 11391 2369
rect 11333 2329 11345 2363
rect 11379 2360 11391 2363
rect 13354 2360 13360 2372
rect 11379 2332 13360 2360
rect 11379 2329 11391 2332
rect 11333 2323 11391 2329
rect 13354 2320 13360 2332
rect 13412 2320 13418 2372
rect 20640 2369 20668 2468
rect 21612 2465 21624 2499
rect 21658 2496 21670 2499
rect 22716 2499 22774 2505
rect 21658 2468 22140 2496
rect 21658 2465 21670 2468
rect 21612 2459 21670 2465
rect 20625 2363 20683 2369
rect 20625 2329 20637 2363
rect 20671 2360 20683 2363
rect 21818 2360 21824 2372
rect 20671 2332 21824 2360
rect 20671 2329 20683 2332
rect 20625 2323 20683 2329
rect 21818 2320 21824 2332
rect 21876 2320 21882 2372
rect 6822 2252 6828 2304
rect 6880 2292 6886 2304
rect 7101 2295 7159 2301
rect 7101 2292 7113 2295
rect 6880 2264 7113 2292
rect 6880 2252 6886 2264
rect 7101 2261 7113 2264
rect 7147 2261 7159 2295
rect 7101 2255 7159 2261
rect 14461 2295 14519 2301
rect 14461 2261 14473 2295
rect 14507 2292 14519 2295
rect 14642 2292 14648 2304
rect 14507 2264 14648 2292
rect 14507 2261 14519 2264
rect 14461 2255 14519 2261
rect 14642 2252 14648 2264
rect 14700 2252 14706 2304
rect 16666 2292 16672 2304
rect 16627 2264 16672 2292
rect 16666 2252 16672 2264
rect 16724 2252 16730 2304
rect 17678 2252 17684 2304
rect 17736 2292 17742 2304
rect 22112 2301 22140 2468
rect 22716 2465 22728 2499
rect 22762 2496 22774 2499
rect 23216 2496 23244 2527
rect 24762 2524 24768 2536
rect 24820 2524 24826 2576
rect 22762 2468 23244 2496
rect 24096 2499 24154 2505
rect 22762 2465 22774 2468
rect 22716 2459 22774 2465
rect 24096 2465 24108 2499
rect 24142 2496 24154 2499
rect 24142 2468 24624 2496
rect 24142 2465 24154 2468
rect 24096 2459 24154 2465
rect 21683 2295 21741 2301
rect 21683 2292 21695 2295
rect 17736 2264 21695 2292
rect 17736 2252 17742 2264
rect 21683 2261 21695 2264
rect 21729 2261 21741 2295
rect 21683 2255 21741 2261
rect 22097 2295 22155 2301
rect 22097 2261 22109 2295
rect 22143 2292 22155 2295
rect 23014 2292 23020 2304
rect 22143 2264 23020 2292
rect 22143 2261 22155 2264
rect 22097 2255 22155 2261
rect 23014 2252 23020 2264
rect 23072 2252 23078 2304
rect 23106 2252 23112 2304
rect 23164 2292 23170 2304
rect 24596 2301 24624 2468
rect 24167 2295 24225 2301
rect 24167 2292 24179 2295
rect 23164 2264 24179 2292
rect 23164 2252 23170 2264
rect 24167 2261 24179 2264
rect 24213 2261 24225 2295
rect 24167 2255 24225 2261
rect 24581 2295 24639 2301
rect 24581 2261 24593 2295
rect 24627 2292 24639 2295
rect 25590 2292 25596 2304
rect 24627 2264 25596 2292
rect 24627 2261 24639 2264
rect 24581 2255 24639 2261
rect 25590 2252 25596 2264
rect 25648 2252 25654 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 18230 416 18236 468
rect 18288 456 18294 468
rect 19334 456 19340 468
rect 18288 428 19340 456
rect 18288 416 18294 428
rect 19334 416 19340 428
rect 19392 416 19398 468
rect 15746 76 15752 128
rect 15804 116 15810 128
rect 17402 116 17408 128
rect 15804 88 17408 116
rect 15804 76 15810 88
rect 17402 76 17408 88
rect 17460 76 17466 128
<< via1 >>
rect 20 27480 72 27532
rect 664 27480 716 27532
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 11612 24828 11664 24880
rect 27620 24828 27672 24880
rect 11244 24556 11296 24608
rect 13176 24556 13228 24608
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 7472 24395 7524 24404
rect 7472 24361 7481 24395
rect 7481 24361 7515 24395
rect 7515 24361 7524 24395
rect 7472 24352 7524 24361
rect 7288 24259 7340 24268
rect 7288 24225 7297 24259
rect 7297 24225 7331 24259
rect 7331 24225 7340 24259
rect 7288 24216 7340 24225
rect 11612 24216 11664 24268
rect 10048 24012 10100 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 9036 23808 9088 23860
rect 11428 23808 11480 23860
rect 11612 23851 11664 23860
rect 11612 23817 11621 23851
rect 11621 23817 11655 23851
rect 11655 23817 11664 23851
rect 11612 23808 11664 23817
rect 20168 23808 20220 23860
rect 11244 23783 11296 23792
rect 11244 23749 11253 23783
rect 11253 23749 11287 23783
rect 11287 23749 11296 23783
rect 11244 23740 11296 23749
rect 1308 23672 1360 23724
rect 7840 23647 7892 23656
rect 7840 23613 7849 23647
rect 7849 23613 7883 23647
rect 7883 23613 7892 23647
rect 7840 23604 7892 23613
rect 11244 23604 11296 23656
rect 16396 23604 16448 23656
rect 16488 23647 16540 23656
rect 16488 23613 16497 23647
rect 16497 23613 16531 23647
rect 16531 23613 16540 23647
rect 18144 23647 18196 23656
rect 16488 23604 16540 23613
rect 18144 23613 18153 23647
rect 18153 23613 18187 23647
rect 18187 23613 18196 23647
rect 18144 23604 18196 23613
rect 21640 23808 21692 23860
rect 23020 23808 23072 23860
rect 22284 23740 22336 23792
rect 19432 23536 19484 23588
rect 27160 23808 27212 23860
rect 25780 23536 25832 23588
rect 1676 23468 1728 23520
rect 7288 23468 7340 23520
rect 7748 23468 7800 23520
rect 19984 23468 20036 23520
rect 22560 23468 22612 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 15660 23239 15712 23248
rect 15660 23205 15669 23239
rect 15669 23205 15703 23239
rect 15703 23205 15712 23239
rect 15660 23196 15712 23205
rect 1216 23128 1268 23180
rect 2228 23128 2280 23180
rect 8484 23128 8536 23180
rect 13636 23171 13688 23180
rect 13636 23137 13645 23171
rect 13645 23137 13679 23171
rect 13679 23137 13688 23171
rect 13636 23128 13688 23137
rect 14096 23171 14148 23180
rect 14096 23137 14105 23171
rect 14105 23137 14139 23171
rect 14139 23137 14148 23171
rect 14096 23128 14148 23137
rect 16304 23128 16356 23180
rect 17316 23128 17368 23180
rect 20996 23171 21048 23180
rect 20996 23137 21014 23171
rect 21014 23137 21048 23171
rect 20996 23128 21048 23137
rect 24124 23128 24176 23180
rect 14280 23103 14332 23112
rect 14280 23069 14289 23103
rect 14289 23069 14323 23103
rect 14323 23069 14332 23103
rect 14280 23060 14332 23069
rect 16396 23060 16448 23112
rect 10968 22992 11020 23044
rect 14372 22992 14424 23044
rect 12440 22924 12492 22976
rect 12716 22967 12768 22976
rect 12716 22933 12725 22967
rect 12725 22933 12759 22967
rect 12759 22933 12768 22967
rect 12716 22924 12768 22933
rect 14648 22967 14700 22976
rect 14648 22933 14657 22967
rect 14657 22933 14691 22967
rect 14691 22933 14700 22967
rect 14648 22924 14700 22933
rect 17408 22924 17460 22976
rect 21180 22924 21232 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 2228 22763 2280 22772
rect 2228 22729 2237 22763
rect 2237 22729 2271 22763
rect 2271 22729 2280 22763
rect 2228 22720 2280 22729
rect 14096 22763 14148 22772
rect 14096 22729 14105 22763
rect 14105 22729 14139 22763
rect 14139 22729 14148 22763
rect 14096 22720 14148 22729
rect 14464 22763 14516 22772
rect 14464 22729 14473 22763
rect 14473 22729 14507 22763
rect 14507 22729 14516 22763
rect 14464 22720 14516 22729
rect 16396 22763 16448 22772
rect 16396 22729 16405 22763
rect 16405 22729 16439 22763
rect 16439 22729 16448 22763
rect 16396 22720 16448 22729
rect 20996 22763 21048 22772
rect 20996 22729 21005 22763
rect 21005 22729 21039 22763
rect 21039 22729 21048 22763
rect 20996 22720 21048 22729
rect 13268 22627 13320 22636
rect 13268 22593 13277 22627
rect 13277 22593 13311 22627
rect 13311 22593 13320 22627
rect 13268 22584 13320 22593
rect 112 22516 164 22568
rect 12716 22559 12768 22568
rect 12716 22525 12725 22559
rect 12725 22525 12759 22559
rect 12759 22525 12768 22559
rect 12716 22516 12768 22525
rect 14096 22516 14148 22568
rect 1768 22380 1820 22432
rect 8484 22380 8536 22432
rect 12256 22423 12308 22432
rect 12256 22389 12265 22423
rect 12265 22389 12299 22423
rect 12299 22389 12308 22423
rect 12256 22380 12308 22389
rect 13636 22380 13688 22432
rect 17316 22516 17368 22568
rect 14464 22448 14516 22500
rect 15660 22448 15712 22500
rect 16120 22491 16172 22500
rect 16120 22457 16129 22491
rect 16129 22457 16163 22491
rect 16163 22457 16172 22491
rect 16120 22448 16172 22457
rect 14648 22380 14700 22432
rect 15384 22380 15436 22432
rect 16948 22380 17000 22432
rect 17776 22380 17828 22432
rect 18420 22380 18472 22432
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 12440 22176 12492 22228
rect 13820 22151 13872 22160
rect 13820 22117 13829 22151
rect 13829 22117 13863 22151
rect 13863 22117 13872 22151
rect 13820 22108 13872 22117
rect 17408 22108 17460 22160
rect 18512 22151 18564 22160
rect 18512 22117 18521 22151
rect 18521 22117 18555 22151
rect 18555 22117 18564 22151
rect 18512 22108 18564 22117
rect 12164 22040 12216 22092
rect 14372 22083 14424 22092
rect 14372 22049 14381 22083
rect 14381 22049 14415 22083
rect 14415 22049 14424 22083
rect 16948 22083 17000 22092
rect 14372 22040 14424 22049
rect 16948 22049 16957 22083
rect 16957 22049 16991 22083
rect 16991 22049 17000 22083
rect 16948 22040 17000 22049
rect 16120 22015 16172 22024
rect 15292 21904 15344 21956
rect 16120 21981 16129 22015
rect 16129 21981 16163 22015
rect 16163 21981 16172 22015
rect 16120 21972 16172 21981
rect 16672 21972 16724 22024
rect 19064 22015 19116 22024
rect 19064 21981 19073 22015
rect 19073 21981 19107 22015
rect 19107 21981 19116 22015
rect 19064 21972 19116 21981
rect 13176 21836 13228 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 12164 21675 12216 21684
rect 12164 21641 12173 21675
rect 12173 21641 12207 21675
rect 12207 21641 12216 21675
rect 12164 21632 12216 21641
rect 16948 21675 17000 21684
rect 16948 21641 16957 21675
rect 16957 21641 16991 21675
rect 16991 21641 17000 21675
rect 16948 21632 17000 21641
rect 17408 21675 17460 21684
rect 17408 21641 17417 21675
rect 17417 21641 17451 21675
rect 17451 21641 17460 21675
rect 17408 21632 17460 21641
rect 24768 21675 24820 21684
rect 24768 21641 24777 21675
rect 24777 21641 24811 21675
rect 24811 21641 24820 21675
rect 24768 21632 24820 21641
rect 14648 21496 14700 21548
rect 16396 21496 16448 21548
rect 18420 21496 18472 21548
rect 12624 21471 12676 21480
rect 12624 21437 12633 21471
rect 12633 21437 12667 21471
rect 12667 21437 12676 21471
rect 12624 21428 12676 21437
rect 12900 21428 12952 21480
rect 23848 21428 23900 21480
rect 12256 21360 12308 21412
rect 13360 21403 13412 21412
rect 13360 21369 13369 21403
rect 13369 21369 13403 21403
rect 13403 21369 13412 21403
rect 13360 21360 13412 21369
rect 13820 21292 13872 21344
rect 14188 21335 14240 21344
rect 14188 21301 14197 21335
rect 14197 21301 14231 21335
rect 14231 21301 14240 21335
rect 15200 21360 15252 21412
rect 14188 21292 14240 21301
rect 15476 21292 15528 21344
rect 16672 21403 16724 21412
rect 16672 21369 16681 21403
rect 16681 21369 16715 21403
rect 16715 21369 16724 21403
rect 16672 21360 16724 21369
rect 18972 21360 19024 21412
rect 19248 21403 19300 21412
rect 19248 21369 19257 21403
rect 19257 21369 19291 21403
rect 19291 21369 19300 21403
rect 19248 21360 19300 21369
rect 17868 21335 17920 21344
rect 17868 21301 17877 21335
rect 17877 21301 17911 21335
rect 17911 21301 17920 21335
rect 17868 21292 17920 21301
rect 19432 21292 19484 21344
rect 20352 21292 20404 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 13360 21088 13412 21140
rect 15292 21088 15344 21140
rect 15384 21088 15436 21140
rect 1216 21020 1268 21072
rect 11520 21063 11572 21072
rect 11520 21029 11529 21063
rect 11529 21029 11563 21063
rect 11563 21029 11572 21063
rect 11520 21020 11572 21029
rect 13176 21020 13228 21072
rect 13728 21063 13780 21072
rect 13728 21029 13737 21063
rect 13737 21029 13771 21063
rect 13771 21029 13780 21063
rect 13728 21020 13780 21029
rect 14464 21020 14516 21072
rect 15476 21063 15528 21072
rect 15476 21029 15485 21063
rect 15485 21029 15519 21063
rect 15519 21029 15528 21063
rect 15476 21020 15528 21029
rect 17868 21020 17920 21072
rect 18512 21063 18564 21072
rect 18512 21029 18521 21063
rect 18521 21029 18555 21063
rect 18555 21029 18564 21063
rect 18512 21020 18564 21029
rect 19248 21020 19300 21072
rect 20076 21020 20128 21072
rect 9588 20952 9640 21004
rect 17408 20952 17460 21004
rect 24676 20995 24728 21004
rect 24676 20961 24694 20995
rect 24694 20961 24728 20995
rect 24676 20952 24728 20961
rect 25136 20952 25188 21004
rect 8300 20927 8352 20936
rect 8300 20893 8309 20927
rect 8309 20893 8343 20927
rect 8343 20893 8352 20927
rect 8300 20884 8352 20893
rect 10048 20884 10100 20936
rect 11060 20884 11112 20936
rect 11796 20884 11848 20936
rect 12808 20884 12860 20936
rect 15384 20927 15436 20936
rect 15384 20893 15393 20927
rect 15393 20893 15427 20927
rect 15427 20893 15436 20927
rect 15384 20884 15436 20893
rect 15292 20816 15344 20868
rect 17776 20884 17828 20936
rect 18052 20816 18104 20868
rect 19984 20816 20036 20868
rect 7656 20748 7708 20800
rect 8852 20791 8904 20800
rect 8852 20757 8861 20791
rect 8861 20757 8895 20791
rect 8895 20757 8904 20791
rect 8852 20748 8904 20757
rect 10048 20748 10100 20800
rect 10324 20791 10376 20800
rect 10324 20757 10333 20791
rect 10333 20757 10367 20791
rect 10367 20757 10376 20791
rect 10324 20748 10376 20757
rect 11612 20748 11664 20800
rect 12624 20791 12676 20800
rect 12624 20757 12633 20791
rect 12633 20757 12667 20791
rect 12667 20757 12676 20791
rect 12624 20748 12676 20757
rect 14648 20791 14700 20800
rect 14648 20757 14657 20791
rect 14657 20757 14691 20791
rect 14691 20757 14700 20791
rect 14648 20748 14700 20757
rect 16396 20791 16448 20800
rect 16396 20757 16405 20791
rect 16405 20757 16439 20791
rect 16439 20757 16448 20791
rect 16396 20748 16448 20757
rect 18604 20748 18656 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 1216 20544 1268 20596
rect 4068 20587 4120 20596
rect 4068 20553 4077 20587
rect 4077 20553 4111 20587
rect 4111 20553 4120 20587
rect 4068 20544 4120 20553
rect 11520 20544 11572 20596
rect 13728 20544 13780 20596
rect 15384 20587 15436 20596
rect 10232 20476 10284 20528
rect 12716 20476 12768 20528
rect 13544 20476 13596 20528
rect 14464 20519 14516 20528
rect 14464 20485 14473 20519
rect 14473 20485 14507 20519
rect 14507 20485 14516 20519
rect 14464 20476 14516 20485
rect 4160 20408 4212 20460
rect 7840 20408 7892 20460
rect 6368 20340 6420 20392
rect 11612 20408 11664 20460
rect 11796 20451 11848 20460
rect 11796 20417 11805 20451
rect 11805 20417 11839 20451
rect 11839 20417 11848 20451
rect 11796 20408 11848 20417
rect 13360 20408 13412 20460
rect 15384 20553 15393 20587
rect 15393 20553 15427 20587
rect 15427 20553 15436 20587
rect 15384 20544 15436 20553
rect 17776 20587 17828 20596
rect 17776 20553 17785 20587
rect 17785 20553 17819 20587
rect 17819 20553 17828 20587
rect 17776 20544 17828 20553
rect 18512 20544 18564 20596
rect 24676 20587 24728 20596
rect 24676 20553 24685 20587
rect 24685 20553 24719 20587
rect 24719 20553 24728 20587
rect 24676 20544 24728 20553
rect 20536 20476 20588 20528
rect 21180 20408 21232 20460
rect 8852 20340 8904 20392
rect 10232 20383 10284 20392
rect 9772 20272 9824 20324
rect 10232 20349 10241 20383
rect 10241 20349 10275 20383
rect 10275 20349 10284 20383
rect 10232 20340 10284 20349
rect 10324 20340 10376 20392
rect 11244 20340 11296 20392
rect 12624 20340 12676 20392
rect 16304 20340 16356 20392
rect 19064 20340 19116 20392
rect 13728 20272 13780 20324
rect 16488 20315 16540 20324
rect 16488 20281 16497 20315
rect 16497 20281 16531 20315
rect 16531 20281 16540 20315
rect 16488 20272 16540 20281
rect 8944 20247 8996 20256
rect 8944 20213 8953 20247
rect 8953 20213 8987 20247
rect 8987 20213 8996 20247
rect 8944 20204 8996 20213
rect 9588 20204 9640 20256
rect 10140 20204 10192 20256
rect 10876 20204 10928 20256
rect 13360 20204 13412 20256
rect 15476 20204 15528 20256
rect 19524 20315 19576 20324
rect 19524 20281 19533 20315
rect 19533 20281 19567 20315
rect 19567 20281 19576 20315
rect 19524 20272 19576 20281
rect 17224 20204 17276 20256
rect 17408 20247 17460 20256
rect 17408 20213 17417 20247
rect 17417 20213 17451 20247
rect 17451 20213 17460 20247
rect 17408 20204 17460 20213
rect 19984 20204 20036 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 7656 20000 7708 20052
rect 4344 19932 4396 19984
rect 7840 20000 7892 20052
rect 8852 20000 8904 20052
rect 14188 20043 14240 20052
rect 14188 20009 14197 20043
rect 14197 20009 14231 20043
rect 14231 20009 14240 20043
rect 14188 20000 14240 20009
rect 14280 20000 14332 20052
rect 16396 20000 16448 20052
rect 18328 20043 18380 20052
rect 18328 20009 18337 20043
rect 18337 20009 18371 20043
rect 18371 20009 18380 20043
rect 18328 20000 18380 20009
rect 18512 20000 18564 20052
rect 19524 20000 19576 20052
rect 24768 20043 24820 20052
rect 24768 20009 24777 20043
rect 24777 20009 24811 20043
rect 24811 20009 24820 20043
rect 24768 20000 24820 20009
rect 8116 19975 8168 19984
rect 8116 19941 8125 19975
rect 8125 19941 8159 19975
rect 8159 19941 8168 19975
rect 8116 19932 8168 19941
rect 10232 19932 10284 19984
rect 13360 19932 13412 19984
rect 13728 19932 13780 19984
rect 15752 19932 15804 19984
rect 6276 19864 6328 19916
rect 10140 19864 10192 19916
rect 11888 19864 11940 19916
rect 13268 19907 13320 19916
rect 13268 19873 13277 19907
rect 13277 19873 13311 19907
rect 13311 19873 13320 19907
rect 13268 19864 13320 19873
rect 17132 19864 17184 19916
rect 19432 19864 19484 19916
rect 20996 19864 21048 19916
rect 24676 19864 24728 19916
rect 3976 19796 4028 19848
rect 3884 19728 3936 19780
rect 5448 19796 5500 19848
rect 6000 19796 6052 19848
rect 8852 19796 8904 19848
rect 5356 19728 5408 19780
rect 15292 19728 15344 19780
rect 16396 19796 16448 19848
rect 17408 19796 17460 19848
rect 17960 19839 18012 19848
rect 17960 19805 17969 19839
rect 17969 19805 18003 19839
rect 18003 19805 18012 19839
rect 17960 19796 18012 19805
rect 16488 19771 16540 19780
rect 16488 19737 16497 19771
rect 16497 19737 16531 19771
rect 16531 19737 16540 19771
rect 16488 19728 16540 19737
rect 5080 19660 5132 19712
rect 6000 19660 6052 19712
rect 11152 19660 11204 19712
rect 11336 19703 11388 19712
rect 11336 19669 11345 19703
rect 11345 19669 11379 19703
rect 11379 19669 11388 19703
rect 11336 19660 11388 19669
rect 12532 19660 12584 19712
rect 20260 19703 20312 19712
rect 20260 19669 20269 19703
rect 20269 19669 20303 19703
rect 20303 19669 20312 19703
rect 20260 19660 20312 19669
rect 21364 19703 21416 19712
rect 21364 19669 21373 19703
rect 21373 19669 21407 19703
rect 21407 19669 21416 19703
rect 21364 19660 21416 19669
rect 21824 19703 21876 19712
rect 21824 19669 21833 19703
rect 21833 19669 21867 19703
rect 21867 19669 21876 19703
rect 21824 19660 21876 19669
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 1584 19499 1636 19508
rect 1584 19465 1593 19499
rect 1593 19465 1627 19499
rect 1627 19465 1636 19499
rect 1584 19456 1636 19465
rect 3976 19456 4028 19508
rect 4160 19499 4212 19508
rect 4160 19465 4169 19499
rect 4169 19465 4203 19499
rect 4203 19465 4212 19499
rect 6276 19499 6328 19508
rect 4160 19456 4212 19465
rect 6276 19465 6285 19499
rect 6285 19465 6319 19499
rect 6319 19465 6328 19499
rect 6276 19456 6328 19465
rect 8300 19499 8352 19508
rect 8300 19465 8309 19499
rect 8309 19465 8343 19499
rect 8343 19465 8352 19499
rect 8300 19456 8352 19465
rect 10140 19456 10192 19508
rect 11520 19499 11572 19508
rect 11520 19465 11529 19499
rect 11529 19465 11563 19499
rect 11563 19465 11572 19499
rect 11520 19456 11572 19465
rect 17224 19456 17276 19508
rect 5080 19363 5132 19372
rect 5080 19329 5089 19363
rect 5089 19329 5123 19363
rect 5123 19329 5132 19363
rect 5080 19320 5132 19329
rect 5356 19363 5408 19372
rect 5356 19329 5365 19363
rect 5365 19329 5399 19363
rect 5399 19329 5408 19363
rect 5356 19320 5408 19329
rect 10232 19388 10284 19440
rect 10876 19388 10928 19440
rect 8852 19363 8904 19372
rect 8852 19329 8861 19363
rect 8861 19329 8895 19363
rect 8895 19329 8904 19363
rect 8852 19320 8904 19329
rect 11888 19431 11940 19440
rect 11888 19397 11897 19431
rect 11897 19397 11931 19431
rect 11931 19397 11940 19431
rect 17132 19431 17184 19440
rect 11888 19388 11940 19397
rect 12532 19363 12584 19372
rect 3884 19184 3936 19236
rect 7196 19295 7248 19304
rect 7196 19261 7205 19295
rect 7205 19261 7239 19295
rect 7239 19261 7248 19295
rect 7196 19252 7248 19261
rect 7472 19295 7524 19304
rect 7472 19261 7481 19295
rect 7481 19261 7515 19295
rect 7515 19261 7524 19295
rect 7472 19252 7524 19261
rect 7840 19252 7892 19304
rect 5172 19227 5224 19236
rect 5172 19193 5181 19227
rect 5181 19193 5215 19227
rect 5215 19193 5224 19227
rect 5172 19184 5224 19193
rect 7656 19227 7708 19236
rect 7656 19193 7665 19227
rect 7665 19193 7699 19227
rect 7699 19193 7708 19227
rect 7656 19184 7708 19193
rect 8576 19184 8628 19236
rect 12532 19329 12541 19363
rect 12541 19329 12575 19363
rect 12575 19329 12584 19363
rect 12532 19320 12584 19329
rect 12808 19363 12860 19372
rect 12808 19329 12817 19363
rect 12817 19329 12851 19363
rect 12851 19329 12860 19363
rect 12808 19320 12860 19329
rect 13452 19363 13504 19372
rect 13452 19329 13461 19363
rect 13461 19329 13495 19363
rect 13495 19329 13504 19363
rect 13452 19320 13504 19329
rect 14280 19363 14332 19372
rect 14280 19329 14289 19363
rect 14289 19329 14323 19363
rect 14323 19329 14332 19363
rect 14280 19320 14332 19329
rect 16396 19363 16448 19372
rect 16396 19329 16405 19363
rect 16405 19329 16439 19363
rect 16439 19329 16448 19363
rect 16396 19320 16448 19329
rect 17132 19397 17141 19431
rect 17141 19397 17175 19431
rect 17175 19397 17184 19431
rect 17132 19388 17184 19397
rect 20996 19388 21048 19440
rect 18788 19320 18840 19372
rect 19432 19320 19484 19372
rect 20260 19320 20312 19372
rect 23388 19320 23440 19372
rect 24676 19320 24728 19372
rect 11336 19252 11388 19304
rect 10876 19227 10928 19236
rect 1952 19159 2004 19168
rect 1952 19125 1961 19159
rect 1961 19125 1995 19159
rect 1995 19125 2004 19159
rect 1952 19116 2004 19125
rect 4344 19116 4396 19168
rect 8116 19116 8168 19168
rect 10140 19159 10192 19168
rect 10140 19125 10149 19159
rect 10149 19125 10183 19159
rect 10183 19125 10192 19159
rect 10140 19116 10192 19125
rect 10876 19193 10885 19227
rect 10885 19193 10919 19227
rect 10919 19193 10928 19227
rect 10876 19184 10928 19193
rect 11152 19184 11204 19236
rect 15752 19184 15804 19236
rect 16120 19227 16172 19236
rect 16120 19193 16129 19227
rect 16129 19193 16163 19227
rect 16163 19193 16172 19227
rect 16120 19184 16172 19193
rect 13452 19116 13504 19168
rect 15476 19116 15528 19168
rect 15660 19116 15712 19168
rect 21364 19252 21416 19304
rect 21824 19295 21876 19304
rect 18328 19184 18380 19236
rect 19984 19227 20036 19236
rect 19984 19193 19993 19227
rect 19993 19193 20027 19227
rect 20027 19193 20036 19227
rect 19984 19184 20036 19193
rect 20076 19184 20128 19236
rect 20812 19184 20864 19236
rect 21824 19261 21833 19295
rect 21833 19261 21867 19295
rect 21867 19261 21876 19295
rect 21824 19252 21876 19261
rect 23480 19184 23532 19236
rect 17408 19159 17460 19168
rect 17408 19125 17417 19159
rect 17417 19125 17451 19159
rect 17451 19125 17460 19159
rect 17408 19116 17460 19125
rect 17776 19159 17828 19168
rect 17776 19125 17785 19159
rect 17785 19125 17819 19159
rect 17819 19125 17828 19159
rect 20996 19159 21048 19168
rect 17776 19116 17828 19125
rect 20996 19125 21005 19159
rect 21005 19125 21039 19159
rect 21039 19125 21048 19159
rect 20996 19116 21048 19125
rect 21456 19159 21508 19168
rect 21456 19125 21465 19159
rect 21465 19125 21499 19159
rect 21499 19125 21508 19159
rect 21456 19116 21508 19125
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 3976 18912 4028 18964
rect 5080 18912 5132 18964
rect 5540 18912 5592 18964
rect 6092 18844 6144 18896
rect 7472 18912 7524 18964
rect 8116 18912 8168 18964
rect 8576 18955 8628 18964
rect 8576 18921 8585 18955
rect 8585 18921 8619 18955
rect 8619 18921 8628 18955
rect 8576 18912 8628 18921
rect 8944 18955 8996 18964
rect 8944 18921 8953 18955
rect 8953 18921 8987 18955
rect 8987 18921 8996 18955
rect 8944 18912 8996 18921
rect 11336 18912 11388 18964
rect 13268 18912 13320 18964
rect 14648 18912 14700 18964
rect 15200 18912 15252 18964
rect 16120 18912 16172 18964
rect 16672 18955 16724 18964
rect 16672 18921 16681 18955
rect 16681 18921 16715 18955
rect 16715 18921 16724 18955
rect 16672 18912 16724 18921
rect 17960 18912 18012 18964
rect 21456 18912 21508 18964
rect 10508 18844 10560 18896
rect 15384 18844 15436 18896
rect 16396 18844 16448 18896
rect 19340 18844 19392 18896
rect 4712 18776 4764 18828
rect 9680 18776 9732 18828
rect 11796 18776 11848 18828
rect 12992 18776 13044 18828
rect 14280 18776 14332 18828
rect 16304 18776 16356 18828
rect 17224 18819 17276 18828
rect 17224 18785 17233 18819
rect 17233 18785 17267 18819
rect 17267 18785 17276 18819
rect 17224 18776 17276 18785
rect 20904 18819 20956 18828
rect 20904 18785 20913 18819
rect 20913 18785 20947 18819
rect 20947 18785 20956 18819
rect 20904 18776 20956 18785
rect 21180 18776 21232 18828
rect 6000 18708 6052 18760
rect 7564 18751 7616 18760
rect 7564 18717 7573 18751
rect 7573 18717 7607 18751
rect 7607 18717 7616 18751
rect 7564 18708 7616 18717
rect 7840 18751 7892 18760
rect 7840 18717 7849 18751
rect 7849 18717 7883 18751
rect 7883 18717 7892 18751
rect 7840 18708 7892 18717
rect 5264 18640 5316 18692
rect 7380 18683 7432 18692
rect 7380 18649 7389 18683
rect 7389 18649 7423 18683
rect 7423 18649 7432 18683
rect 10876 18751 10928 18760
rect 10876 18717 10885 18751
rect 10885 18717 10919 18751
rect 10919 18717 10928 18751
rect 10876 18708 10928 18717
rect 7380 18640 7432 18649
rect 8852 18640 8904 18692
rect 10968 18640 11020 18692
rect 14372 18708 14424 18760
rect 14832 18708 14884 18760
rect 16488 18708 16540 18760
rect 17868 18751 17920 18760
rect 17868 18717 17877 18751
rect 17877 18717 17911 18751
rect 17911 18717 17920 18751
rect 17868 18708 17920 18717
rect 19064 18708 19116 18760
rect 19524 18708 19576 18760
rect 20076 18708 20128 18760
rect 14740 18640 14792 18692
rect 20996 18640 21048 18692
rect 27620 18640 27672 18692
rect 4160 18572 4212 18624
rect 4804 18572 4856 18624
rect 5080 18615 5132 18624
rect 5080 18581 5089 18615
rect 5089 18581 5123 18615
rect 5123 18581 5132 18615
rect 5080 18572 5132 18581
rect 14556 18615 14608 18624
rect 14556 18581 14565 18615
rect 14565 18581 14599 18615
rect 14599 18581 14608 18615
rect 14556 18572 14608 18581
rect 16396 18615 16448 18624
rect 16396 18581 16405 18615
rect 16405 18581 16439 18615
rect 16439 18581 16448 18615
rect 16396 18572 16448 18581
rect 17776 18572 17828 18624
rect 18328 18615 18380 18624
rect 18328 18581 18337 18615
rect 18337 18581 18371 18615
rect 18371 18581 18380 18615
rect 18328 18572 18380 18581
rect 21824 18572 21876 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 6092 18368 6144 18420
rect 8116 18368 8168 18420
rect 9864 18368 9916 18420
rect 10508 18411 10560 18420
rect 10508 18377 10517 18411
rect 10517 18377 10551 18411
rect 10551 18377 10560 18411
rect 10508 18368 10560 18377
rect 10784 18368 10836 18420
rect 14556 18368 14608 18420
rect 7932 18300 7984 18352
rect 9680 18300 9732 18352
rect 4344 18275 4396 18284
rect 4344 18241 4353 18275
rect 4353 18241 4387 18275
rect 4387 18241 4396 18275
rect 4344 18232 4396 18241
rect 5264 18275 5316 18284
rect 5264 18241 5273 18275
rect 5273 18241 5307 18275
rect 5307 18241 5316 18275
rect 5264 18232 5316 18241
rect 5540 18275 5592 18284
rect 5540 18241 5549 18275
rect 5549 18241 5583 18275
rect 5583 18241 5592 18275
rect 5540 18232 5592 18241
rect 7380 18275 7432 18284
rect 7380 18241 7389 18275
rect 7389 18241 7423 18275
rect 7423 18241 7432 18275
rect 7380 18232 7432 18241
rect 7840 18275 7892 18284
rect 7840 18241 7849 18275
rect 7849 18241 7883 18275
rect 7883 18241 7892 18275
rect 7840 18232 7892 18241
rect 8944 18232 8996 18284
rect 10048 18232 10100 18284
rect 10692 18275 10744 18284
rect 10692 18241 10701 18275
rect 10701 18241 10735 18275
rect 10735 18241 10744 18275
rect 10692 18232 10744 18241
rect 12440 18232 12492 18284
rect 12808 18232 12860 18284
rect 4988 18164 5040 18216
rect 12716 18207 12768 18216
rect 12716 18173 12725 18207
rect 12725 18173 12759 18207
rect 12759 18173 12768 18207
rect 12716 18164 12768 18173
rect 12992 18207 13044 18216
rect 12992 18173 13001 18207
rect 13001 18173 13035 18207
rect 13035 18173 13044 18207
rect 12992 18164 13044 18173
rect 18328 18368 18380 18420
rect 18972 18411 19024 18420
rect 18972 18377 18981 18411
rect 18981 18377 19015 18411
rect 19015 18377 19024 18411
rect 18972 18368 19024 18377
rect 20168 18368 20220 18420
rect 20904 18411 20956 18420
rect 20904 18377 20913 18411
rect 20913 18377 20947 18411
rect 20947 18377 20956 18411
rect 20904 18368 20956 18377
rect 24768 18411 24820 18420
rect 24768 18377 24777 18411
rect 24777 18377 24811 18411
rect 24811 18377 24820 18411
rect 24768 18368 24820 18377
rect 17408 18300 17460 18352
rect 20536 18343 20588 18352
rect 20536 18309 20545 18343
rect 20545 18309 20579 18343
rect 20579 18309 20588 18343
rect 20536 18300 20588 18309
rect 16304 18232 16356 18284
rect 16488 18275 16540 18284
rect 16488 18241 16497 18275
rect 16497 18241 16531 18275
rect 16531 18241 16540 18275
rect 16488 18232 16540 18241
rect 17868 18232 17920 18284
rect 5356 18139 5408 18148
rect 5356 18105 5365 18139
rect 5365 18105 5399 18139
rect 5399 18105 5408 18139
rect 5356 18096 5408 18105
rect 8576 18096 8628 18148
rect 8760 18139 8812 18148
rect 8760 18105 8769 18139
rect 8769 18105 8803 18139
rect 8803 18105 8812 18139
rect 8760 18096 8812 18105
rect 10140 18096 10192 18148
rect 10784 18139 10836 18148
rect 10784 18105 10793 18139
rect 10793 18105 10827 18139
rect 10827 18105 10836 18139
rect 10784 18096 10836 18105
rect 4712 18071 4764 18080
rect 4712 18037 4721 18071
rect 4721 18037 4755 18071
rect 4755 18037 4764 18071
rect 4712 18028 4764 18037
rect 7012 18028 7064 18080
rect 11796 18071 11848 18080
rect 11796 18037 11805 18071
rect 11805 18037 11839 18071
rect 11839 18037 11848 18071
rect 11796 18028 11848 18037
rect 12532 18071 12584 18080
rect 12532 18037 12541 18071
rect 12541 18037 12575 18071
rect 12575 18037 12584 18071
rect 12532 18028 12584 18037
rect 13636 18071 13688 18080
rect 13636 18037 13645 18071
rect 13645 18037 13679 18071
rect 13679 18037 13688 18071
rect 24216 18164 24268 18216
rect 15476 18096 15528 18148
rect 19984 18139 20036 18148
rect 13636 18028 13688 18037
rect 14280 18028 14332 18080
rect 15292 18071 15344 18080
rect 15292 18037 15301 18071
rect 15301 18037 15335 18071
rect 15335 18037 15344 18071
rect 15292 18028 15344 18037
rect 17224 18071 17276 18080
rect 17224 18037 17233 18071
rect 17233 18037 17267 18071
rect 17267 18037 17276 18071
rect 17224 18028 17276 18037
rect 17776 18071 17828 18080
rect 17776 18037 17785 18071
rect 17785 18037 17819 18071
rect 17819 18037 17828 18071
rect 19984 18105 19993 18139
rect 19993 18105 20027 18139
rect 20027 18105 20036 18139
rect 19984 18096 20036 18105
rect 20168 18096 20220 18148
rect 19248 18071 19300 18080
rect 17776 18028 17828 18037
rect 19248 18037 19257 18071
rect 19257 18037 19291 18071
rect 19291 18037 19300 18071
rect 19248 18028 19300 18037
rect 21180 18028 21232 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 4804 17867 4856 17876
rect 4804 17833 4813 17867
rect 4813 17833 4847 17867
rect 4847 17833 4856 17867
rect 4804 17824 4856 17833
rect 6000 17824 6052 17876
rect 10692 17867 10744 17876
rect 10692 17833 10701 17867
rect 10701 17833 10735 17867
rect 10735 17833 10744 17867
rect 10692 17824 10744 17833
rect 5356 17756 5408 17808
rect 8208 17799 8260 17808
rect 8208 17765 8217 17799
rect 8217 17765 8251 17799
rect 8251 17765 8260 17799
rect 8208 17756 8260 17765
rect 9864 17799 9916 17808
rect 9864 17765 9873 17799
rect 9873 17765 9907 17799
rect 9907 17765 9916 17799
rect 9864 17756 9916 17765
rect 6092 17688 6144 17740
rect 12532 17824 12584 17876
rect 14832 17824 14884 17876
rect 15292 17824 15344 17876
rect 17868 17824 17920 17876
rect 11612 17756 11664 17808
rect 15476 17756 15528 17808
rect 17776 17756 17828 17808
rect 20536 17799 20588 17808
rect 20536 17765 20545 17799
rect 20545 17765 20579 17799
rect 20579 17765 20588 17799
rect 20536 17756 20588 17765
rect 20812 17756 20864 17808
rect 21456 17756 21508 17808
rect 13636 17731 13688 17740
rect 13636 17697 13645 17731
rect 13645 17697 13679 17731
rect 13679 17697 13688 17731
rect 13636 17688 13688 17697
rect 14188 17731 14240 17740
rect 14188 17697 14197 17731
rect 14197 17697 14231 17731
rect 14231 17697 14240 17731
rect 14188 17688 14240 17697
rect 4252 17620 4304 17672
rect 5540 17620 5592 17672
rect 7564 17620 7616 17672
rect 7840 17620 7892 17672
rect 9772 17663 9824 17672
rect 5080 17552 5132 17604
rect 9772 17629 9781 17663
rect 9781 17629 9815 17663
rect 9815 17629 9824 17663
rect 9772 17620 9824 17629
rect 10048 17663 10100 17672
rect 10048 17629 10057 17663
rect 10057 17629 10091 17663
rect 10091 17629 10100 17663
rect 10048 17620 10100 17629
rect 14832 17620 14884 17672
rect 15292 17663 15344 17672
rect 15292 17629 15301 17663
rect 15301 17629 15335 17663
rect 15335 17629 15344 17663
rect 15292 17620 15344 17629
rect 17684 17620 17736 17672
rect 21272 17663 21324 17672
rect 21272 17629 21281 17663
rect 21281 17629 21315 17663
rect 21315 17629 21324 17663
rect 21272 17620 21324 17629
rect 2044 17484 2096 17536
rect 11152 17552 11204 17604
rect 12348 17527 12400 17536
rect 12348 17493 12357 17527
rect 12357 17493 12391 17527
rect 12391 17493 12400 17527
rect 12348 17484 12400 17493
rect 12992 17484 13044 17536
rect 13360 17484 13412 17536
rect 19524 17527 19576 17536
rect 19524 17493 19533 17527
rect 19533 17493 19567 17527
rect 19567 17493 19576 17527
rect 19524 17484 19576 17493
rect 19984 17527 20036 17536
rect 19984 17493 19993 17527
rect 19993 17493 20027 17527
rect 20027 17493 20036 17527
rect 19984 17484 20036 17493
rect 20260 17484 20312 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 5540 17280 5592 17332
rect 6092 17280 6144 17332
rect 7840 17280 7892 17332
rect 10048 17280 10100 17332
rect 10784 17280 10836 17332
rect 11612 17280 11664 17332
rect 12348 17280 12400 17332
rect 13452 17280 13504 17332
rect 14648 17280 14700 17332
rect 15660 17323 15712 17332
rect 15660 17289 15669 17323
rect 15669 17289 15703 17323
rect 15703 17289 15712 17323
rect 15660 17280 15712 17289
rect 16304 17280 16356 17332
rect 21456 17323 21508 17332
rect 21456 17289 21465 17323
rect 21465 17289 21499 17323
rect 21499 17289 21508 17323
rect 21456 17280 21508 17289
rect 24216 17280 24268 17332
rect 8208 17212 8260 17264
rect 9772 17212 9824 17264
rect 11244 17212 11296 17264
rect 12992 17212 13044 17264
rect 15292 17212 15344 17264
rect 7104 17144 7156 17196
rect 7656 17144 7708 17196
rect 10692 17144 10744 17196
rect 10968 17144 11020 17196
rect 11152 17187 11204 17196
rect 11152 17153 11161 17187
rect 11161 17153 11195 17187
rect 11195 17153 11204 17187
rect 11152 17144 11204 17153
rect 14188 17144 14240 17196
rect 15568 17144 15620 17196
rect 20076 17144 20128 17196
rect 21272 17144 21324 17196
rect 4620 17076 4672 17128
rect 3240 16983 3292 16992
rect 3240 16949 3249 16983
rect 3249 16949 3283 16983
rect 3283 16949 3292 16983
rect 3240 16940 3292 16949
rect 8576 17076 8628 17128
rect 14740 17119 14792 17128
rect 14740 17085 14749 17119
rect 14749 17085 14783 17119
rect 14783 17085 14792 17119
rect 14740 17076 14792 17085
rect 16488 17119 16540 17128
rect 16488 17085 16497 17119
rect 16497 17085 16531 17119
rect 16531 17085 16540 17119
rect 16488 17076 16540 17085
rect 19340 17076 19392 17128
rect 22468 17119 22520 17128
rect 8024 17008 8076 17060
rect 8760 17008 8812 17060
rect 10968 17051 11020 17060
rect 10968 17017 10977 17051
rect 10977 17017 11011 17051
rect 11011 17017 11020 17051
rect 12532 17051 12584 17060
rect 10968 17008 11020 17017
rect 12532 17017 12541 17051
rect 12541 17017 12575 17051
rect 12575 17017 12584 17051
rect 12532 17008 12584 17017
rect 4252 16940 4304 16992
rect 4804 16940 4856 16992
rect 5080 16983 5132 16992
rect 5080 16949 5089 16983
rect 5089 16949 5123 16983
rect 5123 16949 5132 16983
rect 5080 16940 5132 16949
rect 6828 16940 6880 16992
rect 7380 16983 7432 16992
rect 7380 16949 7389 16983
rect 7389 16949 7423 16983
rect 7423 16949 7432 16983
rect 7380 16940 7432 16949
rect 12348 16940 12400 16992
rect 14648 17008 14700 17060
rect 15476 17008 15528 17060
rect 13268 16940 13320 16992
rect 13636 16983 13688 16992
rect 13636 16949 13645 16983
rect 13645 16949 13679 16983
rect 13679 16949 13688 16983
rect 13636 16940 13688 16949
rect 16948 16940 17000 16992
rect 17684 16940 17736 16992
rect 17776 16983 17828 16992
rect 17776 16949 17785 16983
rect 17785 16949 17819 16983
rect 17819 16949 17828 16983
rect 20536 17051 20588 17060
rect 20536 17017 20545 17051
rect 20545 17017 20579 17051
rect 20579 17017 20588 17051
rect 20536 17008 20588 17017
rect 22468 17085 22477 17119
rect 22477 17085 22511 17119
rect 22511 17085 22520 17119
rect 22468 17076 22520 17085
rect 24124 17119 24176 17128
rect 24124 17085 24133 17119
rect 24133 17085 24167 17119
rect 24167 17085 24176 17119
rect 24124 17076 24176 17085
rect 17776 16940 17828 16949
rect 23296 17008 23348 17060
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 5080 16736 5132 16788
rect 8024 16736 8076 16788
rect 8208 16779 8260 16788
rect 8208 16745 8217 16779
rect 8217 16745 8251 16779
rect 8251 16745 8260 16779
rect 8208 16736 8260 16745
rect 10692 16736 10744 16788
rect 12440 16779 12492 16788
rect 12440 16745 12449 16779
rect 12449 16745 12483 16779
rect 12483 16745 12492 16779
rect 12440 16736 12492 16745
rect 14740 16779 14792 16788
rect 14740 16745 14749 16779
rect 14749 16745 14783 16779
rect 14783 16745 14792 16779
rect 14740 16736 14792 16745
rect 15752 16736 15804 16788
rect 16304 16736 16356 16788
rect 19248 16736 19300 16788
rect 19340 16779 19392 16788
rect 19340 16745 19349 16779
rect 19349 16745 19383 16779
rect 19383 16745 19392 16779
rect 19340 16736 19392 16745
rect 21180 16736 21232 16788
rect 22468 16736 22520 16788
rect 5172 16711 5224 16720
rect 5172 16677 5181 16711
rect 5181 16677 5215 16711
rect 5215 16677 5224 16711
rect 5172 16668 5224 16677
rect 7656 16668 7708 16720
rect 11612 16668 11664 16720
rect 15476 16668 15528 16720
rect 17776 16668 17828 16720
rect 20812 16668 20864 16720
rect 2044 16600 2096 16652
rect 7288 16643 7340 16652
rect 7288 16609 7297 16643
rect 7297 16609 7331 16643
rect 7331 16609 7340 16643
rect 7288 16600 7340 16609
rect 9588 16643 9640 16652
rect 9588 16609 9597 16643
rect 9597 16609 9631 16643
rect 9631 16609 9640 16643
rect 9588 16600 9640 16609
rect 10968 16600 11020 16652
rect 12624 16600 12676 16652
rect 13360 16643 13412 16652
rect 13360 16609 13369 16643
rect 13369 16609 13403 16643
rect 13403 16609 13412 16643
rect 13360 16600 13412 16609
rect 15292 16643 15344 16652
rect 15292 16609 15301 16643
rect 15301 16609 15335 16643
rect 15335 16609 15344 16643
rect 15292 16600 15344 16609
rect 4436 16532 4488 16584
rect 5540 16575 5592 16584
rect 5540 16541 5549 16575
rect 5549 16541 5583 16575
rect 5583 16541 5592 16575
rect 5540 16532 5592 16541
rect 11244 16532 11296 16584
rect 17500 16532 17552 16584
rect 20076 16600 20128 16652
rect 21088 16643 21140 16652
rect 21088 16609 21097 16643
rect 21097 16609 21131 16643
rect 21131 16609 21140 16643
rect 21088 16600 21140 16609
rect 21364 16600 21416 16652
rect 21824 16600 21876 16652
rect 22652 16600 22704 16652
rect 22928 16643 22980 16652
rect 22928 16609 22937 16643
rect 22937 16609 22971 16643
rect 22971 16609 22980 16643
rect 22928 16600 22980 16609
rect 1676 16464 1728 16516
rect 9312 16464 9364 16516
rect 12716 16464 12768 16516
rect 15752 16464 15804 16516
rect 1400 16396 1452 16448
rect 4620 16396 4672 16448
rect 7472 16439 7524 16448
rect 7472 16405 7481 16439
rect 7481 16405 7515 16439
rect 7515 16405 7524 16439
rect 7472 16396 7524 16405
rect 10140 16396 10192 16448
rect 13912 16439 13964 16448
rect 13912 16405 13921 16439
rect 13921 16405 13955 16439
rect 13955 16405 13964 16439
rect 13912 16396 13964 16405
rect 16948 16439 17000 16448
rect 16948 16405 16957 16439
rect 16957 16405 16991 16439
rect 16991 16405 17000 16439
rect 16948 16396 17000 16405
rect 19616 16439 19668 16448
rect 19616 16405 19625 16439
rect 19625 16405 19659 16439
rect 19659 16405 19668 16439
rect 19616 16396 19668 16405
rect 20076 16396 20128 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 2044 16235 2096 16244
rect 2044 16201 2053 16235
rect 2053 16201 2087 16235
rect 2087 16201 2096 16235
rect 2044 16192 2096 16201
rect 4436 16235 4488 16244
rect 4436 16201 4445 16235
rect 4445 16201 4479 16235
rect 4479 16201 4488 16235
rect 4436 16192 4488 16201
rect 1400 16031 1452 16040
rect 1400 15997 1409 16031
rect 1409 15997 1443 16031
rect 1443 15997 1452 16031
rect 1400 15988 1452 15997
rect 5172 16192 5224 16244
rect 7104 16235 7156 16244
rect 7104 16201 7113 16235
rect 7113 16201 7147 16235
rect 7147 16201 7156 16235
rect 7104 16192 7156 16201
rect 7472 16235 7524 16244
rect 7472 16201 7481 16235
rect 7481 16201 7515 16235
rect 7515 16201 7524 16235
rect 7472 16192 7524 16201
rect 9588 16192 9640 16244
rect 11612 16192 11664 16244
rect 12900 16192 12952 16244
rect 15292 16192 15344 16244
rect 15476 16192 15528 16244
rect 15936 16235 15988 16244
rect 15936 16201 15945 16235
rect 15945 16201 15979 16235
rect 15979 16201 15988 16235
rect 15936 16192 15988 16201
rect 17500 16235 17552 16244
rect 17500 16201 17509 16235
rect 17509 16201 17543 16235
rect 17543 16201 17552 16235
rect 17500 16192 17552 16201
rect 18972 16235 19024 16244
rect 18972 16201 18981 16235
rect 18981 16201 19015 16235
rect 19015 16201 19024 16235
rect 18972 16192 19024 16201
rect 20168 16235 20220 16244
rect 20168 16201 20177 16235
rect 20177 16201 20211 16235
rect 20211 16201 20220 16235
rect 20168 16192 20220 16201
rect 21364 16235 21416 16244
rect 21364 16201 21373 16235
rect 21373 16201 21407 16235
rect 21407 16201 21416 16235
rect 21364 16192 21416 16201
rect 22652 16235 22704 16244
rect 22652 16201 22661 16235
rect 22661 16201 22695 16235
rect 22695 16201 22704 16235
rect 22652 16192 22704 16201
rect 22928 16192 22980 16244
rect 5540 16167 5592 16176
rect 5540 16133 5549 16167
rect 5549 16133 5583 16167
rect 5583 16133 5592 16167
rect 5540 16124 5592 16133
rect 4988 16099 5040 16108
rect 4988 16065 4997 16099
rect 4997 16065 5031 16099
rect 5031 16065 5040 16099
rect 4988 16056 5040 16065
rect 14188 16124 14240 16176
rect 9312 16099 9364 16108
rect 9312 16065 9321 16099
rect 9321 16065 9355 16099
rect 9355 16065 9364 16099
rect 9312 16056 9364 16065
rect 11060 16056 11112 16108
rect 13360 16056 13412 16108
rect 19524 16124 19576 16176
rect 19616 16056 19668 16108
rect 22192 16056 22244 16108
rect 12348 15988 12400 16040
rect 5264 15920 5316 15972
rect 204 15852 256 15904
rect 7472 15852 7524 15904
rect 8484 15920 8536 15972
rect 9404 15963 9456 15972
rect 9404 15929 9413 15963
rect 9413 15929 9447 15963
rect 9447 15929 9456 15963
rect 9404 15920 9456 15929
rect 12624 15988 12676 16040
rect 14648 15988 14700 16040
rect 16304 15988 16356 16040
rect 16948 16031 17000 16040
rect 16948 15997 16957 16031
rect 16957 15997 16991 16031
rect 16991 15997 17000 16031
rect 16948 15988 17000 15997
rect 18604 16031 18656 16040
rect 18604 15997 18613 16031
rect 18613 15997 18647 16031
rect 18647 15997 18656 16031
rect 18604 15988 18656 15997
rect 10692 15895 10744 15904
rect 10692 15861 10701 15895
rect 10701 15861 10735 15895
rect 10735 15861 10744 15895
rect 13452 15920 13504 15972
rect 13912 15920 13964 15972
rect 14740 15920 14792 15972
rect 18328 15920 18380 15972
rect 18972 15920 19024 15972
rect 21824 15963 21876 15972
rect 21824 15929 21833 15963
rect 21833 15929 21867 15963
rect 21867 15929 21876 15963
rect 21824 15920 21876 15929
rect 22836 15920 22888 15972
rect 10692 15852 10744 15861
rect 15476 15852 15528 15904
rect 15936 15852 15988 15904
rect 17776 15895 17828 15904
rect 17776 15861 17785 15895
rect 17785 15861 17819 15895
rect 17819 15861 17828 15895
rect 17776 15852 17828 15861
rect 21088 15852 21140 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 1400 15648 1452 15700
rect 5264 15691 5316 15700
rect 5264 15657 5273 15691
rect 5273 15657 5307 15691
rect 5307 15657 5316 15691
rect 5264 15648 5316 15657
rect 7288 15691 7340 15700
rect 7288 15657 7297 15691
rect 7297 15657 7331 15691
rect 7331 15657 7340 15691
rect 7288 15648 7340 15657
rect 7840 15648 7892 15700
rect 9220 15691 9272 15700
rect 4436 15623 4488 15632
rect 4436 15589 4445 15623
rect 4445 15589 4479 15623
rect 4479 15589 4488 15623
rect 4436 15580 4488 15589
rect 4988 15623 5040 15632
rect 4988 15589 4997 15623
rect 4997 15589 5031 15623
rect 5031 15589 5040 15623
rect 4988 15580 5040 15589
rect 6276 15580 6328 15632
rect 9220 15657 9229 15691
rect 9229 15657 9263 15691
rect 9263 15657 9272 15691
rect 9220 15648 9272 15657
rect 11244 15691 11296 15700
rect 11244 15657 11253 15691
rect 11253 15657 11287 15691
rect 11287 15657 11296 15691
rect 11244 15648 11296 15657
rect 17684 15691 17736 15700
rect 17684 15657 17693 15691
rect 17693 15657 17727 15691
rect 17727 15657 17736 15691
rect 17684 15648 17736 15657
rect 8484 15623 8536 15632
rect 8484 15589 8493 15623
rect 8493 15589 8527 15623
rect 8527 15589 8536 15623
rect 8484 15580 8536 15589
rect 10140 15623 10192 15632
rect 10140 15589 10149 15623
rect 10149 15589 10183 15623
rect 10183 15589 10192 15623
rect 10140 15580 10192 15589
rect 10600 15580 10652 15632
rect 11060 15580 11112 15632
rect 13176 15623 13228 15632
rect 13176 15589 13185 15623
rect 13185 15589 13219 15623
rect 13219 15589 13228 15623
rect 13176 15580 13228 15589
rect 15936 15580 15988 15632
rect 19524 15648 19576 15700
rect 21824 15648 21876 15700
rect 22284 15691 22336 15700
rect 22284 15657 22293 15691
rect 22293 15657 22327 15691
rect 22327 15657 22336 15691
rect 22284 15648 22336 15657
rect 2964 15555 3016 15564
rect 2964 15521 2973 15555
rect 2973 15521 3007 15555
rect 3007 15521 3016 15555
rect 2964 15512 3016 15521
rect 11888 15512 11940 15564
rect 14832 15512 14884 15564
rect 16304 15512 16356 15564
rect 21456 15580 21508 15632
rect 22560 15623 22612 15632
rect 22560 15589 22569 15623
rect 22569 15589 22603 15623
rect 22603 15589 22612 15623
rect 22560 15580 22612 15589
rect 22652 15623 22704 15632
rect 22652 15589 22661 15623
rect 22661 15589 22695 15623
rect 22695 15589 22704 15623
rect 22652 15580 22704 15589
rect 17684 15512 17736 15564
rect 18328 15512 18380 15564
rect 24676 15512 24728 15564
rect 3148 15351 3200 15360
rect 3148 15317 3157 15351
rect 3157 15317 3191 15351
rect 3191 15317 3200 15351
rect 3148 15308 3200 15317
rect 3424 15308 3476 15360
rect 4344 15308 4396 15360
rect 7472 15444 7524 15496
rect 10416 15487 10468 15496
rect 10416 15453 10425 15487
rect 10425 15453 10459 15487
rect 10459 15453 10468 15487
rect 10416 15444 10468 15453
rect 13084 15487 13136 15496
rect 13084 15453 13093 15487
rect 13093 15453 13127 15487
rect 13127 15453 13136 15487
rect 13084 15444 13136 15453
rect 13452 15444 13504 15496
rect 18788 15487 18840 15496
rect 18788 15453 18797 15487
rect 18797 15453 18831 15487
rect 18831 15453 18840 15487
rect 18788 15444 18840 15453
rect 20996 15487 21048 15496
rect 20996 15453 21005 15487
rect 21005 15453 21039 15487
rect 21039 15453 21048 15487
rect 20996 15444 21048 15453
rect 20536 15376 20588 15428
rect 22836 15487 22888 15496
rect 22836 15453 22845 15487
rect 22845 15453 22879 15487
rect 22879 15453 22888 15487
rect 22836 15444 22888 15453
rect 24768 15419 24820 15428
rect 24768 15385 24777 15419
rect 24777 15385 24811 15419
rect 24811 15385 24820 15419
rect 24768 15376 24820 15385
rect 7564 15351 7616 15360
rect 7564 15317 7573 15351
rect 7573 15317 7607 15351
rect 7607 15317 7616 15351
rect 7564 15308 7616 15317
rect 14004 15351 14056 15360
rect 14004 15317 14013 15351
rect 14013 15317 14047 15351
rect 14047 15317 14056 15351
rect 14004 15308 14056 15317
rect 15660 15351 15712 15360
rect 15660 15317 15669 15351
rect 15669 15317 15703 15351
rect 15703 15317 15712 15351
rect 15660 15308 15712 15317
rect 19064 15351 19116 15360
rect 19064 15317 19073 15351
rect 19073 15317 19107 15351
rect 19107 15317 19116 15351
rect 19064 15308 19116 15317
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 4436 15104 4488 15156
rect 4804 15104 4856 15156
rect 7840 15147 7892 15156
rect 7840 15113 7849 15147
rect 7849 15113 7883 15147
rect 7883 15113 7892 15147
rect 7840 15104 7892 15113
rect 10140 15104 10192 15156
rect 11888 15104 11940 15156
rect 13084 15104 13136 15156
rect 14832 15104 14884 15156
rect 15660 15104 15712 15156
rect 15936 15147 15988 15156
rect 15936 15113 15945 15147
rect 15945 15113 15979 15147
rect 15979 15113 15988 15147
rect 15936 15104 15988 15113
rect 16948 15104 17000 15156
rect 17684 15147 17736 15156
rect 17684 15113 17693 15147
rect 17693 15113 17727 15147
rect 17727 15113 17736 15147
rect 17684 15104 17736 15113
rect 18788 15104 18840 15156
rect 22560 15104 22612 15156
rect 5264 15079 5316 15088
rect 5264 15045 5273 15079
rect 5273 15045 5307 15079
rect 5307 15045 5316 15079
rect 5264 15036 5316 15045
rect 7472 15036 7524 15088
rect 14188 15079 14240 15088
rect 14188 15045 14197 15079
rect 14197 15045 14231 15079
rect 14231 15045 14240 15079
rect 14188 15036 14240 15045
rect 6920 15011 6972 15020
rect 6920 14977 6929 15011
rect 6929 14977 6963 15011
rect 6963 14977 6972 15011
rect 6920 14968 6972 14977
rect 7564 14968 7616 15020
rect 10416 14968 10468 15020
rect 13176 14968 13228 15020
rect 1308 14900 1360 14952
rect 3240 14900 3292 14952
rect 4068 14900 4120 14952
rect 4528 14832 4580 14884
rect 6644 14875 6696 14884
rect 6644 14841 6653 14875
rect 6653 14841 6687 14875
rect 6687 14841 6696 14875
rect 6644 14832 6696 14841
rect 8024 14832 8076 14884
rect 9496 14875 9548 14884
rect 9496 14841 9505 14875
rect 9505 14841 9539 14875
rect 9539 14841 9548 14875
rect 9496 14832 9548 14841
rect 1584 14807 1636 14816
rect 1584 14773 1593 14807
rect 1593 14773 1627 14807
rect 1627 14773 1636 14807
rect 1584 14764 1636 14773
rect 2964 14807 3016 14816
rect 2964 14773 2973 14807
rect 2973 14773 3007 14807
rect 3007 14773 3016 14807
rect 2964 14764 3016 14773
rect 3608 14764 3660 14816
rect 6184 14807 6236 14816
rect 6184 14773 6193 14807
rect 6193 14773 6227 14807
rect 6227 14773 6236 14807
rect 6184 14764 6236 14773
rect 9312 14807 9364 14816
rect 9312 14773 9321 14807
rect 9321 14773 9355 14807
rect 9355 14773 9364 14807
rect 9312 14764 9364 14773
rect 10048 14764 10100 14816
rect 10692 14764 10744 14816
rect 10784 14764 10836 14816
rect 13268 14832 13320 14884
rect 14004 14968 14056 15020
rect 15752 15036 15804 15088
rect 21456 15036 21508 15088
rect 16856 15011 16908 15020
rect 16856 14977 16865 15011
rect 16865 14977 16899 15011
rect 16899 14977 16908 15011
rect 22744 15036 22796 15088
rect 16856 14968 16908 14977
rect 15016 14900 15068 14952
rect 18512 14943 18564 14952
rect 18512 14909 18521 14943
rect 18521 14909 18555 14943
rect 18555 14909 18564 14943
rect 18512 14900 18564 14909
rect 19064 14943 19116 14952
rect 19064 14909 19073 14943
rect 19073 14909 19107 14943
rect 19107 14909 19116 14943
rect 19064 14900 19116 14909
rect 16304 14875 16356 14884
rect 16304 14841 16313 14875
rect 16313 14841 16347 14875
rect 16347 14841 16356 14875
rect 16304 14832 16356 14841
rect 12900 14764 12952 14816
rect 18236 14764 18288 14816
rect 20904 14764 20956 14816
rect 21456 14875 21508 14884
rect 21456 14841 21465 14875
rect 21465 14841 21499 14875
rect 21499 14841 21508 14875
rect 21456 14832 21508 14841
rect 22652 14968 22704 15020
rect 24676 15011 24728 15020
rect 24676 14977 24685 15011
rect 24685 14977 24719 15011
rect 24719 14977 24728 15011
rect 24676 14968 24728 14977
rect 23480 14875 23532 14884
rect 23480 14841 23489 14875
rect 23489 14841 23523 14875
rect 23523 14841 23532 14875
rect 24124 14943 24176 14952
rect 24124 14909 24133 14943
rect 24133 14909 24167 14943
rect 24167 14909 24176 14943
rect 24124 14900 24176 14909
rect 23480 14832 23532 14841
rect 23756 14807 23808 14816
rect 23756 14773 23765 14807
rect 23765 14773 23799 14807
rect 23799 14773 23808 14807
rect 23756 14764 23808 14773
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 940 14560 992 14612
rect 3424 14560 3476 14612
rect 3608 14560 3660 14612
rect 4436 14535 4488 14544
rect 4436 14501 4445 14535
rect 4445 14501 4479 14535
rect 4479 14501 4488 14535
rect 4988 14535 5040 14544
rect 4436 14492 4488 14501
rect 4988 14501 4997 14535
rect 4997 14501 5031 14535
rect 5031 14501 5040 14535
rect 4988 14492 5040 14501
rect 6828 14535 6880 14544
rect 6828 14501 6837 14535
rect 6837 14501 6871 14535
rect 6871 14501 6880 14535
rect 6828 14492 6880 14501
rect 9496 14603 9548 14612
rect 9496 14569 9505 14603
rect 9505 14569 9539 14603
rect 9539 14569 9548 14603
rect 9496 14560 9548 14569
rect 13084 14560 13136 14612
rect 13912 14560 13964 14612
rect 16304 14560 16356 14612
rect 18236 14560 18288 14612
rect 7012 14492 7064 14544
rect 7472 14535 7524 14544
rect 7472 14501 7481 14535
rect 7481 14501 7515 14535
rect 7515 14501 7524 14535
rect 7472 14492 7524 14501
rect 10508 14535 10560 14544
rect 10508 14501 10517 14535
rect 10517 14501 10551 14535
rect 10551 14501 10560 14535
rect 10508 14492 10560 14501
rect 16580 14535 16632 14544
rect 16580 14501 16589 14535
rect 16589 14501 16623 14535
rect 16623 14501 16632 14535
rect 16580 14492 16632 14501
rect 19524 14535 19576 14544
rect 19524 14501 19533 14535
rect 19533 14501 19567 14535
rect 19567 14501 19576 14535
rect 19524 14492 19576 14501
rect 20996 14560 21048 14612
rect 22560 14603 22612 14612
rect 22560 14569 22569 14603
rect 22569 14569 22603 14603
rect 22603 14569 22612 14603
rect 22560 14560 22612 14569
rect 21456 14492 21508 14544
rect 2136 14424 2188 14476
rect 3424 14424 3476 14476
rect 7932 14424 7984 14476
rect 8300 14467 8352 14476
rect 8300 14433 8344 14467
rect 8344 14433 8352 14467
rect 8300 14424 8352 14433
rect 15384 14424 15436 14476
rect 22468 14467 22520 14476
rect 10416 14399 10468 14408
rect 10416 14365 10425 14399
rect 10425 14365 10459 14399
rect 10459 14365 10468 14399
rect 10416 14356 10468 14365
rect 12808 14399 12860 14408
rect 12808 14365 12817 14399
rect 12817 14365 12851 14399
rect 12851 14365 12860 14399
rect 12808 14356 12860 14365
rect 14004 14356 14056 14408
rect 14188 14356 14240 14408
rect 16856 14356 16908 14408
rect 17500 14356 17552 14408
rect 10968 14331 11020 14340
rect 10968 14297 10977 14331
rect 10977 14297 11011 14331
rect 11011 14297 11020 14331
rect 10968 14288 11020 14297
rect 14464 14288 14516 14340
rect 17040 14331 17092 14340
rect 17040 14297 17049 14331
rect 17049 14297 17083 14331
rect 17083 14297 17092 14331
rect 17040 14288 17092 14297
rect 22468 14433 22477 14467
rect 22477 14433 22511 14467
rect 22511 14433 22520 14467
rect 22468 14424 22520 14433
rect 24124 14560 24176 14612
rect 20720 14356 20772 14408
rect 21180 14356 21232 14408
rect 21824 14356 21876 14408
rect 24676 14424 24728 14476
rect 19984 14288 20036 14340
rect 23664 14288 23716 14340
rect 2044 14263 2096 14272
rect 2044 14229 2053 14263
rect 2053 14229 2087 14263
rect 2087 14229 2096 14263
rect 2044 14220 2096 14229
rect 4068 14220 4120 14272
rect 6276 14263 6328 14272
rect 6276 14229 6285 14263
rect 6285 14229 6319 14263
rect 6319 14229 6328 14263
rect 6276 14220 6328 14229
rect 9772 14220 9824 14272
rect 12532 14263 12584 14272
rect 12532 14229 12541 14263
rect 12541 14229 12575 14263
rect 12575 14229 12584 14263
rect 12532 14220 12584 14229
rect 14372 14220 14424 14272
rect 15568 14220 15620 14272
rect 15844 14263 15896 14272
rect 15844 14229 15853 14263
rect 15853 14229 15887 14263
rect 15887 14229 15896 14263
rect 15844 14220 15896 14229
rect 19156 14263 19208 14272
rect 19156 14229 19165 14263
rect 19165 14229 19199 14263
rect 19199 14229 19208 14263
rect 19156 14220 19208 14229
rect 22284 14220 22336 14272
rect 23756 14220 23808 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 4344 14016 4396 14068
rect 4436 14016 4488 14068
rect 5080 14059 5132 14068
rect 5080 14025 5089 14059
rect 5089 14025 5123 14059
rect 5123 14025 5132 14059
rect 5080 14016 5132 14025
rect 6460 14016 6512 14068
rect 7012 14016 7064 14068
rect 8300 14059 8352 14068
rect 8300 14025 8309 14059
rect 8309 14025 8343 14059
rect 8343 14025 8352 14059
rect 8300 14016 8352 14025
rect 10416 14016 10468 14068
rect 11612 14016 11664 14068
rect 2136 13948 2188 14000
rect 2412 13948 2464 14000
rect 4988 13948 5040 14000
rect 6644 13991 6696 14000
rect 6644 13957 6653 13991
rect 6653 13957 6687 13991
rect 6687 13957 6696 13991
rect 6644 13948 6696 13957
rect 8024 13948 8076 14000
rect 112 13812 164 13864
rect 2872 13855 2924 13864
rect 2872 13821 2881 13855
rect 2881 13821 2915 13855
rect 2915 13821 2924 13855
rect 2872 13812 2924 13821
rect 6276 13880 6328 13932
rect 6736 13880 6788 13932
rect 3056 13719 3108 13728
rect 3056 13685 3065 13719
rect 3065 13685 3099 13719
rect 3099 13685 3108 13719
rect 3056 13676 3108 13685
rect 3424 13719 3476 13728
rect 3424 13685 3433 13719
rect 3433 13685 3467 13719
rect 3467 13685 3476 13719
rect 3424 13676 3476 13685
rect 4528 13744 4580 13796
rect 8944 13812 8996 13864
rect 6644 13744 6696 13796
rect 5448 13719 5500 13728
rect 5448 13685 5457 13719
rect 5457 13685 5491 13719
rect 5491 13685 5500 13719
rect 5448 13676 5500 13685
rect 6368 13676 6420 13728
rect 10508 13948 10560 14000
rect 9680 13744 9732 13796
rect 10140 13787 10192 13796
rect 10140 13753 10143 13787
rect 10143 13753 10177 13787
rect 10177 13753 10192 13787
rect 12900 14016 12952 14068
rect 13176 13948 13228 14000
rect 12440 13855 12492 13864
rect 12440 13821 12449 13855
rect 12449 13821 12483 13855
rect 12483 13821 12492 13855
rect 12440 13812 12492 13821
rect 10140 13744 10192 13753
rect 12256 13744 12308 13796
rect 15936 14016 15988 14068
rect 16580 14016 16632 14068
rect 19984 14059 20036 14068
rect 19984 14025 19993 14059
rect 19993 14025 20027 14059
rect 20027 14025 20036 14059
rect 19984 14016 20036 14025
rect 21456 14059 21508 14068
rect 21456 14025 21465 14059
rect 21465 14025 21499 14059
rect 21499 14025 21508 14059
rect 21456 14016 21508 14025
rect 23296 14016 23348 14068
rect 25412 14059 25464 14068
rect 25412 14025 25421 14059
rect 25421 14025 25455 14059
rect 25455 14025 25464 14059
rect 25412 14016 25464 14025
rect 19064 13948 19116 14000
rect 22468 13948 22520 14000
rect 14464 13880 14516 13932
rect 15844 13880 15896 13932
rect 19432 13880 19484 13932
rect 19156 13812 19208 13864
rect 22744 13855 22796 13864
rect 22744 13821 22753 13855
rect 22753 13821 22787 13855
rect 22787 13821 22796 13855
rect 22744 13812 22796 13821
rect 23296 13812 23348 13864
rect 24124 13855 24176 13864
rect 24124 13821 24133 13855
rect 24133 13821 24167 13855
rect 24167 13821 24176 13855
rect 24124 13812 24176 13821
rect 14372 13787 14424 13796
rect 14372 13753 14381 13787
rect 14381 13753 14415 13787
rect 14415 13753 14424 13787
rect 14372 13744 14424 13753
rect 13084 13676 13136 13728
rect 17500 13787 17552 13796
rect 15384 13719 15436 13728
rect 15384 13685 15393 13719
rect 15393 13685 15427 13719
rect 15427 13685 15436 13719
rect 15384 13676 15436 13685
rect 17500 13753 17509 13787
rect 17509 13753 17543 13787
rect 17543 13753 17552 13787
rect 17500 13744 17552 13753
rect 18236 13719 18288 13728
rect 18236 13685 18245 13719
rect 18245 13685 18279 13719
rect 18279 13685 18288 13719
rect 18236 13676 18288 13685
rect 18420 13744 18472 13796
rect 20536 13787 20588 13796
rect 20536 13753 20545 13787
rect 20545 13753 20579 13787
rect 20579 13753 20588 13787
rect 20536 13744 20588 13753
rect 21180 13787 21232 13796
rect 19432 13676 19484 13728
rect 19524 13676 19576 13728
rect 20168 13676 20220 13728
rect 21180 13753 21189 13787
rect 21189 13753 21223 13787
rect 21223 13753 21232 13787
rect 21180 13744 21232 13753
rect 22100 13787 22152 13796
rect 22100 13753 22109 13787
rect 22109 13753 22143 13787
rect 22143 13753 22152 13787
rect 22100 13744 22152 13753
rect 22284 13744 22336 13796
rect 24676 13787 24728 13796
rect 24676 13753 24685 13787
rect 24685 13753 24719 13787
rect 24719 13753 24728 13787
rect 24676 13744 24728 13753
rect 21824 13719 21876 13728
rect 21824 13685 21833 13719
rect 21833 13685 21867 13719
rect 21867 13685 21876 13719
rect 21824 13676 21876 13685
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 3056 13472 3108 13524
rect 4528 13472 4580 13524
rect 5080 13515 5132 13524
rect 5080 13481 5089 13515
rect 5089 13481 5123 13515
rect 5123 13481 5132 13515
rect 5080 13472 5132 13481
rect 6828 13472 6880 13524
rect 4804 13447 4856 13456
rect 4804 13413 4813 13447
rect 4813 13413 4847 13447
rect 4847 13413 4856 13447
rect 4804 13404 4856 13413
rect 2228 13336 2280 13388
rect 2412 13336 2464 13388
rect 10968 13472 11020 13524
rect 12808 13515 12860 13524
rect 12808 13481 12817 13515
rect 12817 13481 12851 13515
rect 12851 13481 12860 13515
rect 12808 13472 12860 13481
rect 6184 13447 6236 13456
rect 6184 13413 6193 13447
rect 6193 13413 6227 13447
rect 6227 13413 6236 13447
rect 6184 13404 6236 13413
rect 10140 13404 10192 13456
rect 10416 13404 10468 13456
rect 6460 13379 6512 13388
rect 6460 13345 6469 13379
rect 6469 13345 6503 13379
rect 6503 13345 6512 13379
rect 6460 13336 6512 13345
rect 8300 13379 8352 13388
rect 8300 13345 8309 13379
rect 8309 13345 8343 13379
rect 8343 13345 8352 13379
rect 8300 13336 8352 13345
rect 8852 13336 8904 13388
rect 11428 13379 11480 13388
rect 11428 13345 11437 13379
rect 11437 13345 11471 13379
rect 11471 13345 11480 13379
rect 11428 13336 11480 13345
rect 11888 13379 11940 13388
rect 11888 13345 11897 13379
rect 11897 13345 11931 13379
rect 11931 13345 11940 13379
rect 11888 13336 11940 13345
rect 12440 13447 12492 13456
rect 12440 13413 12449 13447
rect 12449 13413 12483 13447
rect 12483 13413 12492 13447
rect 12440 13404 12492 13413
rect 13084 13404 13136 13456
rect 14004 13472 14056 13524
rect 14280 13515 14332 13524
rect 14280 13481 14289 13515
rect 14289 13481 14323 13515
rect 14323 13481 14332 13515
rect 14280 13472 14332 13481
rect 16580 13472 16632 13524
rect 16856 13472 16908 13524
rect 20168 13472 20220 13524
rect 20536 13472 20588 13524
rect 20904 13515 20956 13524
rect 20904 13481 20913 13515
rect 20913 13481 20947 13515
rect 20947 13481 20956 13515
rect 20904 13472 20956 13481
rect 22192 13472 22244 13524
rect 23756 13472 23808 13524
rect 18328 13404 18380 13456
rect 19524 13404 19576 13456
rect 22284 13404 22336 13456
rect 15292 13379 15344 13388
rect 15292 13345 15301 13379
rect 15301 13345 15335 13379
rect 15335 13345 15344 13379
rect 15292 13336 15344 13345
rect 15844 13379 15896 13388
rect 15844 13345 15853 13379
rect 15853 13345 15887 13379
rect 15887 13345 15896 13379
rect 15844 13336 15896 13345
rect 17040 13336 17092 13388
rect 21180 13336 21232 13388
rect 10784 13268 10836 13320
rect 13084 13311 13136 13320
rect 13084 13277 13093 13311
rect 13093 13277 13127 13311
rect 13127 13277 13136 13311
rect 13084 13268 13136 13277
rect 16028 13268 16080 13320
rect 18236 13311 18288 13320
rect 18236 13277 18245 13311
rect 18245 13277 18279 13311
rect 18279 13277 18288 13311
rect 18236 13268 18288 13277
rect 18420 13268 18472 13320
rect 21088 13268 21140 13320
rect 21456 13268 21508 13320
rect 22008 13311 22060 13320
rect 22008 13277 22017 13311
rect 22017 13277 22051 13311
rect 22051 13277 22060 13311
rect 22008 13268 22060 13277
rect 8024 13200 8076 13252
rect 12348 13200 12400 13252
rect 14740 13200 14792 13252
rect 17132 13200 17184 13252
rect 20444 13200 20496 13252
rect 20720 13243 20772 13252
rect 20720 13209 20729 13243
rect 20729 13209 20763 13243
rect 20763 13209 20772 13243
rect 22836 13404 22888 13456
rect 23480 13379 23532 13388
rect 23480 13345 23489 13379
rect 23489 13345 23523 13379
rect 23523 13345 23532 13379
rect 23940 13379 23992 13388
rect 23480 13336 23532 13345
rect 23940 13345 23949 13379
rect 23949 13345 23983 13379
rect 23983 13345 23992 13379
rect 23940 13336 23992 13345
rect 25136 13336 25188 13388
rect 24032 13311 24084 13320
rect 24032 13277 24041 13311
rect 24041 13277 24075 13311
rect 24075 13277 24084 13311
rect 24032 13268 24084 13277
rect 20720 13200 20772 13209
rect 1860 13175 1912 13184
rect 1860 13141 1869 13175
rect 1869 13141 1903 13175
rect 1903 13141 1912 13175
rect 1860 13132 1912 13141
rect 2136 13132 2188 13184
rect 2504 13132 2556 13184
rect 2872 13132 2924 13184
rect 5356 13132 5408 13184
rect 7656 13132 7708 13184
rect 9312 13132 9364 13184
rect 14004 13175 14056 13184
rect 14004 13141 14013 13175
rect 14013 13141 14047 13175
rect 14047 13141 14056 13175
rect 14004 13132 14056 13141
rect 15752 13132 15804 13184
rect 16120 13132 16172 13184
rect 18788 13132 18840 13184
rect 19984 13175 20036 13184
rect 19984 13141 19993 13175
rect 19993 13141 20027 13175
rect 20027 13141 20036 13175
rect 19984 13132 20036 13141
rect 21548 13175 21600 13184
rect 21548 13141 21557 13175
rect 21557 13141 21591 13175
rect 21591 13141 21600 13175
rect 21548 13132 21600 13141
rect 24676 13132 24728 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 1952 12928 2004 12980
rect 2412 12971 2464 12980
rect 2412 12937 2421 12971
rect 2421 12937 2455 12971
rect 2455 12937 2464 12971
rect 8852 12971 8904 12980
rect 2412 12928 2464 12937
rect 8852 12937 8861 12971
rect 8861 12937 8895 12971
rect 8895 12937 8904 12971
rect 8852 12928 8904 12937
rect 9312 12971 9364 12980
rect 9312 12937 9321 12971
rect 9321 12937 9355 12971
rect 9355 12937 9364 12971
rect 9312 12928 9364 12937
rect 10140 12928 10192 12980
rect 10784 12971 10836 12980
rect 10784 12937 10793 12971
rect 10793 12937 10827 12971
rect 10827 12937 10836 12971
rect 10784 12928 10836 12937
rect 12256 12971 12308 12980
rect 12256 12937 12265 12971
rect 12265 12937 12299 12971
rect 12299 12937 12308 12971
rect 12256 12928 12308 12937
rect 2872 12860 2924 12912
rect 6828 12860 6880 12912
rect 10416 12903 10468 12912
rect 10416 12869 10425 12903
rect 10425 12869 10459 12903
rect 10459 12869 10468 12903
rect 10416 12860 10468 12869
rect 7932 12792 7984 12844
rect 8116 12835 8168 12844
rect 8116 12801 8125 12835
rect 8125 12801 8159 12835
rect 8159 12801 8168 12835
rect 8116 12792 8168 12801
rect 9496 12792 9548 12844
rect 14004 12971 14056 12980
rect 14004 12937 14013 12971
rect 14013 12937 14047 12971
rect 14047 12937 14056 12971
rect 14004 12928 14056 12937
rect 15292 12971 15344 12980
rect 15292 12937 15301 12971
rect 15301 12937 15335 12971
rect 15335 12937 15344 12971
rect 15292 12928 15344 12937
rect 17132 12928 17184 12980
rect 20076 12928 20128 12980
rect 22192 12928 22244 12980
rect 22284 12928 22336 12980
rect 23480 12928 23532 12980
rect 23940 12928 23992 12980
rect 25136 12971 25188 12980
rect 25136 12937 25145 12971
rect 25145 12937 25179 12971
rect 25179 12937 25188 12971
rect 25136 12928 25188 12937
rect 12624 12860 12676 12912
rect 14280 12835 14332 12844
rect 1584 12724 1636 12776
rect 2596 12767 2648 12776
rect 2596 12733 2605 12767
rect 2605 12733 2639 12767
rect 2639 12733 2648 12767
rect 2596 12724 2648 12733
rect 1768 12656 1820 12708
rect 2964 12656 3016 12708
rect 4528 12724 4580 12776
rect 5356 12767 5408 12776
rect 4344 12656 4396 12708
rect 5356 12733 5365 12767
rect 5365 12733 5399 12767
rect 5399 12733 5408 12767
rect 5356 12724 5408 12733
rect 7656 12767 7708 12776
rect 7656 12733 7665 12767
rect 7665 12733 7699 12767
rect 7699 12733 7708 12767
rect 7656 12724 7708 12733
rect 9312 12656 9364 12708
rect 12532 12724 12584 12776
rect 14280 12801 14289 12835
rect 14289 12801 14323 12835
rect 14323 12801 14332 12835
rect 14280 12792 14332 12801
rect 15752 12767 15804 12776
rect 15752 12733 15761 12767
rect 15761 12733 15795 12767
rect 15795 12733 15804 12767
rect 15752 12724 15804 12733
rect 16304 12767 16356 12776
rect 16304 12733 16313 12767
rect 16313 12733 16347 12767
rect 16347 12733 16356 12767
rect 16304 12724 16356 12733
rect 18328 12860 18380 12912
rect 20536 12903 20588 12912
rect 20536 12869 20545 12903
rect 20545 12869 20579 12903
rect 20579 12869 20588 12903
rect 20536 12860 20588 12869
rect 24768 12903 24820 12912
rect 24768 12869 24777 12903
rect 24777 12869 24811 12903
rect 24811 12869 24820 12903
rect 24768 12860 24820 12869
rect 18604 12835 18656 12844
rect 18604 12801 18613 12835
rect 18613 12801 18647 12835
rect 18647 12801 18656 12835
rect 18604 12792 18656 12801
rect 20076 12792 20128 12844
rect 18420 12724 18472 12776
rect 18788 12724 18840 12776
rect 24676 12724 24728 12776
rect 3884 12588 3936 12640
rect 4252 12631 4304 12640
rect 4252 12597 4261 12631
rect 4261 12597 4295 12631
rect 4295 12597 4304 12631
rect 4252 12588 4304 12597
rect 6000 12631 6052 12640
rect 6000 12597 6009 12631
rect 6009 12597 6043 12631
rect 6043 12597 6052 12631
rect 6000 12588 6052 12597
rect 7196 12631 7248 12640
rect 7196 12597 7205 12631
rect 7205 12597 7239 12631
rect 7239 12597 7248 12631
rect 7196 12588 7248 12597
rect 8300 12588 8352 12640
rect 9036 12588 9088 12640
rect 9680 12588 9732 12640
rect 12716 12656 12768 12708
rect 13176 12656 13228 12708
rect 13728 12656 13780 12708
rect 14924 12699 14976 12708
rect 11428 12588 11480 12640
rect 13544 12588 13596 12640
rect 14004 12588 14056 12640
rect 14924 12665 14933 12699
rect 14933 12665 14967 12699
rect 14967 12665 14976 12699
rect 14924 12656 14976 12665
rect 18236 12656 18288 12708
rect 19984 12699 20036 12708
rect 19984 12665 19993 12699
rect 19993 12665 20027 12699
rect 20027 12665 20036 12699
rect 19984 12656 20036 12665
rect 21548 12699 21600 12708
rect 15844 12631 15896 12640
rect 15844 12597 15853 12631
rect 15853 12597 15887 12631
rect 15887 12597 15896 12631
rect 15844 12588 15896 12597
rect 19524 12588 19576 12640
rect 21548 12665 21557 12699
rect 21557 12665 21591 12699
rect 21591 12665 21600 12699
rect 21548 12656 21600 12665
rect 21088 12588 21140 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 1768 12384 1820 12436
rect 2228 12384 2280 12436
rect 3148 12384 3200 12436
rect 3976 12384 4028 12436
rect 4620 12427 4672 12436
rect 4620 12393 4629 12427
rect 4629 12393 4663 12427
rect 4663 12393 4672 12427
rect 4620 12384 4672 12393
rect 6460 12427 6512 12436
rect 6460 12393 6469 12427
rect 6469 12393 6503 12427
rect 6503 12393 6512 12427
rect 6460 12384 6512 12393
rect 6828 12427 6880 12436
rect 6828 12393 6837 12427
rect 6837 12393 6871 12427
rect 6871 12393 6880 12427
rect 9496 12427 9548 12436
rect 6828 12384 6880 12393
rect 2596 12316 2648 12368
rect 1400 12291 1452 12300
rect 1400 12257 1409 12291
rect 1409 12257 1443 12291
rect 1443 12257 1452 12291
rect 1400 12248 1452 12257
rect 2412 12291 2464 12300
rect 2412 12257 2421 12291
rect 2421 12257 2455 12291
rect 2455 12257 2464 12291
rect 2412 12248 2464 12257
rect 3056 12248 3108 12300
rect 4344 12291 4396 12300
rect 4344 12257 4353 12291
rect 4353 12257 4387 12291
rect 4387 12257 4396 12291
rect 4344 12248 4396 12257
rect 4528 12248 4580 12300
rect 6000 12316 6052 12368
rect 6368 12316 6420 12368
rect 7288 12316 7340 12368
rect 2504 12223 2556 12232
rect 2504 12189 2513 12223
rect 2513 12189 2547 12223
rect 2547 12189 2556 12223
rect 2504 12180 2556 12189
rect 3148 12223 3200 12232
rect 3148 12189 3157 12223
rect 3157 12189 3191 12223
rect 3191 12189 3200 12223
rect 3148 12180 3200 12189
rect 6184 12248 6236 12300
rect 7380 12291 7432 12300
rect 7380 12257 7389 12291
rect 7389 12257 7423 12291
rect 7423 12257 7432 12291
rect 7380 12248 7432 12257
rect 9496 12393 9505 12427
rect 9505 12393 9539 12427
rect 9539 12393 9548 12427
rect 9496 12384 9548 12393
rect 9772 12427 9824 12436
rect 9772 12393 9781 12427
rect 9781 12393 9815 12427
rect 9815 12393 9824 12427
rect 9772 12384 9824 12393
rect 11888 12384 11940 12436
rect 14832 12384 14884 12436
rect 17040 12427 17092 12436
rect 17040 12393 17049 12427
rect 17049 12393 17083 12427
rect 17083 12393 17092 12427
rect 17040 12384 17092 12393
rect 18328 12427 18380 12436
rect 18328 12393 18337 12427
rect 18337 12393 18371 12427
rect 18371 12393 18380 12427
rect 18328 12384 18380 12393
rect 20352 12384 20404 12436
rect 8484 12316 8536 12368
rect 13084 12359 13136 12368
rect 13084 12325 13093 12359
rect 13093 12325 13127 12359
rect 13127 12325 13136 12359
rect 13084 12316 13136 12325
rect 13544 12359 13596 12368
rect 13544 12325 13553 12359
rect 13553 12325 13587 12359
rect 13587 12325 13596 12359
rect 13544 12316 13596 12325
rect 14924 12316 14976 12368
rect 19432 12359 19484 12368
rect 19432 12325 19441 12359
rect 19441 12325 19475 12359
rect 19475 12325 19484 12359
rect 19432 12316 19484 12325
rect 20076 12316 20128 12368
rect 21548 12384 21600 12436
rect 24676 12427 24728 12436
rect 24676 12393 24685 12427
rect 24685 12393 24719 12427
rect 24719 12393 24728 12427
rect 24676 12384 24728 12393
rect 21088 12359 21140 12368
rect 21088 12325 21097 12359
rect 21097 12325 21131 12359
rect 21131 12325 21140 12359
rect 21088 12316 21140 12325
rect 7656 12291 7708 12300
rect 7656 12257 7665 12291
rect 7665 12257 7699 12291
rect 7699 12257 7708 12291
rect 7656 12248 7708 12257
rect 3056 12112 3108 12164
rect 9036 12180 9088 12232
rect 10692 12248 10744 12300
rect 11336 12248 11388 12300
rect 11428 12248 11480 12300
rect 11888 12291 11940 12300
rect 11888 12257 11897 12291
rect 11897 12257 11931 12291
rect 11931 12257 11940 12291
rect 11888 12248 11940 12257
rect 15568 12291 15620 12300
rect 8576 12112 8628 12164
rect 12256 12112 12308 12164
rect 15568 12257 15577 12291
rect 15577 12257 15611 12291
rect 15611 12257 15620 12291
rect 15568 12248 15620 12257
rect 15660 12248 15712 12300
rect 16304 12248 16356 12300
rect 17224 12291 17276 12300
rect 13452 12223 13504 12232
rect 13452 12189 13461 12223
rect 13461 12189 13495 12223
rect 13495 12189 13504 12223
rect 13452 12180 13504 12189
rect 15752 12180 15804 12232
rect 16120 12223 16172 12232
rect 16120 12189 16129 12223
rect 16129 12189 16163 12223
rect 16163 12189 16172 12223
rect 16120 12180 16172 12189
rect 17224 12257 17233 12291
rect 17233 12257 17267 12291
rect 17267 12257 17276 12291
rect 17224 12248 17276 12257
rect 17684 12291 17736 12300
rect 17684 12257 17693 12291
rect 17693 12257 17727 12291
rect 17727 12257 17736 12291
rect 17684 12248 17736 12257
rect 22468 12291 22520 12300
rect 22468 12257 22477 12291
rect 22477 12257 22511 12291
rect 22511 12257 22520 12291
rect 22468 12248 22520 12257
rect 23664 12248 23716 12300
rect 18328 12180 18380 12232
rect 19156 12180 19208 12232
rect 21272 12223 21324 12232
rect 21272 12189 21281 12223
rect 21281 12189 21315 12223
rect 21315 12189 21324 12223
rect 21272 12180 21324 12189
rect 6092 12044 6144 12096
rect 9956 12044 10008 12096
rect 11244 12044 11296 12096
rect 14096 12044 14148 12096
rect 14648 12044 14700 12096
rect 21364 12044 21416 12096
rect 22008 12044 22060 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 2412 11840 2464 11892
rect 4160 11840 4212 11892
rect 6000 11840 6052 11892
rect 7380 11840 7432 11892
rect 8576 11883 8628 11892
rect 4344 11772 4396 11824
rect 1400 11704 1452 11756
rect 3792 11704 3844 11756
rect 7288 11747 7340 11756
rect 7288 11713 7297 11747
rect 7297 11713 7331 11747
rect 7331 11713 7340 11747
rect 7288 11704 7340 11713
rect 1860 11679 1912 11688
rect 1860 11645 1869 11679
rect 1869 11645 1903 11679
rect 1903 11645 1912 11679
rect 1860 11636 1912 11645
rect 3976 11679 4028 11688
rect 3976 11645 3985 11679
rect 3985 11645 4019 11679
rect 4019 11645 4028 11679
rect 3976 11636 4028 11645
rect 4528 11679 4580 11688
rect 4528 11645 4537 11679
rect 4537 11645 4571 11679
rect 4571 11645 4580 11679
rect 4528 11636 4580 11645
rect 5356 11679 5408 11688
rect 4436 11568 4488 11620
rect 5356 11645 5365 11679
rect 5365 11645 5399 11679
rect 5399 11645 5408 11679
rect 5356 11636 5408 11645
rect 7196 11679 7248 11688
rect 7196 11645 7205 11679
rect 7205 11645 7239 11679
rect 7239 11645 7248 11679
rect 7196 11636 7248 11645
rect 7380 11636 7432 11688
rect 8024 11704 8076 11756
rect 8576 11849 8585 11883
rect 8585 11849 8619 11883
rect 8619 11849 8628 11883
rect 8576 11840 8628 11849
rect 9036 11883 9088 11892
rect 9036 11849 9045 11883
rect 9045 11849 9079 11883
rect 9079 11849 9088 11883
rect 9036 11840 9088 11849
rect 9864 11840 9916 11892
rect 12256 11883 12308 11892
rect 12256 11849 12265 11883
rect 12265 11849 12299 11883
rect 12299 11849 12308 11883
rect 12256 11840 12308 11849
rect 13452 11840 13504 11892
rect 14464 11883 14516 11892
rect 14464 11849 14473 11883
rect 14473 11849 14507 11883
rect 14507 11849 14516 11883
rect 14464 11840 14516 11849
rect 14832 11840 14884 11892
rect 17316 11840 17368 11892
rect 18696 11840 18748 11892
rect 22468 11840 22520 11892
rect 23664 11840 23716 11892
rect 8576 11704 8628 11756
rect 7656 11636 7708 11688
rect 11244 11772 11296 11824
rect 11336 11815 11388 11824
rect 11336 11781 11345 11815
rect 11345 11781 11379 11815
rect 11379 11781 11388 11815
rect 11336 11772 11388 11781
rect 15568 11772 15620 11824
rect 17224 11815 17276 11824
rect 10048 11704 10100 11756
rect 13360 11704 13412 11756
rect 14188 11704 14240 11756
rect 17224 11781 17233 11815
rect 17233 11781 17267 11815
rect 17267 11781 17276 11815
rect 17224 11772 17276 11781
rect 18052 11772 18104 11824
rect 21180 11815 21232 11824
rect 16120 11704 16172 11756
rect 18328 11747 18380 11756
rect 18328 11713 18337 11747
rect 18337 11713 18371 11747
rect 18371 11713 18380 11747
rect 18328 11704 18380 11713
rect 21180 11781 21189 11815
rect 21189 11781 21223 11815
rect 21223 11781 21232 11815
rect 21180 11772 21232 11781
rect 20352 11704 20404 11756
rect 21272 11704 21324 11756
rect 21456 11704 21508 11756
rect 9956 11636 10008 11688
rect 10324 11679 10376 11688
rect 10324 11645 10333 11679
rect 10333 11645 10367 11679
rect 10367 11645 10376 11679
rect 10324 11636 10376 11645
rect 10784 11636 10836 11688
rect 4896 11568 4948 11620
rect 6184 11611 6236 11620
rect 2228 11543 2280 11552
rect 2228 11509 2237 11543
rect 2237 11509 2271 11543
rect 2271 11509 2280 11543
rect 2228 11500 2280 11509
rect 4068 11543 4120 11552
rect 4068 11509 4077 11543
rect 4077 11509 4111 11543
rect 4111 11509 4120 11543
rect 4068 11500 4120 11509
rect 6184 11577 6193 11611
rect 6193 11577 6227 11611
rect 6227 11577 6236 11611
rect 6184 11568 6236 11577
rect 8300 11568 8352 11620
rect 8484 11568 8536 11620
rect 13636 11611 13688 11620
rect 13636 11577 13645 11611
rect 13645 11577 13679 11611
rect 13679 11577 13688 11611
rect 13636 11568 13688 11577
rect 14280 11568 14332 11620
rect 10784 11500 10836 11552
rect 11888 11543 11940 11552
rect 11888 11509 11897 11543
rect 11897 11509 11931 11543
rect 11931 11509 11940 11543
rect 11888 11500 11940 11509
rect 12808 11500 12860 11552
rect 13268 11543 13320 11552
rect 13268 11509 13277 11543
rect 13277 11509 13311 11543
rect 13311 11509 13320 11543
rect 13268 11500 13320 11509
rect 13360 11500 13412 11552
rect 17684 11679 17736 11688
rect 17684 11645 17693 11679
rect 17693 11645 17727 11679
rect 17727 11645 17736 11679
rect 17684 11636 17736 11645
rect 18788 11636 18840 11688
rect 20076 11636 20128 11688
rect 15660 11568 15712 11620
rect 15936 11543 15988 11552
rect 15936 11509 15945 11543
rect 15945 11509 15979 11543
rect 15979 11509 15988 11543
rect 15936 11500 15988 11509
rect 16488 11500 16540 11552
rect 18696 11543 18748 11552
rect 18696 11509 18705 11543
rect 18705 11509 18739 11543
rect 18739 11509 18748 11543
rect 18696 11500 18748 11509
rect 19432 11500 19484 11552
rect 21088 11568 21140 11620
rect 21824 11543 21876 11552
rect 21824 11509 21833 11543
rect 21833 11509 21867 11543
rect 21867 11509 21876 11543
rect 21824 11500 21876 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 1860 11339 1912 11348
rect 1860 11305 1869 11339
rect 1869 11305 1903 11339
rect 1903 11305 1912 11339
rect 3056 11339 3108 11348
rect 1860 11296 1912 11305
rect 1952 11228 2004 11280
rect 3056 11305 3065 11339
rect 3065 11305 3099 11339
rect 3099 11305 3108 11339
rect 3056 11296 3108 11305
rect 3976 11296 4028 11348
rect 5448 11339 5500 11348
rect 5448 11305 5457 11339
rect 5457 11305 5491 11339
rect 5491 11305 5500 11339
rect 5448 11296 5500 11305
rect 6828 11296 6880 11348
rect 2780 11228 2832 11280
rect 10140 11296 10192 11348
rect 13544 11339 13596 11348
rect 13544 11305 13553 11339
rect 13553 11305 13587 11339
rect 13587 11305 13596 11339
rect 13544 11296 13596 11305
rect 14188 11339 14240 11348
rect 14188 11305 14197 11339
rect 14197 11305 14231 11339
rect 14231 11305 14240 11339
rect 14188 11296 14240 11305
rect 15568 11339 15620 11348
rect 15568 11305 15577 11339
rect 15577 11305 15611 11339
rect 15611 11305 15620 11339
rect 15568 11296 15620 11305
rect 16120 11339 16172 11348
rect 16120 11305 16129 11339
rect 16129 11305 16163 11339
rect 16163 11305 16172 11339
rect 16120 11296 16172 11305
rect 19984 11296 20036 11348
rect 20352 11339 20404 11348
rect 20352 11305 20361 11339
rect 20361 11305 20395 11339
rect 20395 11305 20404 11339
rect 20352 11296 20404 11305
rect 4528 11203 4580 11212
rect 4528 11169 4537 11203
rect 4537 11169 4571 11203
rect 4571 11169 4580 11203
rect 4528 11160 4580 11169
rect 4896 11203 4948 11212
rect 4896 11169 4905 11203
rect 4905 11169 4939 11203
rect 4939 11169 4948 11203
rect 4896 11160 4948 11169
rect 6184 11160 6236 11212
rect 7380 11203 7432 11212
rect 7380 11169 7389 11203
rect 7389 11169 7423 11203
rect 7423 11169 7432 11203
rect 7380 11160 7432 11169
rect 12716 11228 12768 11280
rect 15476 11228 15528 11280
rect 16304 11271 16356 11280
rect 16304 11237 16313 11271
rect 16313 11237 16347 11271
rect 16347 11237 16356 11271
rect 16304 11228 16356 11237
rect 16488 11228 16540 11280
rect 19156 11271 19208 11280
rect 19156 11237 19165 11271
rect 19165 11237 19199 11271
rect 19199 11237 19208 11271
rect 19156 11228 19208 11237
rect 19800 11228 19852 11280
rect 20076 11228 20128 11280
rect 21088 11271 21140 11280
rect 21088 11237 21097 11271
rect 21097 11237 21131 11271
rect 21131 11237 21140 11271
rect 21088 11228 21140 11237
rect 7656 11160 7708 11212
rect 1584 11092 1636 11144
rect 2320 11092 2372 11144
rect 3424 11092 3476 11144
rect 8300 11160 8352 11212
rect 9588 11160 9640 11212
rect 11336 11203 11388 11212
rect 11336 11169 11345 11203
rect 11345 11169 11379 11203
rect 11379 11169 11388 11203
rect 11336 11160 11388 11169
rect 13268 11160 13320 11212
rect 13636 11160 13688 11212
rect 14004 11203 14056 11212
rect 14004 11169 14013 11203
rect 14013 11169 14047 11203
rect 14047 11169 14056 11203
rect 14004 11160 14056 11169
rect 17960 11160 18012 11212
rect 18696 11203 18748 11212
rect 18696 11169 18705 11203
rect 18705 11169 18739 11203
rect 18739 11169 18748 11203
rect 18696 11160 18748 11169
rect 22744 11160 22796 11212
rect 11796 11092 11848 11144
rect 19432 11092 19484 11144
rect 21732 11092 21784 11144
rect 8208 10956 8260 11008
rect 13728 11024 13780 11076
rect 16672 11024 16724 11076
rect 12624 10956 12676 11008
rect 13452 10956 13504 11008
rect 18144 10999 18196 11008
rect 18144 10965 18153 10999
rect 18153 10965 18187 10999
rect 18187 10965 18196 10999
rect 18144 10956 18196 10965
rect 20996 10956 21048 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 20 10752 72 10804
rect 2044 10684 2096 10736
rect 3240 10752 3292 10804
rect 4988 10795 5040 10804
rect 4988 10761 4997 10795
rect 4997 10761 5031 10795
rect 5031 10761 5040 10795
rect 4988 10752 5040 10761
rect 7380 10752 7432 10804
rect 11336 10795 11388 10804
rect 11336 10761 11345 10795
rect 11345 10761 11379 10795
rect 11379 10761 11388 10795
rect 11336 10752 11388 10761
rect 11796 10795 11848 10804
rect 11796 10761 11805 10795
rect 11805 10761 11839 10795
rect 11839 10761 11848 10795
rect 11796 10752 11848 10761
rect 12716 10795 12768 10804
rect 12716 10761 12725 10795
rect 12725 10761 12759 10795
rect 12759 10761 12768 10795
rect 12716 10752 12768 10761
rect 14004 10795 14056 10804
rect 2136 10659 2188 10668
rect 2136 10625 2145 10659
rect 2145 10625 2179 10659
rect 2179 10625 2188 10659
rect 2136 10616 2188 10625
rect 5356 10684 5408 10736
rect 3884 10616 3936 10668
rect 5172 10591 5224 10600
rect 5172 10557 5181 10591
rect 5181 10557 5215 10591
rect 5215 10557 5224 10591
rect 5172 10548 5224 10557
rect 8484 10616 8536 10668
rect 7380 10591 7432 10600
rect 7380 10557 7389 10591
rect 7389 10557 7423 10591
rect 7423 10557 7432 10591
rect 7380 10548 7432 10557
rect 7656 10591 7708 10600
rect 7656 10557 7665 10591
rect 7665 10557 7699 10591
rect 7699 10557 7708 10591
rect 7656 10548 7708 10557
rect 8208 10591 8260 10600
rect 8208 10557 8217 10591
rect 8217 10557 8251 10591
rect 8251 10557 8260 10591
rect 8208 10548 8260 10557
rect 9588 10684 9640 10736
rect 13084 10684 13136 10736
rect 12900 10616 12952 10668
rect 12992 10616 13044 10668
rect 14004 10761 14013 10795
rect 14013 10761 14047 10795
rect 14047 10761 14056 10795
rect 14004 10752 14056 10761
rect 16028 10752 16080 10804
rect 16304 10752 16356 10804
rect 19340 10752 19392 10804
rect 19800 10795 19852 10804
rect 19800 10761 19809 10795
rect 19809 10761 19843 10795
rect 19843 10761 19852 10795
rect 19800 10752 19852 10761
rect 21088 10752 21140 10804
rect 21732 10795 21784 10804
rect 21732 10761 21741 10795
rect 21741 10761 21775 10795
rect 21775 10761 21784 10795
rect 21732 10752 21784 10761
rect 15844 10616 15896 10668
rect 18604 10659 18656 10668
rect 18604 10625 18613 10659
rect 18613 10625 18647 10659
rect 18647 10625 18656 10659
rect 18604 10616 18656 10625
rect 20444 10659 20496 10668
rect 20444 10625 20453 10659
rect 20453 10625 20487 10659
rect 20487 10625 20496 10659
rect 20444 10616 20496 10625
rect 21272 10616 21324 10668
rect 8760 10548 8812 10600
rect 9312 10548 9364 10600
rect 10140 10548 10192 10600
rect 14556 10591 14608 10600
rect 10692 10523 10744 10532
rect 1952 10455 2004 10464
rect 1952 10421 1961 10455
rect 1961 10421 1995 10455
rect 1995 10421 2004 10455
rect 10692 10489 10701 10523
rect 10701 10489 10735 10523
rect 10735 10489 10744 10523
rect 10692 10480 10744 10489
rect 4068 10455 4120 10464
rect 1952 10412 2004 10421
rect 4068 10421 4077 10455
rect 4077 10421 4111 10455
rect 4111 10421 4120 10455
rect 4068 10412 4120 10421
rect 5172 10412 5224 10464
rect 6552 10412 6604 10464
rect 9312 10412 9364 10464
rect 14556 10557 14565 10591
rect 14565 10557 14599 10591
rect 14599 10557 14608 10591
rect 14556 10548 14608 10557
rect 12716 10480 12768 10532
rect 14004 10480 14056 10532
rect 15936 10480 15988 10532
rect 17960 10480 18012 10532
rect 11336 10412 11388 10464
rect 13636 10412 13688 10464
rect 16856 10455 16908 10464
rect 16856 10421 16865 10455
rect 16865 10421 16899 10455
rect 16899 10421 16908 10455
rect 16856 10412 16908 10421
rect 17408 10412 17460 10464
rect 18144 10412 18196 10464
rect 21640 10548 21692 10600
rect 27620 10616 27672 10668
rect 20904 10480 20956 10532
rect 22744 10455 22796 10464
rect 22744 10421 22753 10455
rect 22753 10421 22787 10455
rect 22787 10421 22796 10455
rect 22744 10412 22796 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 2780 10251 2832 10260
rect 2780 10217 2789 10251
rect 2789 10217 2823 10251
rect 2823 10217 2832 10251
rect 2780 10208 2832 10217
rect 2044 10140 2096 10192
rect 1860 10115 1912 10124
rect 1860 10081 1869 10115
rect 1869 10081 1903 10115
rect 1903 10081 1912 10115
rect 4528 10208 4580 10260
rect 6920 10208 6972 10260
rect 8760 10251 8812 10260
rect 8760 10217 8769 10251
rect 8769 10217 8803 10251
rect 8803 10217 8812 10251
rect 8760 10208 8812 10217
rect 12624 10251 12676 10260
rect 12624 10217 12633 10251
rect 12633 10217 12667 10251
rect 12667 10217 12676 10251
rect 12624 10208 12676 10217
rect 12900 10251 12952 10260
rect 12900 10217 12909 10251
rect 12909 10217 12943 10251
rect 12943 10217 12952 10251
rect 12900 10208 12952 10217
rect 15752 10208 15804 10260
rect 16488 10208 16540 10260
rect 19340 10251 19392 10260
rect 19340 10217 19349 10251
rect 19349 10217 19383 10251
rect 19383 10217 19392 10251
rect 19340 10208 19392 10217
rect 20444 10251 20496 10260
rect 20444 10217 20453 10251
rect 20453 10217 20487 10251
rect 20487 10217 20496 10251
rect 20444 10208 20496 10217
rect 7196 10140 7248 10192
rect 9956 10183 10008 10192
rect 1860 10072 1912 10081
rect 3240 10072 3292 10124
rect 3976 10072 4028 10124
rect 4344 10072 4396 10124
rect 4620 10115 4672 10124
rect 4620 10081 4629 10115
rect 4629 10081 4663 10115
rect 4663 10081 4672 10115
rect 4620 10072 4672 10081
rect 4160 10004 4212 10056
rect 5172 10072 5224 10124
rect 5356 10115 5408 10124
rect 5356 10081 5365 10115
rect 5365 10081 5399 10115
rect 5399 10081 5408 10115
rect 5356 10072 5408 10081
rect 9956 10149 9965 10183
rect 9965 10149 9999 10183
rect 9999 10149 10008 10183
rect 9956 10140 10008 10149
rect 11336 10140 11388 10192
rect 7196 10004 7248 10056
rect 4436 9936 4488 9988
rect 1768 9911 1820 9920
rect 1768 9877 1777 9911
rect 1777 9877 1811 9911
rect 1811 9877 1820 9911
rect 1768 9868 1820 9877
rect 7656 10072 7708 10124
rect 7932 10115 7984 10124
rect 7932 10081 7941 10115
rect 7941 10081 7975 10115
rect 7975 10081 7984 10115
rect 7932 10072 7984 10081
rect 10508 10115 10560 10124
rect 10508 10081 10517 10115
rect 10517 10081 10551 10115
rect 10551 10081 10560 10115
rect 10508 10072 10560 10081
rect 11704 10072 11756 10124
rect 13360 10140 13412 10192
rect 13728 10183 13780 10192
rect 13268 10072 13320 10124
rect 13728 10149 13737 10183
rect 13737 10149 13771 10183
rect 13771 10149 13780 10183
rect 13728 10140 13780 10149
rect 13820 10140 13872 10192
rect 14280 10183 14332 10192
rect 14280 10149 14289 10183
rect 14289 10149 14323 10183
rect 14323 10149 14332 10183
rect 14280 10140 14332 10149
rect 16672 10183 16724 10192
rect 16672 10149 16681 10183
rect 16681 10149 16715 10183
rect 16715 10149 16724 10183
rect 16672 10140 16724 10149
rect 16856 10140 16908 10192
rect 17960 10140 18012 10192
rect 20076 10140 20128 10192
rect 21456 10140 21508 10192
rect 14740 10072 14792 10124
rect 18604 10072 18656 10124
rect 20812 10072 20864 10124
rect 22468 10115 22520 10124
rect 22468 10081 22477 10115
rect 22477 10081 22511 10115
rect 22511 10081 22520 10115
rect 22468 10072 22520 10081
rect 24676 10072 24728 10124
rect 13360 10004 13412 10056
rect 18420 10047 18472 10056
rect 18420 10013 18429 10047
rect 18429 10013 18463 10047
rect 18463 10013 18472 10047
rect 18420 10004 18472 10013
rect 20996 10047 21048 10056
rect 20996 10013 21005 10047
rect 21005 10013 21039 10047
rect 21039 10013 21048 10047
rect 20996 10004 21048 10013
rect 21272 10047 21324 10056
rect 21272 10013 21281 10047
rect 21281 10013 21315 10047
rect 21315 10013 21324 10047
rect 21272 10004 21324 10013
rect 11612 9979 11664 9988
rect 11612 9945 11621 9979
rect 11621 9945 11655 9979
rect 11655 9945 11664 9979
rect 11612 9936 11664 9945
rect 13544 9936 13596 9988
rect 14096 9936 14148 9988
rect 19432 9936 19484 9988
rect 7380 9868 7432 9920
rect 8208 9868 8260 9920
rect 9220 9868 9272 9920
rect 10784 9868 10836 9920
rect 11336 9911 11388 9920
rect 11336 9877 11345 9911
rect 11345 9877 11379 9911
rect 11379 9877 11388 9911
rect 11336 9868 11388 9877
rect 15844 9911 15896 9920
rect 15844 9877 15853 9911
rect 15853 9877 15887 9911
rect 15887 9877 15896 9911
rect 15844 9868 15896 9877
rect 16488 9868 16540 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 2964 9596 3016 9648
rect 4160 9596 4212 9648
rect 2320 9571 2372 9580
rect 2320 9537 2329 9571
rect 2329 9537 2363 9571
rect 2363 9537 2372 9571
rect 2320 9528 2372 9537
rect 3884 9528 3936 9580
rect 4528 9528 4580 9580
rect 7932 9596 7984 9648
rect 3792 9460 3844 9512
rect 4620 9503 4672 9512
rect 2228 9392 2280 9444
rect 2044 9324 2096 9376
rect 4160 9392 4212 9444
rect 4620 9469 4629 9503
rect 4629 9469 4663 9503
rect 4663 9469 4672 9503
rect 4620 9460 4672 9469
rect 5356 9503 5408 9512
rect 5356 9469 5365 9503
rect 5365 9469 5399 9503
rect 5399 9469 5408 9503
rect 5356 9460 5408 9469
rect 7196 9460 7248 9512
rect 7380 9503 7432 9512
rect 7380 9469 7389 9503
rect 7389 9469 7423 9503
rect 7423 9469 7432 9503
rect 7380 9460 7432 9469
rect 7656 9503 7708 9512
rect 7656 9469 7665 9503
rect 7665 9469 7699 9503
rect 7699 9469 7708 9503
rect 7656 9460 7708 9469
rect 9956 9664 10008 9716
rect 13268 9664 13320 9716
rect 16856 9707 16908 9716
rect 16856 9673 16865 9707
rect 16865 9673 16899 9707
rect 16899 9673 16908 9707
rect 16856 9664 16908 9673
rect 18052 9664 18104 9716
rect 18420 9664 18472 9716
rect 10048 9596 10100 9648
rect 11612 9596 11664 9648
rect 13636 9596 13688 9648
rect 13820 9596 13872 9648
rect 14740 9596 14792 9648
rect 16672 9596 16724 9648
rect 17408 9596 17460 9648
rect 20168 9596 20220 9648
rect 20996 9664 21048 9716
rect 21456 9664 21508 9716
rect 24676 9707 24728 9716
rect 24676 9673 24685 9707
rect 24685 9673 24719 9707
rect 24719 9673 24728 9707
rect 24676 9664 24728 9673
rect 22468 9639 22520 9648
rect 12992 9528 13044 9580
rect 13728 9528 13780 9580
rect 16120 9571 16172 9580
rect 16120 9537 16129 9571
rect 16129 9537 16163 9571
rect 16163 9537 16172 9571
rect 16120 9528 16172 9537
rect 17960 9528 18012 9580
rect 10508 9503 10560 9512
rect 4344 9392 4396 9444
rect 10508 9469 10517 9503
rect 10517 9469 10551 9503
rect 10551 9469 10560 9503
rect 10508 9460 10560 9469
rect 10784 9503 10836 9512
rect 10784 9469 10793 9503
rect 10793 9469 10827 9503
rect 10827 9469 10836 9503
rect 10784 9460 10836 9469
rect 12624 9503 12676 9512
rect 12624 9469 12633 9503
rect 12633 9469 12667 9503
rect 12667 9469 12676 9503
rect 12624 9460 12676 9469
rect 12808 9460 12860 9512
rect 3976 9324 4028 9376
rect 5264 9324 5316 9376
rect 6736 9324 6788 9376
rect 7104 9324 7156 9376
rect 9128 9392 9180 9444
rect 10140 9392 10192 9444
rect 9220 9324 9272 9376
rect 9312 9324 9364 9376
rect 10048 9367 10100 9376
rect 10048 9333 10057 9367
rect 10057 9333 10091 9367
rect 10091 9333 10100 9367
rect 10048 9324 10100 9333
rect 11244 9324 11296 9376
rect 12532 9367 12584 9376
rect 12532 9333 12541 9367
rect 12541 9333 12575 9367
rect 12575 9333 12584 9367
rect 12532 9324 12584 9333
rect 13820 9324 13872 9376
rect 15844 9435 15896 9444
rect 15844 9401 15853 9435
rect 15853 9401 15887 9435
rect 15887 9401 15896 9435
rect 15844 9392 15896 9401
rect 18788 9528 18840 9580
rect 22468 9605 22477 9639
rect 22477 9605 22511 9639
rect 22511 9605 22520 9639
rect 22468 9596 22520 9605
rect 20904 9571 20956 9580
rect 20904 9537 20913 9571
rect 20913 9537 20947 9571
rect 20947 9537 20956 9571
rect 20904 9528 20956 9537
rect 15568 9367 15620 9376
rect 15568 9333 15577 9367
rect 15577 9333 15611 9367
rect 15611 9333 15620 9367
rect 15568 9324 15620 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 1860 9120 1912 9172
rect 2044 9120 2096 9172
rect 3792 9163 3844 9172
rect 3792 9129 3801 9163
rect 3801 9129 3835 9163
rect 3835 9129 3844 9163
rect 3792 9120 3844 9129
rect 7288 9120 7340 9172
rect 8392 9120 8444 9172
rect 10140 9120 10192 9172
rect 11704 9120 11756 9172
rect 12808 9163 12860 9172
rect 12808 9129 12817 9163
rect 12817 9129 12851 9163
rect 12851 9129 12860 9163
rect 12808 9120 12860 9129
rect 17960 9120 18012 9172
rect 20168 9163 20220 9172
rect 20168 9129 20177 9163
rect 20177 9129 20211 9163
rect 20211 9129 20220 9163
rect 20168 9120 20220 9129
rect 20996 9120 21048 9172
rect 27620 9120 27672 9172
rect 2872 9052 2924 9104
rect 3424 9095 3476 9104
rect 3424 9061 3433 9095
rect 3433 9061 3467 9095
rect 3467 9061 3476 9095
rect 3424 9052 3476 9061
rect 4252 9095 4304 9104
rect 4252 9061 4261 9095
rect 4261 9061 4295 9095
rect 4295 9061 4304 9095
rect 4252 9052 4304 9061
rect 5356 9052 5408 9104
rect 11336 9052 11388 9104
rect 2044 8984 2096 9036
rect 3976 8984 4028 9036
rect 6000 8984 6052 9036
rect 7196 9027 7248 9036
rect 7196 8993 7205 9027
rect 7205 8993 7239 9027
rect 7239 8993 7248 9027
rect 7196 8984 7248 8993
rect 7380 9027 7432 9036
rect 7380 8993 7389 9027
rect 7389 8993 7423 9027
rect 7423 8993 7432 9027
rect 7380 8984 7432 8993
rect 8300 9027 8352 9036
rect 4160 8959 4212 8968
rect 4160 8925 4169 8959
rect 4169 8925 4203 8959
rect 4203 8925 4212 8959
rect 4436 8959 4488 8968
rect 4160 8916 4212 8925
rect 4436 8925 4445 8959
rect 4445 8925 4479 8959
rect 4479 8925 4488 8959
rect 4436 8916 4488 8925
rect 6092 8916 6144 8968
rect 7012 8916 7064 8968
rect 8300 8993 8309 9027
rect 8309 8993 8343 9027
rect 8343 8993 8352 9027
rect 8300 8984 8352 8993
rect 10784 9027 10836 9036
rect 10784 8993 10793 9027
rect 10793 8993 10827 9027
rect 10827 8993 10836 9027
rect 15568 9052 15620 9104
rect 18052 9095 18104 9104
rect 18052 9061 18061 9095
rect 18061 9061 18095 9095
rect 18095 9061 18104 9095
rect 18052 9052 18104 9061
rect 11704 9027 11756 9036
rect 10784 8984 10836 8993
rect 11704 8993 11713 9027
rect 11713 8993 11747 9027
rect 11747 8993 11756 9027
rect 11704 8984 11756 8993
rect 11888 8984 11940 9036
rect 13820 9027 13872 9036
rect 13820 8993 13829 9027
rect 13829 8993 13863 9027
rect 13863 8993 13872 9027
rect 15384 9027 15436 9036
rect 13820 8984 13872 8993
rect 15384 8993 15393 9027
rect 15393 8993 15427 9027
rect 15427 8993 15436 9027
rect 15384 8984 15436 8993
rect 17316 9027 17368 9036
rect 17316 8993 17325 9027
rect 17325 8993 17359 9027
rect 17359 8993 17368 9027
rect 17316 8984 17368 8993
rect 17684 8984 17736 9036
rect 19800 8984 19852 9036
rect 22192 8984 22244 9036
rect 3516 8848 3568 8900
rect 2780 8823 2832 8832
rect 2780 8789 2789 8823
rect 2789 8789 2823 8823
rect 2823 8789 2832 8823
rect 2780 8780 2832 8789
rect 4344 8848 4396 8900
rect 6644 8848 6696 8900
rect 12348 8916 12400 8968
rect 14556 8916 14608 8968
rect 11704 8848 11756 8900
rect 4620 8780 4672 8832
rect 5080 8823 5132 8832
rect 5080 8789 5089 8823
rect 5089 8789 5123 8823
rect 5123 8789 5132 8823
rect 5080 8780 5132 8789
rect 7196 8780 7248 8832
rect 7564 8780 7616 8832
rect 9220 8780 9272 8832
rect 13360 8780 13412 8832
rect 13728 8780 13780 8832
rect 15752 8823 15804 8832
rect 15752 8789 15761 8823
rect 15761 8789 15795 8823
rect 15795 8789 15804 8823
rect 15752 8780 15804 8789
rect 18788 8823 18840 8832
rect 18788 8789 18797 8823
rect 18797 8789 18831 8823
rect 18831 8789 18840 8823
rect 18788 8780 18840 8789
rect 19984 8780 20036 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 3240 8576 3292 8628
rect 3792 8576 3844 8628
rect 5356 8576 5408 8628
rect 5540 8576 5592 8628
rect 6000 8576 6052 8628
rect 6552 8619 6604 8628
rect 6552 8585 6561 8619
rect 6561 8585 6595 8619
rect 6595 8585 6604 8619
rect 6552 8576 6604 8585
rect 7104 8619 7156 8628
rect 7104 8585 7113 8619
rect 7113 8585 7147 8619
rect 7147 8585 7156 8619
rect 7104 8576 7156 8585
rect 2136 8483 2188 8492
rect 2136 8449 2145 8483
rect 2145 8449 2179 8483
rect 2179 8449 2188 8483
rect 2136 8440 2188 8449
rect 4712 8415 4764 8424
rect 4712 8381 4721 8415
rect 4721 8381 4755 8415
rect 4755 8381 4764 8415
rect 4712 8372 4764 8381
rect 5172 8415 5224 8424
rect 5172 8381 5181 8415
rect 5181 8381 5215 8415
rect 5215 8381 5224 8415
rect 5172 8372 5224 8381
rect 1768 8347 1820 8356
rect 1768 8313 1777 8347
rect 1777 8313 1811 8347
rect 1811 8313 1820 8347
rect 1768 8304 1820 8313
rect 1860 8347 1912 8356
rect 1860 8313 1869 8347
rect 1869 8313 1903 8347
rect 1903 8313 1912 8347
rect 1860 8304 1912 8313
rect 5080 8304 5132 8356
rect 5356 8372 5408 8424
rect 10048 8576 10100 8628
rect 10784 8576 10836 8628
rect 14464 8576 14516 8628
rect 15384 8619 15436 8628
rect 15384 8585 15393 8619
rect 15393 8585 15427 8619
rect 15427 8585 15436 8619
rect 15384 8576 15436 8585
rect 15752 8619 15804 8628
rect 15752 8585 15761 8619
rect 15761 8585 15795 8619
rect 15795 8585 15804 8619
rect 15752 8576 15804 8585
rect 17316 8619 17368 8628
rect 17316 8585 17325 8619
rect 17325 8585 17359 8619
rect 17359 8585 17368 8619
rect 17316 8576 17368 8585
rect 22192 8576 22244 8628
rect 23388 8576 23440 8628
rect 13820 8551 13872 8560
rect 13820 8517 13829 8551
rect 13829 8517 13863 8551
rect 13863 8517 13872 8551
rect 13820 8508 13872 8517
rect 16028 8508 16080 8560
rect 8576 8440 8628 8492
rect 7564 8372 7616 8424
rect 8392 8415 8444 8424
rect 8392 8381 8401 8415
rect 8401 8381 8435 8415
rect 8435 8381 8444 8415
rect 8392 8372 8444 8381
rect 9588 8440 9640 8492
rect 12348 8440 12400 8492
rect 15384 8440 15436 8492
rect 2872 8236 2924 8288
rect 3976 8236 4028 8288
rect 4252 8236 4304 8288
rect 9036 8304 9088 8356
rect 6000 8236 6052 8288
rect 7932 8236 7984 8288
rect 9312 8372 9364 8424
rect 11888 8372 11940 8424
rect 13360 8372 13412 8424
rect 17684 8508 17736 8560
rect 19800 8551 19852 8560
rect 19800 8517 19809 8551
rect 19809 8517 19843 8551
rect 19843 8517 19852 8551
rect 19800 8508 19852 8517
rect 20628 8508 20680 8560
rect 18788 8483 18840 8492
rect 18788 8449 18797 8483
rect 18797 8449 18831 8483
rect 18831 8449 18840 8483
rect 18788 8440 18840 8449
rect 19984 8483 20036 8492
rect 19984 8449 19993 8483
rect 19993 8449 20027 8483
rect 20027 8449 20036 8483
rect 19984 8440 20036 8449
rect 20168 8440 20220 8492
rect 18512 8415 18564 8424
rect 18512 8381 18521 8415
rect 18521 8381 18555 8415
rect 18555 8381 18564 8415
rect 18512 8372 18564 8381
rect 24124 8415 24176 8424
rect 24124 8381 24133 8415
rect 24133 8381 24167 8415
rect 24167 8381 24176 8415
rect 24124 8372 24176 8381
rect 9404 8347 9456 8356
rect 9404 8313 9413 8347
rect 9413 8313 9447 8347
rect 9447 8313 9456 8347
rect 9404 8304 9456 8313
rect 9956 8304 10008 8356
rect 10968 8304 11020 8356
rect 11152 8347 11204 8356
rect 11152 8313 11161 8347
rect 11161 8313 11195 8347
rect 11195 8313 11204 8347
rect 11152 8304 11204 8313
rect 14372 8347 14424 8356
rect 9588 8236 9640 8288
rect 14372 8313 14381 8347
rect 14381 8313 14415 8347
rect 14415 8313 14424 8347
rect 14372 8304 14424 8313
rect 14464 8347 14516 8356
rect 14464 8313 14473 8347
rect 14473 8313 14507 8347
rect 14507 8313 14516 8347
rect 15936 8347 15988 8356
rect 14464 8304 14516 8313
rect 15936 8313 15945 8347
rect 15945 8313 15979 8347
rect 15979 8313 15988 8347
rect 15936 8304 15988 8313
rect 20076 8347 20128 8356
rect 13636 8236 13688 8288
rect 15752 8236 15804 8288
rect 20076 8313 20085 8347
rect 20085 8313 20119 8347
rect 20119 8313 20128 8347
rect 20076 8304 20128 8313
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 2044 8075 2096 8084
rect 2044 8041 2053 8075
rect 2053 8041 2087 8075
rect 2087 8041 2096 8075
rect 2044 8032 2096 8041
rect 3516 8075 3568 8084
rect 3516 8041 3525 8075
rect 3525 8041 3559 8075
rect 3559 8041 3568 8075
rect 3516 8032 3568 8041
rect 3792 8075 3844 8084
rect 3792 8041 3801 8075
rect 3801 8041 3835 8075
rect 3835 8041 3844 8075
rect 3792 8032 3844 8041
rect 1860 7964 1912 8016
rect 2780 7964 2832 8016
rect 2964 8007 3016 8016
rect 2964 7973 2973 8007
rect 2973 7973 3007 8007
rect 3007 7973 3016 8007
rect 2964 7964 3016 7973
rect 4436 7964 4488 8016
rect 5448 7964 5500 8016
rect 4712 7896 4764 7948
rect 5264 7939 5316 7948
rect 5264 7905 5273 7939
rect 5273 7905 5307 7939
rect 5307 7905 5316 7939
rect 5264 7896 5316 7905
rect 6000 7939 6052 7948
rect 3148 7828 3200 7880
rect 4620 7828 4672 7880
rect 5172 7828 5224 7880
rect 6000 7905 6009 7939
rect 6009 7905 6043 7939
rect 6043 7905 6052 7939
rect 6000 7896 6052 7905
rect 7564 7939 7616 7948
rect 7564 7905 7573 7939
rect 7573 7905 7607 7939
rect 7607 7905 7616 7939
rect 7564 7896 7616 7905
rect 6460 7871 6512 7880
rect 3424 7760 3476 7812
rect 4068 7760 4120 7812
rect 5448 7760 5500 7812
rect 6460 7837 6469 7871
rect 6469 7837 6503 7871
rect 6503 7837 6512 7871
rect 6460 7828 6512 7837
rect 6368 7692 6420 7744
rect 7380 7828 7432 7880
rect 7840 7896 7892 7948
rect 12348 8032 12400 8084
rect 15936 8032 15988 8084
rect 16488 8032 16540 8084
rect 18512 8075 18564 8084
rect 18512 8041 18521 8075
rect 18521 8041 18555 8075
rect 18555 8041 18564 8075
rect 18512 8032 18564 8041
rect 20076 8032 20128 8084
rect 9956 7964 10008 8016
rect 11428 7964 11480 8016
rect 11796 7964 11848 8016
rect 13636 8007 13688 8016
rect 13636 7973 13639 8007
rect 13639 7973 13673 8007
rect 13673 7973 13688 8007
rect 13636 7964 13688 7973
rect 14004 7964 14056 8016
rect 15384 8007 15436 8016
rect 15384 7973 15393 8007
rect 15393 7973 15427 8007
rect 15427 7973 15436 8007
rect 15384 7964 15436 7973
rect 15476 8007 15528 8016
rect 15476 7973 15485 8007
rect 15485 7973 15519 8007
rect 15519 7973 15528 8007
rect 15476 7964 15528 7973
rect 8852 7896 8904 7948
rect 10968 7896 11020 7948
rect 11152 7828 11204 7880
rect 12808 7828 12860 7880
rect 13820 7896 13872 7948
rect 16856 7939 16908 7948
rect 16856 7905 16865 7939
rect 16865 7905 16899 7939
rect 16899 7905 16908 7939
rect 16856 7896 16908 7905
rect 16304 7828 16356 7880
rect 9220 7692 9272 7744
rect 10048 7735 10100 7744
rect 10048 7701 10057 7735
rect 10057 7701 10091 7735
rect 10091 7701 10100 7735
rect 10048 7692 10100 7701
rect 10968 7692 11020 7744
rect 12532 7692 12584 7744
rect 14372 7760 14424 7812
rect 15936 7803 15988 7812
rect 15936 7769 15945 7803
rect 15945 7769 15979 7803
rect 15979 7769 15988 7803
rect 15936 7760 15988 7769
rect 18144 7692 18196 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 2780 7531 2832 7540
rect 2780 7497 2789 7531
rect 2789 7497 2823 7531
rect 2823 7497 2832 7531
rect 2780 7488 2832 7497
rect 3516 7488 3568 7540
rect 4160 7488 4212 7540
rect 4620 7531 4672 7540
rect 4620 7497 4629 7531
rect 4629 7497 4663 7531
rect 4663 7497 4672 7531
rect 4620 7488 4672 7497
rect 5264 7488 5316 7540
rect 6552 7488 6604 7540
rect 9956 7488 10008 7540
rect 10968 7488 11020 7540
rect 11704 7531 11756 7540
rect 11704 7497 11713 7531
rect 11713 7497 11747 7531
rect 11747 7497 11756 7531
rect 11704 7488 11756 7497
rect 13452 7488 13504 7540
rect 16304 7531 16356 7540
rect 16304 7497 16313 7531
rect 16313 7497 16347 7531
rect 16347 7497 16356 7531
rect 16304 7488 16356 7497
rect 18604 7531 18656 7540
rect 18604 7497 18613 7531
rect 18613 7497 18647 7531
rect 18647 7497 18656 7531
rect 18604 7488 18656 7497
rect 4344 7420 4396 7472
rect 7840 7420 7892 7472
rect 1952 7352 2004 7404
rect 3976 7352 4028 7404
rect 2780 7284 2832 7336
rect 4712 7327 4764 7336
rect 4712 7293 4721 7327
rect 4721 7293 4755 7327
rect 4755 7293 4764 7327
rect 4712 7284 4764 7293
rect 5356 7284 5408 7336
rect 7748 7352 7800 7404
rect 7564 7284 7616 7336
rect 9220 7420 9272 7472
rect 13820 7463 13872 7472
rect 13820 7429 13829 7463
rect 13829 7429 13863 7463
rect 13863 7429 13872 7463
rect 13820 7420 13872 7429
rect 9404 7352 9456 7404
rect 10784 7352 10836 7404
rect 12808 7395 12860 7404
rect 12808 7361 12817 7395
rect 12817 7361 12851 7395
rect 12851 7361 12860 7395
rect 12808 7352 12860 7361
rect 16856 7420 16908 7472
rect 15936 7395 15988 7404
rect 15936 7361 15945 7395
rect 15945 7361 15979 7395
rect 15979 7361 15988 7395
rect 15936 7352 15988 7361
rect 8392 7327 8444 7336
rect 8392 7293 8401 7327
rect 8401 7293 8435 7327
rect 8435 7293 8444 7327
rect 8392 7284 8444 7293
rect 9128 7327 9180 7336
rect 5080 7216 5132 7268
rect 9128 7293 9137 7327
rect 9137 7293 9171 7327
rect 9171 7293 9180 7327
rect 9128 7284 9180 7293
rect 11428 7284 11480 7336
rect 13544 7284 13596 7336
rect 16120 7284 16172 7336
rect 18604 7284 18656 7336
rect 9312 7259 9364 7268
rect 3148 7191 3200 7200
rect 3148 7157 3157 7191
rect 3157 7157 3191 7191
rect 3191 7157 3200 7191
rect 3148 7148 3200 7157
rect 3516 7191 3568 7200
rect 3516 7157 3525 7191
rect 3525 7157 3559 7191
rect 3559 7157 3568 7191
rect 3516 7148 3568 7157
rect 6368 7148 6420 7200
rect 9312 7225 9321 7259
rect 9321 7225 9355 7259
rect 9355 7225 9364 7259
rect 9312 7216 9364 7225
rect 9588 7191 9640 7200
rect 9588 7157 9597 7191
rect 9597 7157 9631 7191
rect 9631 7157 9640 7191
rect 9588 7148 9640 7157
rect 9956 7191 10008 7200
rect 9956 7157 9965 7191
rect 9965 7157 9999 7191
rect 9999 7157 10008 7191
rect 9956 7148 10008 7157
rect 12164 7191 12216 7200
rect 12164 7157 12173 7191
rect 12173 7157 12207 7191
rect 12207 7157 12216 7191
rect 12164 7148 12216 7157
rect 12440 7148 12492 7200
rect 12624 7259 12676 7268
rect 12624 7225 12633 7259
rect 12633 7225 12667 7259
rect 12667 7225 12676 7259
rect 12624 7216 12676 7225
rect 15384 7259 15436 7268
rect 15384 7225 15393 7259
rect 15393 7225 15427 7259
rect 15427 7225 15436 7259
rect 15384 7216 15436 7225
rect 16948 7216 17000 7268
rect 13452 7191 13504 7200
rect 13452 7157 13461 7191
rect 13461 7157 13495 7191
rect 13495 7157 13504 7191
rect 13452 7148 13504 7157
rect 15476 7148 15528 7200
rect 18604 7148 18656 7200
rect 25136 7191 25188 7200
rect 25136 7157 25145 7191
rect 25145 7157 25179 7191
rect 25179 7157 25188 7191
rect 25136 7148 25188 7157
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 3516 6944 3568 6996
rect 4068 6944 4120 6996
rect 6644 6987 6696 6996
rect 6644 6953 6653 6987
rect 6653 6953 6687 6987
rect 6687 6953 6696 6987
rect 6644 6944 6696 6953
rect 8392 6944 8444 6996
rect 8852 6987 8904 6996
rect 8852 6953 8861 6987
rect 8861 6953 8895 6987
rect 8895 6953 8904 6987
rect 8852 6944 8904 6953
rect 9220 6987 9272 6996
rect 9220 6953 9229 6987
rect 9229 6953 9263 6987
rect 9263 6953 9272 6987
rect 9220 6944 9272 6953
rect 9956 6944 10008 6996
rect 10968 6944 11020 6996
rect 11152 6944 11204 6996
rect 13084 6944 13136 6996
rect 15292 6944 15344 6996
rect 15384 6944 15436 6996
rect 24768 6987 24820 6996
rect 24768 6953 24777 6987
rect 24777 6953 24811 6987
rect 24811 6953 24820 6987
rect 24768 6944 24820 6953
rect 1860 6919 1912 6928
rect 1860 6885 1869 6919
rect 1869 6885 1903 6919
rect 1903 6885 1912 6919
rect 1860 6876 1912 6885
rect 2964 6876 3016 6928
rect 4712 6876 4764 6928
rect 5540 6919 5592 6928
rect 5540 6885 5549 6919
rect 5549 6885 5583 6919
rect 5583 6885 5592 6919
rect 5540 6876 5592 6885
rect 2596 6808 2648 6860
rect 2780 6808 2832 6860
rect 4528 6808 4580 6860
rect 6736 6876 6788 6928
rect 6552 6808 6604 6860
rect 7748 6876 7800 6928
rect 10784 6876 10836 6928
rect 12164 6919 12216 6928
rect 12164 6885 12173 6919
rect 12173 6885 12207 6919
rect 12207 6885 12216 6919
rect 12164 6876 12216 6885
rect 12624 6876 12676 6928
rect 7288 6808 7340 6860
rect 9128 6808 9180 6860
rect 11428 6808 11480 6860
rect 12992 6851 13044 6860
rect 12992 6817 13001 6851
rect 13001 6817 13035 6851
rect 13035 6817 13044 6851
rect 12992 6808 13044 6817
rect 13268 6851 13320 6860
rect 13268 6817 13277 6851
rect 13277 6817 13311 6851
rect 13311 6817 13320 6851
rect 13268 6808 13320 6817
rect 15476 6851 15528 6860
rect 15476 6817 15485 6851
rect 15485 6817 15519 6851
rect 15519 6817 15528 6851
rect 15476 6808 15528 6817
rect 15936 6808 15988 6860
rect 16856 6851 16908 6860
rect 16856 6817 16900 6851
rect 16900 6817 16908 6851
rect 16856 6808 16908 6817
rect 24676 6808 24728 6860
rect 3240 6604 3292 6656
rect 4620 6647 4672 6656
rect 4620 6613 4629 6647
rect 4629 6613 4663 6647
rect 4663 6613 4672 6647
rect 4620 6604 4672 6613
rect 5540 6604 5592 6656
rect 6000 6604 6052 6656
rect 8116 6740 8168 6792
rect 9312 6740 9364 6792
rect 11244 6740 11296 6792
rect 11704 6740 11756 6792
rect 14004 6672 14056 6724
rect 11428 6604 11480 6656
rect 12440 6647 12492 6656
rect 12440 6613 12449 6647
rect 12449 6613 12483 6647
rect 12483 6613 12492 6647
rect 12440 6604 12492 6613
rect 14464 6604 14516 6656
rect 18052 6604 18104 6656
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 1584 6443 1636 6452
rect 1584 6409 1593 6443
rect 1593 6409 1627 6443
rect 1627 6409 1636 6443
rect 1584 6400 1636 6409
rect 6000 6400 6052 6452
rect 6552 6400 6604 6452
rect 10048 6443 10100 6452
rect 10048 6409 10057 6443
rect 10057 6409 10091 6443
rect 10091 6409 10100 6443
rect 10048 6400 10100 6409
rect 11244 6443 11296 6452
rect 11244 6409 11253 6443
rect 11253 6409 11287 6443
rect 11287 6409 11296 6443
rect 11244 6400 11296 6409
rect 14004 6443 14056 6452
rect 14004 6409 14013 6443
rect 14013 6409 14047 6443
rect 14047 6409 14056 6443
rect 14004 6400 14056 6409
rect 15476 6400 15528 6452
rect 16856 6443 16908 6452
rect 16856 6409 16865 6443
rect 16865 6409 16899 6443
rect 16899 6409 16908 6443
rect 16856 6400 16908 6409
rect 23848 6400 23900 6452
rect 3332 6332 3384 6384
rect 4528 6332 4580 6384
rect 6460 6332 6512 6384
rect 1308 6196 1360 6248
rect 2688 6128 2740 6180
rect 3240 6196 3292 6248
rect 3424 6264 3476 6316
rect 5080 6307 5132 6316
rect 5080 6273 5089 6307
rect 5089 6273 5123 6307
rect 5123 6273 5132 6307
rect 5080 6264 5132 6273
rect 6736 6264 6788 6316
rect 4620 6239 4672 6248
rect 3792 6171 3844 6180
rect 2780 6060 2832 6112
rect 3792 6137 3801 6171
rect 3801 6137 3835 6171
rect 3835 6137 3844 6171
rect 3792 6128 3844 6137
rect 4620 6205 4629 6239
rect 4629 6205 4663 6239
rect 4663 6205 4672 6239
rect 4620 6196 4672 6205
rect 4896 6239 4948 6248
rect 4896 6205 4905 6239
rect 4905 6205 4939 6239
rect 4939 6205 4948 6239
rect 4896 6196 4948 6205
rect 10692 6264 10744 6316
rect 11152 6264 11204 6316
rect 15844 6264 15896 6316
rect 7748 6239 7800 6248
rect 7748 6205 7757 6239
rect 7757 6205 7791 6239
rect 7791 6205 7800 6239
rect 7748 6196 7800 6205
rect 8116 6239 8168 6248
rect 8116 6205 8125 6239
rect 8125 6205 8159 6239
rect 8159 6205 8168 6239
rect 8116 6196 8168 6205
rect 8668 6239 8720 6248
rect 8668 6205 8677 6239
rect 8677 6205 8711 6239
rect 8711 6205 8720 6239
rect 8668 6196 8720 6205
rect 14464 6239 14516 6248
rect 4160 6060 4212 6112
rect 6276 6128 6328 6180
rect 7932 6128 7984 6180
rect 7288 6060 7340 6112
rect 7564 6103 7616 6112
rect 7564 6069 7573 6103
rect 7573 6069 7607 6103
rect 7607 6069 7616 6103
rect 7564 6060 7616 6069
rect 8024 6060 8076 6112
rect 9956 6060 10008 6112
rect 10048 6060 10100 6112
rect 12256 6103 12308 6112
rect 12256 6069 12265 6103
rect 12265 6069 12299 6103
rect 12299 6069 12308 6103
rect 13452 6128 13504 6180
rect 14188 6171 14240 6180
rect 14188 6137 14197 6171
rect 14197 6137 14231 6171
rect 14231 6137 14240 6171
rect 14188 6128 14240 6137
rect 14464 6205 14473 6239
rect 14473 6205 14507 6239
rect 14507 6205 14516 6239
rect 14464 6196 14516 6205
rect 18052 6239 18104 6248
rect 18052 6205 18061 6239
rect 18061 6205 18095 6239
rect 18095 6205 18104 6239
rect 18052 6196 18104 6205
rect 24124 6239 24176 6248
rect 24124 6205 24133 6239
rect 24133 6205 24167 6239
rect 24167 6205 24176 6239
rect 24124 6196 24176 6205
rect 15660 6128 15712 6180
rect 16856 6128 16908 6180
rect 18972 6128 19024 6180
rect 24676 6128 24728 6180
rect 12256 6060 12308 6069
rect 13268 6060 13320 6112
rect 14004 6060 14056 6112
rect 18236 6103 18288 6112
rect 18236 6069 18245 6103
rect 18245 6069 18279 6103
rect 18279 6069 18288 6103
rect 18236 6060 18288 6069
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 3424 5899 3476 5908
rect 3424 5865 3433 5899
rect 3433 5865 3467 5899
rect 3467 5865 3476 5899
rect 3424 5856 3476 5865
rect 4896 5856 4948 5908
rect 5448 5856 5500 5908
rect 6736 5856 6788 5908
rect 7748 5856 7800 5908
rect 11428 5899 11480 5908
rect 3240 5788 3292 5840
rect 8024 5788 8076 5840
rect 11428 5865 11437 5899
rect 11437 5865 11471 5899
rect 11471 5865 11480 5899
rect 11428 5856 11480 5865
rect 9864 5831 9916 5840
rect 9864 5797 9873 5831
rect 9873 5797 9907 5831
rect 9907 5797 9916 5831
rect 9864 5788 9916 5797
rect 12256 5788 12308 5840
rect 12992 5788 13044 5840
rect 13728 5856 13780 5908
rect 14464 5788 14516 5840
rect 15476 5831 15528 5840
rect 15476 5797 15485 5831
rect 15485 5797 15519 5831
rect 15519 5797 15528 5831
rect 15476 5788 15528 5797
rect 2780 5763 2832 5772
rect 2780 5729 2789 5763
rect 2789 5729 2823 5763
rect 2823 5729 2832 5763
rect 2780 5720 2832 5729
rect 4160 5763 4212 5772
rect 4160 5729 4169 5763
rect 4169 5729 4203 5763
rect 4203 5729 4212 5763
rect 4160 5720 4212 5729
rect 6276 5720 6328 5772
rect 6552 5720 6604 5772
rect 7564 5720 7616 5772
rect 8392 5720 8444 5772
rect 12164 5763 12216 5772
rect 9312 5652 9364 5704
rect 10968 5652 11020 5704
rect 9036 5584 9088 5636
rect 12164 5729 12173 5763
rect 12173 5729 12207 5763
rect 12207 5729 12216 5763
rect 12164 5720 12216 5729
rect 13176 5720 13228 5772
rect 13728 5720 13780 5772
rect 15384 5695 15436 5704
rect 15384 5661 15393 5695
rect 15393 5661 15427 5695
rect 15427 5661 15436 5695
rect 15384 5652 15436 5661
rect 16028 5695 16080 5704
rect 16028 5661 16037 5695
rect 16037 5661 16071 5695
rect 16071 5661 16080 5695
rect 16028 5652 16080 5661
rect 7196 5516 7248 5568
rect 10692 5559 10744 5568
rect 10692 5525 10701 5559
rect 10701 5525 10735 5559
rect 10735 5525 10744 5559
rect 10692 5516 10744 5525
rect 14464 5559 14516 5568
rect 14464 5525 14473 5559
rect 14473 5525 14507 5559
rect 14507 5525 14516 5559
rect 14464 5516 14516 5525
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 5540 5312 5592 5364
rect 6368 5312 6420 5364
rect 9956 5312 10008 5364
rect 12256 5312 12308 5364
rect 13728 5312 13780 5364
rect 15384 5312 15436 5364
rect 2044 5176 2096 5228
rect 4160 5176 4212 5228
rect 2688 5108 2740 5160
rect 3792 5108 3844 5160
rect 6000 5244 6052 5296
rect 6276 5287 6328 5296
rect 6276 5253 6285 5287
rect 6285 5253 6319 5287
rect 6319 5253 6328 5287
rect 6276 5244 6328 5253
rect 6644 5176 6696 5228
rect 10968 5176 11020 5228
rect 15660 5287 15712 5296
rect 15660 5253 15669 5287
rect 15669 5253 15703 5287
rect 15703 5253 15712 5287
rect 15660 5244 15712 5253
rect 15476 5176 15528 5228
rect 5356 5040 5408 5092
rect 6552 5083 6604 5092
rect 6552 5049 6561 5083
rect 6561 5049 6595 5083
rect 6595 5049 6604 5083
rect 6552 5040 6604 5049
rect 6828 5040 6880 5092
rect 8024 5083 8076 5092
rect 8024 5049 8033 5083
rect 8033 5049 8067 5083
rect 8067 5049 8076 5083
rect 8024 5040 8076 5049
rect 8668 5083 8720 5092
rect 8668 5049 8677 5083
rect 8677 5049 8711 5083
rect 8711 5049 8720 5083
rect 8668 5040 8720 5049
rect 9312 5083 9364 5092
rect 2044 5015 2096 5024
rect 2044 4981 2053 5015
rect 2053 4981 2087 5015
rect 2087 4981 2096 5015
rect 2044 4972 2096 4981
rect 2780 4972 2832 5024
rect 7748 5015 7800 5024
rect 7748 4981 7757 5015
rect 7757 4981 7791 5015
rect 7791 4981 7800 5015
rect 7748 4972 7800 4981
rect 8300 4972 8352 5024
rect 9312 5049 9321 5083
rect 9321 5049 9355 5083
rect 9355 5049 9364 5083
rect 9312 5040 9364 5049
rect 10048 5040 10100 5092
rect 12808 5083 12860 5092
rect 9956 5015 10008 5024
rect 9956 4981 9965 5015
rect 9965 4981 9999 5015
rect 9999 4981 10008 5015
rect 12808 5049 12817 5083
rect 12817 5049 12851 5083
rect 12851 5049 12860 5083
rect 12808 5040 12860 5049
rect 12900 5083 12952 5092
rect 12900 5049 12909 5083
rect 12909 5049 12943 5083
rect 12943 5049 12952 5083
rect 14372 5083 14424 5092
rect 12900 5040 12952 5049
rect 14372 5049 14381 5083
rect 14381 5049 14415 5083
rect 14415 5049 14424 5083
rect 14372 5040 14424 5049
rect 14464 5083 14516 5092
rect 14464 5049 14473 5083
rect 14473 5049 14507 5083
rect 14507 5049 14516 5083
rect 14464 5040 14516 5049
rect 11152 5015 11204 5024
rect 9956 4972 10008 4981
rect 11152 4981 11161 5015
rect 11161 4981 11195 5015
rect 11195 4981 11204 5015
rect 11152 4972 11204 4981
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 6644 4768 6696 4820
rect 8392 4811 8444 4820
rect 8392 4777 8401 4811
rect 8401 4777 8435 4811
rect 8435 4777 8444 4811
rect 8392 4768 8444 4777
rect 9956 4811 10008 4820
rect 9956 4777 9965 4811
rect 9965 4777 9999 4811
rect 9999 4777 10008 4811
rect 9956 4768 10008 4777
rect 12532 4768 12584 4820
rect 14372 4768 14424 4820
rect 14740 4768 14792 4820
rect 2688 4700 2740 4752
rect 7196 4700 7248 4752
rect 7748 4700 7800 4752
rect 9312 4700 9364 4752
rect 12164 4743 12216 4752
rect 12164 4709 12173 4743
rect 12173 4709 12207 4743
rect 12207 4709 12216 4743
rect 12164 4700 12216 4709
rect 14188 4700 14240 4752
rect 15660 4700 15712 4752
rect 16028 4743 16080 4752
rect 16028 4709 16037 4743
rect 16037 4709 16071 4743
rect 16071 4709 16080 4743
rect 16028 4700 16080 4709
rect 27620 4700 27672 4752
rect 1492 4675 1544 4684
rect 1492 4641 1501 4675
rect 1501 4641 1535 4675
rect 1535 4641 1544 4675
rect 1492 4632 1544 4641
rect 5448 4632 5500 4684
rect 9864 4632 9916 4684
rect 10324 4675 10376 4684
rect 10324 4641 10333 4675
rect 10333 4641 10367 4675
rect 10367 4641 10376 4675
rect 10324 4632 10376 4641
rect 11152 4632 11204 4684
rect 11520 4632 11572 4684
rect 11980 4632 12032 4684
rect 24676 4675 24728 4684
rect 24676 4641 24694 4675
rect 24694 4641 24728 4675
rect 24676 4632 24728 4641
rect 8668 4564 8720 4616
rect 13728 4607 13780 4616
rect 13728 4573 13737 4607
rect 13737 4573 13771 4607
rect 13771 4573 13780 4607
rect 13728 4564 13780 4573
rect 14556 4564 14608 4616
rect 1676 4496 1728 4548
rect 2872 4496 2924 4548
rect 6828 4539 6880 4548
rect 6828 4505 6837 4539
rect 6837 4505 6871 4539
rect 6871 4505 6880 4539
rect 6828 4496 6880 4505
rect 12900 4496 12952 4548
rect 14188 4496 14240 4548
rect 2780 4471 2832 4480
rect 2780 4437 2789 4471
rect 2789 4437 2823 4471
rect 2823 4437 2832 4471
rect 2780 4428 2832 4437
rect 21548 4428 21600 4480
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 5448 4224 5500 4276
rect 7748 4224 7800 4276
rect 10692 4224 10744 4276
rect 11520 4224 11572 4276
rect 11980 4224 12032 4276
rect 14188 4224 14240 4276
rect 15660 4224 15712 4276
rect 24676 4267 24728 4276
rect 24676 4233 24685 4267
rect 24685 4233 24719 4267
rect 24719 4233 24728 4267
rect 24676 4224 24728 4233
rect 10324 4156 10376 4208
rect 14464 4156 14516 4208
rect 8300 4088 8352 4140
rect 7748 4020 7800 4072
rect 6552 3952 6604 4004
rect 9864 4088 9916 4140
rect 10048 4088 10100 4140
rect 12440 4088 12492 4140
rect 12808 4088 12860 4140
rect 14556 4131 14608 4140
rect 14556 4097 14565 4131
rect 14565 4097 14599 4131
rect 14599 4097 14608 4131
rect 14556 4088 14608 4097
rect 14280 3995 14332 4004
rect 14280 3961 14289 3995
rect 14289 3961 14323 3995
rect 14323 3961 14332 3995
rect 14280 3952 14332 3961
rect 14464 3952 14516 4004
rect 14740 3952 14792 4004
rect 21548 3952 21600 4004
rect 1492 3884 1544 3936
rect 9588 3927 9640 3936
rect 9588 3893 9597 3927
rect 9597 3893 9631 3927
rect 9631 3893 9640 3927
rect 9588 3884 9640 3893
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 1768 3680 1820 3732
rect 7196 3680 7248 3732
rect 13728 3723 13780 3732
rect 13728 3689 13737 3723
rect 13737 3689 13771 3723
rect 13771 3689 13780 3723
rect 13728 3680 13780 3689
rect 1400 3587 1452 3596
rect 1400 3553 1409 3587
rect 1409 3553 1443 3587
rect 1443 3553 1452 3587
rect 1400 3544 1452 3553
rect 15384 3587 15436 3596
rect 15384 3553 15402 3587
rect 15402 3553 15436 3587
rect 15384 3544 15436 3553
rect 16028 3544 16080 3596
rect 24676 3587 24728 3596
rect 24676 3553 24694 3587
rect 24694 3553 24728 3587
rect 24676 3544 24728 3553
rect 27620 3544 27672 3596
rect 14280 3451 14332 3460
rect 14280 3417 14289 3451
rect 14289 3417 14323 3451
rect 14323 3417 14332 3451
rect 14280 3408 14332 3417
rect 15660 3340 15712 3392
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 112 3068 164 3120
rect 1400 3068 1452 3120
rect 9864 3136 9916 3188
rect 10784 3068 10836 3120
rect 11980 3136 12032 3188
rect 15384 3179 15436 3188
rect 15384 3145 15393 3179
rect 15393 3145 15427 3179
rect 15427 3145 15436 3179
rect 15384 3136 15436 3145
rect 24676 3179 24728 3188
rect 24676 3145 24685 3179
rect 24685 3145 24719 3179
rect 24719 3145 24728 3179
rect 24676 3136 24728 3145
rect 12072 3068 12124 3120
rect 13912 3068 13964 3120
rect 23112 3068 23164 3120
rect 15660 2975 15712 2984
rect 15660 2941 15669 2975
rect 15669 2941 15703 2975
rect 15703 2941 15712 2975
rect 15660 2932 15712 2941
rect 16764 2796 16816 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 848 2592 900 2644
rect 1492 2592 1544 2644
rect 14832 2635 14884 2644
rect 14832 2601 14841 2635
rect 14841 2601 14875 2635
rect 14875 2601 14884 2635
rect 14832 2592 14884 2601
rect 16396 2592 16448 2644
rect 20260 2592 20312 2644
rect 21364 2592 21416 2644
rect 7564 2499 7616 2508
rect 7564 2465 7573 2499
rect 7573 2465 7607 2499
rect 7607 2465 7616 2499
rect 7564 2456 7616 2465
rect 8944 2456 8996 2508
rect 16672 2456 16724 2508
rect 4712 2320 4764 2372
rect 8944 2320 8996 2372
rect 13360 2320 13412 2372
rect 21824 2320 21876 2372
rect 6828 2252 6880 2304
rect 14648 2252 14700 2304
rect 16672 2295 16724 2304
rect 16672 2261 16681 2295
rect 16681 2261 16715 2295
rect 16715 2261 16724 2295
rect 16672 2252 16724 2261
rect 17684 2252 17736 2304
rect 24768 2524 24820 2576
rect 23020 2252 23072 2304
rect 23112 2252 23164 2304
rect 25596 2252 25648 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 18236 416 18288 468
rect 19340 416 19392 468
rect 15752 76 15804 128
rect 17408 76 17460 128
<< metal2 >>
rect 20 27532 72 27538
rect 662 27532 718 28000
rect 662 27520 664 27532
rect 20 27474 72 27480
rect 716 27520 718 27532
rect 2042 27554 2098 28000
rect 2042 27526 2452 27554
rect 2042 27520 2098 27526
rect 664 27474 716 27480
rect 32 10810 60 27474
rect 676 27443 704 27474
rect 1214 26888 1270 26897
rect 1214 26823 1270 26832
rect 110 24576 166 24585
rect 110 24511 166 24520
rect 124 22574 152 24511
rect 1228 23186 1256 26823
rect 1306 25392 1362 25401
rect 1306 25327 1362 25336
rect 1320 23730 1348 25327
rect 1308 23724 1360 23730
rect 1308 23666 1360 23672
rect 1676 23520 1728 23526
rect 1676 23462 1728 23468
rect 1216 23180 1268 23186
rect 1216 23122 1268 23128
rect 1214 22672 1270 22681
rect 1214 22607 1270 22616
rect 112 22568 164 22574
rect 112 22510 164 22516
rect 1228 21078 1256 22607
rect 1216 21072 1268 21078
rect 1216 21014 1268 21020
rect 1228 20602 1256 21014
rect 1216 20596 1268 20602
rect 1216 20538 1268 20544
rect 1582 20088 1638 20097
rect 1582 20023 1638 20032
rect 1596 19514 1624 20023
rect 1584 19508 1636 19514
rect 1584 19450 1636 19456
rect 1306 18728 1362 18737
rect 1306 18663 1362 18672
rect 204 15904 256 15910
rect 204 15846 256 15852
rect 110 13968 166 13977
rect 110 13903 166 13912
rect 124 13870 152 13903
rect 112 13864 164 13870
rect 112 13806 164 13812
rect 20 10804 72 10810
rect 20 10746 72 10752
rect 110 10160 166 10169
rect 110 10095 166 10104
rect 124 9897 152 10095
rect 110 9888 166 9897
rect 110 9823 166 9832
rect 110 8528 166 8537
rect 216 8514 244 15846
rect 1320 15065 1348 18663
rect 1688 16522 1716 23462
rect 2228 23180 2280 23186
rect 2228 23122 2280 23128
rect 2240 22778 2268 23122
rect 2228 22772 2280 22778
rect 2228 22714 2280 22720
rect 1768 22432 1820 22438
rect 1768 22374 1820 22380
rect 1780 21593 1808 22374
rect 1766 21584 1822 21593
rect 1766 21519 1822 21528
rect 1952 19168 2004 19174
rect 1952 19110 2004 19116
rect 1676 16516 1728 16522
rect 1676 16458 1728 16464
rect 1400 16448 1452 16454
rect 1400 16390 1452 16396
rect 1412 16046 1440 16390
rect 1400 16040 1452 16046
rect 1400 15982 1452 15988
rect 1412 15706 1440 15982
rect 1400 15700 1452 15706
rect 1400 15642 1452 15648
rect 1306 15056 1362 15065
rect 1306 14991 1362 15000
rect 1308 14952 1360 14958
rect 1308 14894 1360 14900
rect 938 14784 994 14793
rect 938 14719 994 14728
rect 952 14618 980 14719
rect 940 14612 992 14618
rect 940 14554 992 14560
rect 1320 12345 1348 14894
rect 1584 14816 1636 14822
rect 1584 14758 1636 14764
rect 1596 12782 1624 14758
rect 1860 13184 1912 13190
rect 1860 13126 1912 13132
rect 1584 12776 1636 12782
rect 1584 12718 1636 12724
rect 1306 12336 1362 12345
rect 1306 12271 1362 12280
rect 1400 12300 1452 12306
rect 166 8486 244 8514
rect 110 8463 166 8472
rect 1320 6254 1348 12271
rect 1400 12242 1452 12248
rect 1412 11762 1440 12242
rect 1400 11756 1452 11762
rect 1400 11698 1452 11704
rect 1596 11150 1624 12718
rect 1768 12708 1820 12714
rect 1768 12650 1820 12656
rect 1780 12442 1808 12650
rect 1768 12436 1820 12442
rect 1768 12378 1820 12384
rect 1872 11694 1900 13126
rect 1964 12986 1992 19110
rect 2044 17536 2096 17542
rect 2044 17478 2096 17484
rect 2056 16658 2084 17478
rect 2044 16652 2096 16658
rect 2044 16594 2096 16600
rect 2056 16250 2084 16594
rect 2044 16244 2096 16250
rect 2044 16186 2096 16192
rect 2134 14512 2190 14521
rect 2134 14447 2136 14456
rect 2188 14447 2190 14456
rect 2136 14418 2188 14424
rect 2044 14272 2096 14278
rect 2044 14214 2096 14220
rect 1952 12980 2004 12986
rect 1952 12922 2004 12928
rect 1860 11688 1912 11694
rect 1860 11630 1912 11636
rect 1872 11354 1900 11630
rect 1860 11348 1912 11354
rect 1860 11290 1912 11296
rect 1952 11280 2004 11286
rect 2056 11268 2084 14214
rect 2148 14006 2176 14418
rect 2424 14006 2452 27526
rect 3422 27520 3478 28000
rect 4802 27520 4858 28000
rect 6182 27554 6238 28000
rect 7654 27554 7710 28000
rect 6012 27526 6238 27554
rect 3436 22681 3464 27520
rect 3422 22672 3478 22681
rect 3422 22607 3478 22616
rect 4066 21312 4122 21321
rect 4066 21247 4122 21256
rect 4080 20602 4108 21247
rect 4068 20596 4120 20602
rect 4068 20538 4120 20544
rect 4160 20460 4212 20466
rect 4160 20402 4212 20408
rect 3976 19848 4028 19854
rect 3976 19790 4028 19796
rect 3884 19780 3936 19786
rect 3884 19722 3936 19728
rect 3896 19242 3924 19722
rect 3988 19514 4016 19790
rect 4172 19514 4200 20402
rect 4344 19984 4396 19990
rect 4344 19926 4396 19932
rect 3976 19508 4028 19514
rect 3976 19450 4028 19456
rect 4160 19508 4212 19514
rect 4160 19450 4212 19456
rect 3884 19236 3936 19242
rect 3884 19178 3936 19184
rect 3988 18970 4016 19450
rect 4356 19174 4384 19926
rect 4344 19168 4396 19174
rect 4344 19110 4396 19116
rect 3976 18964 4028 18970
rect 3976 18906 4028 18912
rect 4160 18624 4212 18630
rect 4160 18566 4212 18572
rect 3240 16992 3292 16998
rect 3240 16934 3292 16940
rect 2964 15564 3016 15570
rect 2964 15506 3016 15512
rect 2976 14822 3004 15506
rect 3148 15360 3200 15366
rect 3148 15302 3200 15308
rect 2964 14816 3016 14822
rect 2964 14758 3016 14764
rect 2136 14000 2188 14006
rect 2136 13942 2188 13948
rect 2412 14000 2464 14006
rect 2412 13942 2464 13948
rect 2424 13394 2452 13942
rect 2872 13864 2924 13870
rect 2872 13806 2924 13812
rect 2228 13388 2280 13394
rect 2228 13330 2280 13336
rect 2412 13388 2464 13394
rect 2412 13330 2464 13336
rect 2240 13297 2268 13330
rect 2226 13288 2282 13297
rect 2226 13223 2282 13232
rect 2136 13184 2188 13190
rect 2136 13126 2188 13132
rect 2004 11240 2084 11268
rect 1952 11222 2004 11228
rect 1584 11144 1636 11150
rect 1584 11086 1636 11092
rect 2056 10742 2084 11240
rect 2044 10736 2096 10742
rect 2044 10678 2096 10684
rect 2056 10520 2084 10678
rect 2148 10674 2176 13126
rect 2240 12442 2268 13223
rect 2424 12986 2452 13330
rect 2884 13190 2912 13806
rect 2504 13184 2556 13190
rect 2504 13126 2556 13132
rect 2872 13184 2924 13190
rect 2872 13126 2924 13132
rect 2412 12980 2464 12986
rect 2412 12922 2464 12928
rect 2228 12436 2280 12442
rect 2228 12378 2280 12384
rect 2412 12300 2464 12306
rect 2412 12242 2464 12248
rect 2424 11898 2452 12242
rect 2516 12238 2544 13126
rect 2884 12918 2912 13126
rect 2872 12912 2924 12918
rect 2872 12854 2924 12860
rect 2596 12776 2648 12782
rect 2596 12718 2648 12724
rect 2608 12374 2636 12718
rect 2976 12714 3004 14758
rect 3056 13728 3108 13734
rect 3056 13670 3108 13676
rect 3068 13530 3096 13670
rect 3056 13524 3108 13530
rect 3056 13466 3108 13472
rect 2964 12708 3016 12714
rect 2964 12650 3016 12656
rect 3160 12442 3188 15302
rect 3252 14958 3280 16934
rect 3424 15360 3476 15366
rect 3424 15302 3476 15308
rect 3240 14952 3292 14958
rect 3240 14894 3292 14900
rect 3436 14618 3464 15302
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 3608 14816 3660 14822
rect 3608 14758 3660 14764
rect 3620 14618 3648 14758
rect 3424 14612 3476 14618
rect 3424 14554 3476 14560
rect 3608 14612 3660 14618
rect 3608 14554 3660 14560
rect 3424 14476 3476 14482
rect 3424 14418 3476 14424
rect 3436 13841 3464 14418
rect 4080 14278 4108 14894
rect 4068 14272 4120 14278
rect 4068 14214 4120 14220
rect 3422 13832 3478 13841
rect 3422 13767 3478 13776
rect 3436 13734 3464 13767
rect 3424 13728 3476 13734
rect 3424 13670 3476 13676
rect 3884 12640 3936 12646
rect 3884 12582 3936 12588
rect 3148 12436 3200 12442
rect 3148 12378 3200 12384
rect 2596 12368 2648 12374
rect 2596 12310 2648 12316
rect 3056 12300 3108 12306
rect 3056 12242 3108 12248
rect 2504 12232 2556 12238
rect 2504 12174 2556 12180
rect 3068 12170 3096 12242
rect 3148 12232 3200 12238
rect 3148 12174 3200 12180
rect 3056 12164 3108 12170
rect 3056 12106 3108 12112
rect 2412 11892 2464 11898
rect 2412 11834 2464 11840
rect 2228 11552 2280 11558
rect 2228 11494 2280 11500
rect 2136 10668 2188 10674
rect 2136 10610 2188 10616
rect 2056 10492 2176 10520
rect 1952 10464 2004 10470
rect 1952 10406 2004 10412
rect 1860 10124 1912 10130
rect 1860 10066 1912 10072
rect 1768 9920 1820 9926
rect 1768 9862 1820 9868
rect 1780 8362 1808 9862
rect 1872 9178 1900 10066
rect 1860 9172 1912 9178
rect 1860 9114 1912 9120
rect 1768 8356 1820 8362
rect 1768 8298 1820 8304
rect 1860 8356 1912 8362
rect 1860 8298 1912 8304
rect 1582 6760 1638 6769
rect 1582 6695 1638 6704
rect 1596 6458 1624 6695
rect 1584 6452 1636 6458
rect 1584 6394 1636 6400
rect 1308 6248 1360 6254
rect 1308 6190 1360 6196
rect 1492 4684 1544 4690
rect 1492 4626 1544 4632
rect 1504 3942 1532 4626
rect 1676 4548 1728 4554
rect 1676 4490 1728 4496
rect 1492 3936 1544 3942
rect 1492 3878 1544 3884
rect 1400 3596 1452 3602
rect 1400 3538 1452 3544
rect 110 3224 166 3233
rect 110 3159 166 3168
rect 124 3126 152 3159
rect 1412 3126 1440 3538
rect 112 3120 164 3126
rect 112 3062 164 3068
rect 1400 3120 1452 3126
rect 1400 3062 1452 3068
rect 1504 2650 1532 3878
rect 848 2644 900 2650
rect 848 2586 900 2592
rect 1492 2644 1544 2650
rect 1492 2586 1544 2592
rect 570 82 626 480
rect 860 82 888 2586
rect 570 54 888 82
rect 1688 82 1716 4490
rect 1780 3738 1808 8298
rect 1872 8022 1900 8298
rect 1860 8016 1912 8022
rect 1860 7958 1912 7964
rect 1872 6934 1900 7958
rect 1964 7410 1992 10406
rect 2044 10192 2096 10198
rect 2044 10134 2096 10140
rect 2056 9382 2084 10134
rect 2044 9376 2096 9382
rect 2044 9318 2096 9324
rect 2056 9178 2084 9318
rect 2044 9172 2096 9178
rect 2044 9114 2096 9120
rect 2044 9036 2096 9042
rect 2044 8978 2096 8984
rect 2056 8090 2084 8978
rect 2148 8498 2176 10492
rect 2240 9450 2268 11494
rect 3068 11354 3096 12106
rect 3056 11348 3108 11354
rect 3056 11290 3108 11296
rect 2780 11280 2832 11286
rect 2780 11222 2832 11228
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 2332 9586 2360 11086
rect 2792 10266 2820 11222
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 3160 10169 3188 12174
rect 3792 11756 3844 11762
rect 3896 11744 3924 12582
rect 3976 12436 4028 12442
rect 3976 12378 4028 12384
rect 3844 11716 3924 11744
rect 3792 11698 3844 11704
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 3240 10804 3292 10810
rect 3240 10746 3292 10752
rect 3146 10160 3202 10169
rect 3252 10130 3280 10746
rect 3146 10095 3202 10104
rect 3240 10124 3292 10130
rect 3240 10066 3292 10072
rect 2964 9648 3016 9654
rect 2964 9590 3016 9596
rect 2320 9580 2372 9586
rect 2320 9522 2372 9528
rect 2228 9444 2280 9450
rect 2228 9386 2280 9392
rect 2872 9104 2924 9110
rect 2872 9046 2924 9052
rect 2780 8832 2832 8838
rect 2780 8774 2832 8780
rect 2136 8492 2188 8498
rect 2136 8434 2188 8440
rect 2044 8084 2096 8090
rect 2044 8026 2096 8032
rect 2792 8022 2820 8774
rect 2884 8294 2912 9046
rect 2872 8288 2924 8294
rect 2872 8230 2924 8236
rect 2780 8016 2832 8022
rect 2780 7958 2832 7964
rect 2792 7546 2820 7958
rect 2780 7540 2832 7546
rect 2780 7482 2832 7488
rect 1952 7404 2004 7410
rect 1952 7346 2004 7352
rect 2792 7342 2820 7482
rect 2780 7336 2832 7342
rect 2780 7278 2832 7284
rect 1860 6928 1912 6934
rect 1860 6870 1912 6876
rect 2596 6860 2648 6866
rect 2780 6860 2832 6866
rect 2648 6820 2728 6848
rect 2596 6802 2648 6808
rect 2700 6186 2728 6820
rect 2780 6802 2832 6808
rect 2688 6180 2740 6186
rect 2688 6122 2740 6128
rect 2044 5228 2096 5234
rect 2044 5170 2096 5176
rect 2056 5030 2084 5170
rect 2700 5166 2728 6122
rect 2792 6118 2820 6802
rect 2780 6112 2832 6118
rect 2780 6054 2832 6060
rect 2792 5778 2820 6054
rect 2780 5772 2832 5778
rect 2780 5714 2832 5720
rect 2688 5160 2740 5166
rect 2688 5102 2740 5108
rect 2044 5024 2096 5030
rect 2044 4966 2096 4972
rect 1768 3732 1820 3738
rect 1768 3674 1820 3680
rect 2056 2281 2084 4966
rect 2700 4758 2728 5102
rect 2792 5030 2820 5714
rect 2780 5024 2832 5030
rect 2780 4966 2832 4972
rect 2688 4752 2740 4758
rect 2688 4694 2740 4700
rect 2792 4486 2820 4966
rect 2884 4554 2912 8230
rect 2976 8022 3004 9590
rect 3252 8634 3280 10066
rect 3436 9110 3464 11086
rect 3896 10674 3924 11716
rect 3988 11694 4016 12378
rect 3976 11688 4028 11694
rect 3976 11630 4028 11636
rect 3988 11354 4016 11630
rect 4080 11558 4108 14214
rect 4172 13297 4200 18566
rect 4356 18290 4384 19110
rect 4712 18828 4764 18834
rect 4712 18770 4764 18776
rect 4344 18284 4396 18290
rect 4344 18226 4396 18232
rect 4724 18086 4752 18770
rect 4816 18630 4844 27520
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 6012 19854 6040 27526
rect 6182 27520 6238 27526
rect 7484 27526 7710 27554
rect 7484 24410 7512 27526
rect 7654 27520 7710 27526
rect 9034 27520 9090 28000
rect 10414 27554 10470 28000
rect 11794 27554 11850 28000
rect 9968 27526 10470 27554
rect 7472 24404 7524 24410
rect 7472 24346 7524 24352
rect 7288 24268 7340 24274
rect 7288 24210 7340 24216
rect 7300 23526 7328 24210
rect 9048 23866 9076 27520
rect 9036 23860 9088 23866
rect 9036 23802 9088 23808
rect 7840 23656 7892 23662
rect 7840 23598 7892 23604
rect 7288 23520 7340 23526
rect 7288 23462 7340 23468
rect 7748 23520 7800 23526
rect 7748 23462 7800 23468
rect 7656 20800 7708 20806
rect 7656 20742 7708 20748
rect 6274 20496 6330 20505
rect 6274 20431 6330 20440
rect 6288 19922 6316 20431
rect 6368 20392 6420 20398
rect 6368 20334 6420 20340
rect 6276 19916 6328 19922
rect 6276 19858 6328 19864
rect 5448 19848 5500 19854
rect 5448 19790 5500 19796
rect 6000 19848 6052 19854
rect 6000 19790 6052 19796
rect 5356 19780 5408 19786
rect 5356 19722 5408 19728
rect 5080 19712 5132 19718
rect 5080 19654 5132 19660
rect 5092 19378 5120 19654
rect 5368 19378 5396 19722
rect 5080 19372 5132 19378
rect 5080 19314 5132 19320
rect 5356 19372 5408 19378
rect 5356 19314 5408 19320
rect 5092 18970 5120 19314
rect 5172 19236 5224 19242
rect 5172 19178 5224 19184
rect 5080 18964 5132 18970
rect 5080 18906 5132 18912
rect 4804 18624 4856 18630
rect 4804 18566 4856 18572
rect 5080 18624 5132 18630
rect 5184 18612 5212 19178
rect 5264 18692 5316 18698
rect 5264 18634 5316 18640
rect 5132 18584 5212 18612
rect 5080 18566 5132 18572
rect 4988 18216 5040 18222
rect 5092 18204 5120 18566
rect 5276 18290 5304 18634
rect 5264 18284 5316 18290
rect 5264 18226 5316 18232
rect 5040 18176 5120 18204
rect 4988 18158 5040 18164
rect 4712 18080 4764 18086
rect 4712 18022 4764 18028
rect 4804 17876 4856 17882
rect 4804 17818 4856 17824
rect 4252 17672 4304 17678
rect 4252 17614 4304 17620
rect 4264 16998 4292 17614
rect 4620 17128 4672 17134
rect 4620 17070 4672 17076
rect 4252 16992 4304 16998
rect 4252 16934 4304 16940
rect 4158 13288 4214 13297
rect 4158 13223 4214 13232
rect 4264 12646 4292 16934
rect 4436 16584 4488 16590
rect 4436 16526 4488 16532
rect 4448 16250 4476 16526
rect 4632 16454 4660 17070
rect 4816 16998 4844 17818
rect 5092 17610 5120 18176
rect 5356 18148 5408 18154
rect 5356 18090 5408 18096
rect 5368 17814 5396 18090
rect 5356 17808 5408 17814
rect 5356 17750 5408 17756
rect 5080 17604 5132 17610
rect 5080 17546 5132 17552
rect 4804 16992 4856 16998
rect 4804 16934 4856 16940
rect 5080 16992 5132 16998
rect 5080 16934 5132 16940
rect 5092 16794 5120 16934
rect 5080 16788 5132 16794
rect 5080 16730 5132 16736
rect 5172 16720 5224 16726
rect 5172 16662 5224 16668
rect 4620 16448 4672 16454
rect 4620 16390 4672 16396
rect 4436 16244 4488 16250
rect 4436 16186 4488 16192
rect 4436 15632 4488 15638
rect 4436 15574 4488 15580
rect 4344 15360 4396 15366
rect 4344 15302 4396 15308
rect 4356 14074 4384 15302
rect 4448 15162 4476 15574
rect 4436 15156 4488 15162
rect 4436 15098 4488 15104
rect 4528 14884 4580 14890
rect 4528 14826 4580 14832
rect 4436 14544 4488 14550
rect 4436 14486 4488 14492
rect 4448 14074 4476 14486
rect 4344 14068 4396 14074
rect 4344 14010 4396 14016
rect 4436 14068 4488 14074
rect 4436 14010 4488 14016
rect 4540 13802 4568 14826
rect 4528 13796 4580 13802
rect 4528 13738 4580 13744
rect 4528 13524 4580 13530
rect 4528 13466 4580 13472
rect 4540 12782 4568 13466
rect 4528 12776 4580 12782
rect 4528 12718 4580 12724
rect 4344 12708 4396 12714
rect 4344 12650 4396 12656
rect 4252 12640 4304 12646
rect 4252 12582 4304 12588
rect 4356 12306 4384 12650
rect 4540 12306 4568 12718
rect 4632 12442 4660 16390
rect 5184 16250 5212 16662
rect 5172 16244 5224 16250
rect 5172 16186 5224 16192
rect 4988 16108 5040 16114
rect 4988 16050 5040 16056
rect 5000 15638 5028 16050
rect 5264 15972 5316 15978
rect 5264 15914 5316 15920
rect 5276 15706 5304 15914
rect 5264 15700 5316 15706
rect 5264 15642 5316 15648
rect 4988 15632 5040 15638
rect 4988 15574 5040 15580
rect 4804 15156 4856 15162
rect 4804 15098 4856 15104
rect 4816 13462 4844 15098
rect 5000 14550 5028 15574
rect 5276 15094 5304 15642
rect 5264 15088 5316 15094
rect 5264 15030 5316 15036
rect 4988 14544 5040 14550
rect 5460 14521 5488 19790
rect 6000 19712 6052 19718
rect 6000 19654 6052 19660
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5540 18964 5592 18970
rect 5540 18906 5592 18912
rect 5552 18290 5580 18906
rect 6012 18766 6040 19654
rect 6288 19514 6316 19858
rect 6276 19508 6328 19514
rect 6276 19450 6328 19456
rect 6092 18896 6144 18902
rect 6092 18838 6144 18844
rect 6000 18760 6052 18766
rect 6000 18702 6052 18708
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5540 18284 5592 18290
rect 5540 18226 5592 18232
rect 6012 17882 6040 18702
rect 6104 18426 6132 18838
rect 6092 18420 6144 18426
rect 6092 18362 6144 18368
rect 6000 17876 6052 17882
rect 6000 17818 6052 17824
rect 6104 17746 6132 18362
rect 6092 17740 6144 17746
rect 6092 17682 6144 17688
rect 5540 17672 5592 17678
rect 5540 17614 5592 17620
rect 5552 17338 5580 17614
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 6104 17338 6132 17682
rect 5540 17332 5592 17338
rect 5540 17274 5592 17280
rect 6092 17332 6144 17338
rect 6092 17274 6144 17280
rect 5540 16584 5592 16590
rect 5540 16526 5592 16532
rect 5552 16182 5580 16526
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5540 16176 5592 16182
rect 5540 16118 5592 16124
rect 5552 16017 5580 16118
rect 5538 16008 5594 16017
rect 5538 15943 5594 15952
rect 6276 15632 6328 15638
rect 6196 15592 6276 15620
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 6196 14822 6224 15592
rect 6276 15574 6328 15580
rect 6184 14816 6236 14822
rect 6184 14758 6236 14764
rect 4988 14486 5040 14492
rect 5446 14512 5502 14521
rect 5446 14447 5502 14456
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5080 14068 5132 14074
rect 5080 14010 5132 14016
rect 4988 14000 5040 14006
rect 4988 13942 5040 13948
rect 4804 13456 4856 13462
rect 4804 13398 4856 13404
rect 4620 12436 4672 12442
rect 4620 12378 4672 12384
rect 4344 12300 4396 12306
rect 4344 12242 4396 12248
rect 4528 12300 4580 12306
rect 4528 12242 4580 12248
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 4068 11552 4120 11558
rect 4068 11494 4120 11500
rect 3976 11348 4028 11354
rect 3976 11290 4028 11296
rect 3884 10668 3936 10674
rect 3884 10610 3936 10616
rect 3896 9586 3924 10610
rect 3988 10130 4016 11290
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 3976 10124 4028 10130
rect 3976 10066 4028 10072
rect 3884 9580 3936 9586
rect 3884 9522 3936 9528
rect 3792 9512 3844 9518
rect 3792 9454 3844 9460
rect 3804 9178 3832 9454
rect 3976 9376 4028 9382
rect 3976 9318 4028 9324
rect 3792 9172 3844 9178
rect 3792 9114 3844 9120
rect 3424 9104 3476 9110
rect 3424 9046 3476 9052
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 2964 8016 3016 8022
rect 2964 7958 3016 7964
rect 2976 6934 3004 7958
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 3160 7206 3188 7822
rect 3436 7818 3464 9046
rect 3988 9042 4016 9318
rect 3976 9036 4028 9042
rect 3976 8978 4028 8984
rect 3516 8900 3568 8906
rect 3516 8842 3568 8848
rect 3528 8090 3556 8842
rect 3792 8628 3844 8634
rect 3792 8570 3844 8576
rect 3804 8090 3832 8570
rect 3976 8288 4028 8294
rect 3976 8230 4028 8236
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 3792 8084 3844 8090
rect 3792 8026 3844 8032
rect 3424 7812 3476 7818
rect 3424 7754 3476 7760
rect 3516 7540 3568 7546
rect 3516 7482 3568 7488
rect 3528 7206 3556 7482
rect 3988 7410 4016 8230
rect 4080 7993 4108 10406
rect 4172 10062 4200 11834
rect 4356 11830 4384 12242
rect 4344 11824 4396 11830
rect 4344 11766 4396 11772
rect 4540 11694 4568 12242
rect 4528 11688 4580 11694
rect 4528 11630 4580 11636
rect 4436 11620 4488 11626
rect 4436 11562 4488 11568
rect 4344 10124 4396 10130
rect 4344 10066 4396 10072
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 4172 9654 4200 9998
rect 4160 9648 4212 9654
rect 4160 9590 4212 9596
rect 4172 9450 4200 9590
rect 4356 9450 4384 10066
rect 4448 9994 4476 11562
rect 4540 11218 4568 11630
rect 4896 11620 4948 11626
rect 4896 11562 4948 11568
rect 4908 11218 4936 11562
rect 4528 11212 4580 11218
rect 4528 11154 4580 11160
rect 4896 11212 4948 11218
rect 4896 11154 4948 11160
rect 4540 10266 4568 11154
rect 5000 10810 5028 13942
rect 5092 13530 5120 14010
rect 5448 13728 5500 13734
rect 5448 13670 5500 13676
rect 5080 13524 5132 13530
rect 5080 13466 5132 13472
rect 5356 13184 5408 13190
rect 5356 13126 5408 13132
rect 5368 12782 5396 13126
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 5368 11694 5396 12718
rect 5356 11688 5408 11694
rect 5356 11630 5408 11636
rect 4988 10804 5040 10810
rect 4988 10746 5040 10752
rect 5368 10742 5396 11630
rect 5460 11354 5488 13670
rect 6196 13462 6224 14758
rect 6276 14272 6328 14278
rect 6276 14214 6328 14220
rect 6288 13938 6316 14214
rect 6276 13932 6328 13938
rect 6276 13874 6328 13880
rect 6380 13814 6408 20334
rect 7668 20058 7696 20742
rect 7656 20052 7708 20058
rect 7656 19994 7708 20000
rect 7196 19304 7248 19310
rect 7196 19246 7248 19252
rect 7472 19304 7524 19310
rect 7472 19246 7524 19252
rect 7012 18080 7064 18086
rect 7012 18022 7064 18028
rect 6828 16992 6880 16998
rect 6828 16934 6880 16940
rect 6644 14884 6696 14890
rect 6644 14826 6696 14832
rect 6460 14068 6512 14074
rect 6460 14010 6512 14016
rect 6288 13786 6408 13814
rect 6184 13456 6236 13462
rect 6184 13398 6236 13404
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 6000 12640 6052 12646
rect 6000 12582 6052 12588
rect 6012 12374 6040 12582
rect 6000 12368 6052 12374
rect 6000 12310 6052 12316
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 6012 11898 6040 12310
rect 6184 12300 6236 12306
rect 6184 12242 6236 12248
rect 6092 12096 6144 12102
rect 6092 12038 6144 12044
rect 6000 11892 6052 11898
rect 6000 11834 6052 11840
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5356 10736 5408 10742
rect 5356 10678 5408 10684
rect 5172 10600 5224 10606
rect 5172 10542 5224 10548
rect 5184 10470 5212 10542
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 4528 10260 4580 10266
rect 4528 10202 4580 10208
rect 5184 10130 5212 10406
rect 5368 10130 5396 10678
rect 4620 10124 4672 10130
rect 4620 10066 4672 10072
rect 5172 10124 5224 10130
rect 5172 10066 5224 10072
rect 5356 10124 5408 10130
rect 5408 10084 5488 10112
rect 5356 10066 5408 10072
rect 4436 9988 4488 9994
rect 4436 9930 4488 9936
rect 4160 9444 4212 9450
rect 4160 9386 4212 9392
rect 4344 9444 4396 9450
rect 4344 9386 4396 9392
rect 4252 9104 4304 9110
rect 4448 9058 4476 9930
rect 4528 9580 4580 9586
rect 4528 9522 4580 9528
rect 4252 9046 4304 9052
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 4066 7984 4122 7993
rect 4066 7919 4122 7928
rect 4068 7812 4120 7818
rect 4068 7754 4120 7760
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 3148 7200 3200 7206
rect 3148 7142 3200 7148
rect 3516 7200 3568 7206
rect 3516 7142 3568 7148
rect 2964 6928 3016 6934
rect 2964 6870 3016 6876
rect 3160 5817 3188 7142
rect 3528 7002 3556 7142
rect 4080 7002 4108 7754
rect 4172 7546 4200 8910
rect 4264 8294 4292 9046
rect 4356 9030 4476 9058
rect 4356 8906 4384 9030
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 4344 8900 4396 8906
rect 4344 8842 4396 8848
rect 4252 8288 4304 8294
rect 4252 8230 4304 8236
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 4356 7478 4384 8842
rect 4448 8022 4476 8910
rect 4436 8016 4488 8022
rect 4436 7958 4488 7964
rect 4344 7472 4396 7478
rect 4344 7414 4396 7420
rect 3516 6996 3568 7002
rect 3516 6938 3568 6944
rect 4068 6996 4120 7002
rect 4068 6938 4120 6944
rect 4540 6866 4568 9522
rect 4632 9518 4660 10066
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 4632 8838 4660 9454
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 4712 8424 4764 8430
rect 4712 8366 4764 8372
rect 4724 7954 4752 8366
rect 5092 8362 5120 8774
rect 5172 8424 5224 8430
rect 5172 8366 5224 8372
rect 5080 8356 5132 8362
rect 5080 8298 5132 8304
rect 4712 7948 4764 7954
rect 4712 7890 4764 7896
rect 5184 7886 5212 8366
rect 5276 7954 5304 9318
rect 5368 9110 5396 9454
rect 5356 9104 5408 9110
rect 5356 9046 5408 9052
rect 5368 8634 5396 9046
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 5368 8430 5396 8570
rect 5356 8424 5408 8430
rect 5356 8366 5408 8372
rect 5460 8022 5488 10084
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 6104 9674 6132 12038
rect 6196 11626 6224 12242
rect 6184 11620 6236 11626
rect 6184 11562 6236 11568
rect 6196 11218 6224 11562
rect 6184 11212 6236 11218
rect 6184 11154 6236 11160
rect 6288 10033 6316 13786
rect 6368 13728 6420 13734
rect 6368 13670 6420 13676
rect 6380 12374 6408 13670
rect 6472 13394 6500 14010
rect 6656 14006 6684 14826
rect 6840 14550 6868 16934
rect 6920 15020 6972 15026
rect 6920 14962 6972 14968
rect 6828 14544 6880 14550
rect 6828 14486 6880 14492
rect 6644 14000 6696 14006
rect 6644 13942 6696 13948
rect 6656 13802 6684 13942
rect 6736 13932 6788 13938
rect 6736 13874 6788 13880
rect 6644 13796 6696 13802
rect 6644 13738 6696 13744
rect 6460 13388 6512 13394
rect 6460 13330 6512 13336
rect 6472 12442 6500 13330
rect 6460 12436 6512 12442
rect 6460 12378 6512 12384
rect 6368 12368 6420 12374
rect 6368 12310 6420 12316
rect 6552 10464 6604 10470
rect 6552 10406 6604 10412
rect 6274 10024 6330 10033
rect 6274 9959 6330 9968
rect 6012 9646 6132 9674
rect 6012 9042 6040 9646
rect 6000 9036 6052 9042
rect 6000 8978 6052 8984
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 6012 8634 6040 8978
rect 6092 8968 6144 8974
rect 6092 8910 6144 8916
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 5448 8016 5500 8022
rect 5448 7958 5500 7964
rect 5264 7948 5316 7954
rect 5264 7890 5316 7896
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 4632 7546 4660 7822
rect 5276 7546 5304 7890
rect 5460 7818 5488 7958
rect 5448 7812 5500 7818
rect 5448 7754 5500 7760
rect 4620 7540 4672 7546
rect 4620 7482 4672 7488
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 5356 7336 5408 7342
rect 5356 7278 5408 7284
rect 4724 6934 4752 7278
rect 5080 7268 5132 7274
rect 5080 7210 5132 7216
rect 4712 6928 4764 6934
rect 4712 6870 4764 6876
rect 4528 6860 4580 6866
rect 4528 6802 4580 6808
rect 3240 6656 3292 6662
rect 3240 6598 3292 6604
rect 3252 6254 3280 6598
rect 4540 6390 4568 6802
rect 4620 6656 4672 6662
rect 4620 6598 4672 6604
rect 3332 6384 3384 6390
rect 3332 6326 3384 6332
rect 4528 6384 4580 6390
rect 4528 6326 4580 6332
rect 3240 6248 3292 6254
rect 3240 6190 3292 6196
rect 3252 5846 3280 6190
rect 3240 5840 3292 5846
rect 3146 5808 3202 5817
rect 3240 5782 3292 5788
rect 3146 5743 3202 5752
rect 2872 4548 2924 4554
rect 2872 4490 2924 4496
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 2042 2272 2098 2281
rect 2042 2207 2098 2216
rect 2792 921 2820 4422
rect 3344 4154 3372 6326
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 3436 5914 3464 6258
rect 4632 6254 4660 6598
rect 5092 6322 5120 7210
rect 5080 6316 5132 6322
rect 5080 6258 5132 6264
rect 4620 6248 4672 6254
rect 4620 6190 4672 6196
rect 4896 6248 4948 6254
rect 4896 6190 4948 6196
rect 3792 6180 3844 6186
rect 3792 6122 3844 6128
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 3804 5166 3832 6122
rect 4160 6112 4212 6118
rect 4160 6054 4212 6060
rect 4172 5778 4200 6054
rect 4908 5914 4936 6190
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 4172 5234 4200 5714
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 3792 5160 3844 5166
rect 3792 5102 3844 5108
rect 5368 5098 5396 7278
rect 5460 5914 5488 7754
rect 5552 6934 5580 8570
rect 6000 8288 6052 8294
rect 6000 8230 6052 8236
rect 6012 7954 6040 8230
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5540 6928 5592 6934
rect 5540 6870 5592 6876
rect 6012 6662 6040 7890
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 6000 6656 6052 6662
rect 6000 6598 6052 6604
rect 5448 5908 5500 5914
rect 5448 5850 5500 5856
rect 5446 5672 5502 5681
rect 5446 5607 5502 5616
rect 5356 5092 5408 5098
rect 5356 5034 5408 5040
rect 5460 4690 5488 5607
rect 5552 5370 5580 6598
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 6000 6452 6052 6458
rect 6000 6394 6052 6400
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5540 5364 5592 5370
rect 5540 5306 5592 5312
rect 6012 5302 6040 6394
rect 6000 5296 6052 5302
rect 6000 5238 6052 5244
rect 5448 4684 5500 4690
rect 5448 4626 5500 4632
rect 5460 4282 5488 4626
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5448 4276 5500 4282
rect 5448 4218 5500 4224
rect 3252 4126 3372 4154
rect 2778 912 2834 921
rect 2778 847 2834 856
rect 1766 82 1822 480
rect 1688 54 1822 82
rect 570 0 626 54
rect 1766 0 1822 54
rect 3054 82 3110 480
rect 3252 82 3280 4126
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 4712 2372 4764 2378
rect 4712 2314 4764 2320
rect 3054 54 3280 82
rect 4342 82 4398 480
rect 4724 82 4752 2314
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 4342 54 4752 82
rect 5630 82 5686 480
rect 6104 82 6132 8910
rect 6564 8888 6592 10406
rect 6748 9382 6776 13874
rect 6840 13530 6868 14486
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 6828 12912 6880 12918
rect 6828 12854 6880 12860
rect 6840 12442 6868 12854
rect 6828 12436 6880 12442
rect 6828 12378 6880 12384
rect 6840 11354 6868 12378
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6932 10266 6960 14962
rect 7024 14906 7052 18022
rect 7208 17785 7236 19246
rect 7484 18970 7512 19246
rect 7656 19236 7708 19242
rect 7656 19178 7708 19184
rect 7472 18964 7524 18970
rect 7472 18906 7524 18912
rect 7564 18760 7616 18766
rect 7564 18702 7616 18708
rect 7380 18692 7432 18698
rect 7380 18634 7432 18640
rect 7392 18290 7420 18634
rect 7380 18284 7432 18290
rect 7380 18226 7432 18232
rect 7194 17776 7250 17785
rect 7194 17711 7250 17720
rect 7576 17678 7604 18702
rect 7564 17672 7616 17678
rect 7564 17614 7616 17620
rect 7668 17202 7696 19178
rect 7104 17196 7156 17202
rect 7104 17138 7156 17144
rect 7656 17196 7708 17202
rect 7656 17138 7708 17144
rect 7116 16250 7144 17138
rect 7380 16992 7432 16998
rect 7380 16934 7432 16940
rect 7288 16652 7340 16658
rect 7288 16594 7340 16600
rect 7104 16244 7156 16250
rect 7104 16186 7156 16192
rect 7300 15706 7328 16594
rect 7288 15700 7340 15706
rect 7288 15642 7340 15648
rect 7392 15609 7420 16934
rect 7668 16726 7696 17138
rect 7656 16720 7708 16726
rect 7656 16662 7708 16668
rect 7472 16448 7524 16454
rect 7472 16390 7524 16396
rect 7484 16250 7512 16390
rect 7472 16244 7524 16250
rect 7472 16186 7524 16192
rect 7484 15910 7512 16186
rect 7472 15904 7524 15910
rect 7472 15846 7524 15852
rect 7378 15600 7434 15609
rect 7378 15535 7434 15544
rect 7472 15496 7524 15502
rect 7472 15438 7524 15444
rect 7484 15094 7512 15438
rect 7564 15360 7616 15366
rect 7564 15302 7616 15308
rect 7472 15088 7524 15094
rect 7472 15030 7524 15036
rect 7102 14920 7158 14929
rect 7024 14878 7102 14906
rect 7102 14855 7158 14864
rect 7012 14544 7064 14550
rect 7012 14486 7064 14492
rect 7024 14074 7052 14486
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 7116 13814 7144 14855
rect 7484 14550 7512 15030
rect 7576 15026 7604 15302
rect 7564 15020 7616 15026
rect 7564 14962 7616 14968
rect 7472 14544 7524 14550
rect 7472 14486 7524 14492
rect 7024 13786 7144 13814
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 6736 9376 6788 9382
rect 6736 9318 6788 9324
rect 7024 8974 7052 13786
rect 7656 13184 7708 13190
rect 7656 13126 7708 13132
rect 7668 12782 7696 13126
rect 7656 12776 7708 12782
rect 7656 12718 7708 12724
rect 7196 12640 7248 12646
rect 7196 12582 7248 12588
rect 7208 11694 7236 12582
rect 7288 12368 7340 12374
rect 7288 12310 7340 12316
rect 7300 11762 7328 12310
rect 7668 12306 7696 12718
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 7656 12300 7708 12306
rect 7656 12242 7708 12248
rect 7392 11898 7420 12242
rect 7380 11892 7432 11898
rect 7380 11834 7432 11840
rect 7288 11756 7340 11762
rect 7288 11698 7340 11704
rect 7196 11688 7248 11694
rect 7196 11630 7248 11636
rect 7208 10198 7236 11630
rect 7196 10192 7248 10198
rect 7196 10134 7248 10140
rect 7196 10056 7248 10062
rect 7196 9998 7248 10004
rect 7208 9518 7236 9998
rect 7196 9512 7248 9518
rect 7196 9454 7248 9460
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 7012 8968 7064 8974
rect 7012 8910 7064 8916
rect 6644 8900 6696 8906
rect 6564 8860 6644 8888
rect 6564 8634 6592 8860
rect 6644 8842 6696 8848
rect 7116 8634 7144 9318
rect 7208 9042 7236 9454
rect 7300 9178 7328 11698
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 7656 11688 7708 11694
rect 7656 11630 7708 11636
rect 7392 11218 7420 11630
rect 7668 11529 7696 11630
rect 7654 11520 7710 11529
rect 7654 11455 7710 11464
rect 7380 11212 7432 11218
rect 7380 11154 7432 11160
rect 7656 11212 7708 11218
rect 7656 11154 7708 11160
rect 7392 10810 7420 11154
rect 7380 10804 7432 10810
rect 7380 10746 7432 10752
rect 7392 10606 7420 10746
rect 7668 10606 7696 11154
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 7656 10600 7708 10606
rect 7656 10542 7708 10548
rect 7656 10124 7708 10130
rect 7656 10066 7708 10072
rect 7380 9920 7432 9926
rect 7380 9862 7432 9868
rect 7392 9518 7420 9862
rect 7668 9518 7696 10066
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 7656 9512 7708 9518
rect 7760 9489 7788 23462
rect 7852 20466 7880 23598
rect 8484 23180 8536 23186
rect 8484 23122 8536 23128
rect 8496 22438 8524 23122
rect 8484 22432 8536 22438
rect 8484 22374 8536 22380
rect 8300 20936 8352 20942
rect 8300 20878 8352 20884
rect 7840 20460 7892 20466
rect 7840 20402 7892 20408
rect 7840 20052 7892 20058
rect 7840 19994 7892 20000
rect 7852 19310 7880 19994
rect 8116 19984 8168 19990
rect 8116 19926 8168 19932
rect 7840 19304 7892 19310
rect 7840 19246 7892 19252
rect 8128 19174 8156 19926
rect 8312 19514 8340 20878
rect 8300 19508 8352 19514
rect 8300 19450 8352 19456
rect 8116 19168 8168 19174
rect 8116 19110 8168 19116
rect 8128 18970 8156 19110
rect 8116 18964 8168 18970
rect 8116 18906 8168 18912
rect 7840 18760 7892 18766
rect 7840 18702 7892 18708
rect 7852 18290 7880 18702
rect 8128 18426 8156 18906
rect 8116 18420 8168 18426
rect 8116 18362 8168 18368
rect 7932 18352 7984 18358
rect 7932 18294 7984 18300
rect 7840 18284 7892 18290
rect 7840 18226 7892 18232
rect 7852 17678 7880 18226
rect 7840 17672 7892 17678
rect 7840 17614 7892 17620
rect 7852 17338 7880 17614
rect 7840 17332 7892 17338
rect 7840 17274 7892 17280
rect 7944 16153 7972 18294
rect 8208 17808 8260 17814
rect 8208 17750 8260 17756
rect 8220 17270 8248 17750
rect 8208 17264 8260 17270
rect 8208 17206 8260 17212
rect 8024 17060 8076 17066
rect 8024 17002 8076 17008
rect 8036 16794 8064 17002
rect 8220 16794 8248 17206
rect 8024 16788 8076 16794
rect 8024 16730 8076 16736
rect 8208 16788 8260 16794
rect 8208 16730 8260 16736
rect 7930 16144 7986 16153
rect 7930 16079 7986 16088
rect 7840 15700 7892 15706
rect 7840 15642 7892 15648
rect 7852 15162 7880 15642
rect 7840 15156 7892 15162
rect 7840 15098 7892 15104
rect 7944 14482 7972 16079
rect 8036 14890 8064 16730
rect 8114 16144 8170 16153
rect 8114 16079 8170 16088
rect 8024 14884 8076 14890
rect 8024 14826 8076 14832
rect 7932 14476 7984 14482
rect 7932 14418 7984 14424
rect 8036 14006 8064 14826
rect 8024 14000 8076 14006
rect 8024 13942 8076 13948
rect 8024 13252 8076 13258
rect 8024 13194 8076 13200
rect 7932 12844 7984 12850
rect 7932 12786 7984 12792
rect 7944 12753 7972 12786
rect 7930 12744 7986 12753
rect 7930 12679 7986 12688
rect 8036 11762 8064 13194
rect 8128 12850 8156 16079
rect 8496 15978 8524 22374
rect 9588 21004 9640 21010
rect 9588 20946 9640 20952
rect 8852 20800 8904 20806
rect 8852 20742 8904 20748
rect 8864 20398 8892 20742
rect 8852 20392 8904 20398
rect 8852 20334 8904 20340
rect 8864 20058 8892 20334
rect 9600 20262 9628 20946
rect 9772 20324 9824 20330
rect 9772 20266 9824 20272
rect 8944 20256 8996 20262
rect 8944 20198 8996 20204
rect 9588 20256 9640 20262
rect 9588 20198 9640 20204
rect 8852 20052 8904 20058
rect 8852 19994 8904 20000
rect 8852 19848 8904 19854
rect 8852 19790 8904 19796
rect 8864 19378 8892 19790
rect 8852 19372 8904 19378
rect 8852 19314 8904 19320
rect 8576 19236 8628 19242
rect 8576 19178 8628 19184
rect 8588 18970 8616 19178
rect 8576 18964 8628 18970
rect 8576 18906 8628 18912
rect 8588 18154 8616 18906
rect 8864 18698 8892 19314
rect 8956 18970 8984 20198
rect 8944 18964 8996 18970
rect 8944 18906 8996 18912
rect 8852 18692 8904 18698
rect 8852 18634 8904 18640
rect 8956 18290 8984 18906
rect 8944 18284 8996 18290
rect 8944 18226 8996 18232
rect 9600 18193 9628 20198
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 9692 18358 9720 18770
rect 9680 18352 9732 18358
rect 9680 18294 9732 18300
rect 9586 18184 9642 18193
rect 8576 18148 8628 18154
rect 8576 18090 8628 18096
rect 8760 18148 8812 18154
rect 9586 18119 9642 18128
rect 8760 18090 8812 18096
rect 8576 17128 8628 17134
rect 8576 17070 8628 17076
rect 8484 15972 8536 15978
rect 8484 15914 8536 15920
rect 8496 15638 8524 15914
rect 8484 15632 8536 15638
rect 8484 15574 8536 15580
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 8312 14074 8340 14418
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 8588 13814 8616 17070
rect 8772 17066 8800 18090
rect 8760 17060 8812 17066
rect 8760 17002 8812 17008
rect 9600 16658 9628 18119
rect 9784 17678 9812 20266
rect 9864 18420 9916 18426
rect 9864 18362 9916 18368
rect 9876 17814 9904 18362
rect 9864 17808 9916 17814
rect 9864 17750 9916 17756
rect 9772 17672 9824 17678
rect 9772 17614 9824 17620
rect 9784 17270 9812 17614
rect 9772 17264 9824 17270
rect 9772 17206 9824 17212
rect 9588 16652 9640 16658
rect 9588 16594 9640 16600
rect 9312 16516 9364 16522
rect 9312 16458 9364 16464
rect 9324 16114 9352 16458
rect 9600 16250 9628 16594
rect 9588 16244 9640 16250
rect 9588 16186 9640 16192
rect 9312 16108 9364 16114
rect 9232 16068 9312 16096
rect 9232 15706 9260 16068
rect 9312 16050 9364 16056
rect 9404 15972 9456 15978
rect 9324 15932 9404 15960
rect 9220 15700 9272 15706
rect 9220 15642 9272 15648
rect 9324 14822 9352 15932
rect 9404 15914 9456 15920
rect 9496 14884 9548 14890
rect 9496 14826 9548 14832
rect 9312 14816 9364 14822
rect 9312 14758 9364 14764
rect 8944 13864 8996 13870
rect 8496 13786 8616 13814
rect 8942 13832 8944 13841
rect 8996 13832 8998 13841
rect 8300 13388 8352 13394
rect 8300 13330 8352 13336
rect 8116 12844 8168 12850
rect 8116 12786 8168 12792
rect 8312 12646 8340 13330
rect 8300 12640 8352 12646
rect 8300 12582 8352 12588
rect 8496 12374 8524 13786
rect 8942 13767 8998 13776
rect 8852 13388 8904 13394
rect 8852 13330 8904 13336
rect 8864 12986 8892 13330
rect 8852 12980 8904 12986
rect 8852 12922 8904 12928
rect 8864 12889 8892 12922
rect 8850 12880 8906 12889
rect 8850 12815 8906 12824
rect 8484 12368 8536 12374
rect 8484 12310 8536 12316
rect 8576 12164 8628 12170
rect 8576 12106 8628 12112
rect 8588 11898 8616 12106
rect 8576 11892 8628 11898
rect 8576 11834 8628 11840
rect 8024 11756 8076 11762
rect 8024 11698 8076 11704
rect 8576 11756 8628 11762
rect 8576 11698 8628 11704
rect 8300 11620 8352 11626
rect 8300 11562 8352 11568
rect 8484 11620 8536 11626
rect 8484 11562 8536 11568
rect 8312 11218 8340 11562
rect 8300 11212 8352 11218
rect 8300 11154 8352 11160
rect 8208 11008 8260 11014
rect 8208 10950 8260 10956
rect 8220 10606 8248 10950
rect 8208 10600 8260 10606
rect 8208 10542 8260 10548
rect 7932 10124 7984 10130
rect 7932 10066 7984 10072
rect 7944 9654 7972 10066
rect 8220 9926 8248 10542
rect 8208 9920 8260 9926
rect 8208 9862 8260 9868
rect 7932 9648 7984 9654
rect 7932 9590 7984 9596
rect 7656 9454 7708 9460
rect 7746 9480 7802 9489
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7392 9042 7420 9454
rect 7746 9415 7802 9424
rect 7196 9036 7248 9042
rect 7196 8978 7248 8984
rect 7380 9036 7432 9042
rect 7380 8978 7432 8984
rect 7208 8838 7236 8978
rect 7196 8832 7248 8838
rect 7196 8774 7248 8780
rect 6552 8628 6604 8634
rect 6552 8570 6604 8576
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 6368 7744 6420 7750
rect 6368 7686 6420 7692
rect 6380 7206 6408 7686
rect 6368 7200 6420 7206
rect 6368 7142 6420 7148
rect 6276 6180 6328 6186
rect 6276 6122 6328 6128
rect 6288 5778 6316 6122
rect 6276 5772 6328 5778
rect 6276 5714 6328 5720
rect 6288 5302 6316 5714
rect 6380 5370 6408 7142
rect 6472 6390 6500 7822
rect 6564 7546 6592 8570
rect 7392 7886 7420 8978
rect 7564 8832 7616 8838
rect 7564 8774 7616 8780
rect 7576 8430 7604 8774
rect 7564 8424 7616 8430
rect 7564 8366 7616 8372
rect 7576 7954 7604 8366
rect 7564 7948 7616 7954
rect 7564 7890 7616 7896
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 7576 7342 7604 7890
rect 7760 7410 7788 9415
rect 7944 8294 7972 9590
rect 7932 8288 7984 8294
rect 7932 8230 7984 8236
rect 7840 7948 7892 7954
rect 7840 7890 7892 7896
rect 7852 7478 7880 7890
rect 7840 7472 7892 7478
rect 7840 7414 7892 7420
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 6644 6996 6696 7002
rect 6644 6938 6696 6944
rect 6552 6860 6604 6866
rect 6552 6802 6604 6808
rect 6564 6458 6592 6802
rect 6552 6452 6604 6458
rect 6552 6394 6604 6400
rect 6460 6384 6512 6390
rect 6460 6326 6512 6332
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 6276 5296 6328 5302
rect 6276 5238 6328 5244
rect 6564 5098 6592 5714
rect 6656 5234 6684 6938
rect 6736 6928 6788 6934
rect 6736 6870 6788 6876
rect 7748 6928 7800 6934
rect 7748 6870 7800 6876
rect 6748 6322 6776 6870
rect 7288 6860 7340 6866
rect 7288 6802 7340 6808
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 6748 5914 6776 6258
rect 7300 6118 7328 6802
rect 7760 6254 7788 6870
rect 7748 6248 7800 6254
rect 7748 6190 7800 6196
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 7576 5778 7604 6054
rect 7760 5914 7788 6190
rect 7944 6186 7972 8230
rect 8116 6792 8168 6798
rect 8220 6780 8248 9862
rect 8312 9042 8340 11154
rect 8496 10674 8524 11562
rect 8484 10668 8536 10674
rect 8484 10610 8536 10616
rect 8392 9172 8444 9178
rect 8392 9114 8444 9120
rect 8300 9036 8352 9042
rect 8300 8978 8352 8984
rect 8404 8430 8432 9114
rect 8588 8498 8616 11698
rect 8760 10600 8812 10606
rect 8760 10542 8812 10548
rect 8772 10266 8800 10542
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 8576 8492 8628 8498
rect 8576 8434 8628 8440
rect 8392 8424 8444 8430
rect 8392 8366 8444 8372
rect 8404 7342 8432 8366
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 8392 7336 8444 7342
rect 8392 7278 8444 7284
rect 8404 7002 8432 7278
rect 8864 7002 8892 7890
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8852 6996 8904 7002
rect 8852 6938 8904 6944
rect 8168 6752 8248 6780
rect 8116 6734 8168 6740
rect 8128 6254 8156 6734
rect 8666 6352 8722 6361
rect 8666 6287 8722 6296
rect 8680 6254 8708 6287
rect 8116 6248 8168 6254
rect 8116 6190 8168 6196
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 7932 6180 7984 6186
rect 7932 6122 7984 6128
rect 8024 6112 8076 6118
rect 8024 6054 8076 6060
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 8036 5846 8064 6054
rect 8024 5840 8076 5846
rect 8024 5782 8076 5788
rect 7564 5772 7616 5778
rect 7564 5714 7616 5720
rect 7196 5568 7248 5574
rect 7196 5510 7248 5516
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 6552 5092 6604 5098
rect 6552 5034 6604 5040
rect 6564 5001 6592 5034
rect 6550 4992 6606 5001
rect 6550 4927 6606 4936
rect 6564 4010 6592 4927
rect 6656 4826 6684 5170
rect 6828 5092 6880 5098
rect 6828 5034 6880 5040
rect 6644 4820 6696 4826
rect 6644 4762 6696 4768
rect 6840 4554 6868 5034
rect 7208 4758 7236 5510
rect 8036 5098 8064 5782
rect 8392 5772 8444 5778
rect 8392 5714 8444 5720
rect 8024 5092 8076 5098
rect 8024 5034 8076 5040
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 7760 4758 7788 4966
rect 7196 4752 7248 4758
rect 7196 4694 7248 4700
rect 7748 4752 7800 4758
rect 7748 4694 7800 4700
rect 6828 4548 6880 4554
rect 6828 4490 6880 4496
rect 6552 4004 6604 4010
rect 6552 3946 6604 3952
rect 7208 3738 7236 4694
rect 7760 4282 7788 4694
rect 7748 4276 7800 4282
rect 7748 4218 7800 4224
rect 7760 4078 7788 4218
rect 8312 4146 8340 4966
rect 8404 4826 8432 5714
rect 8668 5092 8720 5098
rect 8668 5034 8720 5040
rect 8392 4820 8444 4826
rect 8392 4762 8444 4768
rect 8680 4622 8708 5034
rect 8668 4616 8720 4622
rect 8668 4558 8720 4564
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 7748 4072 7800 4078
rect 7748 4014 7800 4020
rect 7196 3732 7248 3738
rect 7196 3674 7248 3680
rect 8390 2952 8446 2961
rect 8390 2887 8446 2896
rect 7564 2508 7616 2514
rect 7564 2450 7616 2456
rect 7576 2417 7604 2450
rect 7562 2408 7618 2417
rect 7562 2343 7618 2352
rect 6828 2304 6880 2310
rect 6828 2246 6880 2252
rect 5630 54 6132 82
rect 6840 82 6868 2246
rect 6918 82 6974 480
rect 6840 54 6974 82
rect 3054 0 3110 54
rect 4342 0 4398 54
rect 5630 0 5686 54
rect 6918 0 6974 54
rect 8114 82 8170 480
rect 8404 82 8432 2887
rect 8956 2514 8984 13767
rect 9324 13190 9352 14758
rect 9508 14618 9536 14826
rect 9496 14612 9548 14618
rect 9496 14554 9548 14560
rect 9772 14272 9824 14278
rect 9772 14214 9824 14220
rect 9680 13796 9732 13802
rect 9784 13784 9812 14214
rect 9968 13814 9996 27526
rect 10414 27520 10470 27526
rect 11440 27526 11850 27554
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 11244 24608 11296 24614
rect 11244 24550 11296 24556
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10048 24064 10100 24070
rect 10048 24006 10100 24012
rect 10060 20942 10088 24006
rect 11256 23798 11284 24550
rect 11440 23866 11468 27526
rect 11794 27520 11850 27526
rect 13174 27520 13230 28000
rect 14646 27554 14702 28000
rect 14476 27526 14702 27554
rect 11612 24880 11664 24886
rect 11612 24822 11664 24828
rect 11624 24274 11652 24822
rect 13188 24614 13216 27520
rect 13176 24608 13228 24614
rect 13176 24550 13228 24556
rect 11612 24268 11664 24274
rect 11612 24210 11664 24216
rect 11624 23866 11652 24210
rect 11428 23860 11480 23866
rect 11428 23802 11480 23808
rect 11612 23860 11664 23866
rect 11612 23802 11664 23808
rect 11244 23792 11296 23798
rect 11244 23734 11296 23740
rect 11256 23662 11284 23734
rect 11244 23656 11296 23662
rect 11244 23598 11296 23604
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 11058 23080 11114 23089
rect 10980 23050 11058 23066
rect 10968 23044 11058 23050
rect 11020 23038 11058 23044
rect 11058 23015 11114 23024
rect 10968 22986 11020 22992
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10048 20936 10100 20942
rect 10048 20878 10100 20884
rect 11060 20936 11112 20942
rect 11060 20878 11112 20884
rect 10048 20800 10100 20806
rect 10048 20742 10100 20748
rect 10324 20800 10376 20806
rect 10324 20742 10376 20748
rect 10060 18290 10088 20742
rect 10232 20528 10284 20534
rect 10232 20470 10284 20476
rect 10244 20398 10272 20470
rect 10336 20398 10364 20742
rect 10232 20392 10284 20398
rect 10232 20334 10284 20340
rect 10324 20392 10376 20398
rect 10324 20334 10376 20340
rect 10140 20256 10192 20262
rect 10140 20198 10192 20204
rect 10876 20256 10928 20262
rect 10876 20198 10928 20204
rect 10152 19922 10180 20198
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10232 19984 10284 19990
rect 10232 19926 10284 19932
rect 10140 19916 10192 19922
rect 10140 19858 10192 19864
rect 10152 19514 10180 19858
rect 10140 19508 10192 19514
rect 10140 19450 10192 19456
rect 10244 19446 10272 19926
rect 10888 19446 10916 20198
rect 10232 19440 10284 19446
rect 10232 19382 10284 19388
rect 10876 19440 10928 19446
rect 10876 19382 10928 19388
rect 10244 19334 10272 19382
rect 10152 19306 10272 19334
rect 10152 19174 10180 19306
rect 10888 19242 10916 19382
rect 10876 19236 10928 19242
rect 10876 19178 10928 19184
rect 10140 19168 10192 19174
rect 10140 19110 10192 19116
rect 10048 18284 10100 18290
rect 10048 18226 10100 18232
rect 10152 18154 10180 19110
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10508 18896 10560 18902
rect 10508 18838 10560 18844
rect 10520 18426 10548 18838
rect 10876 18760 10928 18766
rect 10876 18702 10928 18708
rect 10508 18420 10560 18426
rect 10508 18362 10560 18368
rect 10784 18420 10836 18426
rect 10784 18362 10836 18368
rect 10692 18284 10744 18290
rect 10692 18226 10744 18232
rect 10140 18148 10192 18154
rect 10140 18090 10192 18096
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10704 17882 10732 18226
rect 10796 18154 10824 18362
rect 10784 18148 10836 18154
rect 10784 18090 10836 18096
rect 10692 17876 10744 17882
rect 10692 17818 10744 17824
rect 10048 17672 10100 17678
rect 10048 17614 10100 17620
rect 10060 17338 10088 17614
rect 10796 17338 10824 18090
rect 10048 17332 10100 17338
rect 10048 17274 10100 17280
rect 10784 17332 10836 17338
rect 10784 17274 10836 17280
rect 10692 17196 10744 17202
rect 10692 17138 10744 17144
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10704 16794 10732 17138
rect 10692 16788 10744 16794
rect 10692 16730 10744 16736
rect 10140 16448 10192 16454
rect 10140 16390 10192 16396
rect 10152 15638 10180 16390
rect 10692 15904 10744 15910
rect 10692 15846 10744 15852
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10140 15632 10192 15638
rect 10140 15574 10192 15580
rect 10600 15632 10652 15638
rect 10704 15620 10732 15846
rect 10652 15592 10732 15620
rect 10600 15574 10652 15580
rect 10152 15162 10180 15574
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10140 15156 10192 15162
rect 10140 15098 10192 15104
rect 10428 15026 10456 15438
rect 10416 15020 10468 15026
rect 10416 14962 10468 14968
rect 10704 14822 10732 15592
rect 10048 14816 10100 14822
rect 10048 14758 10100 14764
rect 10692 14816 10744 14822
rect 10692 14758 10744 14764
rect 10784 14816 10836 14822
rect 10784 14758 10836 14764
rect 9732 13756 9812 13784
rect 9680 13738 9732 13744
rect 9312 13184 9364 13190
rect 9312 13126 9364 13132
rect 9324 12986 9352 13126
rect 9312 12980 9364 12986
rect 9312 12922 9364 12928
rect 9324 12714 9352 12922
rect 9496 12844 9548 12850
rect 9496 12786 9548 12792
rect 9312 12708 9364 12714
rect 9312 12650 9364 12656
rect 9036 12640 9088 12646
rect 9036 12582 9088 12588
rect 9048 12238 9076 12582
rect 9508 12442 9536 12786
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9496 12436 9548 12442
rect 9496 12378 9548 12384
rect 9036 12232 9088 12238
rect 9036 12174 9088 12180
rect 9048 11898 9076 12174
rect 9036 11892 9088 11898
rect 9036 11834 9088 11840
rect 9588 11212 9640 11218
rect 9588 11154 9640 11160
rect 9600 10742 9628 11154
rect 9588 10736 9640 10742
rect 9588 10678 9640 10684
rect 9312 10600 9364 10606
rect 9312 10542 9364 10548
rect 9324 10470 9352 10542
rect 9312 10464 9364 10470
rect 9312 10406 9364 10412
rect 9220 9920 9272 9926
rect 9220 9862 9272 9868
rect 9128 9444 9180 9450
rect 9128 9386 9180 9392
rect 9036 8356 9088 8362
rect 9036 8298 9088 8304
rect 9048 5642 9076 8298
rect 9140 7342 9168 9386
rect 9232 9382 9260 9862
rect 9324 9382 9352 10406
rect 9220 9376 9272 9382
rect 9220 9318 9272 9324
rect 9312 9376 9364 9382
rect 9312 9318 9364 9324
rect 9232 8838 9260 9318
rect 9220 8832 9272 8838
rect 9220 8774 9272 8780
rect 9232 7750 9260 8774
rect 9324 8430 9352 9318
rect 9588 8492 9640 8498
rect 9588 8434 9640 8440
rect 9312 8424 9364 8430
rect 9312 8366 9364 8372
rect 9404 8356 9456 8362
rect 9404 8298 9456 8304
rect 9220 7744 9272 7750
rect 9220 7686 9272 7692
rect 9232 7478 9260 7686
rect 9220 7472 9272 7478
rect 9220 7414 9272 7420
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 9140 6866 9168 7278
rect 9232 7002 9260 7414
rect 9416 7410 9444 8298
rect 9600 8294 9628 8434
rect 9588 8288 9640 8294
rect 9588 8230 9640 8236
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 9312 7268 9364 7274
rect 9312 7210 9364 7216
rect 9220 6996 9272 7002
rect 9220 6938 9272 6944
rect 9128 6860 9180 6866
rect 9128 6802 9180 6808
rect 9324 6798 9352 7210
rect 9600 7206 9628 8230
rect 9588 7200 9640 7206
rect 9588 7142 9640 7148
rect 9312 6792 9364 6798
rect 9312 6734 9364 6740
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 9036 5636 9088 5642
rect 9036 5578 9088 5584
rect 9324 5098 9352 5646
rect 9312 5092 9364 5098
rect 9312 5034 9364 5040
rect 9324 4758 9352 5034
rect 9312 4752 9364 4758
rect 9312 4694 9364 4700
rect 9692 4154 9720 12582
rect 9784 12442 9812 13756
rect 9876 13786 9996 13814
rect 9772 12436 9824 12442
rect 9772 12378 9824 12384
rect 9876 11898 9904 13786
rect 9956 12096 10008 12102
rect 9956 12038 10008 12044
rect 9864 11892 9916 11898
rect 9864 11834 9916 11840
rect 9968 11694 9996 12038
rect 10060 11762 10088 14758
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10508 14544 10560 14550
rect 10704 14532 10732 14758
rect 10560 14504 10732 14532
rect 10508 14486 10560 14492
rect 10416 14408 10468 14414
rect 10416 14350 10468 14356
rect 10428 14074 10456 14350
rect 10416 14068 10468 14074
rect 10416 14010 10468 14016
rect 10520 14006 10548 14486
rect 10508 14000 10560 14006
rect 10508 13942 10560 13948
rect 10796 13814 10824 14758
rect 10140 13796 10192 13802
rect 10140 13738 10192 13744
rect 10704 13786 10824 13814
rect 10152 13462 10180 13738
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10140 13456 10192 13462
rect 10140 13398 10192 13404
rect 10416 13456 10468 13462
rect 10416 13398 10468 13404
rect 10152 12986 10180 13398
rect 10140 12980 10192 12986
rect 10140 12922 10192 12928
rect 10428 12918 10456 13398
rect 10416 12912 10468 12918
rect 10416 12854 10468 12860
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10704 12306 10732 13786
rect 10784 13320 10836 13326
rect 10784 13262 10836 13268
rect 10796 12986 10824 13262
rect 10784 12980 10836 12986
rect 10784 12922 10836 12928
rect 10692 12300 10744 12306
rect 10692 12242 10744 12248
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 9956 11688 10008 11694
rect 10324 11688 10376 11694
rect 9956 11630 10008 11636
rect 10152 11648 10324 11676
rect 9968 10198 9996 11630
rect 10152 11354 10180 11648
rect 10324 11630 10376 11636
rect 10784 11688 10836 11694
rect 10784 11630 10836 11636
rect 10796 11558 10824 11630
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 10152 10606 10180 11290
rect 10140 10600 10192 10606
rect 10140 10542 10192 10548
rect 9956 10192 10008 10198
rect 9956 10134 10008 10140
rect 9968 9722 9996 10134
rect 9956 9716 10008 9722
rect 10152 9674 10180 10542
rect 10692 10532 10744 10538
rect 10692 10474 10744 10480
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 9956 9658 10008 9664
rect 10060 9654 10180 9674
rect 10048 9648 10180 9654
rect 10100 9646 10180 9648
rect 10048 9590 10100 9596
rect 10520 9518 10548 10066
rect 10704 9761 10732 10474
rect 10796 9926 10824 11494
rect 10784 9920 10836 9926
rect 10784 9862 10836 9868
rect 10690 9752 10746 9761
rect 10690 9687 10746 9696
rect 10796 9518 10824 9862
rect 10508 9512 10560 9518
rect 10508 9454 10560 9460
rect 10784 9512 10836 9518
rect 10784 9454 10836 9460
rect 10140 9444 10192 9450
rect 10140 9386 10192 9392
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 10060 8634 10088 9318
rect 10152 9178 10180 9386
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10796 9042 10824 9454
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 10796 8634 10824 8978
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 9956 8356 10008 8362
rect 9956 8298 10008 8304
rect 9968 8022 9996 8298
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 9956 8016 10008 8022
rect 9956 7958 10008 7964
rect 9968 7546 9996 7958
rect 10048 7744 10100 7750
rect 10048 7686 10100 7692
rect 9956 7540 10008 7546
rect 9956 7482 10008 7488
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 9968 7002 9996 7142
rect 9956 6996 10008 7002
rect 9956 6938 10008 6944
rect 9968 6118 9996 6938
rect 10060 6458 10088 7686
rect 10784 7404 10836 7410
rect 10784 7346 10836 7352
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10796 6934 10824 7346
rect 10784 6928 10836 6934
rect 10784 6870 10836 6876
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 10060 6118 10088 6394
rect 10692 6316 10744 6322
rect 10692 6258 10744 6264
rect 9956 6112 10008 6118
rect 9956 6054 10008 6060
rect 10048 6112 10100 6118
rect 10048 6054 10100 6060
rect 9864 5840 9916 5846
rect 9864 5782 9916 5788
rect 9876 4690 9904 5782
rect 9968 5370 9996 6054
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10704 5574 10732 6258
rect 10692 5568 10744 5574
rect 10692 5510 10744 5516
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 10048 5092 10100 5098
rect 10048 5034 10100 5040
rect 9956 5024 10008 5030
rect 9956 4966 10008 4972
rect 9968 4826 9996 4966
rect 9956 4820 10008 4826
rect 9956 4762 10008 4768
rect 9864 4684 9916 4690
rect 9864 4626 9916 4632
rect 9692 4146 9904 4154
rect 10060 4146 10088 5034
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10324 4684 10376 4690
rect 10324 4626 10376 4632
rect 10336 4214 10364 4626
rect 10704 4282 10732 5510
rect 10692 4276 10744 4282
rect 10692 4218 10744 4224
rect 10324 4208 10376 4214
rect 10324 4150 10376 4156
rect 10888 4154 10916 18702
rect 10968 18692 11020 18698
rect 10968 18634 11020 18640
rect 10980 17202 11008 18634
rect 10968 17196 11020 17202
rect 10968 17138 11020 17144
rect 10968 17060 11020 17066
rect 10968 17002 11020 17008
rect 10980 16658 11008 17002
rect 10968 16652 11020 16658
rect 10968 16594 11020 16600
rect 11072 16114 11100 20878
rect 11256 20505 11284 23598
rect 13636 23180 13688 23186
rect 13636 23122 13688 23128
rect 14096 23180 14148 23186
rect 14096 23122 14148 23128
rect 12440 22976 12492 22982
rect 12440 22918 12492 22924
rect 12716 22976 12768 22982
rect 12716 22918 12768 22924
rect 12162 22672 12218 22681
rect 12162 22607 12218 22616
rect 12176 22098 12204 22607
rect 12256 22432 12308 22438
rect 12256 22374 12308 22380
rect 12164 22092 12216 22098
rect 12164 22034 12216 22040
rect 12176 21690 12204 22034
rect 12164 21684 12216 21690
rect 11992 21644 12164 21672
rect 11520 21072 11572 21078
rect 11520 21014 11572 21020
rect 11532 20602 11560 21014
rect 11796 20936 11848 20942
rect 11796 20878 11848 20884
rect 11612 20800 11664 20806
rect 11612 20742 11664 20748
rect 11520 20596 11572 20602
rect 11520 20538 11572 20544
rect 11242 20496 11298 20505
rect 11242 20431 11298 20440
rect 11244 20392 11296 20398
rect 11244 20334 11296 20340
rect 11152 19712 11204 19718
rect 11152 19654 11204 19660
rect 11164 19242 11192 19654
rect 11152 19236 11204 19242
rect 11152 19178 11204 19184
rect 11152 17604 11204 17610
rect 11152 17546 11204 17552
rect 11164 17202 11192 17546
rect 11256 17270 11284 20334
rect 11336 19712 11388 19718
rect 11336 19654 11388 19660
rect 11348 19310 11376 19654
rect 11532 19514 11560 20538
rect 11624 20466 11652 20742
rect 11808 20466 11836 20878
rect 11612 20460 11664 20466
rect 11612 20402 11664 20408
rect 11796 20460 11848 20466
rect 11796 20402 11848 20408
rect 11808 20369 11836 20402
rect 11794 20360 11850 20369
rect 11794 20295 11850 20304
rect 11888 19916 11940 19922
rect 11888 19858 11940 19864
rect 11520 19508 11572 19514
rect 11520 19450 11572 19456
rect 11900 19446 11928 19858
rect 11888 19440 11940 19446
rect 11888 19382 11940 19388
rect 11336 19304 11388 19310
rect 11336 19246 11388 19252
rect 11348 18970 11376 19246
rect 11336 18964 11388 18970
rect 11336 18906 11388 18912
rect 11794 18864 11850 18873
rect 11794 18799 11796 18808
rect 11848 18799 11850 18808
rect 11796 18770 11848 18776
rect 11808 18086 11836 18770
rect 11796 18080 11848 18086
rect 11796 18022 11848 18028
rect 11612 17808 11664 17814
rect 11612 17750 11664 17756
rect 11624 17338 11652 17750
rect 11612 17332 11664 17338
rect 11612 17274 11664 17280
rect 11244 17264 11296 17270
rect 11244 17206 11296 17212
rect 11152 17196 11204 17202
rect 11152 17138 11204 17144
rect 11624 16726 11652 17274
rect 11612 16720 11664 16726
rect 11612 16662 11664 16668
rect 11244 16584 11296 16590
rect 11244 16526 11296 16532
rect 11060 16108 11112 16114
rect 11060 16050 11112 16056
rect 11072 15638 11100 16050
rect 11256 15706 11284 16526
rect 11624 16250 11652 16662
rect 11612 16244 11664 16250
rect 11612 16186 11664 16192
rect 11244 15700 11296 15706
rect 11244 15642 11296 15648
rect 11060 15632 11112 15638
rect 11060 15574 11112 15580
rect 10968 14340 11020 14346
rect 10968 14282 11020 14288
rect 10980 13530 11008 14282
rect 11624 14074 11652 16186
rect 11612 14068 11664 14074
rect 11612 14010 11664 14016
rect 11808 13814 11836 18022
rect 11900 15570 11928 19382
rect 11888 15564 11940 15570
rect 11888 15506 11940 15512
rect 11900 15162 11928 15506
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 11808 13786 11928 13814
rect 10968 13524 11020 13530
rect 10968 13466 11020 13472
rect 11900 13394 11928 13786
rect 11428 13388 11480 13394
rect 11428 13330 11480 13336
rect 11888 13388 11940 13394
rect 11888 13330 11940 13336
rect 11440 12646 11468 13330
rect 11428 12640 11480 12646
rect 11428 12582 11480 12588
rect 11440 12306 11468 12582
rect 11900 12442 11928 13330
rect 11888 12436 11940 12442
rect 11888 12378 11940 12384
rect 11336 12300 11388 12306
rect 11336 12242 11388 12248
rect 11428 12300 11480 12306
rect 11428 12242 11480 12248
rect 11888 12300 11940 12306
rect 11888 12242 11940 12248
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 11256 11830 11284 12038
rect 11348 11830 11376 12242
rect 11244 11824 11296 11830
rect 11244 11766 11296 11772
rect 11336 11824 11388 11830
rect 11336 11766 11388 11772
rect 11900 11558 11928 12242
rect 11888 11552 11940 11558
rect 11888 11494 11940 11500
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 11348 10810 11376 11154
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 11808 10810 11836 11086
rect 11336 10804 11388 10810
rect 11336 10746 11388 10752
rect 11796 10804 11848 10810
rect 11796 10746 11848 10752
rect 11336 10464 11388 10470
rect 11336 10406 11388 10412
rect 11348 10198 11376 10406
rect 11336 10192 11388 10198
rect 11336 10134 11388 10140
rect 11348 9926 11376 10134
rect 11704 10124 11756 10130
rect 11704 10066 11756 10072
rect 11518 10024 11574 10033
rect 11518 9959 11574 9968
rect 11612 9988 11664 9994
rect 11336 9920 11388 9926
rect 11336 9862 11388 9868
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 11256 8412 11284 9318
rect 11348 9110 11376 9862
rect 11336 9104 11388 9110
rect 11336 9046 11388 9052
rect 11256 8384 11376 8412
rect 10968 8356 11020 8362
rect 10968 8298 11020 8304
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 10980 7954 11008 8298
rect 10968 7948 11020 7954
rect 10968 7890 11020 7896
rect 10980 7750 11008 7890
rect 11164 7886 11192 8298
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 10980 7546 11008 7686
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 10980 7002 11008 7482
rect 11164 7002 11192 7822
rect 10968 6996 11020 7002
rect 10968 6938 11020 6944
rect 11152 6996 11204 7002
rect 11152 6938 11204 6944
rect 11164 6322 11192 6938
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 11256 6458 11284 6734
rect 11244 6452 11296 6458
rect 11244 6394 11296 6400
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 10968 5704 11020 5710
rect 10966 5672 10968 5681
rect 11020 5672 11022 5681
rect 10966 5607 11022 5616
rect 10980 5234 11008 5607
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 11152 5024 11204 5030
rect 11152 4966 11204 4972
rect 11164 4690 11192 4966
rect 11152 4684 11204 4690
rect 11152 4626 11204 4632
rect 9692 4140 9916 4146
rect 9692 4126 9864 4140
rect 9864 4082 9916 4088
rect 10048 4140 10100 4146
rect 10888 4126 11100 4154
rect 10048 4082 10100 4088
rect 9588 3936 9640 3942
rect 9588 3878 9640 3884
rect 8944 2508 8996 2514
rect 8944 2450 8996 2456
rect 8956 2378 8984 2450
rect 8944 2372 8996 2378
rect 8944 2314 8996 2320
rect 8114 54 8432 82
rect 9402 82 9458 480
rect 9600 82 9628 3878
rect 9876 3194 9904 4082
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 10784 3120 10836 3126
rect 10784 3062 10836 3068
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 9402 54 9628 82
rect 10690 82 10746 480
rect 10796 82 10824 3062
rect 11072 1601 11100 4126
rect 11058 1592 11114 1601
rect 11058 1527 11114 1536
rect 11348 241 11376 8384
rect 11428 8016 11480 8022
rect 11428 7958 11480 7964
rect 11440 7342 11468 7958
rect 11428 7336 11480 7342
rect 11428 7278 11480 7284
rect 11440 6866 11468 7278
rect 11428 6860 11480 6866
rect 11428 6802 11480 6808
rect 11440 6662 11468 6802
rect 11428 6656 11480 6662
rect 11428 6598 11480 6604
rect 11440 5914 11468 6598
rect 11428 5908 11480 5914
rect 11428 5850 11480 5856
rect 11532 4690 11560 9959
rect 11612 9930 11664 9936
rect 11624 9654 11652 9930
rect 11612 9648 11664 9654
rect 11612 9590 11664 9596
rect 11716 9178 11744 10066
rect 11704 9172 11756 9178
rect 11704 9114 11756 9120
rect 11716 9042 11744 9114
rect 11704 9036 11756 9042
rect 11888 9036 11940 9042
rect 11756 8996 11836 9024
rect 11704 8978 11756 8984
rect 11704 8900 11756 8906
rect 11704 8842 11756 8848
rect 11716 7993 11744 8842
rect 11808 8022 11836 8996
rect 11888 8978 11940 8984
rect 11900 8430 11928 8978
rect 11888 8424 11940 8430
rect 11888 8366 11940 8372
rect 11796 8016 11848 8022
rect 11702 7984 11758 7993
rect 11796 7958 11848 7964
rect 11702 7919 11758 7928
rect 11716 7546 11744 7919
rect 11704 7540 11756 7546
rect 11704 7482 11756 7488
rect 11716 6798 11744 7482
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 11992 4690 12020 21644
rect 12164 21626 12216 21632
rect 12268 21418 12296 22374
rect 12452 22234 12480 22918
rect 12728 22574 12756 22918
rect 13268 22636 13320 22642
rect 13268 22578 13320 22584
rect 12716 22568 12768 22574
rect 12716 22510 12768 22516
rect 12440 22228 12492 22234
rect 12440 22170 12492 22176
rect 12624 21480 12676 21486
rect 12624 21422 12676 21428
rect 12256 21412 12308 21418
rect 12256 21354 12308 21360
rect 12636 20806 12664 21422
rect 12624 20800 12676 20806
rect 12624 20742 12676 20748
rect 12636 20398 12664 20742
rect 12728 20534 12756 22510
rect 13176 21888 13228 21894
rect 13176 21830 13228 21836
rect 12900 21480 12952 21486
rect 12900 21422 12952 21428
rect 12808 20936 12860 20942
rect 12808 20878 12860 20884
rect 12716 20528 12768 20534
rect 12716 20470 12768 20476
rect 12624 20392 12676 20398
rect 12624 20334 12676 20340
rect 12532 19712 12584 19718
rect 12532 19654 12584 19660
rect 12544 19378 12572 19654
rect 12820 19378 12848 20878
rect 12532 19372 12584 19378
rect 12532 19314 12584 19320
rect 12808 19372 12860 19378
rect 12808 19314 12860 19320
rect 12820 18290 12848 19314
rect 12440 18284 12492 18290
rect 12440 18226 12492 18232
rect 12808 18284 12860 18290
rect 12808 18226 12860 18232
rect 12348 17536 12400 17542
rect 12348 17478 12400 17484
rect 12360 17338 12388 17478
rect 12348 17332 12400 17338
rect 12348 17274 12400 17280
rect 12360 16998 12388 17274
rect 12452 17048 12480 18226
rect 12716 18216 12768 18222
rect 12716 18158 12768 18164
rect 12532 18080 12584 18086
rect 12532 18022 12584 18028
rect 12544 17882 12572 18022
rect 12532 17876 12584 17882
rect 12532 17818 12584 17824
rect 12532 17060 12584 17066
rect 12452 17020 12532 17048
rect 12348 16992 12400 16998
rect 12348 16934 12400 16940
rect 12452 16794 12480 17020
rect 12532 17002 12584 17008
rect 12440 16788 12492 16794
rect 12440 16730 12492 16736
rect 12624 16652 12676 16658
rect 12624 16594 12676 16600
rect 12636 16046 12664 16594
rect 12728 16522 12756 18158
rect 12912 17649 12940 21422
rect 13188 21078 13216 21830
rect 13176 21072 13228 21078
rect 13176 21014 13228 21020
rect 13280 19922 13308 22578
rect 13648 22438 13676 23122
rect 14108 22778 14136 23122
rect 14280 23112 14332 23118
rect 14280 23054 14332 23060
rect 14096 22772 14148 22778
rect 14096 22714 14148 22720
rect 14108 22574 14136 22714
rect 14096 22568 14148 22574
rect 14096 22510 14148 22516
rect 13636 22432 13688 22438
rect 13636 22374 13688 22380
rect 13360 21412 13412 21418
rect 13360 21354 13412 21360
rect 13372 21146 13400 21354
rect 13360 21140 13412 21146
rect 13360 21082 13412 21088
rect 13372 20466 13400 21082
rect 13544 20528 13596 20534
rect 13544 20470 13596 20476
rect 13360 20460 13412 20466
rect 13360 20402 13412 20408
rect 13360 20256 13412 20262
rect 13360 20198 13412 20204
rect 13372 19990 13400 20198
rect 13360 19984 13412 19990
rect 13360 19926 13412 19932
rect 13268 19916 13320 19922
rect 13268 19858 13320 19864
rect 13280 18970 13308 19858
rect 13372 19334 13400 19926
rect 13452 19372 13504 19378
rect 13372 19320 13452 19334
rect 13372 19314 13504 19320
rect 13372 19306 13492 19314
rect 13464 19174 13492 19306
rect 13452 19168 13504 19174
rect 13452 19110 13504 19116
rect 13268 18964 13320 18970
rect 13268 18906 13320 18912
rect 12992 18828 13044 18834
rect 12992 18770 13044 18776
rect 13004 18222 13032 18770
rect 12992 18216 13044 18222
rect 12992 18158 13044 18164
rect 12898 17640 12954 17649
rect 12898 17575 12954 17584
rect 12716 16516 12768 16522
rect 12716 16458 12768 16464
rect 12912 16250 12940 17575
rect 13004 17542 13032 18158
rect 12992 17536 13044 17542
rect 12992 17478 13044 17484
rect 13360 17536 13412 17542
rect 13360 17478 13412 17484
rect 13004 17270 13032 17478
rect 12992 17264 13044 17270
rect 12992 17206 13044 17212
rect 13268 16992 13320 16998
rect 13268 16934 13320 16940
rect 12900 16244 12952 16250
rect 12900 16186 12952 16192
rect 12348 16040 12400 16046
rect 12348 15982 12400 15988
rect 12624 16040 12676 16046
rect 12624 15982 12676 15988
rect 12256 13796 12308 13802
rect 12256 13738 12308 13744
rect 12268 12986 12296 13738
rect 12360 13258 12388 15982
rect 12532 14272 12584 14278
rect 12532 14214 12584 14220
rect 12440 13864 12492 13870
rect 12440 13806 12492 13812
rect 12452 13462 12480 13806
rect 12440 13456 12492 13462
rect 12440 13398 12492 13404
rect 12348 13252 12400 13258
rect 12348 13194 12400 13200
rect 12256 12980 12308 12986
rect 12256 12922 12308 12928
rect 12544 12782 12572 14214
rect 12636 12918 12664 15982
rect 13176 15632 13228 15638
rect 13176 15574 13228 15580
rect 13084 15496 13136 15502
rect 13084 15438 13136 15444
rect 13096 15162 13124 15438
rect 13084 15156 13136 15162
rect 13084 15098 13136 15104
rect 13188 15026 13216 15574
rect 13176 15020 13228 15026
rect 13176 14962 13228 14968
rect 12900 14816 12952 14822
rect 12900 14758 12952 14764
rect 12808 14408 12860 14414
rect 12808 14350 12860 14356
rect 12820 13530 12848 14350
rect 12912 14074 12940 14758
rect 13084 14612 13136 14618
rect 13084 14554 13136 14560
rect 12900 14068 12952 14074
rect 12900 14010 12952 14016
rect 13096 13734 13124 14554
rect 13188 14006 13216 14962
rect 13280 14890 13308 16934
rect 13372 16658 13400 17478
rect 13464 17338 13492 19110
rect 13556 18068 13584 20470
rect 13648 18873 13676 22374
rect 13820 22160 13872 22166
rect 13820 22102 13872 22108
rect 13832 21350 13860 22102
rect 13820 21344 13872 21350
rect 13820 21286 13872 21292
rect 14188 21344 14240 21350
rect 14188 21286 14240 21292
rect 13728 21072 13780 21078
rect 13728 21014 13780 21020
rect 13740 20602 13768 21014
rect 13728 20596 13780 20602
rect 13728 20538 13780 20544
rect 13728 20324 13780 20330
rect 13728 20266 13780 20272
rect 13740 19990 13768 20266
rect 14200 20058 14228 21286
rect 14292 20058 14320 23054
rect 14372 23044 14424 23050
rect 14372 22986 14424 22992
rect 14384 22098 14412 22986
rect 14476 22778 14504 27526
rect 14646 27520 14702 27526
rect 16026 27554 16082 28000
rect 16026 27526 16344 27554
rect 16026 27520 16082 27526
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 15660 23248 15712 23254
rect 15660 23190 15712 23196
rect 14648 22976 14700 22982
rect 14648 22918 14700 22924
rect 14464 22772 14516 22778
rect 14464 22714 14516 22720
rect 14464 22500 14516 22506
rect 14464 22442 14516 22448
rect 14372 22092 14424 22098
rect 14372 22034 14424 22040
rect 14188 20052 14240 20058
rect 14188 19994 14240 20000
rect 14280 20052 14332 20058
rect 14280 19994 14332 20000
rect 13728 19984 13780 19990
rect 13728 19926 13780 19932
rect 14292 19378 14320 19994
rect 14280 19372 14332 19378
rect 14280 19314 14332 19320
rect 13634 18864 13690 18873
rect 13634 18799 13690 18808
rect 14280 18828 14332 18834
rect 14280 18770 14332 18776
rect 14292 18086 14320 18770
rect 14384 18766 14412 22034
rect 14476 21078 14504 22442
rect 14660 22438 14688 22918
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 15672 22506 15700 23190
rect 16316 23186 16344 27526
rect 17406 27520 17462 28000
rect 17512 27526 17816 27554
rect 17420 27418 17448 27520
rect 17512 27418 17540 27526
rect 17420 27390 17540 27418
rect 16486 23760 16542 23769
rect 16486 23695 16542 23704
rect 16500 23662 16528 23695
rect 16396 23656 16448 23662
rect 16396 23598 16448 23604
rect 16488 23656 16540 23662
rect 16488 23598 16540 23604
rect 16304 23180 16356 23186
rect 16304 23122 16356 23128
rect 16408 23118 16436 23598
rect 17316 23180 17368 23186
rect 17316 23122 17368 23128
rect 16396 23112 16448 23118
rect 16396 23054 16448 23060
rect 16408 22778 16436 23054
rect 16396 22772 16448 22778
rect 16396 22714 16448 22720
rect 17328 22574 17356 23122
rect 17408 22976 17460 22982
rect 17408 22918 17460 22924
rect 17316 22568 17368 22574
rect 17316 22510 17368 22516
rect 15660 22500 15712 22506
rect 15660 22442 15712 22448
rect 16120 22500 16172 22506
rect 16120 22442 16172 22448
rect 14648 22432 14700 22438
rect 14648 22374 14700 22380
rect 15384 22432 15436 22438
rect 15384 22374 15436 22380
rect 15292 21956 15344 21962
rect 15292 21898 15344 21904
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 14648 21548 14700 21554
rect 14648 21490 14700 21496
rect 14464 21072 14516 21078
rect 14464 21014 14516 21020
rect 14476 20534 14504 21014
rect 14660 20806 14688 21490
rect 15200 21412 15252 21418
rect 15200 21354 15252 21360
rect 15212 21026 15240 21354
rect 15304 21146 15332 21898
rect 15396 21146 15424 22374
rect 16132 22030 16160 22442
rect 16948 22432 17000 22438
rect 16948 22374 17000 22380
rect 16960 22098 16988 22374
rect 17420 22166 17448 22918
rect 17788 22438 17816 27526
rect 18786 27520 18842 28000
rect 20166 27520 20222 28000
rect 21638 27520 21694 28000
rect 23018 27520 23074 28000
rect 24398 27554 24454 28000
rect 24136 27526 24454 27554
rect 18144 23656 18196 23662
rect 18144 23598 18196 23604
rect 18156 23089 18184 23598
rect 18142 23080 18198 23089
rect 18142 23015 18198 23024
rect 17776 22432 17828 22438
rect 17776 22374 17828 22380
rect 18420 22432 18472 22438
rect 18420 22374 18472 22380
rect 17408 22160 17460 22166
rect 17408 22102 17460 22108
rect 16948 22092 17000 22098
rect 16948 22034 17000 22040
rect 16120 22024 16172 22030
rect 16120 21966 16172 21972
rect 16672 22024 16724 22030
rect 16672 21966 16724 21972
rect 16396 21548 16448 21554
rect 16396 21490 16448 21496
rect 15476 21344 15528 21350
rect 15476 21286 15528 21292
rect 15292 21140 15344 21146
rect 15292 21082 15344 21088
rect 15384 21140 15436 21146
rect 15384 21082 15436 21088
rect 15488 21078 15516 21286
rect 15476 21072 15528 21078
rect 15212 20998 15332 21026
rect 15476 21014 15528 21020
rect 15304 20874 15332 20998
rect 15384 20936 15436 20942
rect 15384 20878 15436 20884
rect 15292 20868 15344 20874
rect 15292 20810 15344 20816
rect 14648 20800 14700 20806
rect 14648 20742 14700 20748
rect 14464 20528 14516 20534
rect 14464 20470 14516 20476
rect 14660 18970 14688 20742
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 15304 19786 15332 20810
rect 15396 20602 15424 20878
rect 15384 20596 15436 20602
rect 15384 20538 15436 20544
rect 15488 20262 15516 21014
rect 16408 20806 16436 21490
rect 16684 21418 16712 21966
rect 16960 21690 16988 22034
rect 17420 21690 17448 22102
rect 16948 21684 17000 21690
rect 16948 21626 17000 21632
rect 17408 21684 17460 21690
rect 17408 21626 17460 21632
rect 17774 21584 17830 21593
rect 18432 21554 18460 22374
rect 18512 22160 18564 22166
rect 18512 22102 18564 22108
rect 17774 21519 17830 21528
rect 18420 21548 18472 21554
rect 16672 21412 16724 21418
rect 16672 21354 16724 21360
rect 16396 20800 16448 20806
rect 16396 20742 16448 20748
rect 16304 20392 16356 20398
rect 16304 20334 16356 20340
rect 15476 20256 15528 20262
rect 15476 20198 15528 20204
rect 15292 19780 15344 19786
rect 15292 19722 15344 19728
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 14648 18964 14700 18970
rect 14648 18906 14700 18912
rect 15200 18964 15252 18970
rect 15304 18952 15332 19722
rect 15488 19174 15516 20198
rect 15752 19984 15804 19990
rect 15752 19926 15804 19932
rect 15764 19242 15792 19926
rect 15752 19236 15804 19242
rect 15752 19178 15804 19184
rect 16120 19236 16172 19242
rect 16120 19178 16172 19184
rect 15476 19168 15528 19174
rect 15476 19110 15528 19116
rect 15660 19168 15712 19174
rect 15660 19110 15712 19116
rect 15252 18924 15332 18952
rect 15200 18906 15252 18912
rect 15384 18896 15436 18902
rect 15304 18856 15384 18884
rect 14372 18760 14424 18766
rect 14372 18702 14424 18708
rect 14832 18760 14884 18766
rect 14832 18702 14884 18708
rect 14740 18692 14792 18698
rect 14740 18634 14792 18640
rect 14556 18624 14608 18630
rect 14556 18566 14608 18572
rect 14568 18426 14596 18566
rect 14556 18420 14608 18426
rect 14556 18362 14608 18368
rect 13636 18080 13688 18086
rect 13556 18040 13636 18068
rect 13636 18022 13688 18028
rect 14280 18080 14332 18086
rect 14280 18022 14332 18028
rect 13648 17746 13676 18022
rect 13636 17740 13688 17746
rect 13636 17682 13688 17688
rect 14188 17740 14240 17746
rect 14188 17682 14240 17688
rect 13452 17332 13504 17338
rect 13452 17274 13504 17280
rect 13648 16998 13676 17682
rect 14200 17202 14228 17682
rect 14188 17196 14240 17202
rect 14188 17138 14240 17144
rect 13636 16992 13688 16998
rect 13636 16934 13688 16940
rect 13360 16652 13412 16658
rect 13360 16594 13412 16600
rect 13372 16114 13400 16594
rect 13912 16448 13964 16454
rect 13912 16390 13964 16396
rect 13360 16108 13412 16114
rect 13360 16050 13412 16056
rect 13924 15978 13952 16390
rect 14188 16176 14240 16182
rect 14188 16118 14240 16124
rect 13452 15972 13504 15978
rect 13452 15914 13504 15920
rect 13912 15972 13964 15978
rect 13912 15914 13964 15920
rect 13464 15502 13492 15914
rect 13452 15496 13504 15502
rect 13452 15438 13504 15444
rect 13268 14884 13320 14890
rect 13268 14826 13320 14832
rect 13924 14618 13952 15914
rect 14004 15360 14056 15366
rect 14004 15302 14056 15308
rect 14016 15026 14044 15302
rect 14200 15094 14228 16118
rect 14188 15088 14240 15094
rect 14188 15030 14240 15036
rect 14004 15020 14056 15026
rect 14004 14962 14056 14968
rect 13912 14612 13964 14618
rect 13912 14554 13964 14560
rect 13726 14512 13782 14521
rect 14016 14498 14044 14962
rect 13726 14447 13782 14456
rect 13924 14470 14044 14498
rect 13176 14000 13228 14006
rect 13176 13942 13228 13948
rect 13084 13728 13136 13734
rect 13084 13670 13136 13676
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 13096 13462 13124 13670
rect 13084 13456 13136 13462
rect 13084 13398 13136 13404
rect 13084 13320 13136 13326
rect 13084 13262 13136 13268
rect 12624 12912 12676 12918
rect 12624 12854 12676 12860
rect 12532 12776 12584 12782
rect 12532 12718 12584 12724
rect 12256 12164 12308 12170
rect 12256 12106 12308 12112
rect 12268 11898 12296 12106
rect 12256 11892 12308 11898
rect 12256 11834 12308 11840
rect 12544 9382 12572 12718
rect 12636 11014 12664 12854
rect 12716 12708 12768 12714
rect 12716 12650 12768 12656
rect 12728 11286 12756 12650
rect 13096 12374 13124 13262
rect 13740 12714 13768 14447
rect 13176 12708 13228 12714
rect 13176 12650 13228 12656
rect 13728 12708 13780 12714
rect 13728 12650 13780 12656
rect 13084 12368 13136 12374
rect 13084 12310 13136 12316
rect 12808 11552 12860 11558
rect 12808 11494 12860 11500
rect 12716 11280 12768 11286
rect 12716 11222 12768 11228
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 12636 10266 12664 10950
rect 12728 10810 12756 11222
rect 12716 10804 12768 10810
rect 12716 10746 12768 10752
rect 12728 10538 12756 10746
rect 12716 10532 12768 10538
rect 12716 10474 12768 10480
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12636 9518 12664 10202
rect 12820 9518 12848 11494
rect 13084 10736 13136 10742
rect 13084 10678 13136 10684
rect 12900 10668 12952 10674
rect 12900 10610 12952 10616
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 12912 10266 12940 10610
rect 12900 10260 12952 10266
rect 12900 10202 12952 10208
rect 13004 9586 13032 10610
rect 12992 9580 13044 9586
rect 12992 9522 13044 9528
rect 12624 9512 12676 9518
rect 12624 9454 12676 9460
rect 12808 9512 12860 9518
rect 12808 9454 12860 9460
rect 12532 9376 12584 9382
rect 12532 9318 12584 9324
rect 12820 9178 12848 9454
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 12360 8498 12388 8910
rect 12348 8492 12400 8498
rect 12348 8434 12400 8440
rect 12360 8090 12388 8434
rect 12348 8084 12400 8090
rect 12348 8026 12400 8032
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12532 7744 12584 7750
rect 12532 7686 12584 7692
rect 12164 7200 12216 7206
rect 12164 7142 12216 7148
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12176 6934 12204 7142
rect 12164 6928 12216 6934
rect 12164 6870 12216 6876
rect 12452 6662 12480 7142
rect 12440 6656 12492 6662
rect 12440 6598 12492 6604
rect 12256 6112 12308 6118
rect 12256 6054 12308 6060
rect 12268 5846 12296 6054
rect 12256 5840 12308 5846
rect 12256 5782 12308 5788
rect 12164 5772 12216 5778
rect 12164 5714 12216 5720
rect 12176 4758 12204 5714
rect 12268 5370 12296 5782
rect 12256 5364 12308 5370
rect 12256 5306 12308 5312
rect 12164 4752 12216 4758
rect 12164 4694 12216 4700
rect 11520 4684 11572 4690
rect 11520 4626 11572 4632
rect 11980 4684 12032 4690
rect 11980 4626 12032 4632
rect 11532 4282 11560 4626
rect 11992 4282 12020 4626
rect 11520 4276 11572 4282
rect 11520 4218 11572 4224
rect 11980 4276 12032 4282
rect 11980 4218 12032 4224
rect 11992 3194 12020 4218
rect 12452 4146 12480 6598
rect 12544 4826 12572 7686
rect 12820 7410 12848 7822
rect 12808 7404 12860 7410
rect 12808 7346 12860 7352
rect 12820 7313 12848 7346
rect 12806 7304 12862 7313
rect 12624 7268 12676 7274
rect 12806 7239 12862 7248
rect 12624 7210 12676 7216
rect 12636 6934 12664 7210
rect 13096 7002 13124 10678
rect 13084 6996 13136 7002
rect 13084 6938 13136 6944
rect 12624 6928 12676 6934
rect 12624 6870 12676 6876
rect 12992 6860 13044 6866
rect 12992 6802 13044 6808
rect 13004 6361 13032 6802
rect 12990 6352 13046 6361
rect 12990 6287 13046 6296
rect 13004 5846 13032 6287
rect 12992 5840 13044 5846
rect 12992 5782 13044 5788
rect 13188 5778 13216 12650
rect 13544 12640 13596 12646
rect 13544 12582 13596 12588
rect 13556 12374 13584 12582
rect 13544 12368 13596 12374
rect 13544 12310 13596 12316
rect 13452 12232 13504 12238
rect 13452 12174 13504 12180
rect 13464 11898 13492 12174
rect 13452 11892 13504 11898
rect 13452 11834 13504 11840
rect 13360 11756 13412 11762
rect 13412 11716 13492 11744
rect 13360 11698 13412 11704
rect 13268 11552 13320 11558
rect 13268 11494 13320 11500
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 13280 11218 13308 11494
rect 13268 11212 13320 11218
rect 13268 11154 13320 11160
rect 13372 10198 13400 11494
rect 13464 11014 13492 11716
rect 13556 11354 13584 12310
rect 13636 11620 13688 11626
rect 13636 11562 13688 11568
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13648 11218 13676 11562
rect 13636 11212 13688 11218
rect 13636 11154 13688 11160
rect 13728 11076 13780 11082
rect 13728 11018 13780 11024
rect 13452 11008 13504 11014
rect 13452 10950 13504 10956
rect 13360 10192 13412 10198
rect 13360 10134 13412 10140
rect 13268 10124 13320 10130
rect 13268 10066 13320 10072
rect 13280 9722 13308 10066
rect 13360 10056 13412 10062
rect 13360 9998 13412 10004
rect 13268 9716 13320 9722
rect 13268 9658 13320 9664
rect 13372 8838 13400 9998
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 13360 8424 13412 8430
rect 13360 8366 13412 8372
rect 13268 6860 13320 6866
rect 13372 6848 13400 8366
rect 13464 7546 13492 10950
rect 13636 10464 13688 10470
rect 13636 10406 13688 10412
rect 13544 9988 13596 9994
rect 13544 9930 13596 9936
rect 13452 7540 13504 7546
rect 13452 7482 13504 7488
rect 13556 7342 13584 9930
rect 13648 9654 13676 10406
rect 13740 10198 13768 11018
rect 13728 10192 13780 10198
rect 13728 10134 13780 10140
rect 13820 10192 13872 10198
rect 13820 10134 13872 10140
rect 13832 10044 13860 10134
rect 13740 10016 13860 10044
rect 13636 9648 13688 9654
rect 13636 9590 13688 9596
rect 13740 9586 13768 10016
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 13832 9382 13860 9590
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 13832 9042 13860 9318
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 13728 8832 13780 8838
rect 13728 8774 13780 8780
rect 13636 8288 13688 8294
rect 13636 8230 13688 8236
rect 13648 8022 13676 8230
rect 13636 8016 13688 8022
rect 13636 7958 13688 7964
rect 13544 7336 13596 7342
rect 13544 7278 13596 7284
rect 13452 7200 13504 7206
rect 13648 7188 13676 7958
rect 13504 7160 13676 7188
rect 13452 7142 13504 7148
rect 13320 6820 13400 6848
rect 13268 6802 13320 6808
rect 13280 6118 13308 6802
rect 13464 6186 13492 7142
rect 13452 6180 13504 6186
rect 13452 6122 13504 6128
rect 13268 6112 13320 6118
rect 13268 6054 13320 6060
rect 13740 5914 13768 8774
rect 13832 8566 13860 8978
rect 13820 8560 13872 8566
rect 13820 8502 13872 8508
rect 13820 7948 13872 7954
rect 13820 7890 13872 7896
rect 13832 7478 13860 7890
rect 13820 7472 13872 7478
rect 13820 7414 13872 7420
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 13176 5772 13228 5778
rect 13176 5714 13228 5720
rect 13728 5772 13780 5778
rect 13728 5714 13780 5720
rect 13740 5370 13768 5714
rect 13728 5364 13780 5370
rect 13728 5306 13780 5312
rect 12808 5092 12860 5098
rect 12808 5034 12860 5040
rect 12900 5092 12952 5098
rect 12900 5034 12952 5040
rect 12532 4820 12584 4826
rect 12532 4762 12584 4768
rect 12820 4146 12848 5034
rect 12912 4554 12940 5034
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 12900 4548 12952 4554
rect 12900 4490 12952 4496
rect 12440 4140 12492 4146
rect 12440 4082 12492 4088
rect 12808 4140 12860 4146
rect 12808 4082 12860 4088
rect 13740 3738 13768 4558
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 11980 3188 12032 3194
rect 11980 3130 12032 3136
rect 13924 3126 13952 14470
rect 14200 14414 14228 15030
rect 14292 14929 14320 18022
rect 14648 17332 14700 17338
rect 14648 17274 14700 17280
rect 14660 17066 14688 17274
rect 14752 17134 14780 18634
rect 14844 17882 14872 18702
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 15304 18086 15332 18856
rect 15384 18838 15436 18844
rect 15488 18154 15516 19110
rect 15476 18148 15528 18154
rect 15476 18090 15528 18096
rect 15292 18080 15344 18086
rect 15292 18022 15344 18028
rect 15304 17882 15332 18022
rect 14832 17876 14884 17882
rect 14832 17818 14884 17824
rect 15292 17876 15344 17882
rect 15292 17818 15344 17824
rect 15476 17808 15528 17814
rect 15476 17750 15528 17756
rect 14832 17672 14884 17678
rect 14832 17614 14884 17620
rect 15292 17672 15344 17678
rect 15292 17614 15344 17620
rect 14740 17128 14792 17134
rect 14740 17070 14792 17076
rect 14648 17060 14700 17066
rect 14648 17002 14700 17008
rect 14752 16794 14780 17070
rect 14740 16788 14792 16794
rect 14740 16730 14792 16736
rect 14648 16040 14700 16046
rect 14648 15982 14700 15988
rect 14278 14920 14334 14929
rect 14278 14855 14334 14864
rect 14004 14408 14056 14414
rect 14004 14350 14056 14356
rect 14188 14408 14240 14414
rect 14188 14350 14240 14356
rect 14016 13530 14044 14350
rect 14464 14340 14516 14346
rect 14464 14282 14516 14288
rect 14372 14272 14424 14278
rect 14372 14214 14424 14220
rect 14384 13802 14412 14214
rect 14476 13938 14504 14282
rect 14464 13932 14516 13938
rect 14464 13874 14516 13880
rect 14372 13796 14424 13802
rect 14372 13738 14424 13744
rect 14004 13524 14056 13530
rect 14004 13466 14056 13472
rect 14280 13524 14332 13530
rect 14280 13466 14332 13472
rect 14004 13184 14056 13190
rect 14004 13126 14056 13132
rect 14016 12986 14044 13126
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 14016 12646 14044 12922
rect 14186 12880 14242 12889
rect 14292 12850 14320 13466
rect 14186 12815 14242 12824
rect 14280 12844 14332 12850
rect 14004 12640 14056 12646
rect 14004 12582 14056 12588
rect 14096 12096 14148 12102
rect 14096 12038 14148 12044
rect 14004 11212 14056 11218
rect 14004 11154 14056 11160
rect 14016 10810 14044 11154
rect 14004 10804 14056 10810
rect 14004 10746 14056 10752
rect 14004 10532 14056 10538
rect 14004 10474 14056 10480
rect 14016 8022 14044 10474
rect 14108 9994 14136 12038
rect 14200 11762 14228 12815
rect 14280 12786 14332 12792
rect 14476 11898 14504 13874
rect 14660 12102 14688 15982
rect 14740 15972 14792 15978
rect 14740 15914 14792 15920
rect 14752 15042 14780 15914
rect 14844 15570 14872 17614
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15304 17270 15332 17614
rect 15292 17264 15344 17270
rect 15292 17206 15344 17212
rect 15488 17066 15516 17750
rect 15672 17338 15700 19110
rect 15660 17332 15712 17338
rect 15660 17274 15712 17280
rect 15568 17196 15620 17202
rect 15568 17138 15620 17144
rect 15476 17060 15528 17066
rect 15476 17002 15528 17008
rect 15488 16726 15516 17002
rect 15476 16720 15528 16726
rect 15476 16662 15528 16668
rect 15292 16652 15344 16658
rect 15292 16594 15344 16600
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15304 16250 15332 16594
rect 15488 16250 15516 16662
rect 15292 16244 15344 16250
rect 15292 16186 15344 16192
rect 15476 16244 15528 16250
rect 15476 16186 15528 16192
rect 15476 15904 15528 15910
rect 15476 15846 15528 15852
rect 14832 15564 14884 15570
rect 14832 15506 14884 15512
rect 14844 15162 14872 15506
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14832 15156 14884 15162
rect 14832 15098 14884 15104
rect 14752 15014 14872 15042
rect 14740 13252 14792 13258
rect 14740 13194 14792 13200
rect 14648 12096 14700 12102
rect 14648 12038 14700 12044
rect 14464 11892 14516 11898
rect 14464 11834 14516 11840
rect 14188 11756 14240 11762
rect 14188 11698 14240 11704
rect 14200 11354 14228 11698
rect 14280 11620 14332 11626
rect 14280 11562 14332 11568
rect 14188 11348 14240 11354
rect 14188 11290 14240 11296
rect 14292 10198 14320 11562
rect 14556 10600 14608 10606
rect 14556 10542 14608 10548
rect 14280 10192 14332 10198
rect 14280 10134 14332 10140
rect 14096 9988 14148 9994
rect 14096 9930 14148 9936
rect 14568 8974 14596 10542
rect 14752 10248 14780 13194
rect 14844 12866 14872 15014
rect 15016 14952 15068 14958
rect 15016 14894 15068 14900
rect 15028 14521 15056 14894
rect 15014 14512 15070 14521
rect 15014 14447 15070 14456
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15396 13734 15424 14418
rect 15384 13728 15436 13734
rect 15384 13670 15436 13676
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15304 12986 15332 13330
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 14922 12880 14978 12889
rect 14844 12838 14922 12866
rect 14922 12815 14978 12824
rect 14936 12714 14964 12815
rect 15396 12753 15424 13670
rect 15382 12744 15438 12753
rect 14924 12708 14976 12714
rect 15382 12679 15438 12688
rect 14924 12650 14976 12656
rect 14832 12436 14884 12442
rect 14832 12378 14884 12384
rect 14844 11898 14872 12378
rect 14936 12374 14964 12650
rect 14924 12368 14976 12374
rect 14924 12310 14976 12316
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 14832 11892 14884 11898
rect 14832 11834 14884 11840
rect 15488 11286 15516 15846
rect 15580 14278 15608 17138
rect 15764 16794 15792 19178
rect 16132 18970 16160 19178
rect 16120 18964 16172 18970
rect 16120 18906 16172 18912
rect 16316 18834 16344 20334
rect 16408 20058 16436 20742
rect 16488 20324 16540 20330
rect 16488 20266 16540 20272
rect 16396 20052 16448 20058
rect 16396 19994 16448 20000
rect 16396 19848 16448 19854
rect 16396 19790 16448 19796
rect 16408 19378 16436 19790
rect 16500 19786 16528 20266
rect 16488 19780 16540 19786
rect 16488 19722 16540 19728
rect 16396 19372 16448 19378
rect 16396 19314 16448 19320
rect 16408 18902 16436 19314
rect 16684 18970 16712 21354
rect 17408 21004 17460 21010
rect 17408 20946 17460 20952
rect 17420 20262 17448 20946
rect 17788 20942 17816 21519
rect 18420 21490 18472 21496
rect 17868 21344 17920 21350
rect 17868 21286 17920 21292
rect 17880 21078 17908 21286
rect 18524 21078 18552 22102
rect 17868 21072 17920 21078
rect 17868 21014 17920 21020
rect 18512 21072 18564 21078
rect 18512 21014 18564 21020
rect 17776 20936 17828 20942
rect 17776 20878 17828 20884
rect 17788 20602 17816 20878
rect 18052 20868 18104 20874
rect 18052 20810 18104 20816
rect 17776 20596 17828 20602
rect 17776 20538 17828 20544
rect 17224 20256 17276 20262
rect 17224 20198 17276 20204
rect 17408 20256 17460 20262
rect 17408 20198 17460 20204
rect 17132 19916 17184 19922
rect 17132 19858 17184 19864
rect 17144 19446 17172 19858
rect 17236 19514 17264 20198
rect 17420 19854 17448 20198
rect 17408 19848 17460 19854
rect 17408 19790 17460 19796
rect 17960 19848 18012 19854
rect 17960 19790 18012 19796
rect 17224 19508 17276 19514
rect 17224 19450 17276 19456
rect 17132 19440 17184 19446
rect 17132 19382 17184 19388
rect 17408 19168 17460 19174
rect 17408 19110 17460 19116
rect 17776 19168 17828 19174
rect 17776 19110 17828 19116
rect 16672 18964 16724 18970
rect 16672 18906 16724 18912
rect 16396 18896 16448 18902
rect 16396 18838 16448 18844
rect 16304 18828 16356 18834
rect 16304 18770 16356 18776
rect 17224 18828 17276 18834
rect 17224 18770 17276 18776
rect 16488 18760 16540 18766
rect 16488 18702 16540 18708
rect 16396 18624 16448 18630
rect 16396 18566 16448 18572
rect 16304 18284 16356 18290
rect 16408 18272 16436 18566
rect 16500 18290 16528 18702
rect 16356 18244 16436 18272
rect 16304 18226 16356 18232
rect 16302 17776 16358 17785
rect 16302 17711 16358 17720
rect 16316 17338 16344 17711
rect 16304 17332 16356 17338
rect 16304 17274 16356 17280
rect 16316 16794 16344 17274
rect 15752 16788 15804 16794
rect 15752 16730 15804 16736
rect 16304 16788 16356 16794
rect 16304 16730 16356 16736
rect 15752 16516 15804 16522
rect 15752 16458 15804 16464
rect 15660 15360 15712 15366
rect 15660 15302 15712 15308
rect 15672 15162 15700 15302
rect 15660 15156 15712 15162
rect 15660 15098 15712 15104
rect 15764 15094 15792 16458
rect 15936 16244 15988 16250
rect 15936 16186 15988 16192
rect 15948 15910 15976 16186
rect 16316 16046 16344 16730
rect 16304 16040 16356 16046
rect 16132 16000 16304 16028
rect 15936 15904 15988 15910
rect 15936 15846 15988 15852
rect 15948 15638 15976 15846
rect 15936 15632 15988 15638
rect 15936 15574 15988 15580
rect 15948 15162 15976 15574
rect 15936 15156 15988 15162
rect 15936 15098 15988 15104
rect 15752 15088 15804 15094
rect 15752 15030 15804 15036
rect 15568 14272 15620 14278
rect 15568 14214 15620 14220
rect 15580 13297 15608 14214
rect 15764 13814 15792 15030
rect 15844 14272 15896 14278
rect 15844 14214 15896 14220
rect 15856 13938 15884 14214
rect 15948 14074 15976 15098
rect 15936 14068 15988 14074
rect 15936 14010 15988 14016
rect 15844 13932 15896 13938
rect 15896 13892 15976 13920
rect 15844 13874 15896 13880
rect 15764 13786 15884 13814
rect 15856 13394 15884 13786
rect 15844 13388 15896 13394
rect 15844 13330 15896 13336
rect 15566 13288 15622 13297
rect 15566 13223 15622 13232
rect 15752 13184 15804 13190
rect 15752 13126 15804 13132
rect 15764 12782 15792 13126
rect 15752 12776 15804 12782
rect 15948 12753 15976 13892
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 15752 12718 15804 12724
rect 15934 12744 15990 12753
rect 15568 12300 15620 12306
rect 15568 12242 15620 12248
rect 15660 12300 15712 12306
rect 15660 12242 15712 12248
rect 15580 11830 15608 12242
rect 15568 11824 15620 11830
rect 15568 11766 15620 11772
rect 15580 11354 15608 11766
rect 15672 11626 15700 12242
rect 15764 12238 15792 12718
rect 15934 12679 15990 12688
rect 15844 12640 15896 12646
rect 15844 12582 15896 12588
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 15660 11620 15712 11626
rect 15660 11562 15712 11568
rect 15568 11348 15620 11354
rect 15568 11290 15620 11296
rect 15476 11280 15528 11286
rect 15476 11222 15528 11228
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15764 10266 15792 12174
rect 15856 10674 15884 12582
rect 15936 11552 15988 11558
rect 15936 11494 15988 11500
rect 15844 10668 15896 10674
rect 15844 10610 15896 10616
rect 15948 10538 15976 11494
rect 16040 10810 16068 13262
rect 16132 13190 16160 16000
rect 16304 15982 16356 15988
rect 16304 15564 16356 15570
rect 16304 15506 16356 15512
rect 16316 14890 16344 15506
rect 16304 14884 16356 14890
rect 16304 14826 16356 14832
rect 16316 14618 16344 14826
rect 16304 14612 16356 14618
rect 16304 14554 16356 14560
rect 16120 13184 16172 13190
rect 16120 13126 16172 13132
rect 16304 12776 16356 12782
rect 16304 12718 16356 12724
rect 16316 12306 16344 12718
rect 16304 12300 16356 12306
rect 16304 12242 16356 12248
rect 16120 12232 16172 12238
rect 16120 12174 16172 12180
rect 16132 11762 16160 12174
rect 16120 11756 16172 11762
rect 16120 11698 16172 11704
rect 16132 11354 16160 11698
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 16304 11280 16356 11286
rect 16304 11222 16356 11228
rect 16316 10810 16344 11222
rect 16028 10804 16080 10810
rect 16028 10746 16080 10752
rect 16304 10804 16356 10810
rect 16304 10746 16356 10752
rect 15936 10532 15988 10538
rect 15936 10474 15988 10480
rect 15752 10260 15804 10266
rect 14752 10220 14872 10248
rect 14740 10124 14792 10130
rect 14740 10066 14792 10072
rect 14752 9761 14780 10066
rect 14738 9752 14794 9761
rect 14738 9687 14794 9696
rect 14752 9654 14780 9687
rect 14740 9648 14792 9654
rect 14740 9590 14792 9596
rect 14556 8968 14608 8974
rect 14556 8910 14608 8916
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14476 8362 14504 8570
rect 14372 8356 14424 8362
rect 14372 8298 14424 8304
rect 14464 8356 14516 8362
rect 14464 8298 14516 8304
rect 14004 8016 14056 8022
rect 14004 7958 14056 7964
rect 14384 7818 14412 8298
rect 14372 7812 14424 7818
rect 14372 7754 14424 7760
rect 14004 6724 14056 6730
rect 14004 6666 14056 6672
rect 14016 6458 14044 6666
rect 14464 6656 14516 6662
rect 14464 6598 14516 6604
rect 14004 6452 14056 6458
rect 14004 6394 14056 6400
rect 14476 6254 14504 6598
rect 14464 6248 14516 6254
rect 14464 6190 14516 6196
rect 14188 6180 14240 6186
rect 14188 6122 14240 6128
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 14016 3641 14044 6054
rect 14200 4758 14228 6122
rect 14476 5846 14504 6190
rect 14464 5840 14516 5846
rect 14464 5782 14516 5788
rect 14476 5574 14504 5782
rect 14464 5568 14516 5574
rect 14464 5510 14516 5516
rect 14476 5098 14504 5510
rect 14372 5092 14424 5098
rect 14372 5034 14424 5040
rect 14464 5092 14516 5098
rect 14464 5034 14516 5040
rect 14384 4826 14412 5034
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 14188 4752 14240 4758
rect 14188 4694 14240 4700
rect 14200 4554 14228 4694
rect 14188 4548 14240 4554
rect 14188 4490 14240 4496
rect 14200 4282 14228 4490
rect 14188 4276 14240 4282
rect 14188 4218 14240 4224
rect 14476 4214 14504 5034
rect 14740 4820 14792 4826
rect 14740 4762 14792 4768
rect 14556 4616 14608 4622
rect 14556 4558 14608 4564
rect 14464 4208 14516 4214
rect 14464 4150 14516 4156
rect 14476 4010 14504 4150
rect 14568 4146 14596 4558
rect 14556 4140 14608 4146
rect 14556 4082 14608 4088
rect 14752 4010 14780 4762
rect 14280 4004 14332 4010
rect 14280 3946 14332 3952
rect 14464 4004 14516 4010
rect 14464 3946 14516 3952
rect 14740 4004 14792 4010
rect 14740 3946 14792 3952
rect 14002 3632 14058 3641
rect 14002 3567 14058 3576
rect 14292 3466 14320 3946
rect 14280 3460 14332 3466
rect 14280 3402 14332 3408
rect 12072 3120 12124 3126
rect 12072 3062 12124 3068
rect 13912 3120 13964 3126
rect 13912 3062 13964 3068
rect 11334 232 11390 241
rect 11334 167 11390 176
rect 10690 54 10824 82
rect 11978 82 12034 480
rect 12084 82 12112 3062
rect 14844 2650 14872 10220
rect 15752 10202 15804 10208
rect 15844 9920 15896 9926
rect 15844 9862 15896 9868
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15856 9450 15884 9862
rect 15844 9444 15896 9450
rect 15844 9386 15896 9392
rect 15568 9376 15620 9382
rect 15568 9318 15620 9324
rect 15580 9110 15608 9318
rect 15568 9104 15620 9110
rect 15568 9046 15620 9052
rect 15384 9036 15436 9042
rect 15384 8978 15436 8984
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15396 8634 15424 8978
rect 15752 8832 15804 8838
rect 15752 8774 15804 8780
rect 15764 8634 15792 8774
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 15384 8492 15436 8498
rect 15384 8434 15436 8440
rect 15396 8022 15424 8434
rect 15764 8294 15792 8570
rect 15752 8288 15804 8294
rect 15752 8230 15804 8236
rect 15384 8016 15436 8022
rect 15304 7976 15384 8004
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 15304 7002 15332 7976
rect 15384 7958 15436 7964
rect 15476 8016 15528 8022
rect 15476 7958 15528 7964
rect 15384 7268 15436 7274
rect 15384 7210 15436 7216
rect 15396 7002 15424 7210
rect 15488 7206 15516 7958
rect 15476 7200 15528 7206
rect 15476 7142 15528 7148
rect 15292 6996 15344 7002
rect 15292 6938 15344 6944
rect 15384 6996 15436 7002
rect 15384 6938 15436 6944
rect 15488 6866 15516 7142
rect 15476 6860 15528 6866
rect 15476 6802 15528 6808
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15488 6458 15516 6802
rect 15476 6452 15528 6458
rect 15476 6394 15528 6400
rect 15856 6322 15884 9386
rect 16040 8566 16068 10746
rect 16120 9580 16172 9586
rect 16120 9522 16172 9528
rect 16028 8560 16080 8566
rect 16028 8502 16080 8508
rect 15936 8356 15988 8362
rect 15936 8298 15988 8304
rect 15948 8090 15976 8298
rect 15936 8084 15988 8090
rect 15936 8026 15988 8032
rect 15936 7812 15988 7818
rect 15936 7754 15988 7760
rect 15948 7410 15976 7754
rect 15936 7404 15988 7410
rect 15936 7346 15988 7352
rect 15948 6866 15976 7346
rect 16132 7342 16160 9522
rect 16304 7880 16356 7886
rect 16304 7822 16356 7828
rect 16316 7546 16344 7822
rect 16304 7540 16356 7546
rect 16304 7482 16356 7488
rect 16120 7336 16172 7342
rect 16120 7278 16172 7284
rect 15936 6860 15988 6866
rect 15936 6802 15988 6808
rect 15844 6316 15896 6322
rect 15844 6258 15896 6264
rect 15660 6180 15712 6186
rect 15660 6122 15712 6128
rect 15476 5840 15528 5846
rect 15476 5782 15528 5788
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 15396 5370 15424 5646
rect 15384 5364 15436 5370
rect 15384 5306 15436 5312
rect 15488 5234 15516 5782
rect 15672 5302 15700 6122
rect 16028 5704 16080 5710
rect 16028 5646 16080 5652
rect 15660 5296 15712 5302
rect 15660 5238 15712 5244
rect 15476 5228 15528 5234
rect 15476 5170 15528 5176
rect 15672 4758 15700 5238
rect 16040 4758 16068 5646
rect 15660 4752 15712 4758
rect 15660 4694 15712 4700
rect 16028 4752 16080 4758
rect 16028 4694 16080 4700
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 15672 4282 15700 4694
rect 15660 4276 15712 4282
rect 15660 4218 15712 4224
rect 16040 3602 16068 4694
rect 15384 3596 15436 3602
rect 15384 3538 15436 3544
rect 16028 3596 16080 3602
rect 16028 3538 16080 3544
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 15396 3194 15424 3538
rect 15660 3392 15712 3398
rect 15660 3334 15712 3340
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 15672 2990 15700 3334
rect 15660 2984 15712 2990
rect 15660 2926 15712 2932
rect 16408 2650 16436 18244
rect 16488 18284 16540 18290
rect 16488 18226 16540 18232
rect 17236 18086 17264 18770
rect 17420 18358 17448 19110
rect 17788 18630 17816 19110
rect 17972 18970 18000 19790
rect 17960 18964 18012 18970
rect 17960 18906 18012 18912
rect 17868 18760 17920 18766
rect 17868 18702 17920 18708
rect 17776 18624 17828 18630
rect 17776 18566 17828 18572
rect 17408 18352 17460 18358
rect 17408 18294 17460 18300
rect 17788 18086 17816 18566
rect 17880 18290 17908 18702
rect 17868 18284 17920 18290
rect 17868 18226 17920 18232
rect 17224 18080 17276 18086
rect 17224 18022 17276 18028
rect 17776 18080 17828 18086
rect 17776 18022 17828 18028
rect 16488 17128 16540 17134
rect 16488 17070 16540 17076
rect 16500 16153 16528 17070
rect 16948 16992 17000 16998
rect 16948 16934 17000 16940
rect 16960 16454 16988 16934
rect 16948 16448 17000 16454
rect 16948 16390 17000 16396
rect 16486 16144 16542 16153
rect 16486 16079 16542 16088
rect 16960 16046 16988 16390
rect 16948 16040 17000 16046
rect 16948 15982 17000 15988
rect 16960 15162 16988 15982
rect 16948 15156 17000 15162
rect 16948 15098 17000 15104
rect 16856 15020 16908 15026
rect 16856 14962 16908 14968
rect 16580 14544 16632 14550
rect 16580 14486 16632 14492
rect 16592 14074 16620 14486
rect 16868 14414 16896 14962
rect 16856 14408 16908 14414
rect 16856 14350 16908 14356
rect 16580 14068 16632 14074
rect 16580 14010 16632 14016
rect 16592 13530 16620 14010
rect 16868 13530 16896 14350
rect 17040 14340 17092 14346
rect 17040 14282 17092 14288
rect 16580 13524 16632 13530
rect 16580 13466 16632 13472
rect 16856 13524 16908 13530
rect 16856 13466 16908 13472
rect 17052 13394 17080 14282
rect 17236 13705 17264 18022
rect 17788 17814 17816 18022
rect 17880 17882 17908 18226
rect 17868 17876 17920 17882
rect 17868 17818 17920 17824
rect 17776 17808 17828 17814
rect 17776 17750 17828 17756
rect 17684 17672 17736 17678
rect 17684 17614 17736 17620
rect 17696 16998 17724 17614
rect 17788 16998 17816 17750
rect 17684 16992 17736 16998
rect 17684 16934 17736 16940
rect 17776 16992 17828 16998
rect 17776 16934 17828 16940
rect 17500 16584 17552 16590
rect 17500 16526 17552 16532
rect 17512 16250 17540 16526
rect 17500 16244 17552 16250
rect 17500 16186 17552 16192
rect 17696 15706 17724 16934
rect 17788 16726 17816 16934
rect 17776 16720 17828 16726
rect 17776 16662 17828 16668
rect 17788 15910 17816 16662
rect 17776 15904 17828 15910
rect 17776 15846 17828 15852
rect 17684 15700 17736 15706
rect 17684 15642 17736 15648
rect 17684 15564 17736 15570
rect 17684 15506 17736 15512
rect 17696 15162 17724 15506
rect 17684 15156 17736 15162
rect 17684 15098 17736 15104
rect 17500 14408 17552 14414
rect 17500 14350 17552 14356
rect 17512 13802 17540 14350
rect 17500 13796 17552 13802
rect 17500 13738 17552 13744
rect 17222 13696 17278 13705
rect 17222 13631 17278 13640
rect 17040 13388 17092 13394
rect 17040 13330 17092 13336
rect 17052 12442 17080 13330
rect 17132 13252 17184 13258
rect 17132 13194 17184 13200
rect 17144 12986 17172 13194
rect 17132 12980 17184 12986
rect 17132 12922 17184 12928
rect 17040 12436 17092 12442
rect 17040 12378 17092 12384
rect 17236 12306 17264 13631
rect 17224 12300 17276 12306
rect 17224 12242 17276 12248
rect 17684 12300 17736 12306
rect 17684 12242 17736 12248
rect 17236 11830 17264 12242
rect 17316 11892 17368 11898
rect 17316 11834 17368 11840
rect 17224 11824 17276 11830
rect 17224 11766 17276 11772
rect 16488 11552 16540 11558
rect 16488 11494 16540 11500
rect 16500 11286 16528 11494
rect 16488 11280 16540 11286
rect 16488 11222 16540 11228
rect 16500 10266 16528 11222
rect 16672 11076 16724 11082
rect 16672 11018 16724 11024
rect 16488 10260 16540 10266
rect 16488 10202 16540 10208
rect 16684 10198 16712 11018
rect 16856 10464 16908 10470
rect 16856 10406 16908 10412
rect 16868 10198 16896 10406
rect 16672 10192 16724 10198
rect 16672 10134 16724 10140
rect 16856 10192 16908 10198
rect 16856 10134 16908 10140
rect 16488 9920 16540 9926
rect 16488 9862 16540 9868
rect 16500 8090 16528 9862
rect 16684 9654 16712 10134
rect 16868 9722 16896 10134
rect 16856 9716 16908 9722
rect 16856 9658 16908 9664
rect 16672 9648 16724 9654
rect 16672 9590 16724 9596
rect 17328 9042 17356 11834
rect 17696 11694 17724 12242
rect 18064 11830 18092 20810
rect 18524 20602 18552 21014
rect 18604 20800 18656 20806
rect 18604 20742 18656 20748
rect 18512 20596 18564 20602
rect 18512 20538 18564 20544
rect 18524 20058 18552 20538
rect 18616 20369 18644 20742
rect 18602 20360 18658 20369
rect 18602 20295 18658 20304
rect 18328 20052 18380 20058
rect 18328 19994 18380 20000
rect 18512 20052 18564 20058
rect 18512 19994 18564 20000
rect 18340 19242 18368 19994
rect 18800 19378 18828 27520
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 20180 23866 20208 27520
rect 21652 23866 21680 27520
rect 23032 23866 23060 27520
rect 20168 23860 20220 23866
rect 20168 23802 20220 23808
rect 21640 23860 21692 23866
rect 21640 23802 21692 23808
rect 23020 23860 23072 23866
rect 23020 23802 23072 23808
rect 22284 23792 22336 23798
rect 22284 23734 22336 23740
rect 19432 23588 19484 23594
rect 19432 23530 19484 23536
rect 19064 22024 19116 22030
rect 19064 21966 19116 21972
rect 18972 21412 19024 21418
rect 18972 21354 19024 21360
rect 18788 19372 18840 19378
rect 18788 19314 18840 19320
rect 18328 19236 18380 19242
rect 18328 19178 18380 19184
rect 18328 18624 18380 18630
rect 18328 18566 18380 18572
rect 18340 18426 18368 18566
rect 18984 18426 19012 21354
rect 19076 20398 19104 21966
rect 19248 21412 19300 21418
rect 19248 21354 19300 21360
rect 19260 21078 19288 21354
rect 19444 21350 19472 23530
rect 19984 23520 20036 23526
rect 19984 23462 20036 23468
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19432 21344 19484 21350
rect 19432 21286 19484 21292
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19248 21072 19300 21078
rect 19248 21014 19300 21020
rect 19996 20874 20024 23462
rect 20996 23180 21048 23186
rect 20996 23122 21048 23128
rect 21008 22778 21036 23122
rect 21180 22976 21232 22982
rect 21180 22918 21232 22924
rect 20996 22772 21048 22778
rect 20996 22714 21048 22720
rect 20352 21344 20404 21350
rect 20352 21286 20404 21292
rect 20076 21072 20128 21078
rect 20076 21014 20128 21020
rect 19984 20868 20036 20874
rect 19984 20810 20036 20816
rect 19430 20496 19486 20505
rect 19430 20431 19486 20440
rect 19064 20392 19116 20398
rect 19064 20334 19116 20340
rect 19076 18766 19104 20334
rect 19444 19922 19472 20431
rect 19524 20324 19576 20330
rect 19524 20266 19576 20272
rect 19536 20058 19564 20266
rect 19984 20256 20036 20262
rect 19984 20198 20036 20204
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19524 20052 19576 20058
rect 19524 19994 19576 20000
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 19444 19378 19472 19858
rect 19432 19372 19484 19378
rect 19432 19314 19484 19320
rect 19996 19242 20024 20198
rect 20088 19242 20116 21014
rect 20260 19712 20312 19718
rect 20260 19654 20312 19660
rect 20272 19378 20300 19654
rect 20260 19372 20312 19378
rect 20260 19314 20312 19320
rect 19984 19236 20036 19242
rect 19984 19178 20036 19184
rect 20076 19236 20128 19242
rect 20076 19178 20128 19184
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19340 18896 19392 18902
rect 19260 18856 19340 18884
rect 19064 18760 19116 18766
rect 19064 18702 19116 18708
rect 18328 18420 18380 18426
rect 18328 18362 18380 18368
rect 18972 18420 19024 18426
rect 18972 18362 19024 18368
rect 18340 15978 18368 18362
rect 18984 16250 19012 18362
rect 19260 18086 19288 18856
rect 19340 18838 19392 18844
rect 19524 18760 19576 18766
rect 19524 18702 19576 18708
rect 20076 18760 20128 18766
rect 20076 18702 20128 18708
rect 19248 18080 19300 18086
rect 19248 18022 19300 18028
rect 19260 16794 19288 18022
rect 19536 17542 19564 18702
rect 19984 18148 20036 18154
rect 19984 18090 20036 18096
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19996 17542 20024 18090
rect 19524 17536 19576 17542
rect 19524 17478 19576 17484
rect 19984 17536 20036 17542
rect 19984 17478 20036 17484
rect 19340 17128 19392 17134
rect 19340 17070 19392 17076
rect 19352 16794 19380 17070
rect 19248 16788 19300 16794
rect 19248 16730 19300 16736
rect 19340 16788 19392 16794
rect 19340 16730 19392 16736
rect 18972 16244 19024 16250
rect 18972 16186 19024 16192
rect 18604 16040 18656 16046
rect 18604 15982 18656 15988
rect 18328 15972 18380 15978
rect 18328 15914 18380 15920
rect 18340 15570 18368 15914
rect 18616 15609 18644 15982
rect 18984 15978 19012 16186
rect 19536 16182 19564 17478
rect 20088 17202 20116 18702
rect 20168 18420 20220 18426
rect 20168 18362 20220 18368
rect 20180 18154 20208 18362
rect 20168 18148 20220 18154
rect 20168 18090 20220 18096
rect 20260 17536 20312 17542
rect 20260 17478 20312 17484
rect 20076 17196 20128 17202
rect 20076 17138 20128 17144
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 20088 16658 20116 17138
rect 20076 16652 20128 16658
rect 20128 16612 20208 16640
rect 20076 16594 20128 16600
rect 19616 16448 19668 16454
rect 19616 16390 19668 16396
rect 20076 16448 20128 16454
rect 20076 16390 20128 16396
rect 19524 16176 19576 16182
rect 19524 16118 19576 16124
rect 19628 16114 19656 16390
rect 19616 16108 19668 16114
rect 19616 16050 19668 16056
rect 18972 15972 19024 15978
rect 18972 15914 19024 15920
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19524 15700 19576 15706
rect 19524 15642 19576 15648
rect 18602 15600 18658 15609
rect 18328 15564 18380 15570
rect 18602 15535 18658 15544
rect 18970 15600 19026 15609
rect 18970 15535 19026 15544
rect 18328 15506 18380 15512
rect 18788 15496 18840 15502
rect 18788 15438 18840 15444
rect 18800 15162 18828 15438
rect 18788 15156 18840 15162
rect 18788 15098 18840 15104
rect 18510 15056 18566 15065
rect 18510 14991 18566 15000
rect 18524 14958 18552 14991
rect 18512 14952 18564 14958
rect 18564 14912 18736 14940
rect 18512 14894 18564 14900
rect 18236 14816 18288 14822
rect 18236 14758 18288 14764
rect 18248 14618 18276 14758
rect 18236 14612 18288 14618
rect 18236 14554 18288 14560
rect 18248 13734 18276 14554
rect 18420 13796 18472 13802
rect 18340 13756 18420 13784
rect 18236 13728 18288 13734
rect 18340 13716 18368 13756
rect 18420 13738 18472 13744
rect 18288 13688 18368 13716
rect 18236 13670 18288 13676
rect 18340 13462 18368 13688
rect 18328 13456 18380 13462
rect 18328 13398 18380 13404
rect 18236 13320 18288 13326
rect 18236 13262 18288 13268
rect 18248 12714 18276 13262
rect 18340 12918 18368 13398
rect 18420 13320 18472 13326
rect 18420 13262 18472 13268
rect 18328 12912 18380 12918
rect 18328 12854 18380 12860
rect 18236 12708 18288 12714
rect 18236 12650 18288 12656
rect 18248 12345 18276 12650
rect 18340 12442 18368 12854
rect 18432 12782 18460 13262
rect 18604 12844 18656 12850
rect 18604 12786 18656 12792
rect 18420 12776 18472 12782
rect 18420 12718 18472 12724
rect 18328 12436 18380 12442
rect 18328 12378 18380 12384
rect 18234 12336 18290 12345
rect 18234 12271 18290 12280
rect 18328 12232 18380 12238
rect 18328 12174 18380 12180
rect 18052 11824 18104 11830
rect 18052 11766 18104 11772
rect 18340 11762 18368 12174
rect 18328 11756 18380 11762
rect 18328 11698 18380 11704
rect 17684 11688 17736 11694
rect 17684 11630 17736 11636
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 17420 9654 17448 10406
rect 17408 9648 17460 9654
rect 17408 9590 17460 9596
rect 17316 9036 17368 9042
rect 17316 8978 17368 8984
rect 17328 8634 17356 8978
rect 17316 8628 17368 8634
rect 17316 8570 17368 8576
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 16856 7948 16908 7954
rect 16856 7890 16908 7896
rect 16868 7478 16896 7890
rect 16856 7472 16908 7478
rect 16856 7414 16908 7420
rect 16948 7268 17000 7274
rect 16948 7210 17000 7216
rect 16856 6860 16908 6866
rect 16856 6802 16908 6808
rect 16868 6458 16896 6802
rect 16856 6452 16908 6458
rect 16856 6394 16908 6400
rect 16856 6180 16908 6186
rect 16856 6122 16908 6128
rect 16868 2961 16896 6122
rect 16854 2952 16910 2961
rect 16854 2887 16910 2896
rect 16764 2848 16816 2854
rect 16764 2790 16816 2796
rect 14832 2644 14884 2650
rect 14832 2586 14884 2592
rect 16396 2644 16448 2650
rect 16396 2586 16448 2592
rect 16672 2508 16724 2514
rect 16672 2450 16724 2456
rect 13360 2372 13412 2378
rect 13360 2314 13412 2320
rect 11978 54 12112 82
rect 13266 82 13322 480
rect 13372 82 13400 2314
rect 16684 2310 16712 2450
rect 14648 2304 14700 2310
rect 14648 2246 14700 2252
rect 16672 2304 16724 2310
rect 16672 2246 16724 2252
rect 13266 54 13400 82
rect 14554 82 14610 480
rect 14660 82 14688 2246
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 16684 1329 16712 2246
rect 16670 1320 16726 1329
rect 16670 1255 16726 1264
rect 14554 54 14688 82
rect 15750 128 15806 480
rect 15750 76 15752 128
rect 15804 76 15806 128
rect 8114 0 8170 54
rect 9402 0 9458 54
rect 10690 0 10746 54
rect 11978 0 12034 54
rect 13266 0 13322 54
rect 14554 0 14610 54
rect 15750 0 15806 76
rect 16776 82 16804 2790
rect 16960 2417 16988 7210
rect 16946 2408 17002 2417
rect 16946 2343 17002 2352
rect 17038 82 17094 480
rect 17420 134 17448 9590
rect 17696 9042 17724 11630
rect 17960 11212 18012 11218
rect 17960 11154 18012 11160
rect 17972 10538 18000 11154
rect 18144 11008 18196 11014
rect 18144 10950 18196 10956
rect 17960 10532 18012 10538
rect 17960 10474 18012 10480
rect 17972 10198 18000 10474
rect 18156 10470 18184 10950
rect 18616 10674 18644 12786
rect 18708 11898 18736 14912
rect 18788 13184 18840 13190
rect 18788 13126 18840 13132
rect 18800 12782 18828 13126
rect 18788 12776 18840 12782
rect 18788 12718 18840 12724
rect 18696 11892 18748 11898
rect 18696 11834 18748 11840
rect 18800 11694 18828 12718
rect 18788 11688 18840 11694
rect 18788 11630 18840 11636
rect 18696 11552 18748 11558
rect 18696 11494 18748 11500
rect 18708 11218 18736 11494
rect 18696 11212 18748 11218
rect 18696 11154 18748 11160
rect 18604 10668 18656 10674
rect 18604 10610 18656 10616
rect 18144 10464 18196 10470
rect 18144 10406 18196 10412
rect 17960 10192 18012 10198
rect 17960 10134 18012 10140
rect 17972 9586 18000 10134
rect 18604 10124 18656 10130
rect 18604 10066 18656 10072
rect 18420 10056 18472 10062
rect 18420 9998 18472 10004
rect 18432 9722 18460 9998
rect 18052 9716 18104 9722
rect 18052 9658 18104 9664
rect 18420 9716 18472 9722
rect 18420 9658 18472 9664
rect 17960 9580 18012 9586
rect 17960 9522 18012 9528
rect 17972 9178 18000 9522
rect 17960 9172 18012 9178
rect 17960 9114 18012 9120
rect 18064 9110 18092 9658
rect 18052 9104 18104 9110
rect 18052 9046 18104 9052
rect 17684 9036 17736 9042
rect 17684 8978 17736 8984
rect 17696 8566 17724 8978
rect 17684 8560 17736 8566
rect 17684 8502 17736 8508
rect 18512 8424 18564 8430
rect 18512 8366 18564 8372
rect 18524 8090 18552 8366
rect 18512 8084 18564 8090
rect 18512 8026 18564 8032
rect 18144 7744 18196 7750
rect 18144 7686 18196 7692
rect 18052 6656 18104 6662
rect 18052 6598 18104 6604
rect 18064 6254 18092 6598
rect 18052 6248 18104 6254
rect 18052 6190 18104 6196
rect 17684 2304 17736 2310
rect 17684 2246 17736 2252
rect 17696 1601 17724 2246
rect 17682 1592 17738 1601
rect 17682 1527 17738 1536
rect 16776 54 17094 82
rect 17408 128 17460 134
rect 17408 70 17460 76
rect 18156 82 18184 7686
rect 18616 7546 18644 10066
rect 18788 9580 18840 9586
rect 18788 9522 18840 9528
rect 18800 8838 18828 9522
rect 18788 8832 18840 8838
rect 18788 8774 18840 8780
rect 18800 8498 18828 8774
rect 18788 8492 18840 8498
rect 18788 8434 18840 8440
rect 18604 7540 18656 7546
rect 18604 7482 18656 7488
rect 18616 7342 18644 7482
rect 18604 7336 18656 7342
rect 18604 7278 18656 7284
rect 18604 7200 18656 7206
rect 18604 7142 18656 7148
rect 18236 6112 18288 6118
rect 18236 6054 18288 6060
rect 18248 474 18276 6054
rect 18616 5817 18644 7142
rect 18984 6186 19012 15535
rect 19064 15360 19116 15366
rect 19064 15302 19116 15308
rect 19076 15065 19104 15302
rect 19062 15056 19118 15065
rect 19062 14991 19118 15000
rect 19076 14958 19104 14991
rect 19064 14952 19116 14958
rect 19064 14894 19116 14900
rect 19536 14550 19564 15642
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19524 14544 19576 14550
rect 19524 14486 19576 14492
rect 19984 14340 20036 14346
rect 19984 14282 20036 14288
rect 19156 14272 19208 14278
rect 19156 14214 19208 14220
rect 19064 14000 19116 14006
rect 19064 13942 19116 13948
rect 19076 13705 19104 13942
rect 19168 13870 19196 14214
rect 19996 14074 20024 14282
rect 19984 14068 20036 14074
rect 19984 14010 20036 14016
rect 19432 13932 19484 13938
rect 19432 13874 19484 13880
rect 19156 13864 19208 13870
rect 19156 13806 19208 13812
rect 19062 13696 19118 13705
rect 19062 13631 19118 13640
rect 19168 13433 19196 13806
rect 19444 13734 19472 13874
rect 19432 13728 19484 13734
rect 19432 13670 19484 13676
rect 19524 13728 19576 13734
rect 19524 13670 19576 13676
rect 19536 13462 19564 13670
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19524 13456 19576 13462
rect 19154 13424 19210 13433
rect 19524 13398 19576 13404
rect 19154 13359 19210 13368
rect 19536 12646 19564 13398
rect 19984 13184 20036 13190
rect 19984 13126 20036 13132
rect 19996 12714 20024 13126
rect 20088 12986 20116 16390
rect 20180 16250 20208 16612
rect 20168 16244 20220 16250
rect 20168 16186 20220 16192
rect 20168 13728 20220 13734
rect 20168 13670 20220 13676
rect 20180 13530 20208 13670
rect 20168 13524 20220 13530
rect 20168 13466 20220 13472
rect 20076 12980 20128 12986
rect 20076 12922 20128 12928
rect 20076 12844 20128 12850
rect 20076 12786 20128 12792
rect 19984 12708 20036 12714
rect 19984 12650 20036 12656
rect 19524 12640 19576 12646
rect 19524 12582 19576 12588
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19432 12368 19484 12374
rect 19432 12310 19484 12316
rect 19156 12232 19208 12238
rect 19156 12174 19208 12180
rect 19168 11286 19196 12174
rect 19444 11558 19472 12310
rect 19432 11552 19484 11558
rect 19432 11494 19484 11500
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19996 11354 20024 12650
rect 20088 12374 20116 12786
rect 20076 12368 20128 12374
rect 20128 12328 20208 12356
rect 20076 12310 20128 12316
rect 20076 11688 20128 11694
rect 20076 11630 20128 11636
rect 19984 11348 20036 11354
rect 19984 11290 20036 11296
rect 20088 11286 20116 11630
rect 19156 11280 19208 11286
rect 19156 11222 19208 11228
rect 19800 11280 19852 11286
rect 19800 11222 19852 11228
rect 20076 11280 20128 11286
rect 20076 11222 20128 11228
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19340 10804 19392 10810
rect 19340 10746 19392 10752
rect 19352 10266 19380 10746
rect 19340 10260 19392 10266
rect 19340 10202 19392 10208
rect 19444 9994 19472 11086
rect 19812 10810 19840 11222
rect 19800 10804 19852 10810
rect 19800 10746 19852 10752
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 20076 10192 20128 10198
rect 20076 10134 20128 10140
rect 19432 9988 19484 9994
rect 19432 9930 19484 9936
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19800 9036 19852 9042
rect 19800 8978 19852 8984
rect 19812 8566 19840 8978
rect 19984 8832 20036 8838
rect 19984 8774 20036 8780
rect 19800 8560 19852 8566
rect 19800 8502 19852 8508
rect 19996 8498 20024 8774
rect 19984 8492 20036 8498
rect 19984 8434 20036 8440
rect 20088 8362 20116 10134
rect 20180 9654 20208 12328
rect 20168 9648 20220 9654
rect 20168 9590 20220 9596
rect 20180 9178 20208 9590
rect 20168 9172 20220 9178
rect 20168 9114 20220 9120
rect 20180 8498 20208 9114
rect 20168 8492 20220 8498
rect 20168 8434 20220 8440
rect 20076 8356 20128 8362
rect 20076 8298 20128 8304
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 20088 8090 20116 8298
rect 20076 8084 20128 8090
rect 20076 8026 20128 8032
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 18972 6180 19024 6186
rect 18972 6122 19024 6128
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 18602 5808 18658 5817
rect 18602 5743 18658 5752
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 20272 2650 20300 17478
rect 20364 12442 20392 21286
rect 20536 20528 20588 20534
rect 20536 20470 20588 20476
rect 20548 18358 20576 20470
rect 21192 20466 21220 22918
rect 21180 20460 21232 20466
rect 21180 20402 21232 20408
rect 20996 19916 21048 19922
rect 20996 19858 21048 19864
rect 21008 19446 21036 19858
rect 21364 19712 21416 19718
rect 21364 19654 21416 19660
rect 21824 19712 21876 19718
rect 21824 19654 21876 19660
rect 20996 19440 21048 19446
rect 20996 19382 21048 19388
rect 20812 19236 20864 19242
rect 20812 19178 20864 19184
rect 20536 18352 20588 18358
rect 20536 18294 20588 18300
rect 20548 17814 20576 18294
rect 20824 17814 20852 19178
rect 21008 19174 21036 19382
rect 21376 19310 21404 19654
rect 21836 19310 21864 19654
rect 21364 19304 21416 19310
rect 21364 19246 21416 19252
rect 21824 19304 21876 19310
rect 21824 19246 21876 19252
rect 20996 19168 21048 19174
rect 20996 19110 21048 19116
rect 20904 18828 20956 18834
rect 20904 18770 20956 18776
rect 20916 18426 20944 18770
rect 21008 18698 21036 19110
rect 21376 18873 21404 19246
rect 21456 19168 21508 19174
rect 21456 19110 21508 19116
rect 21468 18970 21496 19110
rect 21456 18964 21508 18970
rect 21456 18906 21508 18912
rect 21362 18864 21418 18873
rect 21180 18828 21232 18834
rect 21362 18799 21418 18808
rect 21180 18770 21232 18776
rect 20996 18692 21048 18698
rect 20996 18634 21048 18640
rect 20904 18420 20956 18426
rect 20904 18362 20956 18368
rect 20536 17808 20588 17814
rect 20536 17750 20588 17756
rect 20812 17808 20864 17814
rect 20812 17750 20864 17756
rect 20548 17066 20576 17750
rect 20536 17060 20588 17066
rect 20536 17002 20588 17008
rect 20824 16726 20852 17750
rect 20812 16720 20864 16726
rect 20812 16662 20864 16668
rect 20536 15428 20588 15434
rect 20536 15370 20588 15376
rect 20548 13802 20576 15370
rect 20916 14906 20944 18362
rect 21192 18086 21220 18770
rect 21836 18630 21864 19246
rect 21824 18624 21876 18630
rect 21824 18566 21876 18572
rect 21180 18080 21232 18086
rect 21180 18022 21232 18028
rect 21192 17649 21220 18022
rect 21456 17808 21508 17814
rect 21456 17750 21508 17756
rect 21272 17672 21324 17678
rect 21178 17640 21234 17649
rect 21272 17614 21324 17620
rect 21178 17575 21234 17584
rect 21192 16794 21220 17575
rect 21284 17202 21312 17614
rect 21468 17338 21496 17750
rect 21456 17332 21508 17338
rect 21456 17274 21508 17280
rect 21272 17196 21324 17202
rect 21272 17138 21324 17144
rect 21180 16788 21232 16794
rect 21180 16730 21232 16736
rect 21836 16658 21864 18566
rect 21088 16652 21140 16658
rect 21088 16594 21140 16600
rect 21364 16652 21416 16658
rect 21364 16594 21416 16600
rect 21824 16652 21876 16658
rect 21824 16594 21876 16600
rect 21100 15910 21128 16594
rect 21376 16250 21404 16594
rect 21364 16244 21416 16250
rect 21364 16186 21416 16192
rect 22192 16108 22244 16114
rect 22296 16096 22324 23734
rect 22560 23520 22612 23526
rect 22560 23462 22612 23468
rect 22468 17128 22520 17134
rect 22468 17070 22520 17076
rect 22480 16794 22508 17070
rect 22468 16788 22520 16794
rect 22468 16730 22520 16736
rect 22244 16068 22324 16096
rect 22192 16050 22244 16056
rect 21824 15972 21876 15978
rect 21824 15914 21876 15920
rect 21088 15904 21140 15910
rect 21088 15846 21140 15852
rect 20996 15496 21048 15502
rect 20996 15438 21048 15444
rect 20824 14878 20944 14906
rect 20720 14408 20772 14414
rect 20720 14350 20772 14356
rect 20536 13796 20588 13802
rect 20536 13738 20588 13744
rect 20442 13560 20498 13569
rect 20548 13530 20576 13738
rect 20442 13495 20498 13504
rect 20536 13524 20588 13530
rect 20456 13258 20484 13495
rect 20536 13466 20588 13472
rect 20444 13252 20496 13258
rect 20444 13194 20496 13200
rect 20548 12918 20576 13466
rect 20732 13258 20760 14350
rect 20824 13841 20852 14878
rect 20904 14816 20956 14822
rect 20904 14758 20956 14764
rect 20810 13832 20866 13841
rect 20810 13767 20866 13776
rect 20916 13530 20944 14758
rect 21008 14618 21036 15438
rect 20996 14612 21048 14618
rect 20996 14554 21048 14560
rect 20904 13524 20956 13530
rect 20904 13466 20956 13472
rect 21100 13326 21128 15846
rect 21836 15706 21864 15914
rect 22296 15706 22324 16068
rect 21824 15700 21876 15706
rect 21824 15642 21876 15648
rect 22284 15700 22336 15706
rect 22284 15642 22336 15648
rect 22572 15638 22600 23462
rect 24136 23186 24164 27526
rect 24398 27520 24454 27526
rect 25778 27520 25834 28000
rect 27158 27520 27214 28000
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 25134 24304 25190 24313
rect 25134 24239 25190 24248
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24124 23180 24176 23186
rect 24124 23122 24176 23128
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24766 22536 24822 22545
rect 24766 22471 24822 22480
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24780 21690 24808 22471
rect 24768 21684 24820 21690
rect 24768 21626 24820 21632
rect 23848 21480 23900 21486
rect 23848 21422 23900 21428
rect 23388 19372 23440 19378
rect 23388 19314 23440 19320
rect 23296 17060 23348 17066
rect 23296 17002 23348 17008
rect 22652 16652 22704 16658
rect 22652 16594 22704 16600
rect 22928 16652 22980 16658
rect 22928 16594 22980 16600
rect 22664 16250 22692 16594
rect 22940 16250 22968 16594
rect 22652 16244 22704 16250
rect 22652 16186 22704 16192
rect 22928 16244 22980 16250
rect 22928 16186 22980 16192
rect 22836 15972 22888 15978
rect 22836 15914 22888 15920
rect 21456 15632 21508 15638
rect 21456 15574 21508 15580
rect 22560 15632 22612 15638
rect 22560 15574 22612 15580
rect 22652 15632 22704 15638
rect 22652 15574 22704 15580
rect 21468 15094 21496 15574
rect 22572 15162 22600 15574
rect 22560 15156 22612 15162
rect 22560 15098 22612 15104
rect 21456 15088 21508 15094
rect 21456 15030 21508 15036
rect 21468 14890 21496 15030
rect 22664 15026 22692 15574
rect 22848 15502 22876 15914
rect 22836 15496 22888 15502
rect 22836 15438 22888 15444
rect 22744 15088 22796 15094
rect 22744 15030 22796 15036
rect 22652 15020 22704 15026
rect 22652 14962 22704 14968
rect 21456 14884 21508 14890
rect 21456 14826 21508 14832
rect 22560 14612 22612 14618
rect 22560 14554 22612 14560
rect 21456 14544 21508 14550
rect 21456 14486 21508 14492
rect 21180 14408 21232 14414
rect 21180 14350 21232 14356
rect 21192 13802 21220 14350
rect 21468 14074 21496 14486
rect 22468 14476 22520 14482
rect 22468 14418 22520 14424
rect 21824 14408 21876 14414
rect 21824 14350 21876 14356
rect 21456 14068 21508 14074
rect 21456 14010 21508 14016
rect 21180 13796 21232 13802
rect 21180 13738 21232 13744
rect 21192 13394 21220 13738
rect 21836 13734 21864 14350
rect 22284 14272 22336 14278
rect 22284 14214 22336 14220
rect 22296 13802 22324 14214
rect 22480 14006 22508 14418
rect 22468 14000 22520 14006
rect 22468 13942 22520 13948
rect 22100 13796 22152 13802
rect 22100 13738 22152 13744
rect 22284 13796 22336 13802
rect 22284 13738 22336 13744
rect 21824 13728 21876 13734
rect 21824 13670 21876 13676
rect 21180 13388 21232 13394
rect 21180 13330 21232 13336
rect 21088 13320 21140 13326
rect 21456 13320 21508 13326
rect 21088 13262 21140 13268
rect 21178 13288 21234 13297
rect 20720 13252 20772 13258
rect 21836 13297 21864 13670
rect 22112 13512 22140 13738
rect 22192 13524 22244 13530
rect 22112 13484 22192 13512
rect 22192 13466 22244 13472
rect 22296 13462 22324 13738
rect 22284 13456 22336 13462
rect 22572 13433 22600 14554
rect 22756 13870 22784 15030
rect 22744 13864 22796 13870
rect 22744 13806 22796 13812
rect 22848 13462 22876 15438
rect 23308 14074 23336 17002
rect 23296 14068 23348 14074
rect 23296 14010 23348 14016
rect 23308 13870 23336 14010
rect 23296 13864 23348 13870
rect 23296 13806 23348 13812
rect 22836 13456 22888 13462
rect 22284 13398 22336 13404
rect 22558 13424 22614 13433
rect 22008 13320 22060 13326
rect 21456 13262 21508 13268
rect 21822 13288 21878 13297
rect 21178 13223 21234 13232
rect 20720 13194 20772 13200
rect 20536 12912 20588 12918
rect 20536 12854 20588 12860
rect 21088 12640 21140 12646
rect 21088 12582 21140 12588
rect 20352 12436 20404 12442
rect 20352 12378 20404 12384
rect 21100 12374 21128 12582
rect 21088 12368 21140 12374
rect 21008 12328 21088 12356
rect 20352 11756 20404 11762
rect 20352 11698 20404 11704
rect 20364 11354 20392 11698
rect 20352 11348 20404 11354
rect 20352 11290 20404 11296
rect 21008 11014 21036 12328
rect 21088 12310 21140 12316
rect 21192 11830 21220 13223
rect 21272 12232 21324 12238
rect 21272 12174 21324 12180
rect 21180 11824 21232 11830
rect 21180 11766 21232 11772
rect 21284 11762 21312 12174
rect 21364 12096 21416 12102
rect 21364 12038 21416 12044
rect 21272 11756 21324 11762
rect 21272 11698 21324 11704
rect 21088 11620 21140 11626
rect 21088 11562 21140 11568
rect 21100 11286 21128 11562
rect 21088 11280 21140 11286
rect 21088 11222 21140 11228
rect 20996 11008 21048 11014
rect 20996 10950 21048 10956
rect 21100 10810 21128 11222
rect 21088 10804 21140 10810
rect 21088 10746 21140 10752
rect 21284 10674 21312 11698
rect 20444 10668 20496 10674
rect 20444 10610 20496 10616
rect 21272 10668 21324 10674
rect 21272 10610 21324 10616
rect 20456 10266 20484 10610
rect 20904 10532 20956 10538
rect 20904 10474 20956 10480
rect 20444 10260 20496 10266
rect 20444 10202 20496 10208
rect 20812 10124 20864 10130
rect 20916 10112 20944 10474
rect 20864 10084 20944 10112
rect 20812 10066 20864 10072
rect 20916 9586 20944 10084
rect 21284 10062 21312 10610
rect 20996 10056 21048 10062
rect 20996 9998 21048 10004
rect 21272 10056 21324 10062
rect 21272 9998 21324 10004
rect 21008 9722 21036 9998
rect 20996 9716 21048 9722
rect 20996 9658 21048 9664
rect 20904 9580 20956 9586
rect 20904 9522 20956 9528
rect 21008 9178 21036 9658
rect 20996 9172 21048 9178
rect 20996 9114 21048 9120
rect 20628 8560 20680 8566
rect 20628 8502 20680 8508
rect 20260 2644 20312 2650
rect 20260 2586 20312 2592
rect 18236 468 18288 474
rect 18236 410 18288 416
rect 18326 82 18382 480
rect 19340 468 19392 474
rect 19340 410 19392 416
rect 18156 54 18382 82
rect 19352 82 19380 410
rect 19614 82 19670 480
rect 19352 54 19670 82
rect 20640 82 20668 8502
rect 21376 2650 21404 12038
rect 21468 11762 21496 13262
rect 22008 13262 22060 13268
rect 21822 13223 21878 13232
rect 21548 13184 21600 13190
rect 21548 13126 21600 13132
rect 21560 12714 21588 13126
rect 21822 12744 21878 12753
rect 21548 12708 21600 12714
rect 21822 12679 21878 12688
rect 21548 12650 21600 12656
rect 21560 12442 21588 12650
rect 21548 12436 21600 12442
rect 21548 12378 21600 12384
rect 21456 11756 21508 11762
rect 21456 11698 21508 11704
rect 21836 11558 21864 12679
rect 22020 12102 22048 13262
rect 22296 12986 22324 13398
rect 22836 13398 22888 13404
rect 22558 13359 22614 13368
rect 22192 12980 22244 12986
rect 22192 12922 22244 12928
rect 22284 12980 22336 12986
rect 22284 12922 22336 12928
rect 22008 12096 22060 12102
rect 22008 12038 22060 12044
rect 21824 11552 21876 11558
rect 21824 11494 21876 11500
rect 21732 11144 21784 11150
rect 21732 11086 21784 11092
rect 21744 10810 21772 11086
rect 21732 10804 21784 10810
rect 21732 10746 21784 10752
rect 21640 10600 21692 10606
rect 21640 10542 21692 10548
rect 21456 10192 21508 10198
rect 21456 10134 21508 10140
rect 21468 9722 21496 10134
rect 21456 9716 21508 9722
rect 21456 9658 21508 9664
rect 21652 9489 21680 10542
rect 21638 9480 21694 9489
rect 21638 9415 21694 9424
rect 22204 9042 22232 12922
rect 22468 12300 22520 12306
rect 22468 12242 22520 12248
rect 22480 11898 22508 12242
rect 22468 11892 22520 11898
rect 22468 11834 22520 11840
rect 22744 11212 22796 11218
rect 22744 11154 22796 11160
rect 22756 10470 22784 11154
rect 22744 10464 22796 10470
rect 22744 10406 22796 10412
rect 22756 10169 22784 10406
rect 22742 10160 22798 10169
rect 22468 10124 22520 10130
rect 22742 10095 22798 10104
rect 22468 10066 22520 10072
rect 22480 9654 22508 10066
rect 22468 9648 22520 9654
rect 22468 9590 22520 9596
rect 22192 9036 22244 9042
rect 22192 8978 22244 8984
rect 22204 8634 22232 8978
rect 23400 8634 23428 19314
rect 23480 19236 23532 19242
rect 23480 19178 23532 19184
rect 23492 14890 23520 19178
rect 23662 18320 23718 18329
rect 23662 18255 23718 18264
rect 23480 14884 23532 14890
rect 23480 14826 23532 14832
rect 23676 14346 23704 18255
rect 23754 15056 23810 15065
rect 23754 14991 23810 15000
rect 23768 14822 23796 14991
rect 23756 14816 23808 14822
rect 23756 14758 23808 14764
rect 23664 14340 23716 14346
rect 23664 14282 23716 14288
rect 23478 13560 23534 13569
rect 23478 13495 23534 13504
rect 23492 13394 23520 13495
rect 23480 13388 23532 13394
rect 23480 13330 23532 13336
rect 23492 12986 23520 13330
rect 23480 12980 23532 12986
rect 23480 12922 23532 12928
rect 23676 12306 23704 14282
rect 23756 14272 23808 14278
rect 23756 14214 23808 14220
rect 23768 13530 23796 14214
rect 23756 13524 23808 13530
rect 23756 13466 23808 13472
rect 23664 12300 23716 12306
rect 23664 12242 23716 12248
rect 23676 11898 23704 12242
rect 23664 11892 23716 11898
rect 23664 11834 23716 11840
rect 22192 8628 22244 8634
rect 22192 8570 22244 8576
rect 23388 8628 23440 8634
rect 23388 8570 23440 8576
rect 23860 6458 23888 21422
rect 24766 21176 24822 21185
rect 24766 21111 24822 21120
rect 24676 21004 24728 21010
rect 24676 20946 24728 20952
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24688 20602 24716 20946
rect 24676 20596 24728 20602
rect 24676 20538 24728 20544
rect 24780 20058 24808 21111
rect 25148 21010 25176 24239
rect 25792 23594 25820 27520
rect 27172 23866 27200 27520
rect 27618 27296 27674 27305
rect 27618 27231 27674 27240
rect 27632 24886 27660 27231
rect 27620 24880 27672 24886
rect 27620 24822 27672 24828
rect 27160 23860 27212 23866
rect 27160 23802 27212 23808
rect 25780 23588 25832 23594
rect 25780 23530 25832 23536
rect 25136 21004 25188 21010
rect 25136 20946 25188 20952
rect 24768 20052 24820 20058
rect 24768 19994 24820 20000
rect 24676 19916 24728 19922
rect 24676 19858 24728 19864
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24688 19378 24716 19858
rect 24766 19816 24822 19825
rect 24766 19751 24822 19760
rect 24676 19372 24728 19378
rect 24676 19314 24728 19320
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24780 18426 24808 19751
rect 27620 18692 27672 18698
rect 27620 18634 27672 18640
rect 24768 18420 24820 18426
rect 24768 18362 24820 18368
rect 24216 18216 24268 18222
rect 24216 18158 24268 18164
rect 24228 17338 24256 18158
rect 27632 17513 27660 18634
rect 27618 17504 27674 17513
rect 24289 17436 24585 17456
rect 27618 17439 27674 17448
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24216 17332 24268 17338
rect 24216 17274 24268 17280
rect 24124 17128 24176 17134
rect 24124 17070 24176 17076
rect 24136 16017 24164 17070
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24122 16008 24178 16017
rect 24122 15943 24178 15952
rect 24766 15736 24822 15745
rect 24766 15671 24822 15680
rect 24676 15564 24728 15570
rect 24676 15506 24728 15512
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24688 15026 24716 15506
rect 24780 15434 24808 15671
rect 24768 15428 24820 15434
rect 24768 15370 24820 15376
rect 24676 15020 24728 15026
rect 24676 14962 24728 14968
rect 24124 14952 24176 14958
rect 24688 14929 24716 14962
rect 24124 14894 24176 14900
rect 24674 14920 24730 14929
rect 24136 14618 24164 14894
rect 24674 14855 24730 14864
rect 24124 14612 24176 14618
rect 24124 14554 24176 14560
rect 24136 13870 24164 14554
rect 24676 14476 24728 14482
rect 24676 14418 24728 14424
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24124 13864 24176 13870
rect 23952 13824 24124 13852
rect 23952 13394 23980 13824
rect 24124 13806 24176 13812
rect 24688 13802 24716 14418
rect 25410 14240 25466 14249
rect 25410 14175 25466 14184
rect 25424 14074 25452 14175
rect 25412 14068 25464 14074
rect 25412 14010 25464 14016
rect 24676 13796 24728 13802
rect 24676 13738 24728 13744
rect 23940 13388 23992 13394
rect 23940 13330 23992 13336
rect 23952 12986 23980 13330
rect 24032 13320 24084 13326
rect 24688 13297 24716 13738
rect 25136 13388 25188 13394
rect 25136 13330 25188 13336
rect 24032 13262 24084 13268
rect 24674 13288 24730 13297
rect 23940 12980 23992 12986
rect 23940 12922 23992 12928
rect 24044 12345 24072 13262
rect 24674 13223 24730 13232
rect 24676 13184 24728 13190
rect 24676 13126 24728 13132
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24688 12782 24716 13126
rect 24766 13016 24822 13025
rect 25148 12986 25176 13330
rect 24766 12951 24822 12960
rect 25136 12980 25188 12986
rect 24780 12918 24808 12951
rect 25136 12922 25188 12928
rect 24768 12912 24820 12918
rect 25148 12889 25176 12922
rect 24768 12854 24820 12860
rect 25134 12880 25190 12889
rect 25134 12815 25190 12824
rect 24676 12776 24728 12782
rect 24676 12718 24728 12724
rect 24688 12442 24716 12718
rect 24676 12436 24728 12442
rect 24676 12378 24728 12384
rect 24030 12336 24086 12345
rect 24030 12271 24086 12280
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24674 11384 24730 11393
rect 24674 11319 24730 11328
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24688 10130 24716 11319
rect 27620 10668 27672 10674
rect 27620 10610 27672 10616
rect 27632 10577 27660 10610
rect 27618 10568 27674 10577
rect 27618 10503 27674 10512
rect 24676 10124 24728 10130
rect 24676 10066 24728 10072
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24688 9722 24716 10066
rect 24676 9716 24728 9722
rect 24676 9658 24728 9664
rect 27620 9172 27672 9178
rect 27620 9114 27672 9120
rect 27632 9081 27660 9114
rect 27618 9072 27674 9081
rect 27618 9007 27674 9016
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24124 8424 24176 8430
rect 24124 8366 24176 8372
rect 24136 7313 24164 8366
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24122 7304 24178 7313
rect 24122 7239 24178 7248
rect 25136 7200 25188 7206
rect 24766 7168 24822 7177
rect 25136 7142 25188 7148
rect 24766 7103 24822 7112
rect 24780 7002 24808 7103
rect 24768 6996 24820 7002
rect 24768 6938 24820 6944
rect 25148 6905 25176 7142
rect 25134 6896 25190 6905
rect 24676 6860 24728 6866
rect 25134 6831 25190 6840
rect 24676 6802 24728 6808
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 23848 6452 23900 6458
rect 23848 6394 23900 6400
rect 24124 6248 24176 6254
rect 24124 6190 24176 6196
rect 24136 5681 24164 6190
rect 24688 6186 24716 6802
rect 24676 6180 24728 6186
rect 24676 6122 24728 6128
rect 24122 5672 24178 5681
rect 24122 5607 24178 5616
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 27618 4856 27674 4865
rect 27618 4791 27674 4800
rect 27632 4758 27660 4791
rect 27620 4752 27672 4758
rect 27620 4694 27672 4700
rect 24676 4684 24728 4690
rect 24676 4626 24728 4632
rect 21548 4480 21600 4486
rect 21548 4422 21600 4428
rect 21560 4010 21588 4422
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24688 4282 24716 4626
rect 24676 4276 24728 4282
rect 24676 4218 24728 4224
rect 21548 4004 21600 4010
rect 21548 3946 21600 3952
rect 23478 3632 23534 3641
rect 23478 3567 23534 3576
rect 24676 3596 24728 3602
rect 23112 3120 23164 3126
rect 23112 3062 23164 3068
rect 21364 2644 21416 2650
rect 21364 2586 21416 2592
rect 21824 2372 21876 2378
rect 21824 2314 21876 2320
rect 20902 82 20958 480
rect 20640 54 20958 82
rect 21836 82 21864 2314
rect 23124 2310 23152 3062
rect 23492 2689 23520 3567
rect 24676 3538 24728 3544
rect 27620 3596 27672 3602
rect 27620 3538 27672 3544
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24688 3194 24716 3538
rect 27632 3505 27660 3538
rect 27618 3496 27674 3505
rect 27618 3431 27674 3440
rect 24676 3188 24728 3194
rect 24676 3130 24728 3136
rect 23478 2680 23534 2689
rect 23478 2615 23534 2624
rect 24768 2576 24820 2582
rect 24768 2518 24820 2524
rect 23020 2304 23072 2310
rect 23020 2246 23072 2252
rect 23112 2304 23164 2310
rect 23112 2246 23164 2252
rect 22098 82 22154 480
rect 21836 54 22154 82
rect 23032 82 23060 2246
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 23386 82 23442 480
rect 23032 54 23442 82
rect 17038 0 17094 54
rect 18326 0 18382 54
rect 19614 0 19670 54
rect 20902 0 20958 54
rect 22098 0 22154 54
rect 23386 0 23442 54
rect 24674 82 24730 480
rect 24780 82 24808 2518
rect 25596 2304 25648 2310
rect 25596 2246 25648 2252
rect 24674 54 24808 82
rect 25608 82 25636 2246
rect 27342 1320 27398 1329
rect 27342 1255 27398 1264
rect 25962 82 26018 480
rect 25608 54 26018 82
rect 24674 0 24730 54
rect 25962 0 26018 54
rect 27250 82 27306 480
rect 27356 82 27384 1255
rect 27250 54 27384 82
rect 27250 0 27306 54
<< via2 >>
rect 1214 26832 1270 26888
rect 110 24520 166 24576
rect 1306 25336 1362 25392
rect 1214 22616 1270 22672
rect 1582 20032 1638 20088
rect 1306 18672 1362 18728
rect 110 13912 166 13968
rect 110 10104 166 10160
rect 110 9832 166 9888
rect 110 8472 166 8528
rect 1766 21528 1822 21584
rect 1306 15000 1362 15056
rect 938 14728 994 14784
rect 1306 12280 1362 12336
rect 2134 14476 2190 14512
rect 2134 14456 2136 14476
rect 2136 14456 2188 14476
rect 2188 14456 2190 14476
rect 3422 22616 3478 22672
rect 4066 21256 4122 21312
rect 2226 13232 2282 13288
rect 3422 13776 3478 13832
rect 1582 6704 1638 6760
rect 110 3168 166 3224
rect 3146 10104 3202 10160
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 6274 20440 6330 20496
rect 4158 13232 4214 13288
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5538 15952 5594 16008
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5446 14456 5502 14512
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 4066 7928 4122 7984
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 6274 9968 6330 10024
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 3146 5752 3202 5808
rect 2042 2216 2098 2272
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5446 5616 5502 5672
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 2778 856 2834 912
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 7194 17720 7250 17776
rect 7378 15544 7434 15600
rect 7102 14864 7158 14920
rect 7654 11464 7710 11520
rect 7930 16088 7986 16144
rect 8114 16088 8170 16144
rect 7930 12688 7986 12744
rect 9586 18128 9642 18184
rect 8942 13812 8944 13832
rect 8944 13812 8996 13832
rect 8996 13812 8998 13832
rect 8942 13776 8998 13812
rect 8850 12824 8906 12880
rect 7746 9424 7802 9480
rect 8666 6296 8722 6352
rect 6550 4936 6606 4992
rect 8390 2896 8446 2952
rect 7562 2352 7618 2408
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 11058 23024 11114 23080
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10690 9696 10746 9752
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 12162 22616 12218 22672
rect 11242 20440 11298 20496
rect 11794 20304 11850 20360
rect 11794 18828 11850 18864
rect 11794 18808 11796 18828
rect 11796 18808 11848 18828
rect 11848 18808 11850 18828
rect 11518 9968 11574 10024
rect 10966 5652 10968 5672
rect 10968 5652 11020 5672
rect 11020 5652 11022 5672
rect 10966 5616 11022 5652
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 11058 1536 11114 1592
rect 11702 7928 11758 7984
rect 12898 17584 12954 17640
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 13634 18808 13690 18864
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 16486 23704 16542 23760
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 18142 23024 18198 23080
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 17774 21528 17830 21584
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 13726 14456 13782 14512
rect 12806 7248 12862 7304
rect 12990 6296 13046 6352
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14278 14864 14334 14920
rect 14186 12824 14242 12880
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 15014 14456 15070 14512
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14922 12824 14978 12880
rect 15382 12688 15438 12744
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 16302 17720 16358 17776
rect 15566 13232 15622 13288
rect 15934 12688 15990 12744
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14738 9696 14794 9752
rect 14002 3576 14058 3632
rect 11334 176 11390 232
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 16486 16088 16542 16144
rect 17222 13640 17278 13696
rect 18602 20304 18658 20360
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19430 20440 19486 20496
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 18602 15544 18658 15600
rect 18970 15544 19026 15600
rect 18510 15000 18566 15056
rect 18234 12280 18290 12336
rect 16854 2896 16910 2952
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 16670 1264 16726 1320
rect 16946 2352 17002 2408
rect 17682 1536 17738 1592
rect 19062 15000 19118 15056
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19062 13640 19118 13696
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19154 13368 19210 13424
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 18602 5752 18658 5808
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 21362 18808 21418 18864
rect 21178 17584 21234 17640
rect 20442 13504 20498 13560
rect 20810 13776 20866 13832
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 25134 24248 25190 24304
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24766 22480 24822 22536
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 21178 13232 21234 13288
rect 21822 13232 21878 13288
rect 21822 12688 21878 12744
rect 22558 13368 22614 13424
rect 21638 9424 21694 9480
rect 22742 10104 22798 10160
rect 23662 18264 23718 18320
rect 23754 15000 23810 15056
rect 23478 13504 23534 13560
rect 24766 21120 24822 21176
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 27618 27240 27674 27296
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24766 19760 24822 19816
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 27618 17448 27674 17504
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24122 15952 24178 16008
rect 24766 15680 24822 15736
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24674 14864 24730 14920
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 25410 14184 25466 14240
rect 24674 13232 24730 13288
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24766 12960 24822 13016
rect 25134 12824 25190 12880
rect 24030 12280 24086 12336
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24674 11328 24730 11384
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 27618 10512 27674 10568
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 27618 9016 27674 9072
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24122 7248 24178 7304
rect 24766 7112 24822 7168
rect 25134 6840 25190 6896
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24122 5616 24178 5672
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 27618 4800 27674 4856
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 23478 3576 23534 3632
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 27618 3440 27674 3496
rect 23478 2624 23534 2680
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 27342 1264 27398 1320
<< metal3 >>
rect 0 27208 480 27328
rect 27520 27296 28000 27328
rect 27520 27240 27618 27296
rect 27674 27240 28000 27296
rect 27520 27208 28000 27240
rect 62 26890 122 27208
rect 1209 26890 1275 26893
rect 62 26888 1275 26890
rect 62 26832 1214 26888
rect 1270 26832 1275 26888
rect 62 26830 1275 26832
rect 1209 26827 1275 26830
rect 0 25848 480 25968
rect 27520 25940 28000 25968
rect 27520 25876 27660 25940
rect 27724 25876 28000 25940
rect 27520 25848 28000 25876
rect 62 25394 122 25848
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 1301 25394 1367 25397
rect 62 25392 1367 25394
rect 62 25336 1306 25392
rect 1362 25336 1367 25392
rect 62 25334 1367 25336
rect 1301 25331 1367 25334
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 0 24576 480 24608
rect 0 24520 110 24576
rect 166 24520 480 24576
rect 0 24488 480 24520
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 27520 24488 28000 24608
rect 19610 24447 19930 24448
rect 25129 24306 25195 24309
rect 27662 24306 27722 24488
rect 25129 24304 27722 24306
rect 25129 24248 25134 24304
rect 25190 24248 27722 24304
rect 25129 24246 27722 24248
rect 25129 24243 25195 24246
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 16481 23762 16547 23765
rect 27654 23762 27660 23764
rect 16481 23760 27660 23762
rect 16481 23704 16486 23760
rect 16542 23704 27660 23760
rect 16481 23702 27660 23704
rect 16481 23699 16547 23702
rect 27654 23700 27660 23702
rect 27724 23700 27730 23764
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 0 23128 480 23248
rect 62 22674 122 23128
rect 11053 23082 11119 23085
rect 18137 23082 18203 23085
rect 11053 23080 18203 23082
rect 11053 23024 11058 23080
rect 11114 23024 18142 23080
rect 18198 23024 18203 23080
rect 11053 23022 18203 23024
rect 11053 23019 11119 23022
rect 18137 23019 18203 23022
rect 27520 22992 28000 23112
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 1209 22674 1275 22677
rect 62 22672 1275 22674
rect 62 22616 1214 22672
rect 1270 22616 1275 22672
rect 62 22614 1275 22616
rect 1209 22611 1275 22614
rect 3417 22674 3483 22677
rect 12157 22674 12223 22677
rect 3417 22672 12223 22674
rect 3417 22616 3422 22672
rect 3478 22616 12162 22672
rect 12218 22616 12223 22672
rect 3417 22614 12223 22616
rect 3417 22611 3483 22614
rect 12157 22611 12223 22614
rect 24761 22538 24827 22541
rect 27662 22538 27722 22992
rect 24761 22536 27722 22538
rect 24761 22480 24766 22536
rect 24822 22480 27722 22536
rect 24761 22478 27722 22480
rect 24761 22475 24827 22478
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 0 21768 480 21888
rect 5610 21792 5930 21793
rect 62 21314 122 21768
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 27520 21632 28000 21752
rect 1761 21586 1827 21589
rect 17769 21586 17835 21589
rect 1761 21584 17835 21586
rect 1761 21528 1766 21584
rect 1822 21528 17774 21584
rect 17830 21528 17835 21584
rect 1761 21526 17835 21528
rect 1761 21523 1827 21526
rect 17769 21523 17835 21526
rect 4061 21314 4127 21317
rect 62 21312 4127 21314
rect 62 21256 4066 21312
rect 4122 21256 4127 21312
rect 62 21254 4127 21256
rect 4061 21251 4127 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 24761 21178 24827 21181
rect 27662 21178 27722 21632
rect 24761 21176 27722 21178
rect 24761 21120 24766 21176
rect 24822 21120 27722 21176
rect 24761 21118 27722 21120
rect 24761 21115 24827 21118
rect 5610 20704 5930 20705
rect 0 20544 480 20664
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 62 20090 122 20544
rect 6269 20498 6335 20501
rect 11237 20498 11303 20501
rect 19425 20498 19491 20501
rect 6269 20496 19491 20498
rect 6269 20440 6274 20496
rect 6330 20440 11242 20496
rect 11298 20440 19430 20496
rect 19486 20440 19491 20496
rect 6269 20438 19491 20440
rect 6269 20435 6335 20438
rect 11237 20435 11303 20438
rect 19425 20435 19491 20438
rect 11789 20362 11855 20365
rect 18597 20362 18663 20365
rect 11789 20360 18663 20362
rect 11789 20304 11794 20360
rect 11850 20304 18602 20360
rect 18658 20304 18663 20360
rect 11789 20302 18663 20304
rect 11789 20299 11855 20302
rect 18597 20299 18663 20302
rect 27520 20272 28000 20392
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 1577 20090 1643 20093
rect 62 20088 1643 20090
rect 62 20032 1582 20088
rect 1638 20032 1643 20088
rect 62 20030 1643 20032
rect 1577 20027 1643 20030
rect 24761 19818 24827 19821
rect 27662 19818 27722 20272
rect 24761 19816 27722 19818
rect 24761 19760 24766 19816
rect 24822 19760 27722 19816
rect 24761 19758 27722 19760
rect 24761 19755 24827 19758
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 0 19184 480 19304
rect 62 18730 122 19184
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 11789 18866 11855 18869
rect 13629 18866 13695 18869
rect 21357 18866 21423 18869
rect 11789 18864 21423 18866
rect 11789 18808 11794 18864
rect 11850 18808 13634 18864
rect 13690 18808 21362 18864
rect 21418 18808 21423 18864
rect 11789 18806 21423 18808
rect 11789 18803 11855 18806
rect 13629 18803 13695 18806
rect 21357 18803 21423 18806
rect 27520 18776 28000 18896
rect 1301 18730 1367 18733
rect 62 18728 1367 18730
rect 62 18672 1306 18728
rect 1362 18672 1367 18728
rect 62 18670 1367 18672
rect 1301 18667 1367 18670
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 23657 18322 23723 18325
rect 27662 18322 27722 18776
rect 23657 18320 27722 18322
rect 23657 18264 23662 18320
rect 23718 18264 27722 18320
rect 23657 18262 27722 18264
rect 23657 18259 23723 18262
rect 9581 18186 9647 18189
rect 62 18184 9647 18186
rect 62 18128 9586 18184
rect 9642 18128 9647 18184
rect 62 18126 9647 18128
rect 62 17944 122 18126
rect 9581 18123 9647 18126
rect 10277 17984 10597 17985
rect 0 17824 480 17944
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 7189 17778 7255 17781
rect 16297 17778 16363 17781
rect 7189 17776 16363 17778
rect 7189 17720 7194 17776
rect 7250 17720 16302 17776
rect 16358 17720 16363 17776
rect 7189 17718 16363 17720
rect 7189 17715 7255 17718
rect 16297 17715 16363 17718
rect 12893 17642 12959 17645
rect 21173 17642 21239 17645
rect 12893 17640 21239 17642
rect 12893 17584 12898 17640
rect 12954 17584 21178 17640
rect 21234 17584 21239 17640
rect 12893 17582 21239 17584
rect 12893 17579 12959 17582
rect 21173 17579 21239 17582
rect 27520 17504 28000 17536
rect 27520 17448 27618 17504
rect 27674 17448 28000 17504
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 27520 17416 28000 17448
rect 24277 17375 24597 17376
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 0 16464 480 16584
rect 62 16146 122 16464
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 7925 16146 7991 16149
rect 62 16144 7991 16146
rect 62 16088 7930 16144
rect 7986 16088 7991 16144
rect 62 16086 7991 16088
rect 7925 16083 7991 16086
rect 8109 16146 8175 16149
rect 16481 16146 16547 16149
rect 8109 16144 16547 16146
rect 8109 16088 8114 16144
rect 8170 16088 16486 16144
rect 16542 16088 16547 16144
rect 8109 16086 16547 16088
rect 8109 16083 8175 16086
rect 16481 16083 16547 16086
rect 27520 16056 28000 16176
rect 5533 16010 5599 16013
rect 24117 16010 24183 16013
rect 5533 16008 24183 16010
rect 5533 15952 5538 16008
rect 5594 15952 24122 16008
rect 24178 15952 24183 16008
rect 5533 15950 24183 15952
rect 5533 15947 5599 15950
rect 24117 15947 24183 15950
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 24761 15738 24827 15741
rect 27662 15738 27722 16056
rect 24761 15736 27722 15738
rect 24761 15680 24766 15736
rect 24822 15680 27722 15736
rect 24761 15678 27722 15680
rect 24761 15675 24827 15678
rect 7373 15602 7439 15605
rect 18597 15602 18663 15605
rect 18965 15602 19031 15605
rect 7373 15600 19031 15602
rect 7373 15544 7378 15600
rect 7434 15544 18602 15600
rect 18658 15544 18970 15600
rect 19026 15544 19031 15600
rect 7373 15542 19031 15544
rect 7373 15539 7439 15542
rect 18597 15539 18663 15542
rect 18965 15539 19031 15542
rect 5610 15264 5930 15265
rect 0 15104 480 15224
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 62 14786 122 15104
rect 1301 15058 1367 15061
rect 18505 15058 18571 15061
rect 1301 15056 18571 15058
rect 1301 15000 1306 15056
rect 1362 15000 18510 15056
rect 18566 15000 18571 15056
rect 1301 14998 18571 15000
rect 1301 14995 1367 14998
rect 18505 14995 18571 14998
rect 19057 15058 19123 15061
rect 23749 15058 23815 15061
rect 19057 15056 23815 15058
rect 19057 15000 19062 15056
rect 19118 15000 23754 15056
rect 23810 15000 23815 15056
rect 19057 14998 23815 15000
rect 19057 14995 19123 14998
rect 23749 14995 23815 14998
rect 7097 14922 7163 14925
rect 14273 14922 14339 14925
rect 24669 14922 24735 14925
rect 7097 14920 24735 14922
rect 7097 14864 7102 14920
rect 7158 14864 14278 14920
rect 14334 14864 24674 14920
rect 24730 14864 24735 14920
rect 7097 14862 24735 14864
rect 7097 14859 7163 14862
rect 14273 14859 14339 14862
rect 24669 14859 24735 14862
rect 933 14786 999 14789
rect 62 14784 999 14786
rect 62 14728 938 14784
rect 994 14728 999 14784
rect 62 14726 999 14728
rect 933 14723 999 14726
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 27520 14696 28000 14816
rect 19610 14655 19930 14656
rect 2129 14514 2195 14517
rect 5441 14514 5507 14517
rect 13721 14514 13787 14517
rect 15009 14514 15075 14517
rect 2129 14512 15075 14514
rect 2129 14456 2134 14512
rect 2190 14456 5446 14512
rect 5502 14456 13726 14512
rect 13782 14456 15014 14512
rect 15070 14456 15075 14512
rect 2129 14454 15075 14456
rect 2129 14451 2195 14454
rect 5441 14451 5507 14454
rect 13721 14451 13787 14454
rect 15009 14451 15075 14454
rect 25405 14242 25471 14245
rect 27662 14242 27722 14696
rect 25405 14240 27722 14242
rect 25405 14184 25410 14240
rect 25466 14184 27722 14240
rect 25405 14182 27722 14184
rect 25405 14179 25471 14182
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 0 13968 480 14000
rect 0 13912 110 13968
rect 166 13912 480 13968
rect 0 13880 480 13912
rect 3417 13834 3483 13837
rect 8937 13834 9003 13837
rect 20805 13834 20871 13837
rect 3417 13832 9003 13834
rect 3417 13776 3422 13832
rect 3478 13776 8942 13832
rect 8998 13776 9003 13832
rect 3417 13774 9003 13776
rect 3417 13771 3483 13774
rect 8937 13771 9003 13774
rect 20164 13832 20871 13834
rect 20164 13776 20810 13832
rect 20866 13776 20871 13832
rect 20164 13774 20871 13776
rect 17217 13698 17283 13701
rect 19057 13698 19123 13701
rect 17217 13696 19123 13698
rect 17217 13640 17222 13696
rect 17278 13640 19062 13696
rect 19118 13640 19123 13696
rect 17217 13638 19123 13640
rect 17217 13635 17283 13638
rect 19057 13635 19123 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 20164 13562 20224 13774
rect 20805 13771 20871 13774
rect 20437 13562 20503 13565
rect 23473 13562 23539 13565
rect 20164 13560 23539 13562
rect 20164 13504 20442 13560
rect 20498 13504 23478 13560
rect 23534 13504 23539 13560
rect 20164 13502 23539 13504
rect 20437 13499 20503 13502
rect 23473 13499 23539 13502
rect 19149 13426 19215 13429
rect 22553 13426 22619 13429
rect 19149 13424 22619 13426
rect 19149 13368 19154 13424
rect 19210 13368 22558 13424
rect 22614 13368 22619 13424
rect 19149 13366 22619 13368
rect 19149 13363 19215 13366
rect 22553 13363 22619 13366
rect 2221 13290 2287 13293
rect 4153 13292 4219 13293
rect 4102 13290 4108 13292
rect 2221 13288 4108 13290
rect 4172 13288 4219 13292
rect 2221 13232 2226 13288
rect 2282 13232 4108 13288
rect 4214 13232 4219 13288
rect 2221 13230 4108 13232
rect 2221 13227 2287 13230
rect 4102 13228 4108 13230
rect 4172 13228 4219 13232
rect 4153 13227 4219 13228
rect 15561 13290 15627 13293
rect 21173 13290 21239 13293
rect 21817 13290 21883 13293
rect 15561 13288 21883 13290
rect 15561 13232 15566 13288
rect 15622 13232 21178 13288
rect 21234 13232 21822 13288
rect 21878 13232 21883 13288
rect 15561 13230 21883 13232
rect 15561 13227 15627 13230
rect 21173 13227 21239 13230
rect 21817 13227 21883 13230
rect 23422 13228 23428 13292
rect 23492 13290 23498 13292
rect 24669 13290 24735 13293
rect 23492 13288 24735 13290
rect 23492 13232 24674 13288
rect 24730 13232 24735 13288
rect 23492 13230 24735 13232
rect 23492 13228 23498 13230
rect 24669 13227 24735 13230
rect 27520 13200 28000 13320
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 24761 13018 24827 13021
rect 27662 13018 27722 13200
rect 24761 13016 27722 13018
rect 24761 12960 24766 13016
rect 24822 12960 27722 13016
rect 24761 12958 27722 12960
rect 24761 12955 24827 12958
rect 8845 12882 8911 12885
rect 14181 12882 14247 12885
rect 8845 12880 14247 12882
rect 8845 12824 8850 12880
rect 8906 12824 14186 12880
rect 14242 12824 14247 12880
rect 8845 12822 14247 12824
rect 8845 12819 8911 12822
rect 14181 12819 14247 12822
rect 14917 12882 14983 12885
rect 25129 12882 25195 12885
rect 14917 12880 25195 12882
rect 14917 12824 14922 12880
rect 14978 12824 25134 12880
rect 25190 12824 25195 12880
rect 14917 12822 25195 12824
rect 14917 12819 14983 12822
rect 25129 12819 25195 12822
rect 7925 12746 7991 12749
rect 15377 12746 15443 12749
rect 7925 12744 15443 12746
rect 7925 12688 7930 12744
rect 7986 12688 15382 12744
rect 15438 12688 15443 12744
rect 7925 12686 15443 12688
rect 7925 12683 7991 12686
rect 15377 12683 15443 12686
rect 15929 12746 15995 12749
rect 21817 12746 21883 12749
rect 15929 12744 21883 12746
rect 15929 12688 15934 12744
rect 15990 12688 21822 12744
rect 21878 12688 21883 12744
rect 15929 12686 21883 12688
rect 15929 12683 15995 12686
rect 21817 12683 21883 12686
rect 0 12612 480 12640
rect 0 12548 60 12612
rect 124 12548 480 12612
rect 0 12520 480 12548
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 54 12276 60 12340
rect 124 12338 130 12340
rect 1301 12338 1367 12341
rect 124 12336 1367 12338
rect 124 12280 1306 12336
rect 1362 12280 1367 12336
rect 124 12278 1367 12280
rect 124 12276 130 12278
rect 1301 12275 1367 12278
rect 18229 12338 18295 12341
rect 24025 12338 24091 12341
rect 18229 12336 24091 12338
rect 18229 12280 18234 12336
rect 18290 12280 24030 12336
rect 24086 12280 24091 12336
rect 18229 12278 24091 12280
rect 18229 12275 18295 12278
rect 24025 12275 24091 12278
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 27520 11840 28000 11960
rect 7649 11522 7715 11525
rect 62 11520 7715 11522
rect 62 11464 7654 11520
rect 7710 11464 7715 11520
rect 62 11462 7715 11464
rect 62 11280 122 11462
rect 7649 11459 7715 11462
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 24669 11386 24735 11389
rect 27662 11386 27722 11840
rect 24669 11384 27722 11386
rect 24669 11328 24674 11384
rect 24730 11328 27722 11384
rect 24669 11326 27722 11328
rect 24669 11323 24735 11326
rect 0 11160 480 11280
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 27520 10568 28000 10600
rect 27520 10512 27618 10568
rect 27674 10512 28000 10568
rect 27520 10480 28000 10512
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 105 10162 171 10165
rect 3141 10162 3207 10165
rect 22737 10162 22803 10165
rect 105 10160 3066 10162
rect 105 10104 110 10160
rect 166 10104 3066 10160
rect 105 10102 3066 10104
rect 105 10099 171 10102
rect 3006 10026 3066 10102
rect 3141 10160 22803 10162
rect 3141 10104 3146 10160
rect 3202 10104 22742 10160
rect 22798 10104 22803 10160
rect 3141 10102 22803 10104
rect 3141 10099 3207 10102
rect 22737 10099 22803 10102
rect 6269 10026 6335 10029
rect 11513 10026 11579 10029
rect 3006 10024 11579 10026
rect 3006 9968 6274 10024
rect 6330 9968 11518 10024
rect 11574 9968 11579 10024
rect 3006 9966 11579 9968
rect 6269 9963 6335 9966
rect 11513 9963 11579 9966
rect 0 9888 480 9920
rect 0 9832 110 9888
rect 166 9832 480 9888
rect 0 9800 480 9832
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 10685 9754 10751 9757
rect 14733 9754 14799 9757
rect 10685 9752 14799 9754
rect 10685 9696 10690 9752
rect 10746 9696 14738 9752
rect 14794 9696 14799 9752
rect 10685 9694 14799 9696
rect 10685 9691 10751 9694
rect 14733 9691 14799 9694
rect 7741 9482 7807 9485
rect 21633 9482 21699 9485
rect 7741 9480 21699 9482
rect 7741 9424 7746 9480
rect 7802 9424 21638 9480
rect 21694 9424 21699 9480
rect 7741 9422 21699 9424
rect 7741 9419 7807 9422
rect 21633 9419 21699 9422
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 27520 9072 28000 9104
rect 27520 9016 27618 9072
rect 27674 9016 28000 9072
rect 27520 8984 28000 9016
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 0 8528 480 8560
rect 0 8472 110 8528
rect 166 8472 480 8528
rect 0 8440 480 8472
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 4061 7986 4127 7989
rect 11697 7986 11763 7989
rect 4061 7984 11763 7986
rect 4061 7928 4066 7984
rect 4122 7928 11702 7984
rect 11758 7928 11763 7984
rect 4061 7926 11763 7928
rect 4061 7923 4127 7926
rect 11697 7923 11763 7926
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 27520 7624 28000 7744
rect 24277 7583 24597 7584
rect 0 7216 480 7336
rect 12801 7306 12867 7309
rect 24117 7306 24183 7309
rect 12801 7304 24183 7306
rect 12801 7248 12806 7304
rect 12862 7248 24122 7304
rect 24178 7248 24183 7304
rect 12801 7246 24183 7248
rect 12801 7243 12867 7246
rect 24117 7243 24183 7246
rect 62 6762 122 7216
rect 24761 7170 24827 7173
rect 27662 7170 27722 7624
rect 24761 7168 27722 7170
rect 24761 7112 24766 7168
rect 24822 7112 27722 7168
rect 24761 7110 27722 7112
rect 24761 7107 24827 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 25129 6898 25195 6901
rect 25129 6896 27722 6898
rect 25129 6840 25134 6896
rect 25190 6840 27722 6896
rect 25129 6838 27722 6840
rect 25129 6835 25195 6838
rect 1577 6762 1643 6765
rect 62 6760 1643 6762
rect 62 6704 1582 6760
rect 1638 6704 1643 6760
rect 62 6702 1643 6704
rect 1577 6699 1643 6702
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 27662 6384 27722 6838
rect 8661 6354 8727 6357
rect 12985 6354 13051 6357
rect 8661 6352 13051 6354
rect 8661 6296 8666 6352
rect 8722 6296 12990 6352
rect 13046 6296 13051 6352
rect 8661 6294 13051 6296
rect 8661 6291 8727 6294
rect 12985 6291 13051 6294
rect 27520 6264 28000 6384
rect 10277 6016 10597 6017
rect 0 5856 480 5976
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 62 5674 122 5856
rect 3141 5810 3207 5813
rect 18597 5810 18663 5813
rect 3141 5808 18663 5810
rect 3141 5752 3146 5808
rect 3202 5752 18602 5808
rect 18658 5752 18663 5808
rect 3141 5750 18663 5752
rect 3141 5747 3207 5750
rect 18597 5747 18663 5750
rect 5441 5674 5507 5677
rect 62 5672 5507 5674
rect 62 5616 5446 5672
rect 5502 5616 5507 5672
rect 62 5614 5507 5616
rect 5441 5611 5507 5614
rect 10961 5674 11027 5677
rect 24117 5674 24183 5677
rect 10961 5672 24183 5674
rect 10961 5616 10966 5672
rect 11022 5616 24122 5672
rect 24178 5616 24183 5672
rect 10961 5614 24183 5616
rect 10961 5611 11027 5614
rect 24117 5611 24183 5614
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 6545 4994 6611 4997
rect 62 4992 6611 4994
rect 62 4936 6550 4992
rect 6606 4936 6611 4992
rect 62 4934 6611 4936
rect 62 4616 122 4934
rect 6545 4931 6611 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 27520 4856 28000 4888
rect 27520 4800 27618 4856
rect 27674 4800 28000 4856
rect 27520 4768 28000 4800
rect 0 4496 480 4616
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 13997 3634 14063 3637
rect 23473 3634 23539 3637
rect 13997 3632 23539 3634
rect 13997 3576 14002 3632
rect 14058 3576 23478 3632
rect 23534 3576 23539 3632
rect 13997 3574 23539 3576
rect 13997 3571 14063 3574
rect 23473 3571 23539 3574
rect 27520 3496 28000 3528
rect 27520 3440 27618 3496
rect 27674 3440 28000 3496
rect 27520 3408 28000 3440
rect 5610 3296 5930 3297
rect 0 3224 480 3256
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 0 3168 110 3224
rect 166 3168 480 3224
rect 0 3136 480 3168
rect 8385 2954 8451 2957
rect 16849 2954 16915 2957
rect 8385 2952 16915 2954
rect 8385 2896 8390 2952
rect 8446 2896 16854 2952
rect 16910 2896 16915 2952
rect 8385 2894 16915 2896
rect 8385 2891 8451 2894
rect 16849 2891 16915 2894
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 23473 2682 23539 2685
rect 23473 2680 27722 2682
rect 23473 2624 23478 2680
rect 23534 2624 27722 2680
rect 23473 2622 27722 2624
rect 23473 2619 23539 2622
rect 7557 2410 7623 2413
rect 16941 2410 17007 2413
rect 7557 2408 17007 2410
rect 7557 2352 7562 2408
rect 7618 2352 16946 2408
rect 17002 2352 17007 2408
rect 7557 2350 17007 2352
rect 7557 2347 7623 2350
rect 16941 2347 17007 2350
rect 2037 2274 2103 2277
rect 62 2272 2103 2274
rect 62 2216 2042 2272
rect 2098 2216 2103 2272
rect 62 2214 2103 2216
rect 62 1896 122 2214
rect 2037 2211 2103 2214
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 27662 2168 27722 2622
rect 24277 2143 24597 2144
rect 27520 2048 28000 2168
rect 0 1776 480 1896
rect 11053 1594 11119 1597
rect 17677 1594 17743 1597
rect 11053 1592 17743 1594
rect 11053 1536 11058 1592
rect 11114 1536 17682 1592
rect 17738 1536 17743 1592
rect 11053 1534 17743 1536
rect 11053 1531 11119 1534
rect 17677 1531 17743 1534
rect 16665 1322 16731 1325
rect 27337 1322 27403 1325
rect 16665 1320 27403 1322
rect 16665 1264 16670 1320
rect 16726 1264 27342 1320
rect 27398 1264 27403 1320
rect 16665 1262 27403 1264
rect 16665 1259 16731 1262
rect 27337 1259 27403 1262
rect 2773 914 2839 917
rect 62 912 2839 914
rect 62 856 2778 912
rect 2834 856 2839 912
rect 62 854 2839 856
rect 62 672 122 854
rect 2773 851 2839 854
rect 27520 688 28000 808
rect 0 552 480 672
rect 11329 234 11395 237
rect 27662 234 27722 688
rect 11329 232 27722 234
rect 11329 176 11334 232
rect 11390 176 27722 232
rect 11329 174 27722 176
rect 11329 171 11395 174
<< via3 >>
rect 27660 25876 27724 25940
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 27660 23700 27724 23764
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 4108 13288 4172 13292
rect 4108 13232 4158 13288
rect 4158 13232 4172 13288
rect 4108 13228 4172 13232
rect 23428 13228 23492 13292
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 60 12548 124 12612
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 60 12276 124 12340
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 27659 25940 27725 25941
rect 27659 25876 27660 25940
rect 27724 25876 27725 25940
rect 27659 25875 27725 25876
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 59 12612 125 12613
rect 59 12548 60 12612
rect 124 12548 125 12612
rect 59 12547 125 12548
rect 62 12341 122 12547
rect 59 12340 125 12341
rect 59 12276 60 12340
rect 124 12276 125 12340
rect 59 12275 125 12276
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 27662 23765 27722 25875
rect 27659 23764 27725 23765
rect 27659 23700 27660 23764
rect 27724 23700 27725 23764
rect 27659 23699 27725 23700
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
<< via4 >>
rect 4022 13292 4258 13378
rect 4022 13228 4108 13292
rect 4108 13228 4172 13292
rect 4172 13228 4258 13292
rect 4022 13142 4258 13228
rect 23342 13292 23578 13378
rect 23342 13228 23428 13292
rect 23428 13228 23492 13292
rect 23492 13228 23578 13292
rect 23342 13142 23578 13228
<< metal5 >>
rect 3980 13378 23620 13420
rect 3980 13142 4022 13378
rect 4258 13142 23342 13378
rect 23578 13142 23620 13378
rect 3980 13100 23620 13142
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1564 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_7
timestamp 1586364061
transform 1 0 1748 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_19
timestamp 1586364061
transform 1 0 2852 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_31
timestamp 1586364061
transform 1 0 3956 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_43
timestamp 1586364061
transform 1 0 5060 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _228_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__228__A
timestamp 1586364061
transform 1 0 7452 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_67
timestamp 1586364061
transform 1 0 7268 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_71
timestamp 1586364061
transform 1 0 7636 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_1_55
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _236_
timestamp 1586364061
transform 1 0 9108 0 1 2720
box -38 -48 406 592
use scs8hd_decap_8  FILLER_0_83 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8740 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_1_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 130 592
use scs8hd_buf_2  _235_
timestamp 1586364061
transform 1 0 10764 0 1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__236__A
timestamp 1586364061
transform 1 0 9660 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_91
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_91
timestamp 1586364061
transform 1 0 9476 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_1_95
timestamp 1586364061
transform 1 0 9844 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_103
timestamp 1586364061
transform 1 0 10580 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_1_113
timestamp 1586364061
transform 1 0 11500 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_109
timestamp 1586364061
transform 1 0 11132 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_113
timestamp 1586364061
transform 1 0 11500 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__232__A
timestamp 1586364061
transform 1 0 11684 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__235__A
timestamp 1586364061
transform 1 0 11316 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _232_
timestamp 1586364061
transform 1 0 11132 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_121
timestamp 1586364061
transform 1 0 12236 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_123
timestamp 1586364061
transform 1 0 12420 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_117
timestamp 1586364061
transform 1 0 11868 0 -1 2720
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_147
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__229__A
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _229_
timestamp 1586364061
transform 1 0 14260 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_156
timestamp 1586364061
transform 1 0 15456 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_153
timestamp 1586364061
transform 1 0 15180 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_4  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _246_
timestamp 1586364061
transform 1 0 15640 0 1 2720
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_2_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 16100 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__246__A
timestamp 1586364061
transform 1 0 16192 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_162
timestamp 1586364061
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_166
timestamp 1586364061
transform 1 0 16376 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_170
timestamp 1586364061
transform 1 0 16744 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_162
timestamp 1586364061
transform 1 0 16008 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_166
timestamp 1586364061
transform 1 0 16376 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_178
timestamp 1586364061
transform 1 0 17480 0 1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_1_182
timestamp 1586364061
transform 1 0 17848 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20056 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_0_205
timestamp 1586364061
transform 1 0 19964 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_209
timestamp 1586364061
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21528 0 -1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21988 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_225
timestamp 1586364061
transform 1 0 21804 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_229
timestamp 1586364061
transform 1 0 22172 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_0_237
timestamp 1586364061
transform 1 0 22908 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_233
timestamp 1586364061
transform 1 0 22540 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23092 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22632 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 774 592
use scs8hd_fill_1  FILLER_0_247
timestamp 1586364061
transform 1 0 23828 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_241
timestamp 1586364061
transform 1 0 23276 0 -1 2720
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24472 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_252
timestamp 1586364061
transform 1 0 24288 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_256
timestamp 1586364061
transform 1 0 24656 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_253
timestamp 1586364061
transform 1 0 24380 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_257
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_0_268
timestamp 1586364061
transform 1 0 25760 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_1  FILLER_0_276
timestamp 1586364061
transform 1 0 26496 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_6
timestamp 1586364061
transform 1 0 1656 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_18
timestamp 1586364061
transform 1 0 2760 0 -1 3808
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_2_30
timestamp 1586364061
transform 1 0 3864 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_70
timestamp 1586364061
transform 1 0 7544 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_2_82
timestamp 1586364061
transform 1 0 8648 0 -1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_90
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14168 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_2_135
timestamp 1586364061
transform 1 0 13524 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_138
timestamp 1586364061
transform 1 0 13800 0 -1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_144
timestamp 1586364061
transform 1 0 14352 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_152
timestamp 1586364061
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_157
timestamp 1586364061
transform 1 0 15548 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_169
timestamp 1586364061
transform 1 0 16652 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_181
timestamp 1586364061
transform 1 0 17756 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_193
timestamp 1586364061
transform 1 0 18860 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_205
timestamp 1586364061
transform 1 0 19964 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_213
timestamp 1586364061
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_258
timestamp 1586364061
transform 1 0 24840 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_270
timestamp 1586364061
transform 1 0 25944 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_274
timestamp 1586364061
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 1564 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_7
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_19
timestamp 1586364061
transform 1 0 2852 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_31
timestamp 1586364061
transform 1 0 3956 0 1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5704 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_43
timestamp 1586364061
transform 1 0 5060 0 1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_3_49
timestamp 1586364061
transform 1 0 5612 0 1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_3_52
timestamp 1586364061
transform 1 0 5888 0 1 3808
box -38 -48 590 592
use scs8hd_inv_8  _204_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6900 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_58
timestamp 1586364061
transform 1 0 6440 0 1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9108 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_72
timestamp 1586364061
transform 1 0 7728 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_76
timestamp 1586364061
transform 1 0 8096 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_3_84
timestamp 1586364061
transform 1 0 8832 0 1 3808
box -38 -48 314 592
use scs8hd_conb_1  _209_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9568 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 9936 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_90
timestamp 1586364061
transform 1 0 9384 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_94
timestamp 1586364061
transform 1 0 9752 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_101
timestamp 1586364061
transform 1 0 10396 0 1 3808
box -38 -48 774 592
use scs8hd_conb_1  _208_
timestamp 1586364061
transform 1 0 11316 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_109
timestamp 1586364061
transform 1 0 11132 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 222 592
use scs8hd_conb_1  _205_
timestamp 1586364061
transform 1 0 13156 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 14168 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12604 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_127
timestamp 1586364061
transform 1 0 12788 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_134
timestamp 1586364061
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_138
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15640 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_151
timestamp 1586364061
transform 1 0 14996 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_156
timestamp 1586364061
transform 1 0 15456 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_160
timestamp 1586364061
transform 1 0 15824 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_172
timestamp 1586364061
transform 1 0 16928 0 1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_3_180
timestamp 1586364061
transform 1 0 17664 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_220
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_232
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_253
timestamp 1586364061
transform 1 0 24380 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use scs8hd_inv_8  _088_
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_6  FILLER_4_12
timestamp 1586364061
transform 1 0 2208 0 -1 4896
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 2760 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__C
timestamp 1586364061
transform 1 0 3128 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_20
timestamp 1586364061
transform 1 0 2944 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_24
timestamp 1586364061
transform 1 0 3312 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_4_30
timestamp 1586364061
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_6  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 590 592
use scs8hd_decap_8  FILLER_4_53
timestamp 1586364061
transform 1 0 5980 0 -1 4896
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6808 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7176 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_61
timestamp 1586364061
transform 1 0 6716 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_64
timestamp 1586364061
transform 1 0 6992 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8372 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_77
timestamp 1586364061
transform 1 0 8188 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_81
timestamp 1586364061
transform 1 0 8556 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_85
timestamp 1586364061
transform 1 0 8924 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_89
timestamp 1586364061
transform 1 0 9292 0 -1 4896
box -38 -48 130 592
use scs8hd_inv_8  _203_
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_102
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11592 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12144 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_4_122
timestamp 1586364061
transform 1 0 12328 0 -1 4896
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12604 0 -1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13064 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_128
timestamp 1586364061
transform 1 0 12880 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_132
timestamp 1586364061
transform 1 0 13248 0 -1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_145
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_149
timestamp 1586364061
transform 1 0 14812 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_163
timestamp 1586364061
transform 1 0 16100 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_175
timestamp 1586364061
transform 1 0 17204 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_187
timestamp 1586364061
transform 1 0 18308 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_199
timestamp 1586364061
transform 1 0 19412 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_4_211
timestamp 1586364061
transform 1 0 20516 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_239
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_258
timestamp 1586364061
transform 1 0 24840 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_270
timestamp 1586364061
transform 1 0 25944 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_274
timestamp 1586364061
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 2392 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__B
timestamp 1586364061
transform 1 0 2024 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_5_9
timestamp 1586364061
transform 1 0 1932 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_12
timestamp 1586364061
transform 1 0 2208 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_16
timestamp 1586364061
transform 1 0 2576 0 1 4896
box -38 -48 222 592
use scs8hd_or3_4  _089_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2760 0 1 4896
box -38 -48 866 592
use scs8hd_buf_1  _164_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4324 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 4048 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_31
timestamp 1586364061
transform 1 0 3956 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_34
timestamp 1586364061
transform 1 0 4232 0 1 4896
box -38 -48 130 592
use scs8hd_buf_1  _162_
timestamp 1586364061
transform 1 0 5704 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 5520 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_38
timestamp 1586364061
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_42
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 590 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_73
timestamp 1586364061
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_77
timestamp 1586364061
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9568 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_90
timestamp 1586364061
transform 1 0 9384 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_94
timestamp 1586364061
transform 1 0 9752 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_107
timestamp 1586364061
transform 1 0 10948 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11132 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_111
timestamp 1586364061
transform 1 0 11316 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_115
timestamp 1586364061
transform 1 0 11684 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12696 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13892 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_141
timestamp 1586364061
transform 1 0 14076 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _187_
timestamp 1586364061
transform 1 0 15824 0 1 4896
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14260 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_152
timestamp 1586364061
transform 1 0 15088 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_156
timestamp 1586364061
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_169
timestamp 1586364061
transform 1 0 16652 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_173
timestamp 1586364061
transform 1 0 17020 0 1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_181
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_196
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_220
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_232
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_7
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_buf_2  _221_
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_7_16
timestamp 1586364061
transform 1 0 2576 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_7_11
timestamp 1586364061
transform 1 0 2116 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_11
timestamp 1586364061
transform 1 0 2116 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 2208 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__221__A
timestamp 1586364061
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 2392 0 1 5984
box -38 -48 222 592
use scs8hd_inv_8  _113_
timestamp 1586364061
transform 1 0 2392 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 2852 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_34
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_30
timestamp 1586364061
transform 1 0 3864 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__125__C
timestamp 1586364061
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_or3_4  _163_
timestamp 1586364061
transform 1 0 3036 0 1 5984
box -38 -48 866 592
use scs8hd_inv_8  _124_
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_6_41
timestamp 1586364061
transform 1 0 4876 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 5060 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_47
timestamp 1586364061
transform 1 0 5428 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_45
timestamp 1586364061
transform 1 0 5244 0 -1 5984
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__186__B
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 5612 0 1 5984
box -38 -48 222 592
use scs8hd_buf_1  _165_
timestamp 1586364061
transform 1 0 5796 0 -1 5984
box -38 -48 314 592
use scs8hd_or3_4  _114_
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 866 592
use scs8hd_decap_3  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_55
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_59
timestamp 1586364061
transform 1 0 6532 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_6_54
timestamp 1586364061
transform 1 0 6072 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 6348 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__D
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_69
timestamp 1586364061
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_65
timestamp 1586364061
transform 1 0 7084 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 7636 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__185__B
timestamp 1586364061
transform 1 0 7268 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__185__D
timestamp 1586364061
transform 1 0 7084 0 1 5984
box -38 -48 222 592
use scs8hd_nor4_4  _185_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7268 0 1 5984
box -38 -48 1602 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__185__C
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_84
timestamp 1586364061
transform 1 0 8832 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_88
timestamp 1586364061
transform 1 0 9200 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_95
timestamp 1586364061
transform 1 0 9844 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_92
timestamp 1586364061
transform 1 0 9568 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_6  FILLER_6_106
timestamp 1586364061
transform 1 0 10856 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_6_102
timestamp 1586364061
transform 1 0 10488 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 1 5984
box -38 -48 866 592
use scs8hd_decap_4  FILLER_7_112
timestamp 1586364061
transform 1 0 11408 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_108
timestamp 1586364061
transform 1 0 11040 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_114
timestamp 1586364061
transform 1 0 11592 0 -1 5984
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 11408 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12144 0 -1 5984
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_6_131
timestamp 1586364061
transform 1 0 13156 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__C
timestamp 1586364061
transform 1 0 13340 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_138
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_134
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_142
timestamp 1586364061
transform 1 0 14168 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_135
timestamp 1586364061
transform 1 0 13524 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 13984 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13892 0 -1 5984
box -38 -48 314 592
use scs8hd_inv_8  _188_
timestamp 1586364061
transform 1 0 14168 0 1 5984
box -38 -48 866 592
use scs8hd_conb_1  _213_
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14352 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 15272 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_146
timestamp 1586364061
transform 1 0 14536 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_6_152
timestamp 1586364061
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_151
timestamp 1586364061
transform 1 0 14996 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_7_156
timestamp 1586364061
transform 1 0 15456 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_163
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_175
timestamp 1586364061
transform 1 0 17204 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_162
timestamp 1586364061
transform 1 0 16008 0 1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_7_170
timestamp 1586364061
transform 1 0 16744 0 1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_173
timestamp 1586364061
transform 1 0 17020 0 1 5984
box -38 -48 774 592
use scs8hd_buf_2  _241_
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__241__A
timestamp 1586364061
transform 1 0 18584 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_187
timestamp 1586364061
transform 1 0 18308 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_181
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_188
timestamp 1586364061
transform 1 0 18400 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_192
timestamp 1586364061
transform 1 0 18768 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_199
timestamp 1586364061
transform 1 0 19412 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_6_211
timestamp 1586364061
transform 1 0 20516 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_204
timestamp 1586364061
transform 1 0 19872 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_216
timestamp 1586364061
transform 1 0 20976 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_228
timestamp 1586364061
transform 1 0 22080 0 1 5984
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_240
timestamp 1586364061
transform 1 0 23184 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_248
timestamp 1586364061
transform 1 0 23920 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__226__A
timestamp 1586364061
transform 1 0 24564 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_263
timestamp 1586364061
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_7_252
timestamp 1586364061
transform 1 0 24288 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_257
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use scs8hd_or3_4  _125_
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 866 592
use scs8hd_conb_1  _210_
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 1840 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_6
timestamp 1586364061
transform 1 0 1656 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_10
timestamp 1586364061
transform 1 0 2024 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__D
timestamp 1586364061
transform 1 0 4232 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_8  _135_
timestamp 1586364061
transform 1 0 4784 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__114__C
timestamp 1586364061
transform 1 0 4600 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__C
timestamp 1586364061
transform 1 0 5796 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_36
timestamp 1586364061
transform 1 0 4416 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_49
timestamp 1586364061
transform 1 0 5612 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_53
timestamp 1586364061
transform 1 0 5980 0 -1 7072
box -38 -48 222 592
use scs8hd_nor4_4  _186_
timestamp 1586364061
transform 1 0 6348 0 -1 7072
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__186__C
timestamp 1586364061
transform 1 0 6164 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__D
timestamp 1586364061
transform 1 0 8096 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__B
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__D
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_74
timestamp 1586364061
transform 1 0 7912 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_78
timestamp 1586364061
transform 1 0 8280 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_82
timestamp 1586364061
transform 1 0 8648 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_86
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_15.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_90
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_104
timestamp 1586364061
transform 1 0 10672 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_8  _201_
timestamp 1586364061
transform 1 0 11408 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_108
timestamp 1586364061
transform 1 0 11040 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_121
timestamp 1586364061
transform 1 0 12236 0 -1 7072
box -38 -48 222 592
use scs8hd_or3_4  _086_
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 14168 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_125
timestamp 1586364061
transform 1 0 12604 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_138
timestamp 1586364061
transform 1 0 13800 0 -1 7072
box -38 -48 406 592
use scs8hd_inv_8  _197_
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_144
timestamp 1586364061
transform 1 0 14352 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_150
timestamp 1586364061
transform 1 0 14904 0 -1 7072
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_163
timestamp 1586364061
transform 1 0 16100 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_12  FILLER_8_174
timestamp 1586364061
transform 1 0 17112 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_186
timestamp 1586364061
transform 1 0 18216 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_198
timestamp 1586364061
transform 1 0 19320 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_8_210
timestamp 1586364061
transform 1 0 20424 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use scs8hd_buf_2  _226_
timestamp 1586364061
transform 1 0 24564 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_4  FILLER_8_251
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_259
timestamp 1586364061
transform 1 0 24932 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_271
timestamp 1586364061
transform 1 0 26036 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_inv_8  _190_
timestamp 1586364061
transform 1 0 1656 0 1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2668 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 222 592
use scs8hd_buf_1  _115_
timestamp 1586364061
transform 1 0 3680 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 4140 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3496 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3036 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_19
timestamp 1586364061
transform 1 0 2852 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_23
timestamp 1586364061
transform 1 0 3220 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_31
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_35
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use scs8hd_buf_1  _090_
timestamp 1586364061
transform 1 0 5704 0 1 7072
box -38 -48 314 592
use scs8hd_buf_1  _126_
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 5520 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_42
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_46
timestamp 1586364061
transform 1 0 5336 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__C
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__B
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_65
timestamp 1586364061
transform 1 0 7084 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_69
timestamp 1586364061
transform 1 0 7452 0 1 7072
box -38 -48 222 592
use scs8hd_nor4_4  _184_
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 1602 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_15.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__C
timestamp 1586364061
transform 1 0 9568 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_90
timestamp 1586364061
transform 1 0 9384 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_94
timestamp 1586364061
transform 1 0 9752 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 11316 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_109
timestamp 1586364061
transform 1 0 11132 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_113
timestamp 1586364061
transform 1 0 11500 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_117
timestamp 1586364061
transform 1 0 11868 0 1 7072
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13984 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_132
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_136
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15180 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14444 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14996 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_143
timestamp 1586364061
transform 1 0 14260 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_147
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16744 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16192 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16560 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_162
timestamp 1586364061
transform 1 0 16008 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_166
timestamp 1586364061
transform 1 0 16376 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_173
timestamp 1586364061
transform 1 0 17020 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_177
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__242__A
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_181
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_187
timestamp 1586364061
transform 1 0 18308 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_191
timestamp 1586364061
transform 1 0 18676 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_203
timestamp 1586364061
transform 1 0 19780 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_215
timestamp 1586364061
transform 1 0 20884 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_227
timestamp 1586364061
transform 1 0 21988 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_9_239
timestamp 1586364061
transform 1 0 23092 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_243
timestamp 1586364061
transform 1 0 23460 0 1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_253
timestamp 1586364061
transform 1 0 24380 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_258
timestamp 1586364061
transform 1 0 24840 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_262
timestamp 1586364061
transform 1 0 25208 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_9_274
timestamp 1586364061
transform 1 0 26312 0 1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2208 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1656 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2024 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_8
timestamp 1586364061
transform 1 0 1840 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__168__D
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_21
timestamp 1586364061
transform 1 0 3036 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use scs8hd_nor4_4  _166_
timestamp 1586364061
transform 1 0 4968 0 -1 8160
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 4416 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 4784 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_38
timestamp 1586364061
transform 1 0 4600 0 -1 8160
box -38 -48 222 592
use scs8hd_nor4_4  _179_
timestamp 1586364061
transform 1 0 7268 0 -1 8160
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__180__B
timestamp 1586364061
transform 1 0 6900 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_59
timestamp 1586364061
transform 1 0 6532 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_65
timestamp 1586364061
transform 1 0 7084 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_88
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_8  _202_
timestamp 1586364061
transform 1 0 9752 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_103
timestamp 1586364061
transform 1 0 10580 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_107
timestamp 1586364061
transform 1 0 10948 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11316 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__095__C
timestamp 1586364061
transform 1 0 12328 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_120
timestamp 1586364061
transform 1 0 12144 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_124
timestamp 1586364061
transform 1 0 12512 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_11.LATCH_1_.latch
timestamp 1586364061
transform 1 0 13248 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12696 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_128
timestamp 1586364061
transform 1 0 12880 0 -1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_143
timestamp 1586364061
transform 1 0 14260 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_147
timestamp 1586364061
transform 1 0 14628 0 -1 8160
box -38 -48 590 592
use scs8hd_buf_2  _242_
timestamp 1586364061
transform 1 0 16836 0 -1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_163
timestamp 1586364061
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_167
timestamp 1586364061
transform 1 0 16468 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_8  FILLER_10_175
timestamp 1586364061
transform 1 0 17204 0 -1 8160
box -38 -48 774 592
use scs8hd_conb_1  _206_
timestamp 1586364061
transform 1 0 17940 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 18400 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_186
timestamp 1586364061
transform 1 0 18216 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_190
timestamp 1586364061
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19872 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_202
timestamp 1586364061
transform 1 0 19688 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_206
timestamp 1586364061
transform 1 0 20056 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_227
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_239
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_251
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_263
timestamp 1586364061
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1656 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2668 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 222 592
use scs8hd_buf_1  _167_
timestamp 1586364061
transform 1 0 3404 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 3220 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_19
timestamp 1586364061
transform 1 0 2852 0 1 8160
box -38 -48 406 592
use scs8hd_decap_4  FILLER_11_28
timestamp 1586364061
transform 1 0 3680 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_34
timestamp 1586364061
transform 1 0 4232 0 1 8160
box -38 -48 222 592
use scs8hd_nor4_4  _168_
timestamp 1586364061
transform 1 0 4416 0 1 8160
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_buf_1  _094_
timestamp 1586364061
transform 1 0 6900 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 7360 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__180__C
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_66
timestamp 1586364061
transform 1 0 7176 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_70
timestamp 1586364061
transform 1 0 7544 0 1 8160
box -38 -48 222 592
use scs8hd_nor4_4  _183_
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__183__D
timestamp 1586364061
transform 1 0 7728 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 10120 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__C
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_91
timestamp 1586364061
transform 1 0 9476 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_95
timestamp 1586364061
transform 1 0 9844 0 1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_11_100
timestamp 1586364061
transform 1 0 10304 0 1 8160
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_11.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12512 0 1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 11684 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_110
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_11_117
timestamp 1586364061
transform 1 0 11868 0 1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14076 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 13708 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_139
timestamp 1586364061
transform 1 0 13892 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14260 0 1 8160
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15640 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 15272 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_152
timestamp 1586364061
transform 1 0 15088 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_156
timestamp 1586364061
transform 1 0 15456 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 17296 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 16928 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_169
timestamp 1586364061
transform 1 0 16652 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_174
timestamp 1586364061
transform 1 0 17112 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_178
timestamp 1586364061
transform 1 0 17480 0 1 8160
box -38 -48 314 592
use scs8hd_nor2_4  _140_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_193
timestamp 1586364061
transform 1 0 18860 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19872 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19688 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19320 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_197
timestamp 1586364061
transform 1 0 19228 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_200
timestamp 1586364061
transform 1 0 19504 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_213
timestamp 1586364061
transform 1 0 20700 0 1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__224__A
timestamp 1586364061
transform 1 0 22264 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_225
timestamp 1586364061
transform 1 0 21804 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_229
timestamp 1586364061
transform 1 0 22172 0 1 8160
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_232
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_11_248
timestamp 1586364061
transform 1 0 23920 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_252
timestamp 1586364061
transform 1 0 24288 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_264
timestamp 1586364061
transform 1 0 25392 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_11_276
timestamp 1586364061
transform 1 0 26496 0 1 8160
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 1840 0 -1 9248
box -38 -48 1050 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 1656 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__D
timestamp 1586364061
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 3036 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_19
timestamp 1586364061
transform 1 0 2852 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_1  _178_
timestamp 1586364061
transform 1 0 5888 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__168__C
timestamp 1586364061
transform 1 0 5060 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__180__D
timestamp 1586364061
transform 1 0 5704 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_41
timestamp 1586364061
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_45
timestamp 1586364061
transform 1 0 5244 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_49
timestamp 1586364061
transform 1 0 5612 0 -1 9248
box -38 -48 130 592
use scs8hd_nor4_4  _180_
timestamp 1586364061
transform 1 0 6900 0 -1 9248
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__181__C
timestamp 1586364061
transform 1 0 6532 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_55
timestamp 1586364061
transform 1 0 6164 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_61
timestamp 1586364061
transform 1 0 6716 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__B
timestamp 1586364061
transform 1 0 8648 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_88
timestamp 1586364061
transform 1 0 9200 0 -1 9248
box -38 -48 406 592
use scs8hd_inv_8  _098_
timestamp 1586364061
transform 1 0 10120 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_97
timestamp 1586364061
transform 1 0 10028 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_12_107
timestamp 1586364061
transform 1 0 10948 0 -1 9248
box -38 -48 590 592
use scs8hd_or3_4  _095_
timestamp 1586364061
transform 1 0 11684 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__102__C
timestamp 1586364061
transform 1 0 11500 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_124
timestamp 1586364061
transform 1 0 12512 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_8  _195_
timestamp 1586364061
transform 1 0 13616 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 12696 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_128
timestamp 1586364061
transform 1 0 12880 0 -1 9248
box -38 -48 590 592
use scs8hd_inv_8  _198_
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 774 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 17296 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_12  FILLER_12_163
timestamp 1586364061
transform 1 0 16100 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_12_175
timestamp 1586364061
transform 1 0 17204 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 18400 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18768 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_185
timestamp 1586364061
transform 1 0 18124 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_190
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_194
timestamp 1586364061
transform 1 0 18952 0 -1 9248
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19688 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20148 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_205
timestamp 1586364061
transform 1 0 19964 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_209
timestamp 1586364061
transform 1 0 20332 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_213
timestamp 1586364061
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use scs8hd_conb_1  _214_
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 314 592
use scs8hd_buf_2  _224_
timestamp 1586364061
transform 1 0 22264 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_218
timestamp 1586364061
transform 1 0 21160 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_234
timestamp 1586364061
transform 1 0 22632 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_246
timestamp 1586364061
transform 1 0 23736 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_258
timestamp 1586364061
transform 1 0 24840 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_270
timestamp 1586364061
transform 1 0 25944 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_274
timestamp 1586364061
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 1840 0 -1 10336
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1932 0 1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1656 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use scs8hd_decap_3  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_19
timestamp 1586364061
transform 1 0 2852 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_22
timestamp 1586364061
transform 1 0 3128 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_18
timestamp 1586364061
transform 1 0 2760 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__B
timestamp 1586364061
transform 1 0 3036 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__D
timestamp 1586364061
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__C
timestamp 1586364061
transform 1 0 3404 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2944 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__C
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__C
timestamp 1586364061
transform 1 0 3772 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_nor4_4  _171_
timestamp 1586364061
transform 1 0 3956 0 1 9248
box -38 -48 1602 592
use scs8hd_nor4_4  _170_
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 5704 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__181__B
timestamp 1586364061
transform 1 0 5980 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_48
timestamp 1586364061
transform 1 0 5520 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_52
timestamp 1586364061
transform 1 0 5888 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_49
timestamp 1586364061
transform 1 0 5612 0 -1 10336
box -38 -48 406 592
use scs8hd_nor4_4  _181_
timestamp 1586364061
transform 1 0 6532 0 -1 10336
box -38 -48 1602 592
use scs8hd_nor4_4  _182_
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__181__D
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__D
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__B
timestamp 1586364061
transform 1 0 6348 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_55
timestamp 1586364061
transform 1 0 6164 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_76
timestamp 1586364061
transform 1 0 8096 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_79
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__C
timestamp 1586364061
transform 1 0 8280 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__C
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_83
timestamp 1586364061
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__D
timestamp 1586364061
transform 1 0 8648 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_88
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_87
timestamp 1586364061
transform 1 0 9108 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 9292 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_98
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_94
timestamp 1586364061
transform 1 0 9752 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 9936 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_1  _085_
timestamp 1586364061
transform 1 0 9476 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_105
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 10948 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__C
timestamp 1586364061
transform 1 0 10304 0 1 9248
box -38 -48 222 592
use scs8hd_or3_4  _108_
timestamp 1586364061
transform 1 0 10488 0 1 9248
box -38 -48 866 592
use scs8hd_inv_8  _084_
timestamp 1586364061
transform 1 0 9936 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_109
timestamp 1586364061
transform 1 0 11132 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_115
timestamp 1586364061
transform 1 0 11684 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_111
timestamp 1586364061
transform 1 0 11316 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 11316 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 11500 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_122
timestamp 1586364061
transform 1 0 12328 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_119
timestamp 1586364061
transform 1 0 12052 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 12512 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 11868 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_or3_4  _102_
timestamp 1586364061
transform 1 0 11500 0 -1 10336
box -38 -48 866 592
use scs8hd_nor2_4  _093_
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use scs8hd_decap_4  FILLER_14_130
timestamp 1586364061
transform 1 0 13064 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_126
timestamp 1586364061
transform 1 0 12696 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_132
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12880 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_134
timestamp 1586364061
transform 1 0 13432 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_13_137
timestamp 1586364061
transform 1 0 13708 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_4  FILLER_14_148
timestamp 1586364061
transform 1 0 14720 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_144
timestamp 1586364061
transform 1 0 14352 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_151
timestamp 1586364061
transform 1 0 14996 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_157
timestamp 1586364061
transform 1 0 15548 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_152
timestamp 1586364061
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_155
timestamp 1586364061
transform 1 0 15364 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15732 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 15180 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15548 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_1  _100_
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_166
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_161
timestamp 1586364061
transform 1 0 15916 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_168
timestamp 1586364061
transform 1 0 16560 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_177
timestamp 1586364061
transform 1 0 17388 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_4  FILLER_13_176
timestamp 1586364061
transform 1 0 17296 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_172
timestamp 1586364061
transform 1 0 16928 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17112 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16744 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16560 0 -1 10336
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 18400 0 -1 10336
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 18400 0 1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 18216 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_180
timestamp 1586364061
transform 1 0 17664 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_185
timestamp 1586364061
transform 1 0 18124 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20148 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19964 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19596 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20332 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_199
timestamp 1586364061
transform 1 0 19412 0 1 9248
box -38 -48 590 592
use scs8hd_fill_2  FILLER_14_199
timestamp 1586364061
transform 1 0 19412 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_203
timestamp 1586364061
transform 1 0 19780 0 -1 10336
box -38 -48 590 592
use scs8hd_decap_3  FILLER_14_211
timestamp 1586364061
transform 1 0 20516 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21160 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21528 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_216
timestamp 1586364061
transform 1 0 20976 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_220
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_224
timestamp 1586364061
transform 1 0 21712 0 1 9248
box -38 -48 774 592
use scs8hd_decap_8  FILLER_14_224
timestamp 1586364061
transform 1 0 21712 0 -1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_234
timestamp 1586364061
transform 1 0 22632 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_242
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_235
timestamp 1586364061
transform 1 0 22724 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_247
timestamp 1586364061
transform 1 0 23828 0 -1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_253
timestamp 1586364061
transform 1 0 24380 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_257
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_258
timestamp 1586364061
transform 1 0 24840 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use scs8hd_decap_4  FILLER_14_270
timestamp 1586364061
transform 1 0 25944 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_274
timestamp 1586364061
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2024 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1840 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 130 592
use scs8hd_inv_8  _083_
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 3404 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__D
timestamp 1586364061
transform 1 0 3036 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_19
timestamp 1586364061
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_23
timestamp 1586364061
transform 1 0 3220 0 1 10336
box -38 -48 222 592
use scs8hd_or3_4  _091_
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__091__B
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_36
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_40
timestamp 1586364061
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_nor4_4  _176_
timestamp 1586364061
transform 1 0 7176 0 1 10336
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__091__C
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 6992 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_83
timestamp 1586364061
transform 1 0 8740 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_88
timestamp 1586364061
transform 1 0 9200 0 1 10336
box -38 -48 222 592
use scs8hd_or3_4  _099_
timestamp 1586364061
transform 1 0 9936 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 9752 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__C
timestamp 1586364061
transform 1 0 9384 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 10948 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_92
timestamp 1586364061
transform 1 0 9568 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_105
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_109
timestamp 1586364061
transform 1 0 11132 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_113
timestamp 1586364061
transform 1 0 11500 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12788 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12604 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 13984 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_138
timestamp 1586364061
transform 1 0 13800 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_142
timestamp 1586364061
transform 1 0 14168 0 1 10336
box -38 -48 406 592
use scs8hd_buf_1  _096_
timestamp 1586364061
transform 1 0 14536 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 14996 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15364 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_149
timestamp 1586364061
transform 1 0 14812 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_153
timestamp 1586364061
transform 1 0 15180 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_157
timestamp 1586364061
transform 1 0 15548 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 15916 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17112 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_172
timestamp 1586364061
transform 1 0 16928 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_176
timestamp 1586364061
transform 1 0 17296 0 1 10336
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 18584 0 1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18216 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_180
timestamp 1586364061
transform 1 0 17664 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_188
timestamp 1586364061
transform 1 0 18400 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20332 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19780 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20148 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_201
timestamp 1586364061
transform 1 0 19596 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_205
timestamp 1586364061
transform 1 0 19964 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21896 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22356 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21712 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_218
timestamp 1586364061
transform 1 0 21160 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_222
timestamp 1586364061
transform 1 0 21528 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_229
timestamp 1586364061
transform 1 0 22172 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 22724 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_233
timestamp 1586364061
transform 1 0 22540 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_237
timestamp 1586364061
transform 1 0 22908 0 1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_15_243
timestamp 1586364061
transform 1 0 23460 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_257
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2024 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_7
timestamp 1586364061
transform 1 0 1748 0 -1 11424
box -38 -48 130 592
use scs8hd_nor4_4  _173_
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 3036 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__D
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_19
timestamp 1586364061
transform 1 0 2852 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__B
timestamp 1586364061
transform 1 0 5796 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_49
timestamp 1586364061
transform 1 0 5612 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_53
timestamp 1586364061
transform 1 0 5980 0 -1 11424
box -38 -48 222 592
use scs8hd_nor4_4  _177_
timestamp 1586364061
transform 1 0 7084 0 -1 11424
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__177__B
timestamp 1586364061
transform 1 0 6900 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__B
timestamp 1586364061
transform 1 0 6532 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__C
timestamp 1586364061
transform 1 0 6164 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_57
timestamp 1586364061
transform 1 0 6348 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_61
timestamp 1586364061
transform 1 0 6716 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__D
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_82
timestamp 1586364061
transform 1 0 8648 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_86
timestamp 1586364061
transform 1 0 9016 0 -1 11424
box -38 -48 590 592
use scs8hd_buf_1  _087_
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use scs8hd_inv_8  _196_
timestamp 1586364061
transform 1 0 10672 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 10212 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_96
timestamp 1586364061
transform 1 0 9936 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_101
timestamp 1586364061
transform 1 0 10396 0 -1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12236 0 -1 11424
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_16_113
timestamp 1586364061
transform 1 0 11500 0 -1 11424
box -38 -48 774 592
use scs8hd_buf_1  _109_
timestamp 1586364061
transform 1 0 13984 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_132
timestamp 1586364061
transform 1 0 13248 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_136
timestamp 1586364061
transform 1 0 13616 0 -1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 15548 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_143
timestamp 1586364061
transform 1 0 14260 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_151
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_159
timestamp 1586364061
transform 1 0 15732 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16192 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16008 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_173
timestamp 1586364061
transform 1 0 17020 0 -1 11424
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18216 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 18676 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_185
timestamp 1586364061
transform 1 0 18124 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_189
timestamp 1586364061
transform 1 0 18492 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_193
timestamp 1586364061
transform 1 0 18860 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_206
timestamp 1586364061
transform 1 0 20056 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_210
timestamp 1586364061
transform 1 0 20424 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_224
timestamp 1586364061
transform 1 0 21712 0 -1 11424
box -38 -48 774 592
use scs8hd_buf_1  _138_
timestamp 1586364061
transform 1 0 22448 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_235
timestamp 1586364061
transform 1 0 22724 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_247
timestamp 1586364061
transform 1 0 23828 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_259
timestamp 1586364061
transform 1 0 24932 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_271
timestamp 1586364061
transform 1 0 26036 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_inv_8  _189_
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_16
timestamp 1586364061
transform 1 0 2576 0 1 11424
box -38 -48 222 592
use scs8hd_nor4_4  _172_
timestamp 1586364061
transform 1 0 3956 0 1 11424
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__137__C
timestamp 1586364061
transform 1 0 2760 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 3772 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__C
timestamp 1586364061
transform 1 0 3404 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_20
timestamp 1586364061
transform 1 0 2944 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_24
timestamp 1586364061
transform 1 0 3312 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__C
timestamp 1586364061
transform 1 0 5704 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_48
timestamp 1586364061
transform 1 0 5520 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_52
timestamp 1586364061
transform 1 0 5888 0 1 11424
box -38 -48 222 592
use scs8hd_or3_4  _116_
timestamp 1586364061
transform 1 0 7176 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 6992 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__C
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__D
timestamp 1586364061
transform 1 0 6072 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_56
timestamp 1586364061
transform 1 0 6256 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use scs8hd_buf_2  _223_
timestamp 1586364061
transform 1 0 9108 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 8924 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__C
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 8556 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_75
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_79
timestamp 1586364061
transform 1 0 8372 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_83
timestamp 1586364061
transform 1 0 8740 0 1 11424
box -38 -48 222 592
use scs8hd_or3_4  _105_
timestamp 1586364061
transform 1 0 10212 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__223__A
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_91
timestamp 1586364061
transform 1 0 9476 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_95
timestamp 1586364061
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use scs8hd_buf_1  _092_
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__B
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_108
timestamp 1586364061
transform 1 0 11040 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_112
timestamp 1586364061
transform 1 0 11408 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13432 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 12880 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_126
timestamp 1586364061
transform 1 0 12696 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_130
timestamp 1586364061
transform 1 0 13064 0 1 11424
box -38 -48 222 592
use scs8hd_buf_1  _103_
timestamp 1586364061
transform 1 0 14996 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15824 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 15456 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 14812 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14444 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_143
timestamp 1586364061
transform 1 0 14260 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_147
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_154
timestamp 1586364061
transform 1 0 15272 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_158
timestamp 1586364061
transform 1 0 15640 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16008 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_173
timestamp 1586364061
transform 1 0 17020 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_177
timestamp 1586364061
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18308 0 1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_181
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20148 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19964 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19504 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_198
timestamp 1586364061
transform 1 0 19320 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_202
timestamp 1586364061
transform 1 0 19688 0 1 11424
box -38 -48 314 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 21712 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 21528 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 21160 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_216
timestamp 1586364061
transform 1 0 20976 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_220
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22724 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_233
timestamp 1586364061
transform 1 0 22540 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_237
timestamp 1586364061
transform 1 0 22908 0 1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_17_243
timestamp 1586364061
transform 1 0 23460 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_249
timestamp 1586364061
transform 1 0 24012 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_261
timestamp 1586364061
transform 1 0 25116 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_17_273
timestamp 1586364061
transform 1 0 26220 0 1 11424
box -38 -48 406 592
use scs8hd_buf_1  _111_
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use scs8hd_or3_4  _137_
timestamp 1586364061
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_6
timestamp 1586364061
transform 1 0 1656 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_10
timestamp 1586364061
transform 1 0 2024 0 -1 12512
box -38 -48 222 592
use scs8hd_nor4_4  _175_
timestamp 1586364061
transform 1 0 4324 0 -1 12512
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__127__C
timestamp 1586364061
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_52
timestamp 1586364061
transform 1 0 5888 0 -1 12512
box -38 -48 222 592
use scs8hd_or3_4  _153_
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 7176 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__B
timestamp 1586364061
transform 1 0 6072 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 6440 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_60
timestamp 1586364061
transform 1 0 6624 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_64
timestamp 1586364061
transform 1 0 6992 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_77
timestamp 1586364061
transform 1 0 8188 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_18_89
timestamp 1586364061
transform 1 0 9292 0 -1 12512
box -38 -48 130 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__105__C
timestamp 1586364061
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_106
timestamp 1586364061
transform 1 0 10856 0 -1 12512
box -38 -48 590 592
use scs8hd_nor2_4  _101_
timestamp 1586364061
transform 1 0 11776 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 11408 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_114
timestamp 1586364061
transform 1 0 11592 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13340 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13064 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_125
timestamp 1586364061
transform 1 0 12604 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_129
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_132
timestamp 1586364061
transform 1 0 13248 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_142
timestamp 1586364061
transform 1 0 14168 0 -1 12512
box -38 -48 774 592
use scs8hd_nor2_4  _143_
timestamp 1586364061
transform 1 0 15548 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_18_150
timestamp 1586364061
transform 1 0 14904 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 17204 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 16560 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16928 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_166
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_170
timestamp 1586364061
transform 1 0 16744 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_174
timestamp 1586364061
transform 1 0 17112 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 18308 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18676 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_184
timestamp 1586364061
transform 1 0 18032 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_189
timestamp 1586364061
transform 1 0 18492 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_193
timestamp 1586364061
transform 1 0 18860 0 -1 12512
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_206
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_224
timestamp 1586364061
transform 1 0 21712 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_228
timestamp 1586364061
transform 1 0 22080 0 -1 12512
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 -1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23460 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_235
timestamp 1586364061
transform 1 0 22724 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_8  FILLER_18_246
timestamp 1586364061
transform 1 0 23736 0 -1 12512
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__237__A
timestamp 1586364061
transform 1 0 24564 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_254
timestamp 1586364061
transform 1 0 24472 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_257
timestamp 1586364061
transform 1 0 24748 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_18_269
timestamp 1586364061
transform 1 0 25852 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_6
timestamp 1586364061
transform 1 0 1656 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 1840 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1472 0 1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_10
timestamp 1586364061
transform 1 0 2024 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_12
timestamp 1586364061
transform 1 0 2208 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 2024 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 2392 0 1 12512
box -38 -48 222 592
use scs8hd_inv_8  _136_
timestamp 1586364061
transform 1 0 2392 0 -1 13600
box -38 -48 866 592
use scs8hd_or3_4  _127_
timestamp 1586364061
transform 1 0 2576 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_25
timestamp 1586364061
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__B
timestamp 1586364061
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_29
timestamp 1586364061
transform 1 0 3772 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__D
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 3956 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_inv_8  _192_
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use scs8hd_nor4_4  _174_
timestamp 1586364061
transform 1 0 4140 0 1 12512
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__174__C
timestamp 1586364061
transform 1 0 5888 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 5060 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5980 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_50
timestamp 1586364061
transform 1 0 5704 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_41
timestamp 1586364061
transform 1 0 4876 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_45
timestamp 1586364061
transform 1 0 5244 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_4  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_58
timestamp 1586364061
transform 1 0 6440 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_54
timestamp 1586364061
transform 1 0 6072 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_70
timestamp 1586364061
transform 1 0 7544 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_4  FILLER_20_64
timestamp 1586364061
transform 1 0 6992 0 -1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__C
timestamp 1586364061
transform 1 0 7176 0 1 12512
box -38 -48 222 592
use scs8hd_inv_8  _200_
timestamp 1586364061
transform 1 0 6164 0 -1 13600
box -38 -48 866 592
use scs8hd_or3_4  _145_
timestamp 1586364061
transform 1 0 7360 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _110_
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 8740 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9200 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_77
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_81
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_85
timestamp 1586364061
transform 1 0 8924 0 1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_74
timestamp 1586364061
transform 1 0 7912 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9568 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10764 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_90
timestamp 1586364061
transform 1 0 9384 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_103
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_107
timestamp 1586364061
transform 1 0 10948 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_104
timestamp 1586364061
transform 1 0 10672 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 11132 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_121
timestamp 1586364061
transform 1 0 12236 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1050 592
use scs8hd_nor2_4  _104_
timestamp 1586364061
transform 1 0 11408 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_1  FILLER_20_129
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_125
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12788 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_141
timestamp 1586364061
transform 1 0 14076 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_138
timestamp 1586364061
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_134
timestamp 1586364061
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 13064 0 -1 13600
box -38 -48 1050 592
use scs8hd_nor2_4  _097_
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14260 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_151
timestamp 1586364061
transform 1 0 14996 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_156
timestamp 1586364061
transform 1 0 15456 0 1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_20_167
timestamp 1586364061
transform 1 0 16468 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_163
timestamp 1586364061
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 16284 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_174
timestamp 1586364061
transform 1 0 17112 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_172
timestamp 1586364061
transform 1 0 16928 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_168
timestamp 1586364061
transform 1 0 16560 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16652 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 16744 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_6  FILLER_20_178
timestamp 1586364061
transform 1 0 17480 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_19_176
timestamp 1586364061
transform 1 0 17296 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17296 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _139_
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 18032 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_179
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_193
timestamp 1586364061
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_203
timestamp 1586364061
transform 1 0 19780 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_20_197
timestamp 1586364061
transform 1 0 19228 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_19_201
timestamp 1586364061
transform 1 0 19596 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_197
timestamp 1586364061
transform 1 0 19228 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19872 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19688 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_210
timestamp 1586364061
transform 1 0 20424 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_206
timestamp 1586364061
transform 1 0 20056 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_213
timestamp 1586364061
transform 1 0 20700 0 1 12512
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19872 0 1 12512
box -38 -48 866 592
use scs8hd_conb_1  _218_
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21436 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21896 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21252 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21436 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_230
timestamp 1586364061
transform 1 0 22264 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_218
timestamp 1586364061
transform 1 0 21160 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_223
timestamp 1586364061
transform 1 0 21620 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_239
timestamp 1586364061
transform 1 0 23092 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_235
timestamp 1586364061
transform 1 0 22724 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_234
timestamp 1586364061
transform 1 0 22632 0 1 12512
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22908 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_249
timestamp 1586364061
transform 1 0 24012 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_242
timestamp 1586364061
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 23828 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_nor2_4  _130_
timestamp 1586364061
transform 1 0 23460 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_4  FILLER_20_256
timestamp 1586364061
transform 1 0 24656 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_252
timestamp 1586364061
transform 1 0 24288 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_253
timestamp 1586364061
transform 1 0 24380 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 24196 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 24472 0 -1 13600
box -38 -48 222 592
use scs8hd_buf_2  _237_
timestamp 1586364061
transform 1 0 24564 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_259
timestamp 1586364061
transform 1 0 24932 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25116 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25024 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_263
timestamp 1586364061
transform 1 0 25300 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_263
timestamp 1586364061
transform 1 0 25300 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_275
timestamp 1586364061
transform 1 0 26404 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__230__A
timestamp 1586364061
transform 1 0 1840 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 2668 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_6
timestamp 1586364061
transform 1 0 1656 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_10
timestamp 1586364061
transform 1 0 2024 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_14
timestamp 1586364061
transform 1 0 2392 0 1 13600
box -38 -48 314 592
use scs8hd_buf_1  _169_
timestamp 1586364061
transform 1 0 2852 0 1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 3864 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3312 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3680 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_22
timestamp 1586364061
transform 1 0 3128 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_26
timestamp 1586364061
transform 1 0 3496 0 1 13600
box -38 -48 222 592
use scs8hd_buf_1  _112_
timestamp 1586364061
transform 1 0 5704 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5060 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5428 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_41
timestamp 1586364061
transform 1 0 4876 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_45
timestamp 1586364061
transform 1 0 5244 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_49
timestamp 1586364061
transform 1 0 5612 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_13.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8740 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9200 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8280 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_73
timestamp 1586364061
transform 1 0 7820 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_77
timestamp 1586364061
transform 1 0 8188 0 1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_21_80
timestamp 1586364061
transform 1 0 8464 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_86
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9752 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9568 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10948 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_90
timestamp 1586364061
transform 1 0 9384 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_105
timestamp 1586364061
transform 1 0 10764 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11316 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_109
timestamp 1586364061
transform 1 0 11132 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_113
timestamp 1586364061
transform 1 0 11500 0 1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_21_119
timestamp 1586364061
transform 1 0 12052 0 1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_134
timestamp 1586364061
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_138
timestamp 1586364061
transform 1 0 13800 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 15732 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 15272 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_151
timestamp 1586364061
transform 1 0 14996 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_21_156
timestamp 1586364061
transform 1 0 15456 0 1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 15916 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_172
timestamp 1586364061
transform 1 0 16928 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_176
timestamp 1586364061
transform 1 0 17296 0 1 13600
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18676 0 1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 18216 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_179
timestamp 1586364061
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_188
timestamp 1586364061
transform 1 0 18400 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20424 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19872 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_202
timestamp 1586364061
transform 1 0 19688 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_206
timestamp 1586364061
transform 1 0 20056 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21988 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 21804 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21436 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_219
timestamp 1586364061
transform 1 0 21252 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_223
timestamp 1586364061
transform 1 0 21620 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_236
timestamp 1586364061
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_240
timestamp 1586364061
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use scs8hd_buf_2  _234_
timestamp 1586364061
transform 1 0 25208 0 1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24656 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_254
timestamp 1586364061
transform 1 0 24472 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_258
timestamp 1586364061
transform 1 0 24840 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_266
timestamp 1586364061
transform 1 0 25576 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__234__A
timestamp 1586364061
transform 1 0 25760 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_270
timestamp 1586364061
transform 1 0 25944 0 1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_21_276
timestamp 1586364061
transform 1 0 26496 0 1 13600
box -38 -48 130 592
use scs8hd_buf_2  _230_
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2024 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_7
timestamp 1586364061
transform 1 0 1748 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_12
timestamp 1586364061
transform 1 0 2208 0 -1 14688
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4232 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_23
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_43
timestamp 1586364061
transform 1 0 5060 0 -1 14688
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6716 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_57
timestamp 1586364061
transform 1 0 6348 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_70
timestamp 1586364061
transform 1 0 7544 0 -1 14688
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8280 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_81
timestamp 1586364061
transform 1 0 8556 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_22_89
timestamp 1586364061
transform 1 0 9292 0 -1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9844 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_97
timestamp 1586364061
transform 1 0 10028 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12420 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_109
timestamp 1586364061
transform 1 0 11132 0 -1 14688
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_22_121
timestamp 1586364061
transform 1 0 12236 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 12788 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14168 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_125
timestamp 1586364061
transform 1 0 12604 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_138
timestamp 1586364061
transform 1 0 13800 0 -1 14688
box -38 -48 406 592
use scs8hd_buf_1  _128_
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15732 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_144
timestamp 1586364061
transform 1 0 14352 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_22_152
timestamp 1586364061
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_157
timestamp 1586364061
transform 1 0 15548 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16100 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_161
timestamp 1586364061
transform 1 0 15916 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_165
timestamp 1586364061
transform 1 0 16284 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_175
timestamp 1586364061
transform 1 0 17204 0 -1 14688
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 17940 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19136 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_194
timestamp 1586364061
transform 1 0 18952 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19504 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_198
timestamp 1586364061
transform 1 0 19320 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_202
timestamp 1586364061
transform 1 0 19688 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_6  FILLER_22_206
timestamp 1586364061
transform 1 0 20056 0 -1 14688
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21988 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_224
timestamp 1586364061
transform 1 0 21712 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_22_229
timestamp 1586364061
transform 1 0 22172 0 -1 14688
box -38 -48 314 592
use scs8hd_nor2_4  _134_
timestamp 1586364061
transform 1 0 22448 0 -1 14688
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24012 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 23644 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_241
timestamp 1586364061
transform 1 0 23276 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_247
timestamp 1586364061
transform 1 0 23828 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_252
timestamp 1586364061
transform 1 0 24288 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_22_264
timestamp 1586364061
transform 1 0 25392 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_22_272
timestamp 1586364061
transform 1 0 26128 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_7
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4324 0 1 14688
box -38 -48 1050 592
use scs8hd_inv_1  mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3312 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3772 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4140 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 2944 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_19
timestamp 1586364061
transform 1 0 2852 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_22
timestamp 1586364061
transform 1 0 3128 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_31
timestamp 1586364061
transform 1 0 3956 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5520 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_46
timestamp 1586364061
transform 1 0 5336 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_50
timestamp 1586364061
transform 1 0 5704 0 1 14688
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_13.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6900 0 1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_54
timestamp 1586364061
transform 1 0 6072 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8096 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9200 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8464 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_74
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_78
timestamp 1586364061
transform 1 0 8280 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_82
timestamp 1586364061
transform 1 0 8648 0 1 14688
box -38 -48 590 592
use scs8hd_buf_1  _106_
timestamp 1586364061
transform 1 0 10948 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9384 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_99
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_103
timestamp 1586364061
transform 1 0 10580 0 1 14688
box -38 -48 222 592
use scs8hd_conb_1  _217_
timestamp 1586364061
transform 1 0 12512 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_110
timestamp 1586364061
transform 1 0 11224 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_114
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_120
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12972 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13340 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_127
timestamp 1586364061
transform 1 0 12788 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_131
timestamp 1586364061
transform 1 0 13156 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15088 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15548 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14904 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_144
timestamp 1586364061
transform 1 0 14352 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_148
timestamp 1586364061
transform 1 0 14720 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_155
timestamp 1586364061
transform 1 0 15364 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_159
timestamp 1586364061
transform 1 0 15732 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15916 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_172
timestamp 1586364061
transform 1 0 16928 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_177
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_2_.latch
timestamp 1586364061
transform 1 0 19044 0 1 14688
box -38 -48 1050 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_181
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_187
timestamp 1586364061
transform 1 0 18308 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_191
timestamp 1586364061
transform 1 0 18676 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20700 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20332 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_206
timestamp 1586364061
transform 1 0 20056 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_211
timestamp 1586364061
transform 1 0 20516 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21252 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21068 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_215
timestamp 1586364061
transform 1 0 20884 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_228
timestamp 1586364061
transform 1 0 22080 0 1 14688
box -38 -48 406 592
use scs8hd_nor2_4  _132_
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22448 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22816 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_234
timestamp 1586364061
transform 1 0 22632 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_238
timestamp 1586364061
transform 1 0 23000 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__231__A
timestamp 1586364061
transform 1 0 24656 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_254
timestamp 1586364061
transform 1 0 24472 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_258
timestamp 1586364061
transform 1 0 24840 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_decap_6  FILLER_23_270
timestamp 1586364061
transform 1 0 25944 0 1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_23_276
timestamp 1586364061
transform 1 0 26496 0 1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__220__A
timestamp 1586364061
transform 1 0 1564 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_7
timestamp 1586364061
transform 1 0 1748 0 -1 15776
box -38 -48 1142 592
use scs8hd_buf_1  _161_
timestamp 1586364061
transform 1 0 2944 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4232 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_19
timestamp 1586364061
transform 1 0 2852 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_6  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_2  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5244 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5980 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_43
timestamp 1586364061
transform 1 0 5060 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_47
timestamp 1586364061
transform 1 0 5428 0 -1 15776
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6164 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 7176 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7544 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_64
timestamp 1586364061
transform 1 0 6992 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_68
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7728 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_81
timestamp 1586364061
transform 1 0 8556 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_87
timestamp 1586364061
transform 1 0 9108 0 -1 15776
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10028 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_90
timestamp 1586364061
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_3  FILLER_24_106
timestamp 1586364061
transform 1 0 10856 0 -1 15776
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11960 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11132 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11500 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_111
timestamp 1586364061
transform 1 0 11316 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_115
timestamp 1586364061
transform 1 0 11684 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_121
timestamp 1586364061
transform 1 0 12236 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_138
timestamp 1586364061
transform 1 0 13800 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_142
timestamp 1586364061
transform 1 0 14168 0 -1 15776
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15824 0 -1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15640 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_150
timestamp 1586364061
transform 1 0 14904 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_4  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_8  FILLER_24_171
timestamp 1586364061
transform 1 0 16836 0 -1 15776
box -38 -48 774 592
use scs8hd_nor2_4  _148_
timestamp 1586364061
transform 1 0 17572 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19044 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18676 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_188
timestamp 1586364061
transform 1 0 18400 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_193
timestamp 1586364061
transform 1 0 18860 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_206
timestamp 1586364061
transform 1 0 20056 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21896 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22264 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_224
timestamp 1586364061
transform 1 0 21712 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_228
timestamp 1586364061
transform 1 0 22080 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22448 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_12  FILLER_24_241
timestamp 1586364061
transform 1 0 23276 0 -1 15776
box -38 -48 1142 592
use scs8hd_buf_2  _231_
timestamp 1586364061
transform 1 0 24564 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_253
timestamp 1586364061
transform 1 0 24380 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_259
timestamp 1586364061
transform 1 0 24932 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_271
timestamp 1586364061
transform 1 0 26036 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_buf_2  _220_
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_7
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_11
timestamp 1586364061
transform 1 0 2116 0 1 15776
box -38 -48 774 592
use scs8hd_inv_8  _191_
timestamp 1586364061
transform 1 0 3312 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4324 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 3128 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_19
timestamp 1586364061
transform 1 0 2852 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_33
timestamp 1586364061
transform 1 0 4140 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4876 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5888 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_37
timestamp 1586364061
transform 1 0 4508 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_50
timestamp 1586364061
transform 1 0 5704 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7452 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7084 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_54
timestamp 1586364061
transform 1 0 6072 0 1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_25_60
timestamp 1586364061
transform 1 0 6624 0 1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_67
timestamp 1586364061
transform 1 0 7268 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9200 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_80
timestamp 1586364061
transform 1 0 8464 0 1 15776
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10212 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_97
timestamp 1586364061
transform 1 0 10028 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_101
timestamp 1586364061
transform 1 0 10396 0 1 15776
box -38 -48 222 592
use scs8hd_buf_1  _117_
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__B
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_114
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_118
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 12880 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_126
timestamp 1586364061
transform 1 0 12696 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_130
timestamp 1586364061
transform 1 0 13064 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_134
timestamp 1586364061
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15088 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15548 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14904 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_144
timestamp 1586364061
transform 1 0 14352 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_148
timestamp 1586364061
transform 1 0 14720 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_155
timestamp 1586364061
transform 1 0 15364 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_159
timestamp 1586364061
transform 1 0 15732 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _149_
timestamp 1586364061
transform 1 0 16376 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 15916 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_163
timestamp 1586364061
transform 1 0 16100 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_175
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_179
timestamp 1586364061
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18124 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_192
timestamp 1586364061
transform 1 0 18768 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_188
timestamp 1586364061
transform 1 0 18400 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18952 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18584 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19136 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20148 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_205
timestamp 1586364061
transform 1 0 19964 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_209
timestamp 1586364061
transform 1 0 20332 0 1 15776
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21620 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 20884 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 21252 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_217
timestamp 1586364061
transform 1 0 21068 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_221
timestamp 1586364061
transform 1 0 21436 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 22632 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_232
timestamp 1586364061
transform 1 0 22448 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_236
timestamp 1586364061
transform 1 0 22816 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_240
timestamp 1586364061
transform 1 0 23184 0 1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_257
timestamp 1586364061
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_25_269
timestamp 1586364061
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2668 0 1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1656 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_8  FILLER_26_9
timestamp 1586364061
transform 1 0 1932 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_26_17
timestamp 1586364061
transform 1 0 2668 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_24
timestamp 1586364061
transform 1 0 3312 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_20
timestamp 1586364061
transform 1 0 2944 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3496 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3128 0 1 16864
box -38 -48 222 592
use scs8hd_conb_1  _211_
timestamp 1586364061
transform 1 0 2944 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_27_35
timestamp 1586364061
transform 1 0 4324 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_31
timestamp 1586364061
transform 1 0 3956 0 1 16864
box -38 -48 406 592
use scs8hd_decap_3  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4324 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_conb_1  _207_
timestamp 1586364061
transform 1 0 3680 0 1 16864
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4968 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4416 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4692 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_37
timestamp 1586364061
transform 1 0 4508 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_41
timestamp 1586364061
transform 1 0 4876 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_51
timestamp 1586364061
transform 1 0 5796 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_27_38
timestamp 1586364061
transform 1 0 4600 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_50
timestamp 1586364061
transform 1 0 5704 0 1 16864
box -38 -48 406 592
use scs8hd_decap_4  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_54
timestamp 1586364061
transform 1 0 6072 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_27_69
timestamp 1586364061
transform 1 0 7452 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_65
timestamp 1586364061
transform 1 0 7084 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_63
timestamp 1586364061
transform 1 0 6900 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 16864
box -38 -48 222 592
use scs8hd_inv_8  _199_
timestamp 1586364061
transform 1 0 7176 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_26_79
timestamp 1586364061
transform 1 0 8372 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_75
timestamp 1586364061
transform 1 0 8004 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 7728 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_89
timestamp 1586364061
transform 1 0 9292 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_85
timestamp 1586364061
transform 1 0 8924 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_83
timestamp 1586364061
transform 1 0 8740 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8556 0 -1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_27_96
timestamp 1586364061
transform 1 0 9936 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_96
timestamp 1586364061
transform 1 0 9936 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_91
timestamp 1586364061
transform 1 0 9476 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9476 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 314 592
use scs8hd_buf_1  _154_
timestamp 1586364061
transform 1 0 9660 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_27_104
timestamp 1586364061
transform 1 0 10672 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_100
timestamp 1586364061
transform 1 0 10304 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_107
timestamp 1586364061
transform 1 0 10948 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_103
timestamp 1586364061
transform 1 0 10580 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_100
timestamp 1586364061
transform 1 0 10304 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10396 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_5_.latch
timestamp 1586364061
transform 1 0 11132 0 -1 16864
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_120
timestamp 1586364061
transform 1 0 12144 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_132
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 406 592
use scs8hd_decap_3  FILLER_26_125
timestamp 1586364061
transform 1 0 12604 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_27_142
timestamp 1586364061
transform 1 0 14168 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_138
timestamp 1586364061
transform 1 0 13800 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_141
timestamp 1586364061
transform 1 0 14076 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_26_137
timestamp 1586364061
transform 1 0 13708 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13892 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 13984 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 13616 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _155_
timestamp 1586364061
transform 1 0 12880 0 -1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_4_.latch
timestamp 1586364061
transform 1 0 14720 0 1 16864
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_5_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 14536 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14720 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_147
timestamp 1586364061
transform 1 0 14628 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_26_150
timestamp 1586364061
transform 1 0 14904 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_159
timestamp 1586364061
transform 1 0 15732 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_163
timestamp 1586364061
transform 1 0 16100 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_169
timestamp 1586364061
transform 1 0 16652 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_165
timestamp 1586364061
transform 1 0 16284 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16284 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 16468 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 15916 0 1 16864
box -38 -48 222 592
use scs8hd_buf_1  _146_
timestamp 1586364061
transform 1 0 16468 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_27_174
timestamp 1586364061
transform 1 0 17112 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_170
timestamp 1586364061
transform 1 0 16744 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_173
timestamp 1586364061
transform 1 0 17020 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 16836 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 16928 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_179
timestamp 1586364061
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_181
timestamp 1586364061
transform 1 0 17756 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_27_188
timestamp 1586364061
transform 1 0 18400 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_195
timestamp 1586364061
transform 1 0 19044 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 18492 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_5_.latch
timestamp 1586364061
transform 1 0 18676 0 1 16864
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_3_.latch
timestamp 1586364061
transform 1 0 18032 0 -1 16864
box -38 -48 1050 592
use scs8hd_decap_6  FILLER_27_202
timestamp 1586364061
transform 1 0 19688 0 1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_26_199
timestamp 1586364061
transform 1 0 19412 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19596 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19228 0 -1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_6  FILLER_26_206
timestamp 1586364061
transform 1 0 20056 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20424 0 1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 21988 0 1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _147_
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 21804 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21436 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_224
timestamp 1586364061
transform 1 0 21712 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_26_229
timestamp 1586364061
transform 1 0 22172 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_219
timestamp 1586364061
transform 1 0 21252 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_223
timestamp 1586364061
transform 1 0 21620 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _118_
timestamp 1586364061
transform 1 0 22448 0 -1 16864
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_241
timestamp 1586364061
transform 1 0 23276 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_236
timestamp 1586364061
transform 1 0 22816 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_248
timestamp 1586364061
transform 1 0 23920 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_253
timestamp 1586364061
transform 1 0 24380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_26_265
timestamp 1586364061
transform 1 0 25484 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_12  FILLER_27_252
timestamp 1586364061
transform 1 0 24288 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_264
timestamp 1586364061
transform 1 0 25392 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_273
timestamp 1586364061
transform 1 0 26220 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_27_276
timestamp 1586364061
transform 1 0 26496 0 1 16864
box -38 -48 130 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_4  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4416 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_47
timestamp 1586364061
transform 1 0 5428 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_51
timestamp 1586364061
transform 1 0 5796 0 -1 17952
box -38 -48 406 592
use scs8hd_inv_8  _194_
timestamp 1586364061
transform 1 0 6164 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_64
timestamp 1586364061
transform 1 0 6992 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_71
timestamp 1586364061
transform 1 0 7636 0 -1 17952
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_8  FILLER_28_84
timestamp 1586364061
transform 1 0 8832 0 -1 17952
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_102
timestamp 1586364061
transform 1 0 10488 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_106
timestamp 1586364061
transform 1 0 10856 0 -1 17952
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_4_.latch
timestamp 1586364061
transform 1 0 11408 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11224 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_123
timestamp 1586364061
transform 1 0 12420 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 13616 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 12604 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_127
timestamp 1586364061
transform 1 0 12788 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_131
timestamp 1586364061
transform 1 0 13156 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_135
timestamp 1586364061
transform 1 0 13524 0 -1 17952
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_3_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_145
timestamp 1586364061
transform 1 0 14444 0 -1 17952
box -38 -48 590 592
use scs8hd_decap_12  FILLER_28_165
timestamp 1586364061
transform 1 0 16284 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_28_177
timestamp 1586364061
transform 1 0 17388 0 -1 17952
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_4_.latch
timestamp 1586364061
transform 1 0 18308 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18032 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_183
timestamp 1586364061
transform 1 0 17940 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_186
timestamp 1586364061
transform 1 0 18216 0 -1 17952
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19872 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19504 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20424 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_198
timestamp 1586364061
transform 1 0 19320 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_202
timestamp 1586364061
transform 1 0 19688 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_206
timestamp 1586364061
transform 1 0 20056 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_212
timestamp 1586364061
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_12  FILLER_28_224
timestamp 1586364061
transform 1 0 21712 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_236
timestamp 1586364061
transform 1 0 22816 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_248
timestamp 1586364061
transform 1 0 23920 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_260
timestamp 1586364061
transform 1 0 25024 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_28_272
timestamp 1586364061
transform 1 0 26128 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 774 592
use scs8hd_inv_8  _193_
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 3404 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_23
timestamp 1586364061
transform 1 0 3220 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_36
timestamp 1586364061
transform 1 0 4416 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_40
timestamp 1586364061
transform 1 0 4784 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_53
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_57
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 406 592
use scs8hd_decap_3  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8832 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8648 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8280 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_76
timestamp 1586364061
transform 1 0 8096 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_80
timestamp 1586364061
transform 1 0 8464 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10028 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_95
timestamp 1586364061
transform 1 0 9844 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_99
timestamp 1586364061
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _156_
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_112
timestamp 1586364061
transform 1 0 11408 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 14168 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13984 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_132
timestamp 1586364061
transform 1 0 13248 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_138
timestamp 1586364061
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15548 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15180 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_151
timestamp 1586364061
transform 1 0 14996 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_155
timestamp 1586364061
transform 1 0 15364 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 17112 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 16744 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_168
timestamp 1586364061
transform 1 0 16560 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_172
timestamp 1586364061
transform 1 0 16928 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_176
timestamp 1586364061
transform 1 0 17296 0 1 17952
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_180
timestamp 1586364061
transform 1 0 17664 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_195
timestamp 1586364061
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19872 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19688 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_199
timestamp 1586364061
transform 1 0 19412 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_213
timestamp 1586364061
transform 1 0 20700 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 20884 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 21252 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_217
timestamp 1586364061
transform 1 0 21068 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_221
timestamp 1586364061
transform 1 0 21436 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_29_233
timestamp 1586364061
transform 1 0 22540 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  FILLER_29_241
timestamp 1586364061
transform 1 0 23276 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 774 592
use scs8hd_buf_2  _244_
timestamp 1586364061
transform 1 0 24564 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__244__A
timestamp 1586364061
transform 1 0 25116 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_253
timestamp 1586364061
transform 1 0 24380 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_259
timestamp 1586364061
transform 1 0 24932 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_263
timestamp 1586364061
transform 1 0 25300 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_275
timestamp 1586364061
transform 1 0 26404 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 406 592
use scs8hd_conb_1  _212_
timestamp 1586364061
transform 1 0 2944 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_19
timestamp 1586364061
transform 1 0 2852 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_23
timestamp 1586364061
transform 1 0 3220 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_4  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4508 0 -1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5520 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5336 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_36
timestamp 1586364061
transform 1 0 4416 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_40
timestamp 1586364061
transform 1 0 4784 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 6900 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_57
timestamp 1586364061
transform 1 0 6348 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_2  FILLER_30_65
timestamp 1586364061
transform 1 0 7084 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8832 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_78
timestamp 1586364061
transform 1 0 8280 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_82
timestamp 1586364061
transform 1 0 8648 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_86
timestamp 1586364061
transform 1 0 9016 0 -1 19040
box -38 -48 590 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_96
timestamp 1586364061
transform 1 0 9936 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_101
timestamp 1586364061
transform 1 0 10396 0 -1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _158_
timestamp 1586364061
transform 1 0 12328 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_8  FILLER_30_114
timestamp 1586364061
transform 1 0 11592 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13984 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13340 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_131
timestamp 1586364061
transform 1 0 13156 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_135
timestamp 1586364061
transform 1 0 13524 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_139
timestamp 1586364061
transform 1 0 13892 0 -1 19040
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 14444 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_143
timestamp 1586364061
transform 1 0 14260 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_147
timestamp 1586364061
transform 1 0 14628 0 -1 19040
box -38 -48 406 592
use scs8hd_nor2_4  _152_
timestamp 1586364061
transform 1 0 17112 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16652 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_163
timestamp 1586364061
transform 1 0 16100 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_167
timestamp 1586364061
transform 1 0 16468 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_171
timestamp 1586364061
transform 1 0 16836 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 18124 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18492 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_183
timestamp 1586364061
transform 1 0 17940 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_187
timestamp 1586364061
transform 1 0 18308 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_191
timestamp 1586364061
transform 1 0 18676 0 -1 19040
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_206
timestamp 1586364061
transform 1 0 20056 0 -1 19040
box -38 -48 774 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_12  FILLER_30_224
timestamp 1586364061
transform 1 0 21712 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_236
timestamp 1586364061
transform 1 0 22816 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_248
timestamp 1586364061
transform 1 0 23920 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_260
timestamp 1586364061
transform 1 0 25024 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  FILLER_30_272
timestamp 1586364061
transform 1 0 26128 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_buf_2  _245_
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__245__A
timestamp 1586364061
transform 1 0 1932 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_7
timestamp 1586364061
transform 1 0 1748 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_11
timestamp 1586364061
transform 1 0 2116 0 1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3956 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3404 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_23
timestamp 1586364061
transform 1 0 3220 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_34
timestamp 1586364061
transform 1 0 4232 0 1 19040
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4968 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_40
timestamp 1586364061
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 406 592
use scs8hd_nor2_4  _157_
timestamp 1586364061
transform 1 0 6900 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_57
timestamp 1586364061
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8464 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8280 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_72
timestamp 1586364061
transform 1 0 7728 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_76
timestamp 1586364061
transform 1 0 8096 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_89
timestamp 1586364061
transform 1 0 9292 0 1 19040
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_2_.latch
timestamp 1586364061
transform 1 0 10580 0 1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10028 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9660 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_95
timestamp 1586364061
transform 1 0 9844 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_99
timestamp 1586364061
transform 1 0 10212 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_114
timestamp 1586364061
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_118
timestamp 1586364061
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 14076 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_132
timestamp 1586364061
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_136
timestamp 1586364061
transform 1 0 13616 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_140
timestamp 1586364061
transform 1 0 13984 0 1 19040
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_2_.latch
timestamp 1586364061
transform 1 0 14260 0 1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15456 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_154
timestamp 1586364061
transform 1 0 15272 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_158
timestamp 1586364061
transform 1 0 15640 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16008 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17020 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_171
timestamp 1586364061
transform 1 0 16836 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_175
timestamp 1586364061
transform 1 0 17204 0 1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_179
timestamp 1586364061
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_195
timestamp 1586364061
transform 1 0 19044 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19780 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19596 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_199
timestamp 1586364061
transform 1 0 19412 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_212
timestamp 1586364061
transform 1 0 20608 0 1 19040
box -38 -48 314 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_217
timestamp 1586364061
transform 1 0 21068 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_229
timestamp 1586364061
transform 1 0 22172 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_3  FILLER_31_241
timestamp 1586364061
transform 1 0 23276 0 1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__239__A
timestamp 1586364061
transform 1 0 24564 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_253
timestamp 1586364061
transform 1 0 24380 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_257
timestamp 1586364061
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_31_269
timestamp 1586364061
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_6  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4600 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_47
timestamp 1586364061
transform 1 0 5428 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_51
timestamp 1586364061
transform 1 0 5796 0 -1 20128
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6164 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_58
timestamp 1586364061
transform 1 0 6440 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_32_70
timestamp 1586364061
transform 1 0 7544 0 -1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7912 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7728 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_83
timestamp 1586364061
transform 1 0 8740 0 -1 20128
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10028 0 -1 20128
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_91
timestamp 1586364061
transform 1 0 9476 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11776 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11224 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_108
timestamp 1586364061
transform 1 0 11040 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_112
timestamp 1586364061
transform 1 0 11408 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_4  FILLER_32_119
timestamp 1586364061
transform 1 0 12052 0 -1 20128
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 13248 0 -1 20128
box -38 -48 1050 592
use scs8hd_decap_6  FILLER_32_125
timestamp 1586364061
transform 1 0 12604 0 -1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_32_131
timestamp 1586364061
transform 1 0 13156 0 -1 20128
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14444 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_143
timestamp 1586364061
transform 1 0 14260 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_147
timestamp 1586364061
transform 1 0 14628 0 -1 20128
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_163
timestamp 1586364061
transform 1 0 16100 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  FILLER_32_168
timestamp 1586364061
transform 1 0 16560 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_32_174
timestamp 1586364061
transform 1 0 17112 0 -1 20128
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_2_.latch
timestamp 1586364061
transform 1 0 17940 0 -1 20128
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_32_182
timestamp 1586364061
transform 1 0 17848 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_194
timestamp 1586364061
transform 1 0 18952 0 -1 20128
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19320 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20148 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_200
timestamp 1586364061
transform 1 0 19504 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_205
timestamp 1586364061
transform 1 0 19964 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_209
timestamp 1586364061
transform 1 0 20332 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_213
timestamp 1586364061
transform 1 0 20700 0 -1 20128
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 21344 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 21712 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_218
timestamp 1586364061
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_222
timestamp 1586364061
transform 1 0 21528 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_226
timestamp 1586364061
transform 1 0 21896 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_238
timestamp 1586364061
transform 1 0 23000 0 -1 20128
box -38 -48 1142 592
use scs8hd_buf_2  _239_
timestamp 1586364061
transform 1 0 24564 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_4  FILLER_32_250
timestamp 1586364061
transform 1 0 24104 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_254
timestamp 1586364061
transform 1 0 24472 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_259
timestamp 1586364061
transform 1 0 24932 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_271
timestamp 1586364061
transform 1 0 26036 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_7
timestamp 1586364061
transform 1 0 1748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_6
timestamp 1586364061
transform 1 0 1656 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_2  _243_
timestamp 1586364061
transform 1 0 3864 0 1 20128
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_19
timestamp 1586364061
transform 1 0 2852 0 1 20128
box -38 -48 774 592
use scs8hd_decap_3  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_34
timestamp 1586364061
transform 1 0 4232 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_18
timestamp 1586364061
transform 1 0 2760 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_34_30
timestamp 1586364061
transform 1 0 3864 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__243__A
timestamp 1586364061
transform 1 0 4416 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_38
timestamp 1586364061
transform 1 0 4600 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_50
timestamp 1586364061
transform 1 0 5704 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7636 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_33_58
timestamp 1586364061
transform 1 0 6440 0 1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_33_70
timestamp 1586364061
transform 1 0 7544 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_34_76
timestamp 1586364061
transform 1 0 8096 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_78
timestamp 1586364061
transform 1 0 8280 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 8464 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8096 0 1 20128
box -38 -48 222 592
use scs8hd_conb_1  _215_
timestamp 1586364061
transform 1 0 8280 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_6  FILLER_34_85
timestamp 1586364061
transform 1 0 8924 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_2  FILLER_34_81
timestamp 1586364061
transform 1 0 8556 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 8740 0 -1 21216
box -38 -48 222 592
use scs8hd_nor2_4  _160_
timestamp 1586364061
transform 1 0 8648 0 1 20128
box -38 -48 866 592
use scs8hd_decap_3  FILLER_34_96
timestamp 1586364061
transform 1 0 9936 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_1  FILLER_34_91
timestamp 1586364061
transform 1 0 9476 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_95
timestamp 1586364061
transform 1 0 9844 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_91
timestamp 1586364061
transform 1 0 9476 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 10028 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_34_101
timestamp 1586364061
transform 1 0 10396 0 -1 21216
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 10212 0 -1 21216
box -38 -48 222 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 10212 0 1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_109
timestamp 1586364061
transform 1 0 11132 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_113
timestamp 1586364061
transform 1 0 11500 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_108
timestamp 1586364061
transform 1 0 11040 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11316 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_124
timestamp 1586364061
transform 1 0 12512 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_34_120
timestamp 1586364061
transform 1 0 12144 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_6  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_33_121
timestamp 1586364061
transform 1 0 12236 0 1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_117
timestamp 1586364061
transform 1 0 11868 0 1 20128
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11316 0 -1 21216
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13156 0 1 20128
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12972 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 12604 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13156 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_142
timestamp 1586364061
transform 1 0 14168 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_127
timestamp 1586364061
transform 1 0 12788 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_3  FILLER_34_133
timestamp 1586364061
transform 1 0 13340 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_149
timestamp 1586364061
transform 1 0 14812 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_145
timestamp 1586364061
transform 1 0 14444 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_146
timestamp 1586364061
transform 1 0 14536 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14720 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14352 0 1 20128
box -38 -48 222 592
use scs8hd_conb_1  _219_
timestamp 1586364061
transform 1 0 14904 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_157
timestamp 1586364061
transform 1 0 15548 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_153
timestamp 1586364061
transform 1 0 15180 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15364 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 866 592
use scs8hd_decap_4  FILLER_34_167
timestamp 1586364061
transform 1 0 16468 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_163
timestamp 1586364061
transform 1 0 16100 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_161
timestamp 1586364061
transform 1 0 15916 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_175
timestamp 1586364061
transform 1 0 17204 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_34_174
timestamp 1586364061
transform 1 0 17112 0 -1 21216
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 20128
box -38 -48 866 592
use scs8hd_fill_1  FILLER_34_186
timestamp 1586364061
transform 1 0 18216 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_179
timestamp 1586364061
transform 1 0 17572 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_conb_1  _216_
timestamp 1586364061
transform 1 0 18308 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_194
timestamp 1586364061
transform 1 0 18952 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_190
timestamp 1586364061
transform 1 0 18584 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18768 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_196
timestamp 1586364061
transform 1 0 19136 0 -1 21216
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18308 0 -1 21216
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19320 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20700 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20332 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_207
timestamp 1586364061
transform 1 0 20148 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_211
timestamp 1586364061
transform 1 0 20516 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_34_208
timestamp 1586364061
transform 1 0 20240 0 -1 21216
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 1 20128
box -38 -48 866 592
use scs8hd_decap_12  FILLER_33_224
timestamp 1586364061
transform 1 0 21712 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_236
timestamp 1586364061
transform 1 0 22816 0 1 20128
box -38 -48 774 592
use scs8hd_decap_8  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_253
timestamp 1586364061
transform 1 0 24380 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_258
timestamp 1586364061
transform 1 0 24840 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_decap_4  FILLER_34_270
timestamp 1586364061
transform 1 0 25944 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_274
timestamp 1586364061
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_86
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_110
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 590 592
use scs8hd_fill_2  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 222 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 12604 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14168 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_134
timestamp 1586364061
transform 1 0 13432 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_138
timestamp 1586364061
transform 1 0 13800 0 1 21216
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14352 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15364 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_153
timestamp 1586364061
transform 1 0 15180 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_157
timestamp 1586364061
transform 1 0 15548 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16928 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_170
timestamp 1586364061
transform 1 0 16744 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_174
timestamp 1586364061
transform 1 0 17112 0 1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18492 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18308 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_179
timestamp 1586364061
transform 1 0 17572 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19504 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_198
timestamp 1586364061
transform 1 0 19320 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_202
timestamp 1586364061
transform 1 0 19688 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_214
timestamp 1586364061
transform 1 0 20792 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_226
timestamp 1586364061
transform 1 0 21896 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_238
timestamp 1586364061
transform 1 0 23000 0 1 21216
box -38 -48 590 592
use scs8hd_decap_8  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 774 592
use scs8hd_buf_2  _238_
timestamp 1586364061
transform 1 0 24564 0 1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__238__A
timestamp 1586364061
transform 1 0 25116 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_253
timestamp 1586364061
transform 1 0 24380 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_259
timestamp 1586364061
transform 1 0 24932 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_263
timestamp 1586364061
transform 1 0 25300 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_275
timestamp 1586364061
transform 1 0 26404 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_36_117
timestamp 1586364061
transform 1 0 11868 0 -1 22304
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12604 0 -1 22304
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_128
timestamp 1586364061
transform 1 0 12880 0 -1 22304
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15364 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_36_145
timestamp 1586364061
transform 1 0 14444 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_1  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_36_164
timestamp 1586364061
transform 1 0 16192 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_12  FILLER_36_175
timestamp 1586364061
transform 1 0 17204 0 -1 22304
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18308 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_12  FILLER_36_196
timestamp 1586364061
transform 1 0 19136 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_6  FILLER_36_208
timestamp 1586364061
transform 1 0 20240 0 -1 22304
box -38 -48 590 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_6
timestamp 1586364061
transform 1 0 1656 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_10
timestamp 1586364061
transform 1 0 2024 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_14
timestamp 1586364061
transform 1 0 2392 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_26
timestamp 1586364061
transform 1 0 3496 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_38
timestamp 1586364061
transform 1 0 4600 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_50
timestamp 1586364061
transform 1 0 5704 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_37_58
timestamp 1586364061
transform 1 0 6440 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_37_80
timestamp 1586364061
transform 1 0 8464 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_83
timestamp 1586364061
transform 1 0 8740 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_95
timestamp 1586364061
transform 1 0 9844 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_107
timestamp 1586364061
transform 1 0 10948 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_119
timestamp 1586364061
transform 1 0 12052 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 314 592
use scs8hd_nor2_4  _122_
timestamp 1586364061
transform 1 0 12696 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 13708 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 14076 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_139
timestamp 1586364061
transform 1 0 13892 0 1 22304
box -38 -48 222 592
use scs8hd_buf_2  _233_
timestamp 1586364061
transform 1 0 14260 0 1 22304
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15364 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15180 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14812 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_147
timestamp 1586364061
transform 1 0 14628 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_151
timestamp 1586364061
transform 1 0 14996 0 1 22304
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_164
timestamp 1586364061
transform 1 0 16192 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_168
timestamp 1586364061
transform 1 0 16560 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_175
timestamp 1586364061
transform 1 0 17204 0 1 22304
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_179
timestamp 1586364061
transform 1 0 17572 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_187
timestamp 1586364061
transform 1 0 18308 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_191
timestamp 1586364061
transform 1 0 18676 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_203
timestamp 1586364061
transform 1 0 19780 0 1 22304
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_217
timestamp 1586364061
transform 1 0 21068 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_229
timestamp 1586364061
transform 1 0 22172 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_37_241
timestamp 1586364061
transform 1 0 23276 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_6
timestamp 1586364061
transform 1 0 1656 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_18
timestamp 1586364061
transform 1 0 2760 0 -1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_38_30
timestamp 1586364061
transform 1 0 3864 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_84
timestamp 1586364061
transform 1 0 8832 0 -1 23392
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_105
timestamp 1586364061
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_38_117
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 774 592
use scs8hd_nor2_4  _121_
timestamp 1586364061
transform 1 0 13524 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 12696 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_125
timestamp 1586364061
transform 1 0 12604 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_6  FILLER_38_128
timestamp 1586364061
transform 1 0 12880 0 -1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_38_134
timestamp 1586364061
transform 1 0 13432 0 -1 23392
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__233__A
timestamp 1586364061
transform 1 0 14536 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_144
timestamp 1586364061
transform 1 0 14352 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_148
timestamp 1586364061
transform 1 0 14720 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_152
timestamp 1586364061
transform 1 0 15088 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17020 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_38_165
timestamp 1586364061
transform 1 0 16284 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_38_176
timestamp 1586364061
transform 1 0 17296 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_188
timestamp 1586364061
transform 1 0 18400 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_200
timestamp 1586364061
transform 1 0 19504 0 -1 23392
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_38_212
timestamp 1586364061
transform 1 0 20608 0 -1 23392
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_218
timestamp 1586364061
transform 1 0 21160 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_230
timestamp 1586364061
transform 1 0 22264 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_242
timestamp 1586364061
transform 1 0 23368 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_254
timestamp 1586364061
transform 1 0 24472 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_38_266
timestamp 1586364061
transform 1 0 25576 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_274
timestamp 1586364061
transform 1 0 26312 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_6
timestamp 1586364061
transform 1 0 1656 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_10
timestamp 1586364061
transform 1 0 2024 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_22
timestamp 1586364061
transform 1 0 3128 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_34
timestamp 1586364061
transform 1 0 4232 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_46
timestamp 1586364061
transform 1 0 5336 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_4  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 406 592
use scs8hd_decap_3  FILLER_39_58
timestamp 1586364061
transform 1 0 6440 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_decap_3  FILLER_40_64
timestamp 1586364061
transform 1 0 6992 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_4  FILLER_39_69
timestamp 1586364061
transform 1 0 7452 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_66
timestamp 1586364061
transform 1 0 7176 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__227__A
timestamp 1586364061
transform 1 0 7268 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _227_
timestamp 1586364061
transform 1 0 7268 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_71
timestamp 1586364061
transform 1 0 7636 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _225_
timestamp 1586364061
transform 1 0 7820 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__225__A
timestamp 1586364061
transform 1 0 8372 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_77
timestamp 1586364061
transform 1 0 8188 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_81
timestamp 1586364061
transform 1 0 8556 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_40_83
timestamp 1586364061
transform 1 0 8740 0 -1 24480
box -38 -48 774 592
use scs8hd_buf_2  _222_
timestamp 1586364061
transform 1 0 10580 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_93
timestamp 1586364061
transform 1 0 9660 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_101
timestamp 1586364061
transform 1 0 10396 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_107
timestamp 1586364061
transform 1 0 10948 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_91
timestamp 1586364061
transform 1 0 9476 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11500 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__222__A
timestamp 1586364061
transform 1 0 11132 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11500 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_111
timestamp 1586364061
transform 1 0 11316 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_115
timestamp 1586364061
transform 1 0 11684 0 1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_39_121
timestamp 1586364061
transform 1 0 12236 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_116
timestamp 1586364061
transform 1 0 11776 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_135
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_128
timestamp 1586364061
transform 1 0 12880 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_140
timestamp 1586364061
transform 1 0 13984 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_147
timestamp 1586364061
transform 1 0 14628 0 1 23392
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_39_159
timestamp 1586364061
transform 1 0 15732 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_152
timestamp 1586364061
transform 1 0 15088 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15916 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16376 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_164
timestamp 1586364061
transform 1 0 16192 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_168
timestamp 1586364061
transform 1 0 16560 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_166
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_178
timestamp 1586364061
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _240_
timestamp 1586364061
transform 1 0 18124 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__240__A
timestamp 1586364061
transform 1 0 18676 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_180
timestamp 1586364061
transform 1 0 17664 0 1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_189
timestamp 1586364061
transform 1 0 18492 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_193
timestamp 1586364061
transform 1 0 18860 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_190
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20148 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20608 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_205
timestamp 1586364061
transform 1 0 19964 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_210
timestamp 1586364061
transform 1 0 20424 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_214
timestamp 1586364061
transform 1 0 20792 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_202
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_221
timestamp 1586364061
transform 1 0 21436 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_225
timestamp 1586364061
transform 1 0 21804 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_decap_6  FILLER_39_237
timestamp 1586364061
transform 1 0 22908 0 1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_39_243
timestamp 1586364061
transform 1 0 23460 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_248
timestamp 1586364061
transform 1 0 23920 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24656 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25116 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_252
timestamp 1586364061
transform 1 0 24288 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_259
timestamp 1586364061
transform 1 0 24932 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_263
timestamp 1586364061
transform 1 0 25300 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_251
timestamp 1586364061
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_263
timestamp 1586364061
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_275
timestamp 1586364061
transform 1 0 26404 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal3 s 27520 688 28000 808 6 address[0]
port 0 nsew default input
rlabel metal3 s 27520 2048 28000 2168 6 address[1]
port 1 nsew default input
rlabel metal2 s 662 27520 718 28000 6 address[2]
port 2 nsew default input
rlabel metal3 s 0 552 480 672 6 address[3]
port 3 nsew default input
rlabel metal3 s 0 1776 480 1896 6 address[4]
port 4 nsew default input
rlabel metal2 s 2042 27520 2098 28000 6 address[5]
port 5 nsew default input
rlabel metal2 s 3054 0 3110 480 6 address[6]
port 6 nsew default input
rlabel metal3 s 0 3136 480 3256 6 bottom_left_grid_pin_13_
port 7 nsew default input
rlabel metal3 s 27520 3408 28000 3528 6 bottom_right_grid_pin_11_
port 8 nsew default input
rlabel metal3 s 0 4496 480 4616 6 chanx_left_in[0]
port 9 nsew default input
rlabel metal2 s 3422 27520 3478 28000 6 chanx_left_in[1]
port 10 nsew default input
rlabel metal2 s 4802 27520 4858 28000 6 chanx_left_in[2]
port 11 nsew default input
rlabel metal3 s 0 5856 480 5976 6 chanx_left_in[3]
port 12 nsew default input
rlabel metal2 s 4342 0 4398 480 6 chanx_left_in[4]
port 13 nsew default input
rlabel metal2 s 5630 0 5686 480 6 chanx_left_in[5]
port 14 nsew default input
rlabel metal2 s 6182 27520 6238 28000 6 chanx_left_in[6]
port 15 nsew default input
rlabel metal3 s 27520 4768 28000 4888 6 chanx_left_in[7]
port 16 nsew default input
rlabel metal3 s 27520 6264 28000 6384 6 chanx_left_in[8]
port 17 nsew default input
rlabel metal2 s 6918 0 6974 480 6 chanx_left_out[0]
port 18 nsew default tristate
rlabel metal2 s 7654 27520 7710 28000 6 chanx_left_out[1]
port 19 nsew default tristate
rlabel metal3 s 27520 7624 28000 7744 6 chanx_left_out[2]
port 20 nsew default tristate
rlabel metal2 s 9034 27520 9090 28000 6 chanx_left_out[3]
port 21 nsew default tristate
rlabel metal3 s 27520 8984 28000 9104 6 chanx_left_out[4]
port 22 nsew default tristate
rlabel metal2 s 10414 27520 10470 28000 6 chanx_left_out[5]
port 23 nsew default tristate
rlabel metal2 s 11794 27520 11850 28000 6 chanx_left_out[6]
port 24 nsew default tristate
rlabel metal3 s 0 7216 480 7336 6 chanx_left_out[7]
port 25 nsew default tristate
rlabel metal3 s 0 8440 480 8560 6 chanx_left_out[8]
port 26 nsew default tristate
rlabel metal3 s 27520 10480 28000 10600 6 chanx_right_in[0]
port 27 nsew default input
rlabel metal2 s 8114 0 8170 480 6 chanx_right_in[1]
port 28 nsew default input
rlabel metal3 s 0 9800 480 9920 6 chanx_right_in[2]
port 29 nsew default input
rlabel metal2 s 9402 0 9458 480 6 chanx_right_in[3]
port 30 nsew default input
rlabel metal3 s 0 11160 480 11280 6 chanx_right_in[4]
port 31 nsew default input
rlabel metal2 s 13174 27520 13230 28000 6 chanx_right_in[5]
port 32 nsew default input
rlabel metal3 s 0 12520 480 12640 6 chanx_right_in[6]
port 33 nsew default input
rlabel metal3 s 0 13880 480 14000 6 chanx_right_in[7]
port 34 nsew default input
rlabel metal3 s 27520 11840 28000 11960 6 chanx_right_in[8]
port 35 nsew default input
rlabel metal3 s 27520 13200 28000 13320 6 chanx_right_out[0]
port 36 nsew default tristate
rlabel metal2 s 10690 0 10746 480 6 chanx_right_out[1]
port 37 nsew default tristate
rlabel metal2 s 11978 0 12034 480 6 chanx_right_out[2]
port 38 nsew default tristate
rlabel metal3 s 27520 14696 28000 14816 6 chanx_right_out[3]
port 39 nsew default tristate
rlabel metal2 s 14646 27520 14702 28000 6 chanx_right_out[4]
port 40 nsew default tristate
rlabel metal2 s 13266 0 13322 480 6 chanx_right_out[5]
port 41 nsew default tristate
rlabel metal3 s 27520 16056 28000 16176 6 chanx_right_out[6]
port 42 nsew default tristate
rlabel metal3 s 0 15104 480 15224 6 chanx_right_out[7]
port 43 nsew default tristate
rlabel metal2 s 14554 0 14610 480 6 chanx_right_out[8]
port 44 nsew default tristate
rlabel metal2 s 16026 27520 16082 28000 6 chany_bottom_in[0]
port 45 nsew default input
rlabel metal3 s 0 16464 480 16584 6 chany_bottom_in[1]
port 46 nsew default input
rlabel metal2 s 15750 0 15806 480 6 chany_bottom_in[2]
port 47 nsew default input
rlabel metal2 s 17406 27520 17462 28000 6 chany_bottom_in[3]
port 48 nsew default input
rlabel metal3 s 0 17824 480 17944 6 chany_bottom_in[4]
port 49 nsew default input
rlabel metal3 s 0 19184 480 19304 6 chany_bottom_in[5]
port 50 nsew default input
rlabel metal3 s 27520 17416 28000 17536 6 chany_bottom_in[6]
port 51 nsew default input
rlabel metal2 s 18786 27520 18842 28000 6 chany_bottom_in[7]
port 52 nsew default input
rlabel metal3 s 27520 18776 28000 18896 6 chany_bottom_in[8]
port 53 nsew default input
rlabel metal2 s 17038 0 17094 480 6 chany_bottom_out[0]
port 54 nsew default tristate
rlabel metal3 s 0 20544 480 20664 6 chany_bottom_out[1]
port 55 nsew default tristate
rlabel metal3 s 27520 20272 28000 20392 6 chany_bottom_out[2]
port 56 nsew default tristate
rlabel metal3 s 0 21768 480 21888 6 chany_bottom_out[3]
port 57 nsew default tristate
rlabel metal2 s 18326 0 18382 480 6 chany_bottom_out[4]
port 58 nsew default tristate
rlabel metal2 s 19614 0 19670 480 6 chany_bottom_out[5]
port 59 nsew default tristate
rlabel metal2 s 20166 27520 20222 28000 6 chany_bottom_out[6]
port 60 nsew default tristate
rlabel metal3 s 27520 21632 28000 21752 6 chany_bottom_out[7]
port 61 nsew default tristate
rlabel metal3 s 27520 22992 28000 23112 6 chany_bottom_out[8]
port 62 nsew default tristate
rlabel metal2 s 1766 0 1822 480 6 data_in
port 63 nsew default input
rlabel metal2 s 570 0 626 480 6 enable
port 64 nsew default input
rlabel metal3 s 0 23128 480 23248 6 left_bottom_grid_pin_12_
port 65 nsew default input
rlabel metal2 s 23386 0 23442 480 6 left_top_grid_pin_11_
port 66 nsew default input
rlabel metal2 s 23018 27520 23074 28000 6 left_top_grid_pin_13_
port 67 nsew default input
rlabel metal2 s 24398 27520 24454 28000 6 left_top_grid_pin_15_
port 68 nsew default input
rlabel metal2 s 20902 0 20958 480 6 left_top_grid_pin_1_
port 69 nsew default input
rlabel metal3 s 0 24488 480 24608 6 left_top_grid_pin_3_
port 70 nsew default input
rlabel metal3 s 27520 24488 28000 24608 6 left_top_grid_pin_5_
port 71 nsew default input
rlabel metal2 s 21638 27520 21694 28000 6 left_top_grid_pin_7_
port 72 nsew default input
rlabel metal2 s 22098 0 22154 480 6 left_top_grid_pin_9_
port 73 nsew default input
rlabel metal2 s 25778 27520 25834 28000 6 right_bottom_grid_pin_12_
port 74 nsew default input
rlabel metal2 s 27158 27520 27214 28000 6 right_top_grid_pin_11_
port 75 nsew default input
rlabel metal2 s 25962 0 26018 480 6 right_top_grid_pin_13_
port 76 nsew default input
rlabel metal2 s 27250 0 27306 480 6 right_top_grid_pin_15_
port 77 nsew default input
rlabel metal3 s 0 25848 480 25968 6 right_top_grid_pin_1_
port 78 nsew default input
rlabel metal3 s 27520 25848 28000 25968 6 right_top_grid_pin_3_
port 79 nsew default input
rlabel metal2 s 24674 0 24730 480 6 right_top_grid_pin_5_
port 80 nsew default input
rlabel metal3 s 27520 27208 28000 27328 6 right_top_grid_pin_7_
port 81 nsew default input
rlabel metal3 s 0 27208 480 27328 6 right_top_grid_pin_9_
port 82 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 83 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 84 nsew default input
<< end >>
