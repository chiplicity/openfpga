magic
tech EFS8A
magscale 1 2
timestamp 1603801159
<< locali >>
rect 9873 18207 9907 18377
rect 8493 13175 8527 13413
rect 2237 12155 2271 12325
<< viali >>
rect 16405 24361 16439 24395
rect 1444 24225 1478 24259
rect 16221 24225 16255 24259
rect 17392 24225 17426 24259
rect 1547 24021 1581 24055
rect 16773 24021 16807 24055
rect 17463 24021 17497 24055
rect 2237 23817 2271 23851
rect 13001 23817 13035 23851
rect 15485 23817 15519 23851
rect 17417 23817 17451 23851
rect 18245 23817 18279 23851
rect 23857 23817 23891 23851
rect 25329 23817 25363 23851
rect 1444 23613 1478 23647
rect 1869 23613 1903 23647
rect 12817 23613 12851 23647
rect 13369 23613 13403 23647
rect 15209 23613 15243 23647
rect 15301 23613 15335 23647
rect 18061 23613 18095 23647
rect 22512 23613 22546 23647
rect 22615 23613 22649 23647
rect 23673 23613 23707 23647
rect 24225 23613 24259 23647
rect 24844 23613 24878 23647
rect 1547 23545 1581 23579
rect 15945 23545 15979 23579
rect 16497 23545 16531 23579
rect 16589 23545 16623 23579
rect 17141 23545 17175 23579
rect 22937 23545 22971 23579
rect 16221 23477 16255 23511
rect 18705 23477 18739 23511
rect 24915 23477 24949 23511
rect 15623 23273 15657 23307
rect 21097 23273 21131 23307
rect 22661 23273 22695 23307
rect 16681 23205 16715 23239
rect 15520 23137 15554 23171
rect 18128 23137 18162 23171
rect 20913 23137 20947 23171
rect 22477 23137 22511 23171
rect 16589 23069 16623 23103
rect 16865 23069 16899 23103
rect 18199 23001 18233 23035
rect 17509 22729 17543 22763
rect 18613 22729 18647 22763
rect 16497 22593 16531 22627
rect 16773 22593 16807 22627
rect 14749 22525 14783 22559
rect 15485 22525 15519 22559
rect 15577 22457 15611 22491
rect 16589 22457 16623 22491
rect 20913 22457 20947 22491
rect 15853 22389 15887 22423
rect 16221 22389 16255 22423
rect 18061 22389 18095 22423
rect 22477 22389 22511 22423
rect 15485 22185 15519 22219
rect 17325 22185 17359 22219
rect 13369 22117 13403 22151
rect 16405 22117 16439 22151
rect 17969 22117 18003 22151
rect 19349 22049 19383 22083
rect 21833 22049 21867 22083
rect 13277 21981 13311 22015
rect 13921 21981 13955 22015
rect 16313 21981 16347 22015
rect 16589 21981 16623 22015
rect 17877 21981 17911 22015
rect 18153 21981 18187 22015
rect 16129 21913 16163 21947
rect 19533 21913 19567 21947
rect 22017 21913 22051 21947
rect 13093 21641 13127 21675
rect 15945 21641 15979 21675
rect 17509 21641 17543 21675
rect 19441 21641 19475 21675
rect 15255 21573 15289 21607
rect 13921 21505 13955 21539
rect 14933 21505 14967 21539
rect 16221 21505 16255 21539
rect 16497 21505 16531 21539
rect 1476 21437 1510 21471
rect 1869 21437 1903 21471
rect 15152 21437 15186 21471
rect 18153 21437 18187 21471
rect 19073 21437 19107 21471
rect 21833 21437 21867 21471
rect 13645 21369 13679 21403
rect 13737 21369 13771 21403
rect 15669 21369 15703 21403
rect 16313 21369 16347 21403
rect 1547 21301 1581 21335
rect 13461 21301 13495 21335
rect 17785 21301 17819 21335
rect 18337 21301 18371 21335
rect 13277 21097 13311 21131
rect 13645 21097 13679 21131
rect 13737 21097 13771 21131
rect 19395 21097 19429 21131
rect 10793 21029 10827 21063
rect 12357 21029 12391 21063
rect 12909 21029 12943 21063
rect 16313 21029 16347 21063
rect 17785 20961 17819 20995
rect 19324 20961 19358 20995
rect 10701 20893 10735 20927
rect 12265 20893 12299 20927
rect 16221 20893 16255 20927
rect 11253 20825 11287 20859
rect 16037 20825 16071 20859
rect 16773 20825 16807 20859
rect 14933 20757 14967 20791
rect 17969 20757 18003 20791
rect 18797 20757 18831 20791
rect 11897 20553 11931 20587
rect 13645 20553 13679 20587
rect 15853 20553 15887 20587
rect 16221 20553 16255 20587
rect 16589 20553 16623 20587
rect 16819 20553 16853 20587
rect 17877 20553 17911 20587
rect 10701 20417 10735 20451
rect 10793 20417 10827 20451
rect 18337 20417 18371 20451
rect 18613 20417 18647 20451
rect 19257 20417 19291 20451
rect 20821 20417 20855 20451
rect 10333 20349 10367 20383
rect 11437 20349 11471 20383
rect 12725 20349 12759 20383
rect 14933 20349 14967 20383
rect 16716 20349 16750 20383
rect 17141 20349 17175 20383
rect 19844 20349 19878 20383
rect 20269 20349 20303 20383
rect 12173 20281 12207 20315
rect 13046 20281 13080 20315
rect 14749 20281 14783 20315
rect 15254 20281 15288 20315
rect 18429 20281 18463 20315
rect 13921 20213 13955 20247
rect 19947 20213 19981 20247
rect 10701 20009 10735 20043
rect 12817 20009 12851 20043
rect 13461 20009 13495 20043
rect 13921 20009 13955 20043
rect 16221 20009 16255 20043
rect 17785 20009 17819 20043
rect 12218 19941 12252 19975
rect 15622 19941 15656 19975
rect 18038 19941 18072 19975
rect 18613 19941 18647 19975
rect 9908 19873 9942 19907
rect 10885 19873 10919 19907
rect 13737 19873 13771 19907
rect 19508 19873 19542 19907
rect 11897 19805 11931 19839
rect 15301 19805 15335 19839
rect 17417 19805 17451 19839
rect 17969 19805 18003 19839
rect 11069 19737 11103 19771
rect 10011 19669 10045 19703
rect 11437 19669 11471 19703
rect 13093 19669 13127 19703
rect 14749 19669 14783 19703
rect 16589 19669 16623 19703
rect 19579 19669 19613 19703
rect 9873 19465 9907 19499
rect 11989 19465 12023 19499
rect 15485 19465 15519 19499
rect 16037 19465 16071 19499
rect 17141 19465 17175 19499
rect 17509 19465 17543 19499
rect 14841 19397 14875 19431
rect 18429 19329 18463 19363
rect 1444 19261 1478 19295
rect 1869 19261 1903 19295
rect 7088 19261 7122 19295
rect 8284 19261 8318 19295
rect 8677 19261 8711 19295
rect 9137 19261 9171 19295
rect 9296 19261 9330 19295
rect 11345 19261 11379 19295
rect 12484 19261 12518 19295
rect 14197 19261 14231 19295
rect 14473 19261 14507 19295
rect 14841 19261 14875 19295
rect 16221 19261 16255 19295
rect 19165 19261 19199 19295
rect 19717 19261 19751 19295
rect 21224 19261 21258 19295
rect 21649 19261 21683 19295
rect 24660 19261 24694 19295
rect 25053 19261 25087 19295
rect 13001 19193 13035 19227
rect 13921 19193 13955 19227
rect 16542 19193 16576 19227
rect 18153 19193 18187 19227
rect 18245 19193 18279 19227
rect 19625 19193 19659 19227
rect 1547 19125 1581 19159
rect 7159 19125 7193 19159
rect 7573 19125 7607 19159
rect 8355 19125 8389 19159
rect 9367 19125 9401 19159
rect 10333 19125 10367 19159
rect 10977 19125 11011 19159
rect 11529 19125 11563 19159
rect 12587 19125 12621 19159
rect 13553 19125 13587 19159
rect 17877 19125 17911 19159
rect 19533 19125 19567 19159
rect 21327 19125 21361 19159
rect 24731 19125 24765 19159
rect 12127 18921 12161 18955
rect 16681 18921 16715 18955
rect 18613 18921 18647 18955
rect 21833 18921 21867 18955
rect 7573 18853 7607 18887
rect 10517 18853 10551 18887
rect 10609 18853 10643 18887
rect 16082 18853 16116 18887
rect 17417 18853 17451 18887
rect 17601 18853 17635 18887
rect 17693 18853 17727 18887
rect 18245 18853 18279 18887
rect 24731 18853 24765 18887
rect 6412 18785 6446 18819
rect 12056 18785 12090 18819
rect 13553 18785 13587 18819
rect 13921 18785 13955 18819
rect 14105 18785 14139 18819
rect 19073 18785 19107 18819
rect 19533 18785 19567 18819
rect 20948 18785 20982 18819
rect 24628 18785 24662 18819
rect 6515 18717 6549 18751
rect 7481 18717 7515 18751
rect 7757 18717 7791 18751
rect 10793 18717 10827 18751
rect 14381 18717 14415 18751
rect 15761 18717 15795 18751
rect 19625 18717 19659 18751
rect 10333 18581 10367 18615
rect 11897 18581 11931 18615
rect 12449 18581 12483 18615
rect 12909 18581 12943 18615
rect 14749 18581 14783 18615
rect 15485 18581 15519 18615
rect 20085 18581 20119 18615
rect 21051 18581 21085 18615
rect 21465 18581 21499 18615
rect 5641 18377 5675 18411
rect 6469 18377 6503 18411
rect 8401 18377 8435 18411
rect 9781 18377 9815 18411
rect 9873 18377 9907 18411
rect 14565 18377 14599 18411
rect 16129 18377 16163 18411
rect 16497 18377 16531 18411
rect 19165 18377 19199 18411
rect 24685 18377 24719 18411
rect 7481 18241 7515 18275
rect 8769 18241 8803 18275
rect 15485 18309 15519 18343
rect 10333 18241 10367 18275
rect 11897 18241 11931 18275
rect 20913 18241 20947 18275
rect 21465 18241 21499 18275
rect 21741 18241 21775 18275
rect 5800 18173 5834 18207
rect 9229 18173 9263 18207
rect 9873 18173 9907 18207
rect 10977 18173 11011 18207
rect 12449 18173 12483 18207
rect 12909 18173 12943 18207
rect 13461 18173 13495 18207
rect 13645 18173 13679 18207
rect 14749 18173 14783 18207
rect 15209 18173 15243 18207
rect 15577 18173 15611 18207
rect 16681 18173 16715 18207
rect 17141 18173 17175 18207
rect 18337 18173 18371 18207
rect 18521 18173 18555 18207
rect 18797 18173 18831 18207
rect 19625 18173 19659 18207
rect 7297 18105 7331 18139
rect 7573 18105 7607 18139
rect 8125 18105 8159 18139
rect 10425 18105 10459 18139
rect 19946 18105 19980 18139
rect 21557 18105 21591 18139
rect 5871 18037 5905 18071
rect 9413 18037 9447 18071
rect 10149 18037 10183 18071
rect 11529 18037 11563 18071
rect 12265 18037 12299 18071
rect 12725 18037 12759 18071
rect 14289 18037 14323 18071
rect 16865 18037 16899 18071
rect 17877 18037 17911 18071
rect 19533 18037 19567 18071
rect 20545 18037 20579 18071
rect 8125 17833 8159 17867
rect 10793 17833 10827 17867
rect 11069 17833 11103 17867
rect 12449 17833 12483 17867
rect 13921 17833 13955 17867
rect 16957 17833 16991 17867
rect 17509 17833 17543 17867
rect 18889 17833 18923 17867
rect 19993 17833 20027 17867
rect 5641 17765 5675 17799
rect 5733 17765 5767 17799
rect 7205 17765 7239 17799
rect 7297 17765 7331 17799
rect 7849 17765 7883 17799
rect 9781 17765 9815 17799
rect 9873 17765 9907 17799
rect 10425 17765 10459 17799
rect 16358 17765 16392 17799
rect 19394 17765 19428 17799
rect 21097 17765 21131 17799
rect 2120 17697 2154 17731
rect 4604 17697 4638 17731
rect 12265 17697 12299 17731
rect 12909 17697 12943 17731
rect 13185 17697 13219 17731
rect 13553 17697 13587 17731
rect 17785 17697 17819 17731
rect 16037 17629 16071 17663
rect 19073 17629 19107 17663
rect 20729 17629 20763 17663
rect 21005 17629 21039 17663
rect 22477 17629 22511 17663
rect 1685 17561 1719 17595
rect 6193 17561 6227 17595
rect 20361 17561 20395 17595
rect 21557 17561 21591 17595
rect 2191 17493 2225 17527
rect 4675 17493 4709 17527
rect 5273 17493 5307 17527
rect 6929 17493 6963 17527
rect 12081 17493 12115 17527
rect 14289 17493 14323 17527
rect 14749 17493 14783 17527
rect 15853 17493 15887 17527
rect 17969 17493 18003 17527
rect 18337 17493 18371 17527
rect 4077 17289 4111 17323
rect 4629 17289 4663 17323
rect 6285 17289 6319 17323
rect 7757 17289 7791 17323
rect 8033 17289 8067 17323
rect 10793 17289 10827 17323
rect 11529 17289 11563 17323
rect 11805 17289 11839 17323
rect 13645 17289 13679 17323
rect 15209 17289 15243 17323
rect 15945 17289 15979 17323
rect 18613 17289 18647 17323
rect 18981 17289 19015 17323
rect 20729 17289 20763 17323
rect 22293 17289 22327 17323
rect 23029 17289 23063 17323
rect 20085 17221 20119 17255
rect 12817 17153 12851 17187
rect 21005 17153 21039 17187
rect 21649 17153 21683 17187
rect 1409 17085 1443 17119
rect 3592 17085 3626 17119
rect 5181 17085 5215 17119
rect 5641 17085 5675 17119
rect 6837 17085 6871 17119
rect 8861 17085 8895 17119
rect 9873 17085 9907 17119
rect 14013 17085 14047 17119
rect 14381 17085 14415 17119
rect 14565 17085 14599 17119
rect 14933 17085 14967 17119
rect 16037 17085 16071 17119
rect 18061 17085 18095 17119
rect 19165 17085 19199 17119
rect 22544 17085 22578 17119
rect 23708 17085 23742 17119
rect 24720 17085 24754 17119
rect 25145 17085 25179 17119
rect 5917 17017 5951 17051
rect 6653 17017 6687 17051
rect 7199 17017 7233 17051
rect 10194 17017 10228 17051
rect 12541 17017 12575 17051
rect 12633 17017 12667 17051
rect 16358 17017 16392 17051
rect 17509 17017 17543 17051
rect 19486 17017 19520 17051
rect 21097 17017 21131 17051
rect 24133 17017 24167 17051
rect 1593 16949 1627 16983
rect 2145 16949 2179 16983
rect 2513 16949 2547 16983
rect 3663 16949 3697 16983
rect 5089 16949 5123 16983
rect 9045 16949 9079 16983
rect 9413 16949 9447 16983
rect 9781 16949 9815 16983
rect 11069 16949 11103 16983
rect 12173 16949 12207 16983
rect 15577 16949 15611 16983
rect 16957 16949 16991 16983
rect 17785 16949 17819 16983
rect 18245 16949 18279 16983
rect 20453 16949 20487 16983
rect 21925 16949 21959 16983
rect 22615 16949 22649 16983
rect 23811 16949 23845 16983
rect 24823 16949 24857 16983
rect 1593 16745 1627 16779
rect 3341 16745 3375 16779
rect 5917 16745 5951 16779
rect 7021 16745 7055 16779
rect 7665 16745 7699 16779
rect 9413 16745 9447 16779
rect 10333 16745 10367 16779
rect 12081 16745 12115 16779
rect 13093 16745 13127 16779
rect 16037 16745 16071 16779
rect 19901 16745 19935 16779
rect 22661 16745 22695 16779
rect 24685 16745 24719 16779
rect 2651 16677 2685 16711
rect 6463 16677 6497 16711
rect 8211 16677 8245 16711
rect 11482 16677 11516 16711
rect 12725 16677 12759 16711
rect 14381 16677 14415 16711
rect 16681 16677 16715 16711
rect 19302 16677 19336 16711
rect 20177 16677 20211 16711
rect 20729 16677 20763 16711
rect 21005 16677 21039 16711
rect 21097 16677 21131 16711
rect 21649 16677 21683 16711
rect 1409 16609 1443 16643
rect 2548 16609 2582 16643
rect 2973 16609 3007 16643
rect 4537 16609 4571 16643
rect 5089 16609 5123 16643
rect 5273 16609 5307 16643
rect 7849 16609 7883 16643
rect 8769 16609 8803 16643
rect 10149 16609 10183 16643
rect 12449 16609 12483 16643
rect 13645 16609 13679 16643
rect 13921 16609 13955 16643
rect 15301 16609 15335 16643
rect 22477 16609 22511 16643
rect 23489 16609 23523 16643
rect 24501 16609 24535 16643
rect 6101 16541 6135 16575
rect 11161 16541 11195 16575
rect 16589 16541 16623 16575
rect 18981 16541 19015 16575
rect 13737 16473 13771 16507
rect 17141 16473 17175 16507
rect 5549 16405 5583 16439
rect 7297 16405 7331 16439
rect 9965 16405 9999 16439
rect 10701 16405 10735 16439
rect 15485 16405 15519 16439
rect 18337 16405 18371 16439
rect 1593 16201 1627 16235
rect 2421 16201 2455 16235
rect 4077 16201 4111 16235
rect 6285 16201 6319 16235
rect 8309 16201 8343 16235
rect 10701 16201 10735 16235
rect 11529 16201 11563 16235
rect 15301 16201 15335 16235
rect 16773 16201 16807 16235
rect 17233 16201 17267 16235
rect 19349 16201 19383 16235
rect 21189 16201 21223 16235
rect 24777 16201 24811 16235
rect 6561 16133 6595 16167
rect 9321 16133 9355 16167
rect 20821 16133 20855 16167
rect 2605 16065 2639 16099
rect 7941 16065 7975 16099
rect 9689 16065 9723 16099
rect 9781 16065 9815 16099
rect 14841 16065 14875 16099
rect 18981 16065 19015 16099
rect 20177 16065 20211 16099
rect 23121 16065 23155 16099
rect 23765 16065 23799 16099
rect 25375 16065 25409 16099
rect 1409 15997 1443 16031
rect 4236 15997 4270 16031
rect 4629 15997 4663 16031
rect 5089 15997 5123 16031
rect 5181 15997 5215 16031
rect 5641 15997 5675 16031
rect 6837 15997 6871 16031
rect 7389 15997 7423 16031
rect 8769 15997 8803 16031
rect 12541 15997 12575 16031
rect 13645 15997 13679 16031
rect 14197 15997 14231 16031
rect 14657 15997 14691 16031
rect 15761 15997 15795 16031
rect 16221 15997 16255 16031
rect 18245 15997 18279 16031
rect 18705 15997 18739 16031
rect 21373 15997 21407 16031
rect 21833 15997 21867 16031
rect 22477 15997 22511 16031
rect 25272 15997 25306 16031
rect 25697 15997 25731 16031
rect 2697 15929 2731 15963
rect 3249 15929 3283 15963
rect 3709 15929 3743 15963
rect 5917 15929 5951 15963
rect 10102 15929 10136 15963
rect 11161 15929 11195 15963
rect 13185 15929 13219 15963
rect 15577 15929 15611 15963
rect 17785 15929 17819 15963
rect 19901 15929 19935 15963
rect 19993 15929 20027 15963
rect 23857 15929 23891 15963
rect 24409 15929 24443 15963
rect 2053 15861 2087 15895
rect 4307 15861 4341 15895
rect 6929 15861 6963 15895
rect 8677 15861 8711 15895
rect 8953 15861 8987 15895
rect 12173 15861 12207 15895
rect 14105 15861 14139 15895
rect 15853 15861 15887 15895
rect 19717 15861 19751 15895
rect 21465 15861 21499 15895
rect 23489 15861 23523 15895
rect 4721 15657 4755 15691
rect 6009 15657 6043 15691
rect 6561 15657 6595 15691
rect 7481 15657 7515 15691
rect 8309 15657 8343 15691
rect 9137 15657 9171 15691
rect 9965 15657 9999 15691
rect 10793 15657 10827 15691
rect 11529 15657 11563 15691
rect 14657 15657 14691 15691
rect 15761 15657 15795 15691
rect 16957 15657 16991 15691
rect 20729 15657 20763 15691
rect 24133 15657 24167 15691
rect 24777 15657 24811 15691
rect 2605 15589 2639 15623
rect 3157 15589 3191 15623
rect 6377 15589 6411 15623
rect 18245 15589 18279 15623
rect 18889 15589 18923 15623
rect 19435 15589 19469 15623
rect 21281 15589 21315 15623
rect 23121 15589 23155 15623
rect 23213 15589 23247 15623
rect 23765 15589 23799 15623
rect 1476 15521 1510 15555
rect 4813 15521 4847 15555
rect 5089 15521 5123 15555
rect 6561 15521 6595 15555
rect 7021 15521 7055 15555
rect 8033 15521 8067 15555
rect 8585 15521 8619 15555
rect 9781 15521 9815 15555
rect 10241 15521 10275 15555
rect 11253 15521 11287 15555
rect 11713 15521 11747 15555
rect 13277 15521 13311 15555
rect 13369 15521 13403 15555
rect 13553 15521 13587 15555
rect 16037 15521 16071 15555
rect 16405 15521 16439 15555
rect 17509 15521 17543 15555
rect 17969 15521 18003 15555
rect 19073 15521 19107 15555
rect 24593 15521 24627 15555
rect 2513 15453 2547 15487
rect 13829 15453 13863 15487
rect 16497 15453 16531 15487
rect 21189 15453 21223 15487
rect 21833 15453 21867 15487
rect 1547 15385 1581 15419
rect 1869 15317 1903 15351
rect 14381 15317 14415 15351
rect 18613 15317 18647 15351
rect 19993 15317 20027 15351
rect 22109 15317 22143 15351
rect 1777 15113 1811 15147
rect 8493 15113 8527 15147
rect 8953 15113 8987 15147
rect 10057 15113 10091 15147
rect 11713 15113 11747 15147
rect 14473 15113 14507 15147
rect 15669 15113 15703 15147
rect 17509 15113 17543 15147
rect 18245 15113 18279 15147
rect 19533 15113 19567 15147
rect 19901 15113 19935 15147
rect 21005 15113 21039 15147
rect 21281 15113 21315 15147
rect 23121 15113 23155 15147
rect 23489 15113 23523 15147
rect 24961 15113 24995 15147
rect 8033 15045 8067 15079
rect 9689 15045 9723 15079
rect 15025 15045 15059 15079
rect 19165 15045 19199 15079
rect 2329 14977 2363 15011
rect 2973 14977 3007 15011
rect 3893 14977 3927 15011
rect 4169 14977 4203 15011
rect 6929 14977 6963 15011
rect 9137 14977 9171 15011
rect 11161 14977 11195 15011
rect 13185 14977 13219 15011
rect 18613 14977 18647 15011
rect 20085 14977 20119 15011
rect 24041 14977 24075 15011
rect 5432 14909 5466 14943
rect 10517 14909 10551 14943
rect 10793 14909 10827 14943
rect 11069 14909 11103 14943
rect 12725 14909 12759 14943
rect 14105 14909 14139 14943
rect 16037 14909 16071 14943
rect 16681 14909 16715 14943
rect 16865 14909 16899 14943
rect 21833 14909 21867 14943
rect 25513 14909 25547 14943
rect 26065 14909 26099 14943
rect 2421 14841 2455 14875
rect 3709 14841 3743 14875
rect 3985 14841 4019 14875
rect 5917 14841 5951 14875
rect 7021 14841 7055 14875
rect 7573 14841 7607 14875
rect 9229 14841 9263 14875
rect 17141 14841 17175 14875
rect 18705 14841 18739 14875
rect 20406 14841 20440 14875
rect 22154 14841 22188 14875
rect 24133 14841 24167 14875
rect 24685 14841 24719 14875
rect 2145 14773 2179 14807
rect 3249 14773 3283 14807
rect 4813 14773 4847 14807
rect 5181 14773 5215 14807
rect 5503 14773 5537 14807
rect 6561 14773 6595 14807
rect 12173 14773 12207 14807
rect 13553 14773 13587 14807
rect 13921 14773 13955 14807
rect 21741 14773 21775 14807
rect 22753 14773 22787 14807
rect 25697 14773 25731 14807
rect 1869 14569 1903 14603
rect 2329 14569 2363 14603
rect 3893 14569 3927 14603
rect 5365 14569 5399 14603
rect 7481 14569 7515 14603
rect 9045 14569 9079 14603
rect 10609 14569 10643 14603
rect 11345 14569 11379 14603
rect 12541 14569 12575 14603
rect 13369 14569 13403 14603
rect 15025 14569 15059 14603
rect 18521 14569 18555 14603
rect 19809 14569 19843 14603
rect 20177 14569 20211 14603
rect 21189 14569 21223 14603
rect 22385 14569 22419 14603
rect 2605 14501 2639 14535
rect 4786 14501 4820 14535
rect 6647 14501 6681 14535
rect 10051 14501 10085 14535
rect 11989 14501 12023 14535
rect 14381 14501 14415 14535
rect 14657 14501 14691 14535
rect 16221 14501 16255 14535
rect 18975 14501 19009 14535
rect 21786 14501 21820 14535
rect 23397 14501 23431 14535
rect 24869 14501 24903 14535
rect 24961 14501 24995 14535
rect 1460 14433 1494 14467
rect 4445 14433 4479 14467
rect 6285 14433 6319 14467
rect 8217 14433 8251 14467
rect 8493 14433 8527 14467
rect 9689 14433 9723 14467
rect 12081 14433 12115 14467
rect 12357 14433 12391 14467
rect 13645 14433 13679 14467
rect 13921 14433 13955 14467
rect 15669 14433 15703 14467
rect 16037 14433 16071 14467
rect 17325 14433 17359 14467
rect 17601 14433 17635 14467
rect 18613 14433 18647 14467
rect 2513 14365 2547 14399
rect 3157 14365 3191 14399
rect 3433 14365 3467 14399
rect 8769 14365 8803 14399
rect 16589 14365 16623 14399
rect 17785 14365 17819 14399
rect 21465 14365 21499 14399
rect 23305 14365 23339 14399
rect 23673 14365 23707 14399
rect 25145 14365 25179 14399
rect 12173 14297 12207 14331
rect 13737 14297 13771 14331
rect 16865 14297 16899 14331
rect 1547 14229 1581 14263
rect 4353 14229 4387 14263
rect 7205 14229 7239 14263
rect 19533 14229 19567 14263
rect 23121 14229 23155 14263
rect 1593 14025 1627 14059
rect 2513 14025 2547 14059
rect 3893 14025 3927 14059
rect 5917 14025 5951 14059
rect 6653 14025 6687 14059
rect 7757 14025 7791 14059
rect 8125 14025 8159 14059
rect 8769 14025 8803 14059
rect 14013 14025 14047 14059
rect 15301 14025 15335 14059
rect 16129 14025 16163 14059
rect 18705 14025 18739 14059
rect 20545 14025 20579 14059
rect 22109 14025 22143 14059
rect 22477 14025 22511 14059
rect 23213 14025 23247 14059
rect 25053 14025 25087 14059
rect 2053 13957 2087 13991
rect 5273 13957 5307 13991
rect 6193 13957 6227 13991
rect 9137 13957 9171 13991
rect 11529 13957 11563 13991
rect 12725 13957 12759 13991
rect 14381 13957 14415 13991
rect 15761 13957 15795 13991
rect 17877 13957 17911 13991
rect 19901 13957 19935 13991
rect 20177 13957 20211 13991
rect 24685 13957 24719 13991
rect 25421 13957 25455 13991
rect 2881 13889 2915 13923
rect 6837 13889 6871 13923
rect 9321 13889 9355 13923
rect 13093 13889 13127 13923
rect 14749 13889 14783 13923
rect 16497 13889 16531 13923
rect 20821 13889 20855 13923
rect 21189 13889 21223 13923
rect 25743 13889 25777 13923
rect 1409 13821 1443 13855
rect 3525 13821 3559 13855
rect 4353 13821 4387 13855
rect 8493 13821 8527 13855
rect 10517 13821 10551 13855
rect 11345 13821 11379 13855
rect 12633 13821 12667 13855
rect 12909 13821 12943 13855
rect 13645 13821 13679 13855
rect 14289 13821 14323 13855
rect 14565 13821 14599 13855
rect 18337 13821 18371 13855
rect 18981 13821 19015 13855
rect 22293 13821 22327 13855
rect 22753 13821 22787 13855
rect 23857 13821 23891 13855
rect 25640 13821 25674 13855
rect 26065 13821 26099 13855
rect 2973 13753 3007 13787
rect 4261 13753 4295 13787
rect 4715 13753 4749 13787
rect 7158 13753 7192 13787
rect 9683 13753 9717 13787
rect 16589 13753 16623 13787
rect 17141 13753 17175 13787
rect 19302 13753 19336 13787
rect 20913 13753 20947 13787
rect 24133 13753 24167 13787
rect 24225 13753 24259 13787
rect 10241 13685 10275 13719
rect 11161 13685 11195 13719
rect 12081 13685 12115 13719
rect 17509 13685 17543 13719
rect 21741 13685 21775 13719
rect 1593 13481 1627 13515
rect 3065 13481 3099 13515
rect 3525 13481 3559 13515
rect 4721 13481 4755 13515
rect 6745 13481 6779 13515
rect 8769 13481 8803 13515
rect 9321 13481 9355 13515
rect 12081 13481 12115 13515
rect 13093 13481 13127 13515
rect 14289 13481 14323 13515
rect 15025 13481 15059 13515
rect 15853 13481 15887 13515
rect 19165 13481 19199 13515
rect 21097 13481 21131 13515
rect 23029 13481 23063 13515
rect 2237 13413 2271 13447
rect 4445 13413 4479 13447
rect 7113 13413 7147 13447
rect 7665 13413 7699 13447
rect 8493 13413 8527 13447
rect 9873 13413 9907 13447
rect 12633 13413 12667 13447
rect 16773 13413 16807 13447
rect 17325 13413 17359 13447
rect 18337 13413 18371 13447
rect 18889 13413 18923 13447
rect 21649 13413 21683 13447
rect 23305 13413 23339 13447
rect 23857 13413 23891 13447
rect 24777 13413 24811 13447
rect 24869 13413 24903 13447
rect 25421 13413 25455 13447
rect 4905 13345 4939 13379
rect 5181 13345 5215 13379
rect 2145 13277 2179 13311
rect 7021 13277 7055 13311
rect 2697 13209 2731 13243
rect 8585 13345 8619 13379
rect 11161 13345 11195 13379
rect 11621 13345 11655 13379
rect 11897 13345 11931 13379
rect 13185 13345 13219 13379
rect 13461 13345 13495 13379
rect 15301 13345 15335 13379
rect 19860 13345 19894 13379
rect 9781 13277 9815 13311
rect 10057 13277 10091 13311
rect 13921 13277 13955 13311
rect 16681 13277 16715 13311
rect 18245 13277 18279 13311
rect 19947 13277 19981 13311
rect 21557 13277 21591 13311
rect 22201 13277 22235 13311
rect 23213 13277 23247 13311
rect 11713 13209 11747 13243
rect 13277 13209 13311 13243
rect 8493 13141 8527 13175
rect 11529 13141 11563 13175
rect 14657 13141 14691 13175
rect 15485 13141 15519 13175
rect 16497 13141 16531 13175
rect 17969 13141 18003 13175
rect 24133 13141 24167 13175
rect 1961 12937 1995 12971
rect 7849 12937 7883 12971
rect 8585 12937 8619 12971
rect 10241 12937 10275 12971
rect 15209 12937 15243 12971
rect 16589 12937 16623 12971
rect 17233 12937 17267 12971
rect 19809 12937 19843 12971
rect 23213 12937 23247 12971
rect 23857 12937 23891 12971
rect 24501 12937 24535 12971
rect 25513 12937 25547 12971
rect 2697 12869 2731 12903
rect 4445 12869 4479 12903
rect 5549 12869 5583 12903
rect 12909 12869 12943 12903
rect 15577 12869 15611 12903
rect 2145 12801 2179 12835
rect 3065 12801 3099 12835
rect 4905 12801 4939 12835
rect 9597 12801 9631 12835
rect 18613 12801 18647 12835
rect 20637 12801 20671 12835
rect 21373 12801 21407 12835
rect 21557 12801 21591 12835
rect 22201 12801 22235 12835
rect 5365 12733 5399 12767
rect 6653 12733 6687 12767
rect 7113 12733 7147 12767
rect 7389 12733 7423 12767
rect 10701 12733 10735 12767
rect 11437 12733 11471 12767
rect 12817 12733 12851 12767
rect 14105 12733 14139 12767
rect 14657 12733 14691 12767
rect 14841 12733 14875 12767
rect 15669 12733 15703 12767
rect 16865 12733 16899 12767
rect 20269 12733 20303 12767
rect 20913 12733 20947 12767
rect 24593 12733 24627 12767
rect 25145 12733 25179 12767
rect 2237 12665 2271 12699
rect 3893 12665 3927 12699
rect 3985 12665 4019 12699
rect 9321 12665 9355 12699
rect 9413 12665 9447 12699
rect 11529 12665 11563 12699
rect 13553 12665 13587 12699
rect 15990 12665 16024 12699
rect 17877 12665 17911 12699
rect 18705 12665 18739 12699
rect 19257 12665 19291 12699
rect 20085 12665 20119 12699
rect 21649 12665 21683 12699
rect 22569 12665 22603 12699
rect 3709 12597 3743 12631
rect 5273 12597 5307 12631
rect 6193 12597 6227 12631
rect 7113 12597 7147 12631
rect 8217 12597 8251 12631
rect 9137 12597 9171 12631
rect 11805 12597 11839 12631
rect 12173 12597 12207 12631
rect 13829 12597 13863 12631
rect 18245 12597 18279 12631
rect 24777 12597 24811 12631
rect 2145 12393 2179 12427
rect 3893 12393 3927 12427
rect 5733 12393 5767 12427
rect 9045 12393 9079 12427
rect 18797 12393 18831 12427
rect 20269 12393 20303 12427
rect 20729 12393 20763 12427
rect 2237 12325 2271 12359
rect 2513 12325 2547 12359
rect 3065 12325 3099 12359
rect 4261 12325 4295 12359
rect 7481 12325 7515 12359
rect 8033 12325 8067 12359
rect 9873 12325 9907 12359
rect 12817 12325 12851 12359
rect 15485 12325 15519 12359
rect 15990 12325 16024 12359
rect 18239 12325 18273 12359
rect 19073 12325 19107 12359
rect 21373 12325 21407 12359
rect 22937 12325 22971 12359
rect 23489 12325 23523 12359
rect 24501 12325 24535 12359
rect 5917 12257 5951 12291
rect 6193 12257 6227 12291
rect 12081 12257 12115 12291
rect 12633 12257 12667 12291
rect 13921 12257 13955 12291
rect 14197 12257 14231 12291
rect 15669 12257 15703 12291
rect 16589 12257 16623 12291
rect 19876 12257 19910 12291
rect 2421 12189 2455 12223
rect 4169 12189 4203 12223
rect 4445 12189 4479 12223
rect 7389 12189 7423 12223
rect 9781 12189 9815 12223
rect 10057 12189 10091 12223
rect 14381 12189 14415 12223
rect 17877 12189 17911 12223
rect 21281 12189 21315 12223
rect 21557 12189 21591 12223
rect 22845 12189 22879 12223
rect 24409 12189 24443 12223
rect 24685 12189 24719 12223
rect 2237 12121 2271 12155
rect 11713 12121 11747 12155
rect 19947 12121 19981 12155
rect 23857 12121 23891 12155
rect 1685 12053 1719 12087
rect 5365 12053 5399 12087
rect 6837 12053 6871 12087
rect 9321 12053 9355 12087
rect 13093 12053 13127 12087
rect 13553 12053 13587 12087
rect 14749 12053 14783 12087
rect 16865 12053 16899 12087
rect 22293 12053 22327 12087
rect 4445 11849 4479 11883
rect 6561 11849 6595 11883
rect 8861 11849 8895 11883
rect 10241 11849 10275 11883
rect 10793 11849 10827 11883
rect 11529 11849 11563 11883
rect 12725 11849 12759 11883
rect 16865 11849 16899 11883
rect 19809 11849 19843 11883
rect 23029 11849 23063 11883
rect 24685 11849 24719 11883
rect 25421 11849 25455 11883
rect 4077 11781 4111 11815
rect 5457 11781 5491 11815
rect 9137 11781 9171 11815
rect 11253 11781 11287 11815
rect 17417 11781 17451 11815
rect 17877 11781 17911 11815
rect 25053 11781 25087 11815
rect 2421 11713 2455 11747
rect 3065 11713 3099 11747
rect 3709 11713 3743 11747
rect 4537 11713 4571 11747
rect 8033 11713 8067 11747
rect 9321 11713 9355 11747
rect 12817 11713 12851 11747
rect 21649 11713 21683 11747
rect 23765 11713 23799 11747
rect 24041 11713 24075 11747
rect 5825 11645 5859 11679
rect 6837 11645 6871 11679
rect 11345 11645 11379 11679
rect 11805 11645 11839 11679
rect 12596 11645 12630 11679
rect 14657 11645 14691 11679
rect 14933 11645 14967 11679
rect 15117 11645 15151 11679
rect 15945 11645 15979 11679
rect 18337 11645 18371 11679
rect 18521 11645 18555 11679
rect 19901 11645 19935 11679
rect 21833 11645 21867 11679
rect 22753 11645 22787 11679
rect 23397 11645 23431 11679
rect 25237 11645 25271 11679
rect 25789 11645 25823 11679
rect 2237 11577 2271 11611
rect 2513 11577 2547 11611
rect 4858 11577 4892 11611
rect 7159 11577 7193 11611
rect 9683 11577 9717 11611
rect 12449 11577 12483 11611
rect 13921 11577 13955 11611
rect 14289 11577 14323 11611
rect 15485 11577 15519 11611
rect 15853 11577 15887 11611
rect 16307 11577 16341 11611
rect 20222 11577 20256 11611
rect 22154 11577 22188 11611
rect 23857 11577 23891 11611
rect 1869 11509 1903 11543
rect 6101 11509 6135 11543
rect 7757 11509 7791 11543
rect 8493 11509 8527 11543
rect 12173 11509 12207 11543
rect 13093 11509 13127 11543
rect 13553 11509 13587 11543
rect 18337 11509 18371 11543
rect 19349 11509 19383 11543
rect 20821 11509 20855 11543
rect 21281 11509 21315 11543
rect 1869 11305 1903 11339
rect 2973 11305 3007 11339
rect 3893 11305 3927 11339
rect 5457 11305 5491 11339
rect 7389 11305 7423 11339
rect 10609 11305 10643 11339
rect 14381 11305 14415 11339
rect 14749 11305 14783 11339
rect 16681 11305 16715 11339
rect 17509 11305 17543 11339
rect 18153 11305 18187 11339
rect 18429 11305 18463 11339
rect 20729 11305 20763 11339
rect 21925 11305 21959 11339
rect 22615 11305 22649 11339
rect 25237 11305 25271 11339
rect 2145 11237 2179 11271
rect 4858 11237 4892 11271
rect 6790 11237 6824 11271
rect 8769 11237 8803 11271
rect 10051 11237 10085 11271
rect 11805 11237 11839 11271
rect 15577 11237 15611 11271
rect 15853 11237 15887 11271
rect 19349 11237 19383 11271
rect 21097 11237 21131 11271
rect 22937 11237 22971 11271
rect 23673 11237 23707 11271
rect 8217 11169 8251 11203
rect 8401 11169 8435 11203
rect 11621 11169 11655 11203
rect 12035 11169 12069 11203
rect 13185 11169 13219 11203
rect 13369 11169 13403 11203
rect 13645 11169 13679 11203
rect 17233 11169 17267 11203
rect 17417 11169 17451 11203
rect 18613 11169 18647 11203
rect 19073 11169 19107 11203
rect 22512 11169 22546 11203
rect 25053 11169 25087 11203
rect 2053 11101 2087 11135
rect 2513 11101 2547 11135
rect 4537 11101 4571 11135
rect 6469 11101 6503 11135
rect 7665 11101 7699 11135
rect 9689 11101 9723 11135
rect 12173 11101 12207 11135
rect 12541 11101 12575 11135
rect 13461 11101 13495 11135
rect 13921 11101 13955 11135
rect 15761 11101 15795 11135
rect 16221 11101 16255 11135
rect 21005 11101 21039 11135
rect 21281 11101 21315 11135
rect 23581 11101 23615 11135
rect 23857 11101 23891 11135
rect 3341 11033 3375 11067
rect 4445 11033 4479 11067
rect 9505 11033 9539 11067
rect 10977 11033 11011 11067
rect 17049 11033 17083 11067
rect 8033 10965 8067 10999
rect 9137 10965 9171 10999
rect 11943 10965 11977 10999
rect 12909 10965 12943 10999
rect 19901 10965 19935 10999
rect 4629 10761 4663 10795
rect 6561 10761 6595 10795
rect 7113 10761 7147 10795
rect 8401 10761 8435 10795
rect 8769 10761 8803 10795
rect 12725 10761 12759 10795
rect 13829 10761 13863 10795
rect 15669 10761 15703 10795
rect 17785 10761 17819 10795
rect 19533 10761 19567 10795
rect 21833 10761 21867 10795
rect 22385 10761 22419 10795
rect 22707 10761 22741 10795
rect 23489 10761 23523 10795
rect 25421 10761 25455 10795
rect 1961 10693 1995 10727
rect 2697 10693 2731 10727
rect 8033 10693 8067 10727
rect 21465 10693 21499 10727
rect 3157 10625 3191 10659
rect 4169 10625 4203 10659
rect 5733 10625 5767 10659
rect 9597 10625 9631 10659
rect 12265 10625 12299 10659
rect 12814 10625 12848 10659
rect 15853 10625 15887 10659
rect 16221 10625 16255 10659
rect 19257 10625 19291 10659
rect 20545 10625 20579 10659
rect 21189 10625 21223 10659
rect 24041 10625 24075 10659
rect 5181 10557 5215 10591
rect 5641 10557 5675 10591
rect 9229 10557 9263 10591
rect 9413 10557 9447 10591
rect 10425 10557 10459 10591
rect 10793 10557 10827 10591
rect 11069 10557 11103 10591
rect 12596 10557 12630 10591
rect 13185 10557 13219 10591
rect 14289 10557 14323 10591
rect 14749 10557 14783 10591
rect 18521 10557 18555 10591
rect 18981 10557 19015 10591
rect 22636 10557 22670 10591
rect 25237 10557 25271 10591
rect 25789 10557 25823 10591
rect 2145 10489 2179 10523
rect 2237 10489 2271 10523
rect 3709 10489 3743 10523
rect 3801 10489 3835 10523
rect 7481 10489 7515 10523
rect 7573 10489 7607 10523
rect 12449 10489 12483 10523
rect 14933 10489 14967 10523
rect 15945 10489 15979 10523
rect 20269 10489 20303 10523
rect 20637 10489 20671 10523
rect 23765 10489 23799 10523
rect 23857 10489 23891 10523
rect 3433 10421 3467 10455
rect 4997 10421 5031 10455
rect 10057 10421 10091 10455
rect 10609 10421 10643 10455
rect 11897 10421 11931 10455
rect 13553 10421 13587 10455
rect 15209 10421 15243 10455
rect 16865 10421 16899 10455
rect 17233 10421 17267 10455
rect 18429 10421 18463 10455
rect 23029 10421 23063 10455
rect 24685 10421 24719 10455
rect 25053 10421 25087 10455
rect 3709 10217 3743 10251
rect 5273 10217 5307 10251
rect 7481 10217 7515 10251
rect 9045 10217 9079 10251
rect 9505 10217 9539 10251
rect 11897 10217 11931 10251
rect 13553 10217 13587 10251
rect 13921 10217 13955 10251
rect 14289 10217 14323 10251
rect 16313 10217 16347 10251
rect 16589 10217 16623 10251
rect 18613 10217 18647 10251
rect 19993 10217 20027 10251
rect 22477 10217 22511 10251
rect 24777 10217 24811 10251
rect 25145 10217 25179 10251
rect 2145 10149 2179 10183
rect 4261 10149 4295 10183
rect 6745 10149 6779 10183
rect 7757 10149 7791 10183
rect 9873 10149 9907 10183
rect 14933 10149 14967 10183
rect 15755 10149 15789 10183
rect 17693 10149 17727 10183
rect 19435 10149 19469 10183
rect 21097 10149 21131 10183
rect 23719 10149 23753 10183
rect 6285 10081 6319 10115
rect 6561 10081 6595 10115
rect 12081 10081 12115 10115
rect 12449 10081 12483 10115
rect 13093 10081 13127 10115
rect 14105 10081 14139 10115
rect 14565 10081 14599 10115
rect 23616 10081 23650 10115
rect 24593 10081 24627 10115
rect 2053 10013 2087 10047
rect 2513 10013 2547 10047
rect 4169 10013 4203 10047
rect 4629 10013 4663 10047
rect 7665 10013 7699 10047
rect 9781 10013 9815 10047
rect 10057 10013 10091 10047
rect 13277 10013 13311 10047
rect 15393 10013 15427 10047
rect 17601 10013 17635 10047
rect 19073 10013 19107 10047
rect 21005 10013 21039 10047
rect 21281 10013 21315 10047
rect 8217 9945 8251 9979
rect 8677 9945 8711 9979
rect 18153 9945 18187 9979
rect 24041 9945 24075 9979
rect 1685 9877 1719 9911
rect 2973 9877 3007 9911
rect 10793 9877 10827 9911
rect 11529 9877 11563 9911
rect 16957 9877 16991 9911
rect 20453 9877 20487 9911
rect 21925 9877 21959 9911
rect 2421 9673 2455 9707
rect 6101 9673 6135 9707
rect 6469 9673 6503 9707
rect 10149 9673 10183 9707
rect 10609 9673 10643 9707
rect 24409 9673 24443 9707
rect 5549 9605 5583 9639
rect 11897 9605 11931 9639
rect 12173 9605 12207 9639
rect 12541 9605 12575 9639
rect 13461 9605 13495 9639
rect 13829 9605 13863 9639
rect 16681 9605 16715 9639
rect 18245 9605 18279 9639
rect 22293 9605 22327 9639
rect 24777 9605 24811 9639
rect 25237 9605 25271 9639
rect 3709 9537 3743 9571
rect 4905 9537 4939 9571
rect 8309 9537 8343 9571
rect 9229 9537 9263 9571
rect 9689 9537 9723 9571
rect 12909 9537 12943 9571
rect 21373 9537 21407 9571
rect 21649 9537 21683 9571
rect 1685 9469 1719 9503
rect 1961 9469 1995 9503
rect 10793 9469 10827 9503
rect 11253 9469 11287 9503
rect 12449 9469 12483 9503
rect 12725 9469 12759 9503
rect 14013 9469 14047 9503
rect 15117 9469 15151 9503
rect 16313 9469 16347 9503
rect 16900 9469 16934 9503
rect 17325 9469 17359 9503
rect 19533 9469 19567 9503
rect 20453 9469 20487 9503
rect 21097 9469 21131 9503
rect 24593 9469 24627 9503
rect 2145 9401 2179 9435
rect 3065 9401 3099 9435
rect 3157 9401 3191 9435
rect 4629 9401 4663 9435
rect 4721 9401 4755 9435
rect 7389 9401 7423 9435
rect 7665 9401 7699 9435
rect 7757 9401 7791 9435
rect 9045 9401 9079 9435
rect 9321 9401 9355 9435
rect 14565 9401 14599 9435
rect 15025 9401 15059 9435
rect 15479 9401 15513 9435
rect 17003 9401 17037 9435
rect 19165 9401 19199 9435
rect 19895 9401 19929 9435
rect 21465 9401 21499 9435
rect 2881 9333 2915 9367
rect 4077 9333 4111 9367
rect 7021 9333 7055 9367
rect 8585 9333 8619 9367
rect 10793 9333 10827 9367
rect 14197 9333 14231 9367
rect 16037 9333 16071 9367
rect 17785 9333 17819 9367
rect 18521 9333 18555 9367
rect 20821 9333 20855 9367
rect 22661 9333 22695 9367
rect 23857 9333 23891 9367
rect 1547 9129 1581 9163
rect 1869 9129 1903 9163
rect 3893 9129 3927 9163
rect 7757 9129 7791 9163
rect 8723 9129 8757 9163
rect 10609 9129 10643 9163
rect 13277 9129 13311 9163
rect 16221 9129 16255 9163
rect 18429 9129 18463 9163
rect 19073 9129 19107 9163
rect 19349 9129 19383 9163
rect 21925 9129 21959 9163
rect 2605 9061 2639 9095
rect 3157 9061 3191 9095
rect 5175 9061 5209 9095
rect 7199 9061 7233 9095
rect 10051 9061 10085 9095
rect 14381 9061 14415 9095
rect 15663 9061 15697 9095
rect 17871 9061 17905 9095
rect 21005 9061 21039 9095
rect 21097 9061 21131 9095
rect 22661 9061 22695 9095
rect 1476 8993 1510 9027
rect 4629 8993 4663 9027
rect 5733 8993 5767 9027
rect 8620 8993 8654 9027
rect 12541 8993 12575 9027
rect 13645 8993 13679 9027
rect 14197 8993 14231 9027
rect 15301 8993 15335 9027
rect 19349 8993 19383 9027
rect 19717 8993 19751 9027
rect 24593 8993 24627 9027
rect 2237 8925 2271 8959
rect 2513 8925 2547 8959
rect 4813 8925 4847 8959
rect 6837 8925 6871 8959
rect 9689 8925 9723 8959
rect 17509 8925 17543 8959
rect 21281 8925 21315 8959
rect 22569 8925 22603 8959
rect 22845 8925 22879 8959
rect 12173 8857 12207 8891
rect 20269 8857 20303 8891
rect 3433 8789 3467 8823
rect 8033 8789 8067 8823
rect 9137 8789 9171 8823
rect 9505 8789 9539 8823
rect 11805 8789 11839 8823
rect 13001 8789 13035 8823
rect 14749 8789 14783 8823
rect 24777 8789 24811 8823
rect 1593 8585 1627 8619
rect 7757 8585 7791 8619
rect 8585 8585 8619 8619
rect 10241 8585 10275 8619
rect 10701 8585 10735 8619
rect 11345 8585 11379 8619
rect 13461 8585 13495 8619
rect 15393 8585 15427 8619
rect 16589 8585 16623 8619
rect 17601 8585 17635 8619
rect 19625 8585 19659 8619
rect 20223 8585 20257 8619
rect 21005 8585 21039 8619
rect 22109 8585 22143 8619
rect 22569 8585 22603 8619
rect 25513 8585 25547 8619
rect 10931 8517 10965 8551
rect 11897 8517 11931 8551
rect 16221 8517 16255 8551
rect 19257 8517 19291 8551
rect 20545 8517 20579 8551
rect 2789 8449 2823 8483
rect 3433 8449 3467 8483
rect 12449 8449 12483 8483
rect 13921 8449 13955 8483
rect 14749 8449 14783 8483
rect 15669 8449 15703 8483
rect 18981 8449 19015 8483
rect 21465 8449 21499 8483
rect 22937 8449 22971 8483
rect 24731 8449 24765 8483
rect 1409 8381 1443 8415
rect 3985 8381 4019 8415
rect 4813 8381 4847 8415
rect 5733 8381 5767 8415
rect 6837 8381 6871 8415
rect 9045 8381 9079 8415
rect 9965 8381 9999 8415
rect 10860 8381 10894 8415
rect 12265 8381 12299 8415
rect 13093 8381 13127 8415
rect 14289 8381 14323 8415
rect 14565 8381 14599 8415
rect 18245 8381 18279 8415
rect 18797 8381 18831 8415
rect 20152 8381 20186 8415
rect 24644 8381 24678 8415
rect 2881 8313 2915 8347
rect 4353 8313 4387 8347
rect 4721 8313 4755 8347
rect 5175 8313 5209 8347
rect 6285 8313 6319 8347
rect 6653 8313 6687 8347
rect 7199 8313 7233 8347
rect 9407 8313 9441 8347
rect 15761 8313 15795 8347
rect 21189 8313 21223 8347
rect 21281 8313 21315 8347
rect 25053 8313 25087 8347
rect 2237 8245 2271 8279
rect 2605 8245 2639 8279
rect 8033 8245 8067 8279
rect 17141 8245 17175 8279
rect 1547 8041 1581 8075
rect 1961 8041 1995 8075
rect 2329 8041 2363 8075
rect 3801 8041 3835 8075
rect 5641 8041 5675 8075
rect 7987 8041 8021 8075
rect 9137 8041 9171 8075
rect 9781 8041 9815 8075
rect 12173 8041 12207 8075
rect 14565 8041 14599 8075
rect 15531 8041 15565 8075
rect 15945 8041 15979 8075
rect 16313 8041 16347 8075
rect 17141 8041 17175 8075
rect 18245 8041 18279 8075
rect 18705 8041 18739 8075
rect 19947 8041 19981 8075
rect 20729 8041 20763 8075
rect 24731 8041 24765 8075
rect 2605 7973 2639 8007
rect 3157 7973 3191 8007
rect 4813 7973 4847 8007
rect 7021 7973 7055 8007
rect 7297 7973 7331 8007
rect 13645 7973 13679 8007
rect 14197 7973 14231 8007
rect 21281 7973 21315 8007
rect 21833 7973 21867 8007
rect 23627 7973 23661 8007
rect 1444 7905 1478 7939
rect 6285 7905 6319 7939
rect 6745 7905 6779 7939
rect 7916 7905 7950 7939
rect 9965 7905 9999 7939
rect 10241 7905 10275 7939
rect 11897 7905 11931 7939
rect 12081 7905 12115 7939
rect 13829 7905 13863 7939
rect 15428 7905 15462 7939
rect 17049 7905 17083 7939
rect 17601 7905 17635 7939
rect 19876 7905 19910 7939
rect 23540 7905 23574 7939
rect 24660 7905 24694 7939
rect 2513 7837 2547 7871
rect 4721 7837 4755 7871
rect 4997 7837 5031 7871
rect 21189 7837 21223 7871
rect 3525 7701 3559 7735
rect 2329 7497 2363 7531
rect 2789 7497 2823 7531
rect 4445 7497 4479 7531
rect 4813 7497 4847 7531
rect 6561 7497 6595 7531
rect 7941 7497 7975 7531
rect 8539 7497 8573 7531
rect 9781 7497 9815 7531
rect 10195 7497 10229 7531
rect 11253 7497 11287 7531
rect 11989 7497 12023 7531
rect 12633 7497 12667 7531
rect 13553 7497 13587 7531
rect 13921 7497 13955 7531
rect 17049 7497 17083 7531
rect 17509 7497 17543 7531
rect 19901 7497 19935 7531
rect 21189 7497 21223 7531
rect 23857 7497 23891 7531
rect 24685 7497 24719 7531
rect 1593 7429 1627 7463
rect 2053 7429 2087 7463
rect 6285 7429 6319 7463
rect 9413 7429 9447 7463
rect 11621 7429 11655 7463
rect 14289 7429 14323 7463
rect 3893 7361 3927 7395
rect 7573 7361 7607 7395
rect 1409 7293 1443 7327
rect 4905 7293 4939 7327
rect 5457 7293 5491 7327
rect 6837 7293 6871 7327
rect 7389 7293 7423 7327
rect 8436 7293 8470 7327
rect 8861 7293 8895 7327
rect 10092 7293 10126 7327
rect 10517 7293 10551 7327
rect 11069 7293 11103 7327
rect 12449 7293 12483 7327
rect 12909 7293 12943 7327
rect 13737 7293 13771 7327
rect 14565 7293 14599 7327
rect 15393 7293 15427 7327
rect 3249 7225 3283 7259
rect 3433 7225 3467 7259
rect 3525 7225 3559 7259
rect 4997 7157 5031 7191
rect 21557 7157 21591 7191
rect 2973 6953 3007 6987
rect 4215 6953 4249 6987
rect 4629 6953 4663 6987
rect 4997 6953 5031 6987
rect 6377 6953 6411 6987
rect 6837 6953 6871 6987
rect 11897 6953 11931 6987
rect 1409 6817 1443 6851
rect 3525 6817 3559 6851
rect 4144 6817 4178 6851
rect 5124 6817 5158 6851
rect 5227 6817 5261 6851
rect 7364 6817 7398 6851
rect 8344 6817 8378 6851
rect 10308 6817 10342 6851
rect 11380 6817 11414 6851
rect 11483 6817 11517 6851
rect 1593 6681 1627 6715
rect 7435 6681 7469 6715
rect 8447 6681 8481 6715
rect 10379 6681 10413 6715
rect 2421 6613 2455 6647
rect 1593 6409 1627 6443
rect 2053 6409 2087 6443
rect 3663 6409 3697 6443
rect 4169 6409 4203 6443
rect 5089 6409 5123 6443
rect 7389 6409 7423 6443
rect 8309 6409 8343 6443
rect 10333 6409 10367 6443
rect 11345 6409 11379 6443
rect 2329 6273 2363 6307
rect 2513 6273 2547 6307
rect 1409 6205 1443 6239
rect 3560 6205 3594 6239
rect 3341 6069 3375 6103
rect 1547 5865 1581 5899
rect 2559 5865 2593 5899
rect 1444 5729 1478 5763
rect 2488 5729 2522 5763
rect 1869 5321 1903 5355
rect 2605 5321 2639 5355
rect 1547 5253 1581 5287
rect 1476 5117 1510 5151
rect 2237 5117 2271 5151
rect 1547 4777 1581 4811
rect 1444 4641 1478 4675
rect 1593 4233 1627 4267
rect 1547 3145 1581 3179
rect 24731 3145 24765 3179
rect 1476 2941 1510 2975
rect 1869 2941 1903 2975
rect 24660 2941 24694 2975
rect 25145 2805 25179 2839
rect 1547 2601 1581 2635
rect 2559 2601 2593 2635
rect 24179 2601 24213 2635
rect 25191 2601 25225 2635
rect 1444 2465 1478 2499
rect 1869 2465 1903 2499
rect 2488 2465 2522 2499
rect 2881 2465 2915 2499
rect 24108 2465 24142 2499
rect 25120 2465 25154 2499
rect 24593 2261 24627 2295
rect 25605 2261 25639 2295
<< metal1 >>
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 16390 24392 16396 24404
rect 16351 24364 16396 24392
rect 16390 24352 16396 24364
rect 16448 24352 16454 24404
rect 658 24216 664 24268
rect 716 24256 722 24268
rect 1432 24259 1490 24265
rect 1432 24256 1444 24259
rect 716 24228 1444 24256
rect 716 24216 722 24228
rect 1432 24225 1444 24228
rect 1478 24256 1490 24259
rect 2222 24256 2228 24268
rect 1478 24228 2228 24256
rect 1478 24225 1490 24228
rect 1432 24219 1490 24225
rect 2222 24216 2228 24228
rect 2280 24216 2286 24268
rect 16114 24216 16120 24268
rect 16172 24256 16178 24268
rect 17402 24265 17408 24268
rect 16209 24259 16267 24265
rect 16209 24256 16221 24259
rect 16172 24228 16221 24256
rect 16172 24216 16178 24228
rect 16209 24225 16221 24228
rect 16255 24225 16267 24259
rect 16209 24219 16267 24225
rect 17380 24259 17408 24265
rect 17380 24225 17392 24259
rect 17380 24219 17408 24225
rect 17402 24216 17408 24219
rect 17460 24216 17466 24268
rect 1535 24055 1593 24061
rect 1535 24021 1547 24055
rect 1581 24052 1593 24055
rect 2682 24052 2688 24064
rect 1581 24024 2688 24052
rect 1581 24021 1593 24024
rect 1535 24015 1593 24021
rect 2682 24012 2688 24024
rect 2740 24012 2746 24064
rect 16482 24012 16488 24064
rect 16540 24052 16546 24064
rect 17494 24061 17500 24064
rect 16761 24055 16819 24061
rect 16761 24052 16773 24055
rect 16540 24024 16773 24052
rect 16540 24012 16546 24024
rect 16761 24021 16773 24024
rect 16807 24021 16819 24055
rect 16761 24015 16819 24021
rect 17451 24055 17500 24061
rect 17451 24021 17463 24055
rect 17497 24021 17500 24055
rect 17451 24015 17500 24021
rect 17494 24012 17500 24015
rect 17552 24012 17558 24064
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 2222 23848 2228 23860
rect 2183 23820 2228 23848
rect 2222 23808 2228 23820
rect 2280 23808 2286 23860
rect 12986 23848 12992 23860
rect 12947 23820 12992 23848
rect 12986 23808 12992 23820
rect 13044 23808 13050 23860
rect 15473 23851 15531 23857
rect 15473 23817 15485 23851
rect 15519 23848 15531 23851
rect 16022 23848 16028 23860
rect 15519 23820 16028 23848
rect 15519 23817 15531 23820
rect 15473 23811 15531 23817
rect 16022 23808 16028 23820
rect 16080 23808 16086 23860
rect 17402 23848 17408 23860
rect 17363 23820 17408 23848
rect 17402 23808 17408 23820
rect 17460 23808 17466 23860
rect 18233 23851 18291 23857
rect 18233 23817 18245 23851
rect 18279 23848 18291 23851
rect 18782 23848 18788 23860
rect 18279 23820 18788 23848
rect 18279 23817 18291 23820
rect 18233 23811 18291 23817
rect 18782 23808 18788 23820
rect 18840 23808 18846 23860
rect 23842 23848 23848 23860
rect 23803 23820 23848 23848
rect 23842 23808 23848 23820
rect 23900 23808 23906 23860
rect 25314 23848 25320 23860
rect 25275 23820 25320 23848
rect 25314 23808 25320 23820
rect 25372 23808 25378 23860
rect 1394 23604 1400 23656
rect 1452 23653 1458 23656
rect 1452 23647 1490 23653
rect 1478 23644 1490 23647
rect 1857 23647 1915 23653
rect 1857 23644 1869 23647
rect 1478 23616 1869 23644
rect 1478 23613 1490 23616
rect 1452 23607 1490 23613
rect 1857 23613 1869 23616
rect 1903 23613 1915 23647
rect 1857 23607 1915 23613
rect 1452 23604 1458 23607
rect 12434 23604 12440 23656
rect 12492 23644 12498 23656
rect 12805 23647 12863 23653
rect 12805 23644 12817 23647
rect 12492 23616 12817 23644
rect 12492 23604 12498 23616
rect 12805 23613 12817 23616
rect 12851 23644 12863 23647
rect 13357 23647 13415 23653
rect 13357 23644 13369 23647
rect 12851 23616 13369 23644
rect 12851 23613 12863 23616
rect 12805 23607 12863 23613
rect 13357 23613 13369 23616
rect 13403 23613 13415 23647
rect 13357 23607 13415 23613
rect 15197 23647 15255 23653
rect 15197 23613 15209 23647
rect 15243 23644 15255 23647
rect 15286 23644 15292 23656
rect 15243 23616 15292 23644
rect 15243 23613 15255 23616
rect 15197 23607 15255 23613
rect 15286 23604 15292 23616
rect 15344 23604 15350 23656
rect 18049 23647 18107 23653
rect 18049 23613 18061 23647
rect 18095 23644 18107 23647
rect 18095 23616 18736 23644
rect 18095 23613 18107 23616
rect 18049 23607 18107 23613
rect 1535 23579 1593 23585
rect 1535 23545 1547 23579
rect 1581 23576 1593 23579
rect 2682 23576 2688 23588
rect 1581 23548 2688 23576
rect 1581 23545 1593 23548
rect 1535 23539 1593 23545
rect 2682 23536 2688 23548
rect 2740 23536 2746 23588
rect 15933 23579 15991 23585
rect 15933 23545 15945 23579
rect 15979 23576 15991 23579
rect 16482 23576 16488 23588
rect 15979 23548 16344 23576
rect 16443 23548 16488 23576
rect 15979 23545 15991 23548
rect 15933 23539 15991 23545
rect 16114 23468 16120 23520
rect 16172 23508 16178 23520
rect 16209 23511 16267 23517
rect 16209 23508 16221 23511
rect 16172 23480 16221 23508
rect 16172 23468 16178 23480
rect 16209 23477 16221 23480
rect 16255 23477 16267 23511
rect 16316 23508 16344 23548
rect 16482 23536 16488 23548
rect 16540 23536 16546 23588
rect 16577 23579 16635 23585
rect 16577 23545 16589 23579
rect 16623 23576 16635 23579
rect 16942 23576 16948 23588
rect 16623 23548 16948 23576
rect 16623 23545 16635 23548
rect 16577 23539 16635 23545
rect 16592 23508 16620 23539
rect 16942 23536 16948 23548
rect 17000 23536 17006 23588
rect 17126 23576 17132 23588
rect 17087 23548 17132 23576
rect 17126 23536 17132 23548
rect 17184 23536 17190 23588
rect 18708 23520 18736 23616
rect 22462 23604 22468 23656
rect 22520 23653 22526 23656
rect 22520 23647 22558 23653
rect 22546 23613 22558 23647
rect 22520 23607 22558 23613
rect 22603 23647 22661 23653
rect 22603 23613 22615 23647
rect 22649 23644 22661 23647
rect 23661 23647 23719 23653
rect 23661 23644 23673 23647
rect 22649 23616 23673 23644
rect 22649 23613 22661 23616
rect 22603 23607 22661 23613
rect 23661 23613 23673 23616
rect 23707 23644 23719 23647
rect 24213 23647 24271 23653
rect 24213 23644 24225 23647
rect 23707 23616 24225 23644
rect 23707 23613 23719 23616
rect 23661 23607 23719 23613
rect 24213 23613 24225 23616
rect 24259 23613 24271 23647
rect 24213 23607 24271 23613
rect 24832 23647 24890 23653
rect 24832 23613 24844 23647
rect 24878 23644 24890 23647
rect 25314 23644 25320 23656
rect 24878 23616 25320 23644
rect 24878 23613 24890 23616
rect 24832 23607 24890 23613
rect 22520 23604 22526 23607
rect 25314 23604 25320 23616
rect 25372 23604 25378 23656
rect 22480 23576 22508 23604
rect 22925 23579 22983 23585
rect 22925 23576 22937 23579
rect 22480 23548 22937 23576
rect 22925 23545 22937 23548
rect 22971 23545 22983 23579
rect 22925 23539 22983 23545
rect 18690 23508 18696 23520
rect 16316 23480 16620 23508
rect 18651 23480 18696 23508
rect 16209 23471 16267 23477
rect 18690 23468 18696 23480
rect 18748 23468 18754 23520
rect 24854 23468 24860 23520
rect 24912 23517 24918 23520
rect 24912 23511 24961 23517
rect 24912 23477 24915 23511
rect 24949 23477 24961 23511
rect 24912 23471 24961 23477
rect 24912 23468 24918 23471
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 15286 23264 15292 23316
rect 15344 23304 15350 23316
rect 15611 23307 15669 23313
rect 15611 23304 15623 23307
rect 15344 23276 15623 23304
rect 15344 23264 15350 23276
rect 15611 23273 15623 23276
rect 15657 23273 15669 23307
rect 15611 23267 15669 23273
rect 21085 23307 21143 23313
rect 21085 23273 21097 23307
rect 21131 23304 21143 23307
rect 21634 23304 21640 23316
rect 21131 23276 21640 23304
rect 21131 23273 21143 23276
rect 21085 23267 21143 23273
rect 21634 23264 21640 23276
rect 21692 23264 21698 23316
rect 22646 23304 22652 23316
rect 22607 23276 22652 23304
rect 22646 23264 22652 23276
rect 22704 23264 22710 23316
rect 16574 23196 16580 23248
rect 16632 23236 16638 23248
rect 16669 23239 16727 23245
rect 16669 23236 16681 23239
rect 16632 23208 16681 23236
rect 16632 23196 16638 23208
rect 16669 23205 16681 23208
rect 16715 23205 16727 23239
rect 16669 23199 16727 23205
rect 15470 23128 15476 23180
rect 15528 23177 15534 23180
rect 15528 23171 15566 23177
rect 15554 23137 15566 23171
rect 15528 23131 15566 23137
rect 18116 23171 18174 23177
rect 18116 23137 18128 23171
rect 18162 23168 18174 23171
rect 18598 23168 18604 23180
rect 18162 23140 18604 23168
rect 18162 23137 18174 23140
rect 18116 23131 18174 23137
rect 15528 23128 15534 23131
rect 18598 23128 18604 23140
rect 18656 23128 18662 23180
rect 20898 23168 20904 23180
rect 20859 23140 20904 23168
rect 20898 23128 20904 23140
rect 20956 23128 20962 23180
rect 22462 23168 22468 23180
rect 22423 23140 22468 23168
rect 22462 23128 22468 23140
rect 22520 23128 22526 23180
rect 16577 23103 16635 23109
rect 16577 23069 16589 23103
rect 16623 23069 16635 23103
rect 16577 23063 16635 23069
rect 16592 23032 16620 23063
rect 16666 23060 16672 23112
rect 16724 23100 16730 23112
rect 16853 23103 16911 23109
rect 16853 23100 16865 23103
rect 16724 23072 16865 23100
rect 16724 23060 16730 23072
rect 16853 23069 16865 23072
rect 16899 23069 16911 23103
rect 16853 23063 16911 23069
rect 17310 23032 17316 23044
rect 16592 23004 17316 23032
rect 17310 22992 17316 23004
rect 17368 23032 17374 23044
rect 18187 23035 18245 23041
rect 18187 23032 18199 23035
rect 17368 23004 18199 23032
rect 17368 22992 17374 23004
rect 18187 23001 18199 23004
rect 18233 23001 18245 23035
rect 18187 22995 18245 23001
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 17494 22760 17500 22772
rect 17455 22732 17500 22760
rect 17494 22720 17500 22732
rect 17552 22720 17558 22772
rect 18598 22760 18604 22772
rect 18559 22732 18604 22760
rect 18598 22720 18604 22732
rect 18656 22720 18662 22772
rect 17512 22692 17540 22720
rect 16500 22664 17540 22692
rect 16500 22633 16528 22664
rect 16485 22627 16543 22633
rect 16485 22593 16497 22627
rect 16531 22593 16543 22627
rect 16758 22624 16764 22636
rect 16719 22596 16764 22624
rect 16485 22587 16543 22593
rect 16758 22584 16764 22596
rect 16816 22584 16822 22636
rect 14737 22559 14795 22565
rect 14737 22525 14749 22559
rect 14783 22556 14795 22559
rect 15473 22559 15531 22565
rect 15473 22556 15485 22559
rect 14783 22528 15485 22556
rect 14783 22525 14795 22528
rect 14737 22519 14795 22525
rect 15473 22525 15485 22528
rect 15519 22556 15531 22559
rect 15654 22556 15660 22568
rect 15519 22528 15660 22556
rect 15519 22525 15531 22528
rect 15473 22519 15531 22525
rect 15654 22516 15660 22528
rect 15712 22516 15718 22568
rect 15562 22488 15568 22500
rect 15523 22460 15568 22488
rect 15562 22448 15568 22460
rect 15620 22448 15626 22500
rect 16574 22488 16580 22500
rect 16487 22460 16580 22488
rect 16574 22448 16580 22460
rect 16632 22448 16638 22500
rect 20898 22488 20904 22500
rect 20859 22460 20904 22488
rect 20898 22448 20904 22460
rect 20956 22448 20962 22500
rect 15746 22380 15752 22432
rect 15804 22420 15810 22432
rect 15841 22423 15899 22429
rect 15841 22420 15853 22423
rect 15804 22392 15853 22420
rect 15804 22380 15810 22392
rect 15841 22389 15853 22392
rect 15887 22420 15899 22423
rect 16209 22423 16267 22429
rect 16209 22420 16221 22423
rect 15887 22392 16221 22420
rect 15887 22389 15899 22392
rect 15841 22383 15899 22389
rect 16209 22389 16221 22392
rect 16255 22420 16267 22423
rect 16592 22420 16620 22448
rect 16255 22392 16620 22420
rect 16255 22389 16267 22392
rect 16209 22383 16267 22389
rect 17862 22380 17868 22432
rect 17920 22420 17926 22432
rect 18049 22423 18107 22429
rect 18049 22420 18061 22423
rect 17920 22392 18061 22420
rect 17920 22380 17926 22392
rect 18049 22389 18061 22392
rect 18095 22389 18107 22423
rect 22462 22420 22468 22432
rect 22423 22392 22468 22420
rect 18049 22383 18107 22389
rect 22462 22380 22468 22392
rect 22520 22380 22526 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 15470 22216 15476 22228
rect 15383 22188 15476 22216
rect 15470 22176 15476 22188
rect 15528 22216 15534 22228
rect 17310 22216 17316 22228
rect 15528 22188 16528 22216
rect 17271 22188 17316 22216
rect 15528 22176 15534 22188
rect 16500 22160 16528 22188
rect 17310 22176 17316 22188
rect 17368 22176 17374 22228
rect 13262 22108 13268 22160
rect 13320 22148 13326 22160
rect 13357 22151 13415 22157
rect 13357 22148 13369 22151
rect 13320 22120 13369 22148
rect 13320 22108 13326 22120
rect 13357 22117 13369 22120
rect 13403 22117 13415 22151
rect 13357 22111 13415 22117
rect 15562 22108 15568 22160
rect 15620 22148 15626 22160
rect 15930 22148 15936 22160
rect 15620 22120 15936 22148
rect 15620 22108 15626 22120
rect 15930 22108 15936 22120
rect 15988 22148 15994 22160
rect 16393 22151 16451 22157
rect 16393 22148 16405 22151
rect 15988 22120 16405 22148
rect 15988 22108 15994 22120
rect 16393 22117 16405 22120
rect 16439 22117 16451 22151
rect 16393 22111 16451 22117
rect 16482 22108 16488 22160
rect 16540 22108 16546 22160
rect 17954 22148 17960 22160
rect 17915 22120 17960 22148
rect 17954 22108 17960 22120
rect 18012 22108 18018 22160
rect 19337 22083 19395 22089
rect 19337 22049 19349 22083
rect 19383 22080 19395 22083
rect 19426 22080 19432 22092
rect 19383 22052 19432 22080
rect 19383 22049 19395 22052
rect 19337 22043 19395 22049
rect 19426 22040 19432 22052
rect 19484 22040 19490 22092
rect 21818 22080 21824 22092
rect 21779 22052 21824 22080
rect 21818 22040 21824 22052
rect 21876 22040 21882 22092
rect 13262 22012 13268 22024
rect 13223 21984 13268 22012
rect 13262 21972 13268 21984
rect 13320 21972 13326 22024
rect 13906 22012 13912 22024
rect 13867 21984 13912 22012
rect 13906 21972 13912 21984
rect 13964 21972 13970 22024
rect 16298 22012 16304 22024
rect 16259 21984 16304 22012
rect 16298 21972 16304 21984
rect 16356 21972 16362 22024
rect 16482 21972 16488 22024
rect 16540 22012 16546 22024
rect 16577 22015 16635 22021
rect 16577 22012 16589 22015
rect 16540 21984 16589 22012
rect 16540 21972 16546 21984
rect 16577 21981 16589 21984
rect 16623 21981 16635 22015
rect 17862 22012 17868 22024
rect 17823 21984 17868 22012
rect 16577 21975 16635 21981
rect 17862 21972 17868 21984
rect 17920 21972 17926 22024
rect 18138 22012 18144 22024
rect 18099 21984 18144 22012
rect 18138 21972 18144 21984
rect 18196 21972 18202 22024
rect 16117 21947 16175 21953
rect 16117 21913 16129 21947
rect 16163 21944 16175 21947
rect 16206 21944 16212 21956
rect 16163 21916 16212 21944
rect 16163 21913 16175 21916
rect 16117 21907 16175 21913
rect 16206 21904 16212 21916
rect 16264 21944 16270 21956
rect 16758 21944 16764 21956
rect 16264 21916 16764 21944
rect 16264 21904 16270 21916
rect 16758 21904 16764 21916
rect 16816 21904 16822 21956
rect 19521 21947 19579 21953
rect 19521 21913 19533 21947
rect 19567 21944 19579 21947
rect 20162 21944 20168 21956
rect 19567 21916 20168 21944
rect 19567 21913 19579 21916
rect 19521 21907 19579 21913
rect 20162 21904 20168 21916
rect 20220 21904 20226 21956
rect 22002 21944 22008 21956
rect 21963 21916 22008 21944
rect 22002 21904 22008 21916
rect 22060 21904 22066 21956
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 13081 21675 13139 21681
rect 13081 21641 13093 21675
rect 13127 21672 13139 21675
rect 13170 21672 13176 21684
rect 13127 21644 13176 21672
rect 13127 21641 13139 21644
rect 13081 21635 13139 21641
rect 13170 21632 13176 21644
rect 13228 21632 13234 21684
rect 15930 21672 15936 21684
rect 15891 21644 15936 21672
rect 15930 21632 15936 21644
rect 15988 21632 15994 21684
rect 17497 21675 17555 21681
rect 17497 21641 17509 21675
rect 17543 21672 17555 21675
rect 17862 21672 17868 21684
rect 17543 21644 17868 21672
rect 17543 21641 17555 21644
rect 17497 21635 17555 21641
rect 17862 21632 17868 21644
rect 17920 21632 17926 21684
rect 19426 21672 19432 21684
rect 19387 21644 19432 21672
rect 19426 21632 19432 21644
rect 19484 21632 19490 21684
rect 15243 21607 15301 21613
rect 15243 21573 15255 21607
rect 15289 21604 15301 21607
rect 16390 21604 16396 21616
rect 15289 21576 16396 21604
rect 15289 21573 15301 21576
rect 15243 21567 15301 21573
rect 16390 21564 16396 21576
rect 16448 21564 16454 21616
rect 13906 21536 13912 21548
rect 13867 21508 13912 21536
rect 13906 21496 13912 21508
rect 13964 21536 13970 21548
rect 14921 21539 14979 21545
rect 14921 21536 14933 21539
rect 13964 21508 14933 21536
rect 13964 21496 13970 21508
rect 14921 21505 14933 21508
rect 14967 21505 14979 21539
rect 16206 21536 16212 21548
rect 16167 21508 16212 21536
rect 14921 21499 14979 21505
rect 1486 21477 1492 21480
rect 1464 21471 1492 21477
rect 1464 21437 1476 21471
rect 1544 21468 1550 21480
rect 1857 21471 1915 21477
rect 1857 21468 1869 21471
rect 1544 21440 1869 21468
rect 1464 21431 1492 21437
rect 1486 21428 1492 21431
rect 1544 21428 1550 21440
rect 1857 21437 1869 21440
rect 1903 21437 1915 21471
rect 14936 21468 14964 21499
rect 16206 21496 16212 21508
rect 16264 21496 16270 21548
rect 16482 21536 16488 21548
rect 16443 21508 16488 21536
rect 16482 21496 16488 21508
rect 16540 21496 16546 21548
rect 15140 21471 15198 21477
rect 15140 21468 15152 21471
rect 14936 21440 15152 21468
rect 1857 21431 1915 21437
rect 15140 21437 15152 21440
rect 15186 21437 15198 21471
rect 15140 21431 15198 21437
rect 18046 21428 18052 21480
rect 18104 21468 18110 21480
rect 18141 21471 18199 21477
rect 18141 21468 18153 21471
rect 18104 21440 18153 21468
rect 18104 21428 18110 21440
rect 18141 21437 18153 21440
rect 18187 21468 18199 21471
rect 19061 21471 19119 21477
rect 19061 21468 19073 21471
rect 18187 21440 19073 21468
rect 18187 21437 18199 21440
rect 18141 21431 18199 21437
rect 19061 21437 19073 21440
rect 19107 21437 19119 21471
rect 21818 21468 21824 21480
rect 21779 21440 21824 21468
rect 19061 21431 19119 21437
rect 21818 21428 21824 21440
rect 21876 21428 21882 21480
rect 13630 21400 13636 21412
rect 13591 21372 13636 21400
rect 13630 21360 13636 21372
rect 13688 21360 13694 21412
rect 13722 21360 13728 21412
rect 13780 21400 13786 21412
rect 15654 21400 15660 21412
rect 13780 21372 13825 21400
rect 15567 21372 15660 21400
rect 13780 21360 13786 21372
rect 15654 21360 15660 21372
rect 15712 21400 15718 21412
rect 16206 21400 16212 21412
rect 15712 21372 16212 21400
rect 15712 21360 15718 21372
rect 16206 21360 16212 21372
rect 16264 21400 16270 21412
rect 16301 21403 16359 21409
rect 16301 21400 16313 21403
rect 16264 21372 16313 21400
rect 16264 21360 16270 21372
rect 16301 21369 16313 21372
rect 16347 21369 16359 21403
rect 16301 21363 16359 21369
rect 1535 21335 1593 21341
rect 1535 21301 1547 21335
rect 1581 21332 1593 21335
rect 1762 21332 1768 21344
rect 1581 21304 1768 21332
rect 1581 21301 1593 21304
rect 1535 21295 1593 21301
rect 1762 21292 1768 21304
rect 1820 21292 1826 21344
rect 13449 21335 13507 21341
rect 13449 21301 13461 21335
rect 13495 21332 13507 21335
rect 13740 21332 13768 21360
rect 13495 21304 13768 21332
rect 13495 21301 13507 21304
rect 13449 21295 13507 21301
rect 16390 21292 16396 21344
rect 16448 21332 16454 21344
rect 17773 21335 17831 21341
rect 17773 21332 17785 21335
rect 16448 21304 17785 21332
rect 16448 21292 16454 21304
rect 17773 21301 17785 21304
rect 17819 21332 17831 21335
rect 17954 21332 17960 21344
rect 17819 21304 17960 21332
rect 17819 21301 17831 21304
rect 17773 21295 17831 21301
rect 17954 21292 17960 21304
rect 18012 21332 18018 21344
rect 18325 21335 18383 21341
rect 18325 21332 18337 21335
rect 18012 21304 18337 21332
rect 18012 21292 18018 21304
rect 18325 21301 18337 21304
rect 18371 21301 18383 21335
rect 18325 21295 18383 21301
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 13262 21128 13268 21140
rect 12912 21100 13268 21128
rect 10778 21060 10784 21072
rect 10739 21032 10784 21060
rect 10778 21020 10784 21032
rect 10836 21020 10842 21072
rect 11882 21020 11888 21072
rect 11940 21060 11946 21072
rect 12912 21069 12940 21100
rect 13262 21088 13268 21100
rect 13320 21088 13326 21140
rect 13630 21128 13636 21140
rect 13591 21100 13636 21128
rect 13630 21088 13636 21100
rect 13688 21128 13694 21140
rect 19426 21137 19432 21140
rect 13725 21131 13783 21137
rect 13725 21128 13737 21131
rect 13688 21100 13737 21128
rect 13688 21088 13694 21100
rect 13725 21097 13737 21100
rect 13771 21097 13783 21131
rect 13725 21091 13783 21097
rect 19383 21131 19432 21137
rect 19383 21097 19395 21131
rect 19429 21097 19432 21131
rect 19383 21091 19432 21097
rect 19426 21088 19432 21091
rect 19484 21088 19490 21140
rect 12345 21063 12403 21069
rect 12345 21060 12357 21063
rect 11940 21032 12357 21060
rect 11940 21020 11946 21032
rect 12345 21029 12357 21032
rect 12391 21029 12403 21063
rect 12345 21023 12403 21029
rect 12897 21063 12955 21069
rect 12897 21029 12909 21063
rect 12943 21029 12955 21063
rect 12897 21023 12955 21029
rect 16301 21063 16359 21069
rect 16301 21029 16313 21063
rect 16347 21060 16359 21063
rect 16390 21060 16396 21072
rect 16347 21032 16396 21060
rect 16347 21029 16359 21032
rect 16301 21023 16359 21029
rect 10686 20924 10692 20936
rect 10647 20896 10692 20924
rect 10686 20884 10692 20896
rect 10744 20884 10750 20936
rect 12253 20927 12311 20933
rect 12253 20893 12265 20927
rect 12299 20924 12311 20927
rect 12526 20924 12532 20936
rect 12299 20896 12532 20924
rect 12299 20893 12311 20896
rect 12253 20887 12311 20893
rect 12526 20884 12532 20896
rect 12584 20884 12590 20936
rect 11241 20859 11299 20865
rect 11241 20825 11253 20859
rect 11287 20856 11299 20859
rect 12912 20856 12940 21023
rect 16390 21020 16396 21032
rect 16448 21020 16454 21072
rect 17770 20992 17776 21004
rect 17731 20964 17776 20992
rect 17770 20952 17776 20964
rect 17828 20952 17834 21004
rect 19334 21001 19340 21004
rect 19312 20995 19340 21001
rect 19312 20961 19324 20995
rect 19312 20955 19340 20961
rect 19334 20952 19340 20955
rect 19392 20952 19398 21004
rect 16209 20927 16267 20933
rect 16209 20893 16221 20927
rect 16255 20924 16267 20927
rect 16574 20924 16580 20936
rect 16255 20896 16580 20924
rect 16255 20893 16267 20896
rect 16209 20887 16267 20893
rect 16574 20884 16580 20896
rect 16632 20884 16638 20936
rect 11287 20828 12940 20856
rect 16025 20859 16083 20865
rect 11287 20825 11299 20828
rect 11241 20819 11299 20825
rect 16025 20825 16037 20859
rect 16071 20856 16083 20859
rect 16298 20856 16304 20868
rect 16071 20828 16304 20856
rect 16071 20825 16083 20828
rect 16025 20819 16083 20825
rect 16298 20816 16304 20828
rect 16356 20816 16362 20868
rect 16758 20856 16764 20868
rect 16719 20828 16764 20856
rect 16758 20816 16764 20828
rect 16816 20816 16822 20868
rect 14826 20748 14832 20800
rect 14884 20788 14890 20800
rect 14921 20791 14979 20797
rect 14921 20788 14933 20791
rect 14884 20760 14933 20788
rect 14884 20748 14890 20760
rect 14921 20757 14933 20760
rect 14967 20757 14979 20791
rect 17954 20788 17960 20800
rect 17915 20760 17960 20788
rect 14921 20751 14979 20757
rect 17954 20748 17960 20760
rect 18012 20748 18018 20800
rect 18782 20788 18788 20800
rect 18743 20760 18788 20788
rect 18782 20748 18788 20760
rect 18840 20748 18846 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 11882 20584 11888 20596
rect 11843 20556 11888 20584
rect 11882 20544 11888 20556
rect 11940 20544 11946 20596
rect 13170 20544 13176 20596
rect 13228 20584 13234 20596
rect 13633 20587 13691 20593
rect 13633 20584 13645 20587
rect 13228 20556 13645 20584
rect 13228 20544 13234 20556
rect 13633 20553 13645 20556
rect 13679 20553 13691 20587
rect 13633 20547 13691 20553
rect 15746 20544 15752 20596
rect 15804 20584 15810 20596
rect 15841 20587 15899 20593
rect 15841 20584 15853 20587
rect 15804 20556 15853 20584
rect 15804 20544 15810 20556
rect 15841 20553 15853 20556
rect 15887 20553 15899 20587
rect 15841 20547 15899 20553
rect 16209 20587 16267 20593
rect 16209 20553 16221 20587
rect 16255 20584 16267 20587
rect 16390 20584 16396 20596
rect 16255 20556 16396 20584
rect 16255 20553 16267 20556
rect 16209 20547 16267 20553
rect 16390 20544 16396 20556
rect 16448 20544 16454 20596
rect 16574 20584 16580 20596
rect 16535 20556 16580 20584
rect 16574 20544 16580 20556
rect 16632 20584 16638 20596
rect 16807 20587 16865 20593
rect 16807 20584 16819 20587
rect 16632 20556 16819 20584
rect 16632 20544 16638 20556
rect 16807 20553 16819 20556
rect 16853 20553 16865 20587
rect 16807 20547 16865 20553
rect 17865 20587 17923 20593
rect 17865 20553 17877 20587
rect 17911 20584 17923 20587
rect 17954 20584 17960 20596
rect 17911 20556 17960 20584
rect 17911 20553 17923 20556
rect 17865 20547 17923 20553
rect 17954 20544 17960 20556
rect 18012 20544 18018 20596
rect 18782 20516 18788 20528
rect 18340 20488 18788 20516
rect 10689 20451 10747 20457
rect 10689 20417 10701 20451
rect 10735 20448 10747 20451
rect 10778 20448 10784 20460
rect 10735 20420 10784 20448
rect 10735 20417 10747 20420
rect 10689 20411 10747 20417
rect 10778 20408 10784 20420
rect 10836 20408 10842 20460
rect 18340 20457 18368 20488
rect 18782 20476 18788 20488
rect 18840 20476 18846 20528
rect 18325 20451 18383 20457
rect 18325 20417 18337 20451
rect 18371 20417 18383 20451
rect 18598 20448 18604 20460
rect 18559 20420 18604 20448
rect 18325 20411 18383 20417
rect 18598 20408 18604 20420
rect 18656 20448 18662 20460
rect 19245 20451 19303 20457
rect 19245 20448 19257 20451
rect 18656 20420 19257 20448
rect 18656 20408 18662 20420
rect 19245 20417 19257 20420
rect 19291 20448 19303 20451
rect 19334 20448 19340 20460
rect 19291 20420 19340 20448
rect 19291 20417 19303 20420
rect 19245 20411 19303 20417
rect 19334 20408 19340 20420
rect 19392 20408 19398 20460
rect 20806 20448 20812 20460
rect 20767 20420 20812 20448
rect 20806 20408 20812 20420
rect 20864 20408 20870 20460
rect 10321 20383 10379 20389
rect 10321 20349 10333 20383
rect 10367 20380 10379 20383
rect 11425 20383 11483 20389
rect 11425 20380 11437 20383
rect 10367 20352 11437 20380
rect 10367 20349 10379 20352
rect 10321 20343 10379 20349
rect 11425 20349 11437 20352
rect 11471 20380 11483 20383
rect 11882 20380 11888 20392
rect 11471 20352 11888 20380
rect 11471 20349 11483 20352
rect 11425 20343 11483 20349
rect 11882 20340 11888 20352
rect 11940 20340 11946 20392
rect 12710 20380 12716 20392
rect 12671 20352 12716 20380
rect 12710 20340 12716 20352
rect 12768 20340 12774 20392
rect 14826 20340 14832 20392
rect 14884 20380 14890 20392
rect 14921 20383 14979 20389
rect 14921 20380 14933 20383
rect 14884 20352 14933 20380
rect 14884 20340 14890 20352
rect 14921 20349 14933 20352
rect 14967 20349 14979 20383
rect 14921 20343 14979 20349
rect 16666 20340 16672 20392
rect 16724 20389 16730 20392
rect 16724 20383 16762 20389
rect 16750 20380 16762 20383
rect 17129 20383 17187 20389
rect 17129 20380 17141 20383
rect 16750 20352 17141 20380
rect 16750 20349 16762 20352
rect 16724 20343 16762 20349
rect 17129 20349 17141 20352
rect 17175 20349 17187 20383
rect 17129 20343 17187 20349
rect 16724 20340 16730 20343
rect 19794 20340 19800 20392
rect 19852 20389 19858 20392
rect 19852 20383 19890 20389
rect 19878 20380 19890 20383
rect 20254 20380 20260 20392
rect 19878 20352 20260 20380
rect 19878 20349 19890 20352
rect 19852 20343 19890 20349
rect 19852 20340 19858 20343
rect 20254 20340 20260 20352
rect 20312 20340 20318 20392
rect 11974 20272 11980 20324
rect 12032 20312 12038 20324
rect 12161 20315 12219 20321
rect 12161 20312 12173 20315
rect 12032 20284 12173 20312
rect 12032 20272 12038 20284
rect 12161 20281 12173 20284
rect 12207 20312 12219 20315
rect 13034 20315 13092 20321
rect 13034 20312 13046 20315
rect 12207 20284 13046 20312
rect 12207 20281 12219 20284
rect 12161 20275 12219 20281
rect 13034 20281 13046 20284
rect 13080 20312 13092 20315
rect 14737 20315 14795 20321
rect 14737 20312 14749 20315
rect 13080 20284 14749 20312
rect 13080 20281 13092 20284
rect 13034 20275 13092 20281
rect 14737 20281 14749 20284
rect 14783 20312 14795 20315
rect 15242 20315 15300 20321
rect 15242 20312 15254 20315
rect 14783 20284 15254 20312
rect 14783 20281 14795 20284
rect 14737 20275 14795 20281
rect 15242 20281 15254 20284
rect 15288 20312 15300 20315
rect 15562 20312 15568 20324
rect 15288 20284 15568 20312
rect 15288 20281 15300 20284
rect 15242 20275 15300 20281
rect 15562 20272 15568 20284
rect 15620 20272 15626 20324
rect 18417 20315 18475 20321
rect 18417 20281 18429 20315
rect 18463 20281 18475 20315
rect 18417 20275 18475 20281
rect 13446 20204 13452 20256
rect 13504 20244 13510 20256
rect 13909 20247 13967 20253
rect 13909 20244 13921 20247
rect 13504 20216 13921 20244
rect 13504 20204 13510 20216
rect 13909 20213 13921 20216
rect 13955 20213 13967 20247
rect 13909 20207 13967 20213
rect 17954 20204 17960 20256
rect 18012 20244 18018 20256
rect 18432 20244 18460 20275
rect 18012 20216 18460 20244
rect 18012 20204 18018 20216
rect 19426 20204 19432 20256
rect 19484 20244 19490 20256
rect 19935 20247 19993 20253
rect 19935 20244 19947 20247
rect 19484 20216 19947 20244
rect 19484 20204 19490 20216
rect 19935 20213 19947 20216
rect 19981 20213 19993 20247
rect 19935 20207 19993 20213
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 10686 20040 10692 20052
rect 10647 20012 10692 20040
rect 10686 20000 10692 20012
rect 10744 20000 10750 20052
rect 11882 20000 11888 20052
rect 11940 20040 11946 20052
rect 12805 20043 12863 20049
rect 12805 20040 12817 20043
rect 11940 20012 12817 20040
rect 11940 20000 11946 20012
rect 12805 20009 12817 20012
rect 12851 20009 12863 20043
rect 12805 20003 12863 20009
rect 13170 20000 13176 20052
rect 13228 20040 13234 20052
rect 13449 20043 13507 20049
rect 13449 20040 13461 20043
rect 13228 20012 13461 20040
rect 13228 20000 13234 20012
rect 13449 20009 13461 20012
rect 13495 20009 13507 20043
rect 13449 20003 13507 20009
rect 11974 19932 11980 19984
rect 12032 19972 12038 19984
rect 12206 19975 12264 19981
rect 12206 19972 12218 19975
rect 12032 19944 12218 19972
rect 12032 19932 12038 19944
rect 12206 19941 12218 19944
rect 12252 19941 12264 19975
rect 12206 19935 12264 19941
rect 9858 19864 9864 19916
rect 9916 19913 9922 19916
rect 9916 19907 9954 19913
rect 9942 19873 9954 19907
rect 9916 19867 9954 19873
rect 10873 19907 10931 19913
rect 10873 19873 10885 19907
rect 10919 19904 10931 19907
rect 10962 19904 10968 19916
rect 10919 19876 10968 19904
rect 10919 19873 10931 19876
rect 10873 19867 10931 19873
rect 9916 19864 9922 19867
rect 10962 19864 10968 19876
rect 11020 19864 11026 19916
rect 13464 19904 13492 20003
rect 13814 20000 13820 20052
rect 13872 20040 13878 20052
rect 13909 20043 13967 20049
rect 13909 20040 13921 20043
rect 13872 20012 13921 20040
rect 13872 20000 13878 20012
rect 13909 20009 13921 20012
rect 13955 20009 13967 20043
rect 16206 20040 16212 20052
rect 16167 20012 16212 20040
rect 13909 20003 13967 20009
rect 16206 20000 16212 20012
rect 16264 20000 16270 20052
rect 17770 20040 17776 20052
rect 17731 20012 17776 20040
rect 17770 20000 17776 20012
rect 17828 20000 17834 20052
rect 15562 19932 15568 19984
rect 15620 19981 15626 19984
rect 15620 19975 15668 19981
rect 15620 19941 15622 19975
rect 15656 19941 15668 19975
rect 17788 19972 17816 20000
rect 18026 19975 18084 19981
rect 18026 19972 18038 19975
rect 17788 19944 18038 19972
rect 15620 19935 15668 19941
rect 18026 19941 18038 19944
rect 18072 19941 18084 19975
rect 18598 19972 18604 19984
rect 18559 19944 18604 19972
rect 18026 19935 18084 19941
rect 15620 19932 15626 19935
rect 18598 19932 18604 19944
rect 18656 19932 18662 19984
rect 19518 19913 19524 19916
rect 13725 19907 13783 19913
rect 13725 19904 13737 19907
rect 13464 19876 13737 19904
rect 13725 19873 13737 19876
rect 13771 19873 13783 19907
rect 13725 19867 13783 19873
rect 19496 19907 19524 19913
rect 19496 19873 19508 19907
rect 19496 19867 19524 19873
rect 19518 19864 19524 19867
rect 19576 19864 19582 19916
rect 11882 19836 11888 19848
rect 11843 19808 11888 19836
rect 11882 19796 11888 19808
rect 11940 19796 11946 19848
rect 15289 19839 15347 19845
rect 15289 19805 15301 19839
rect 15335 19836 15347 19839
rect 15470 19836 15476 19848
rect 15335 19808 15476 19836
rect 15335 19805 15347 19808
rect 15289 19799 15347 19805
rect 15470 19796 15476 19808
rect 15528 19796 15534 19848
rect 17405 19839 17463 19845
rect 17405 19805 17417 19839
rect 17451 19836 17463 19839
rect 17957 19839 18015 19845
rect 17957 19836 17969 19839
rect 17451 19808 17969 19836
rect 17451 19805 17463 19808
rect 17405 19799 17463 19805
rect 17957 19805 17969 19808
rect 18003 19836 18015 19839
rect 18414 19836 18420 19848
rect 18003 19808 18420 19836
rect 18003 19805 18015 19808
rect 17957 19799 18015 19805
rect 18414 19796 18420 19808
rect 18472 19796 18478 19848
rect 11057 19771 11115 19777
rect 11057 19737 11069 19771
rect 11103 19768 11115 19771
rect 11330 19768 11336 19780
rect 11103 19740 11336 19768
rect 11103 19737 11115 19740
rect 11057 19731 11115 19737
rect 11330 19728 11336 19740
rect 11388 19728 11394 19780
rect 10042 19709 10048 19712
rect 9999 19703 10048 19709
rect 9999 19669 10011 19703
rect 10045 19669 10048 19703
rect 9999 19663 10048 19669
rect 10042 19660 10048 19663
rect 10100 19660 10106 19712
rect 11422 19700 11428 19712
rect 11383 19672 11428 19700
rect 11422 19660 11428 19672
rect 11480 19660 11486 19712
rect 12710 19660 12716 19712
rect 12768 19700 12774 19712
rect 13081 19703 13139 19709
rect 13081 19700 13093 19703
rect 12768 19672 13093 19700
rect 12768 19660 12774 19672
rect 13081 19669 13093 19672
rect 13127 19669 13139 19703
rect 14734 19700 14740 19712
rect 14695 19672 14740 19700
rect 13081 19663 13139 19669
rect 14734 19660 14740 19672
rect 14792 19660 14798 19712
rect 16577 19703 16635 19709
rect 16577 19669 16589 19703
rect 16623 19700 16635 19703
rect 16666 19700 16672 19712
rect 16623 19672 16672 19700
rect 16623 19669 16635 19672
rect 16577 19663 16635 19669
rect 16666 19660 16672 19672
rect 16724 19660 16730 19712
rect 19334 19660 19340 19712
rect 19392 19700 19398 19712
rect 19567 19703 19625 19709
rect 19567 19700 19579 19703
rect 19392 19672 19579 19700
rect 19392 19660 19398 19672
rect 19567 19669 19579 19672
rect 19613 19669 19625 19703
rect 19567 19663 19625 19669
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 9858 19496 9864 19508
rect 9819 19468 9864 19496
rect 9858 19456 9864 19468
rect 9916 19456 9922 19508
rect 11974 19496 11980 19508
rect 11935 19468 11980 19496
rect 11974 19456 11980 19468
rect 12032 19456 12038 19508
rect 15473 19499 15531 19505
rect 15473 19465 15485 19499
rect 15519 19496 15531 19499
rect 15562 19496 15568 19508
rect 15519 19468 15568 19496
rect 15519 19465 15531 19468
rect 15473 19459 15531 19465
rect 15562 19456 15568 19468
rect 15620 19496 15626 19508
rect 16022 19496 16028 19508
rect 15620 19468 16028 19496
rect 15620 19456 15626 19468
rect 16022 19456 16028 19468
rect 16080 19456 16086 19508
rect 17129 19499 17187 19505
rect 17129 19465 17141 19499
rect 17175 19496 17187 19499
rect 17497 19499 17555 19505
rect 17497 19496 17509 19499
rect 17175 19468 17509 19496
rect 17175 19465 17187 19468
rect 17129 19459 17187 19465
rect 17497 19465 17509 19468
rect 17543 19496 17555 19499
rect 17770 19496 17776 19508
rect 17543 19468 17776 19496
rect 17543 19465 17555 19468
rect 17497 19459 17555 19465
rect 17770 19456 17776 19468
rect 17828 19456 17834 19508
rect 14826 19428 14832 19440
rect 14787 19400 14832 19428
rect 14826 19388 14832 19400
rect 14884 19388 14890 19440
rect 16666 19320 16672 19372
rect 16724 19320 16730 19372
rect 18414 19360 18420 19372
rect 18375 19332 18420 19360
rect 18414 19320 18420 19332
rect 18472 19320 18478 19372
rect 1394 19252 1400 19304
rect 1452 19301 1458 19304
rect 1452 19295 1490 19301
rect 1478 19292 1490 19295
rect 1857 19295 1915 19301
rect 1857 19292 1869 19295
rect 1478 19264 1869 19292
rect 1478 19261 1490 19264
rect 1452 19255 1490 19261
rect 1857 19261 1869 19264
rect 1903 19261 1915 19295
rect 1857 19255 1915 19261
rect 7076 19295 7134 19301
rect 7076 19261 7088 19295
rect 7122 19292 7134 19295
rect 8272 19295 8330 19301
rect 7122 19264 7604 19292
rect 7122 19261 7134 19264
rect 7076 19255 7134 19261
rect 1452 19252 1458 19255
rect 1535 19159 1593 19165
rect 1535 19125 1547 19159
rect 1581 19156 1593 19159
rect 1762 19156 1768 19168
rect 1581 19128 1768 19156
rect 1581 19125 1593 19128
rect 1535 19119 1593 19125
rect 1762 19116 1768 19128
rect 1820 19116 1826 19168
rect 7147 19159 7205 19165
rect 7147 19125 7159 19159
rect 7193 19156 7205 19159
rect 7282 19156 7288 19168
rect 7193 19128 7288 19156
rect 7193 19125 7205 19128
rect 7147 19119 7205 19125
rect 7282 19116 7288 19128
rect 7340 19116 7346 19168
rect 7576 19165 7604 19264
rect 8272 19261 8284 19295
rect 8318 19292 8330 19295
rect 8386 19292 8392 19304
rect 8318 19264 8392 19292
rect 8318 19261 8330 19264
rect 8272 19255 8330 19261
rect 8386 19252 8392 19264
rect 8444 19292 8450 19304
rect 8665 19295 8723 19301
rect 8665 19292 8677 19295
rect 8444 19264 8677 19292
rect 8444 19252 8450 19264
rect 8665 19261 8677 19264
rect 8711 19292 8723 19295
rect 9030 19292 9036 19304
rect 8711 19264 9036 19292
rect 8711 19261 8723 19264
rect 8665 19255 8723 19261
rect 9030 19252 9036 19264
rect 9088 19252 9094 19304
rect 9125 19295 9183 19301
rect 9125 19261 9137 19295
rect 9171 19292 9183 19295
rect 9284 19295 9342 19301
rect 9284 19292 9296 19295
rect 9171 19264 9296 19292
rect 9171 19261 9183 19264
rect 9125 19255 9183 19261
rect 9284 19261 9296 19264
rect 9330 19292 9342 19295
rect 9582 19292 9588 19304
rect 9330 19264 9588 19292
rect 9330 19261 9342 19264
rect 9284 19255 9342 19261
rect 9582 19252 9588 19264
rect 9640 19252 9646 19304
rect 11333 19295 11391 19301
rect 11333 19261 11345 19295
rect 11379 19292 11391 19295
rect 11422 19292 11428 19304
rect 11379 19264 11428 19292
rect 11379 19261 11391 19264
rect 11333 19255 11391 19261
rect 11422 19252 11428 19264
rect 11480 19292 11486 19304
rect 12250 19292 12256 19304
rect 11480 19264 12256 19292
rect 11480 19252 11486 19264
rect 12250 19252 12256 19264
rect 12308 19252 12314 19304
rect 12434 19252 12440 19304
rect 12492 19301 12498 19304
rect 12492 19295 12530 19301
rect 12518 19292 12530 19295
rect 14182 19292 14188 19304
rect 12518 19264 12585 19292
rect 14143 19264 14188 19292
rect 12518 19261 12530 19264
rect 12492 19255 12530 19261
rect 12492 19252 12498 19255
rect 14182 19252 14188 19264
rect 14240 19252 14246 19304
rect 14461 19295 14519 19301
rect 14461 19261 14473 19295
rect 14507 19261 14519 19295
rect 14461 19255 14519 19261
rect 12452 19224 12480 19252
rect 12989 19227 13047 19233
rect 12989 19224 13001 19227
rect 12452 19196 13001 19224
rect 12989 19193 13001 19196
rect 13035 19224 13047 19227
rect 13630 19224 13636 19236
rect 13035 19196 13636 19224
rect 13035 19193 13047 19196
rect 12989 19187 13047 19193
rect 13630 19184 13636 19196
rect 13688 19184 13694 19236
rect 13906 19224 13912 19236
rect 13819 19196 13912 19224
rect 13906 19184 13912 19196
rect 13964 19224 13970 19236
rect 14476 19224 14504 19255
rect 14734 19252 14740 19304
rect 14792 19292 14798 19304
rect 14829 19295 14887 19301
rect 14829 19292 14841 19295
rect 14792 19264 14841 19292
rect 14792 19252 14798 19264
rect 14829 19261 14841 19264
rect 14875 19261 14887 19295
rect 14829 19255 14887 19261
rect 15746 19252 15752 19304
rect 15804 19292 15810 19304
rect 16209 19295 16267 19301
rect 16209 19292 16221 19295
rect 15804 19264 16221 19292
rect 15804 19252 15810 19264
rect 16209 19261 16221 19264
rect 16255 19292 16267 19295
rect 16684 19292 16712 19320
rect 19153 19295 19211 19301
rect 19153 19292 19165 19295
rect 16255 19264 16712 19292
rect 18800 19264 19165 19292
rect 16255 19261 16267 19264
rect 16209 19255 16267 19261
rect 13964 19196 14504 19224
rect 13964 19184 13970 19196
rect 16022 19184 16028 19236
rect 16080 19224 16086 19236
rect 16530 19227 16588 19233
rect 16530 19224 16542 19227
rect 16080 19196 16542 19224
rect 16080 19184 16086 19196
rect 16530 19193 16542 19196
rect 16576 19193 16588 19227
rect 18138 19224 18144 19236
rect 18099 19196 18144 19224
rect 16530 19187 16588 19193
rect 18138 19184 18144 19196
rect 18196 19184 18202 19236
rect 18233 19227 18291 19233
rect 18233 19193 18245 19227
rect 18279 19193 18291 19227
rect 18233 19187 18291 19193
rect 7561 19159 7619 19165
rect 7561 19125 7573 19159
rect 7607 19156 7619 19159
rect 7650 19156 7656 19168
rect 7607 19128 7656 19156
rect 7607 19125 7619 19128
rect 7561 19119 7619 19125
rect 7650 19116 7656 19128
rect 7708 19116 7714 19168
rect 8343 19159 8401 19165
rect 8343 19125 8355 19159
rect 8389 19156 8401 19159
rect 8938 19156 8944 19168
rect 8389 19128 8944 19156
rect 8389 19125 8401 19128
rect 8343 19119 8401 19125
rect 8938 19116 8944 19128
rect 8996 19116 9002 19168
rect 9122 19116 9128 19168
rect 9180 19156 9186 19168
rect 9355 19159 9413 19165
rect 9355 19156 9367 19159
rect 9180 19128 9367 19156
rect 9180 19116 9186 19128
rect 9355 19125 9367 19128
rect 9401 19125 9413 19159
rect 9355 19119 9413 19125
rect 10134 19116 10140 19168
rect 10192 19156 10198 19168
rect 10321 19159 10379 19165
rect 10321 19156 10333 19159
rect 10192 19128 10333 19156
rect 10192 19116 10198 19128
rect 10321 19125 10333 19128
rect 10367 19125 10379 19159
rect 10962 19156 10968 19168
rect 10923 19128 10968 19156
rect 10321 19119 10379 19125
rect 10962 19116 10968 19128
rect 11020 19116 11026 19168
rect 11422 19116 11428 19168
rect 11480 19156 11486 19168
rect 11517 19159 11575 19165
rect 11517 19156 11529 19159
rect 11480 19128 11529 19156
rect 11480 19116 11486 19128
rect 11517 19125 11529 19128
rect 11563 19125 11575 19159
rect 12526 19156 12532 19168
rect 12485 19128 12532 19156
rect 11517 19119 11575 19125
rect 12526 19116 12532 19128
rect 12584 19165 12590 19168
rect 12584 19159 12633 19165
rect 12584 19125 12587 19159
rect 12621 19156 12633 19159
rect 13446 19156 13452 19168
rect 12621 19128 13452 19156
rect 12621 19125 12633 19128
rect 12584 19119 12633 19125
rect 12584 19116 12590 19119
rect 13446 19116 13452 19128
rect 13504 19116 13510 19168
rect 13541 19159 13599 19165
rect 13541 19125 13553 19159
rect 13587 19156 13599 19159
rect 14182 19156 14188 19168
rect 13587 19128 14188 19156
rect 13587 19125 13599 19128
rect 13541 19119 13599 19125
rect 14182 19116 14188 19128
rect 14240 19116 14246 19168
rect 17865 19159 17923 19165
rect 17865 19125 17877 19159
rect 17911 19156 17923 19159
rect 18248 19156 18276 19187
rect 18322 19184 18328 19236
rect 18380 19224 18386 19236
rect 18800 19224 18828 19264
rect 19153 19261 19165 19264
rect 19199 19292 19211 19295
rect 19705 19295 19763 19301
rect 19705 19292 19717 19295
rect 19199 19264 19717 19292
rect 19199 19261 19211 19264
rect 19153 19255 19211 19261
rect 19705 19261 19717 19264
rect 19751 19261 19763 19295
rect 19705 19255 19763 19261
rect 21174 19252 21180 19304
rect 21232 19301 21238 19304
rect 21232 19295 21270 19301
rect 21258 19292 21270 19295
rect 21637 19295 21695 19301
rect 21637 19292 21649 19295
rect 21258 19264 21649 19292
rect 21258 19261 21270 19264
rect 21232 19255 21270 19261
rect 21637 19261 21649 19264
rect 21683 19261 21695 19295
rect 21637 19255 21695 19261
rect 24648 19295 24706 19301
rect 24648 19261 24660 19295
rect 24694 19292 24706 19295
rect 24762 19292 24768 19304
rect 24694 19264 24768 19292
rect 24694 19261 24706 19264
rect 24648 19255 24706 19261
rect 21232 19252 21238 19255
rect 24762 19252 24768 19264
rect 24820 19292 24826 19304
rect 25041 19295 25099 19301
rect 25041 19292 25053 19295
rect 24820 19264 25053 19292
rect 24820 19252 24826 19264
rect 25041 19261 25053 19264
rect 25087 19261 25099 19295
rect 25041 19255 25099 19261
rect 19613 19227 19671 19233
rect 19613 19224 19625 19227
rect 18380 19196 18828 19224
rect 18892 19196 19625 19224
rect 18380 19184 18386 19196
rect 18892 19156 18920 19196
rect 19613 19193 19625 19196
rect 19659 19193 19671 19227
rect 19613 19187 19671 19193
rect 19518 19156 19524 19168
rect 17911 19128 18920 19156
rect 19479 19128 19524 19156
rect 17911 19125 17923 19128
rect 17865 19119 17923 19125
rect 19518 19116 19524 19128
rect 19576 19116 19582 19168
rect 20990 19116 20996 19168
rect 21048 19156 21054 19168
rect 21315 19159 21373 19165
rect 21315 19156 21327 19159
rect 21048 19128 21327 19156
rect 21048 19116 21054 19128
rect 21315 19125 21327 19128
rect 21361 19125 21373 19159
rect 21315 19119 21373 19125
rect 23474 19116 23480 19168
rect 23532 19156 23538 19168
rect 24719 19159 24777 19165
rect 24719 19156 24731 19159
rect 23532 19128 24731 19156
rect 23532 19116 23538 19128
rect 24719 19125 24731 19128
rect 24765 19125 24777 19159
rect 24719 19119 24777 19125
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 12115 18955 12173 18961
rect 12115 18921 12127 18955
rect 12161 18952 12173 18955
rect 12342 18952 12348 18964
rect 12161 18924 12348 18952
rect 12161 18921 12173 18924
rect 12115 18915 12173 18921
rect 12342 18912 12348 18924
rect 12400 18912 12406 18964
rect 16669 18955 16727 18961
rect 16669 18921 16681 18955
rect 16715 18952 16727 18955
rect 17494 18952 17500 18964
rect 16715 18924 17500 18952
rect 16715 18921 16727 18924
rect 16669 18915 16727 18921
rect 17494 18912 17500 18924
rect 17552 18952 17558 18964
rect 17552 18924 17724 18952
rect 17552 18912 17558 18924
rect 7558 18884 7564 18896
rect 7519 18856 7564 18884
rect 7558 18844 7564 18856
rect 7616 18844 7622 18896
rect 10502 18884 10508 18896
rect 10463 18856 10508 18884
rect 10502 18844 10508 18856
rect 10560 18844 10566 18896
rect 10597 18887 10655 18893
rect 10597 18853 10609 18887
rect 10643 18884 10655 18887
rect 10778 18884 10784 18896
rect 10643 18856 10784 18884
rect 10643 18853 10655 18856
rect 10597 18847 10655 18853
rect 10778 18844 10784 18856
rect 10836 18844 10842 18896
rect 16022 18844 16028 18896
rect 16080 18893 16086 18896
rect 16080 18887 16128 18893
rect 16080 18853 16082 18887
rect 16116 18853 16128 18887
rect 16080 18847 16128 18853
rect 17405 18887 17463 18893
rect 17405 18853 17417 18887
rect 17451 18884 17463 18887
rect 17586 18884 17592 18896
rect 17451 18856 17592 18884
rect 17451 18853 17463 18856
rect 17405 18847 17463 18853
rect 16080 18844 16086 18847
rect 17586 18844 17592 18856
rect 17644 18844 17650 18896
rect 17696 18893 17724 18924
rect 18138 18912 18144 18964
rect 18196 18952 18202 18964
rect 18601 18955 18659 18961
rect 18601 18952 18613 18955
rect 18196 18924 18613 18952
rect 18196 18912 18202 18924
rect 18601 18921 18613 18924
rect 18647 18952 18659 18955
rect 19242 18952 19248 18964
rect 18647 18924 19248 18952
rect 18647 18921 18659 18924
rect 18601 18915 18659 18921
rect 19242 18912 19248 18924
rect 19300 18912 19306 18964
rect 21818 18952 21824 18964
rect 21779 18924 21824 18952
rect 21818 18912 21824 18924
rect 21876 18912 21882 18964
rect 17681 18887 17739 18893
rect 17681 18853 17693 18887
rect 17727 18884 17739 18887
rect 18046 18884 18052 18896
rect 17727 18856 18052 18884
rect 17727 18853 17739 18856
rect 17681 18847 17739 18853
rect 18046 18844 18052 18856
rect 18104 18844 18110 18896
rect 18233 18887 18291 18893
rect 18233 18853 18245 18887
rect 18279 18884 18291 18887
rect 18414 18884 18420 18896
rect 18279 18856 18420 18884
rect 18279 18853 18291 18856
rect 18233 18847 18291 18853
rect 18414 18844 18420 18856
rect 18472 18844 18478 18896
rect 23474 18844 23480 18896
rect 23532 18884 23538 18896
rect 24719 18887 24777 18893
rect 24719 18884 24731 18887
rect 23532 18856 24731 18884
rect 23532 18844 23538 18856
rect 24719 18853 24731 18856
rect 24765 18853 24777 18887
rect 24719 18847 24777 18853
rect 6362 18776 6368 18828
rect 6420 18825 6426 18828
rect 6420 18819 6458 18825
rect 6446 18785 6458 18819
rect 6420 18779 6458 18785
rect 12044 18819 12102 18825
rect 12044 18785 12056 18819
rect 12090 18816 12102 18819
rect 12158 18816 12164 18828
rect 12090 18788 12164 18816
rect 12090 18785 12102 18788
rect 12044 18779 12102 18785
rect 6420 18776 6426 18779
rect 12158 18776 12164 18788
rect 12216 18776 12222 18828
rect 13538 18816 13544 18828
rect 13499 18788 13544 18816
rect 13538 18776 13544 18788
rect 13596 18776 13602 18828
rect 13906 18816 13912 18828
rect 13867 18788 13912 18816
rect 13906 18776 13912 18788
rect 13964 18776 13970 18828
rect 14093 18819 14151 18825
rect 14093 18785 14105 18819
rect 14139 18816 14151 18819
rect 14734 18816 14740 18828
rect 14139 18788 14740 18816
rect 14139 18785 14151 18788
rect 14093 18779 14151 18785
rect 6503 18751 6561 18757
rect 6503 18717 6515 18751
rect 6549 18748 6561 18751
rect 7466 18748 7472 18760
rect 6549 18720 7472 18748
rect 6549 18717 6561 18720
rect 6503 18711 6561 18717
rect 7466 18708 7472 18720
rect 7524 18708 7530 18760
rect 7742 18748 7748 18760
rect 7703 18720 7748 18748
rect 7742 18708 7748 18720
rect 7800 18708 7806 18760
rect 10318 18708 10324 18760
rect 10376 18748 10382 18760
rect 10781 18751 10839 18757
rect 10781 18748 10793 18751
rect 10376 18720 10793 18748
rect 10376 18708 10382 18720
rect 10781 18717 10793 18720
rect 10827 18717 10839 18751
rect 10781 18711 10839 18717
rect 13814 18708 13820 18760
rect 13872 18748 13878 18760
rect 14108 18748 14136 18779
rect 14734 18776 14740 18788
rect 14792 18776 14798 18828
rect 18874 18776 18880 18828
rect 18932 18816 18938 18828
rect 19061 18819 19119 18825
rect 19061 18816 19073 18819
rect 18932 18788 19073 18816
rect 18932 18776 18938 18788
rect 19061 18785 19073 18788
rect 19107 18785 19119 18819
rect 19518 18816 19524 18828
rect 19479 18788 19524 18816
rect 19061 18779 19119 18785
rect 19518 18776 19524 18788
rect 19576 18776 19582 18828
rect 20714 18776 20720 18828
rect 20772 18816 20778 18828
rect 20936 18819 20994 18825
rect 20936 18816 20948 18819
rect 20772 18788 20948 18816
rect 20772 18776 20778 18788
rect 20936 18785 20948 18788
rect 20982 18785 20994 18819
rect 20936 18779 20994 18785
rect 24578 18776 24584 18828
rect 24636 18825 24642 18828
rect 24636 18819 24674 18825
rect 24662 18785 24674 18819
rect 24636 18779 24674 18785
rect 24636 18776 24642 18779
rect 13872 18720 14136 18748
rect 14369 18751 14427 18757
rect 13872 18708 13878 18720
rect 14369 18717 14381 18751
rect 14415 18748 14427 18751
rect 15749 18751 15807 18757
rect 15749 18748 15761 18751
rect 14415 18720 15761 18748
rect 14415 18717 14427 18720
rect 14369 18711 14427 18717
rect 15749 18717 15761 18720
rect 15795 18748 15807 18751
rect 16482 18748 16488 18760
rect 15795 18720 16488 18748
rect 15795 18717 15807 18720
rect 15749 18711 15807 18717
rect 16482 18708 16488 18720
rect 16540 18708 16546 18760
rect 19334 18708 19340 18760
rect 19392 18748 19398 18760
rect 19613 18751 19671 18757
rect 19613 18748 19625 18751
rect 19392 18720 19625 18748
rect 19392 18708 19398 18720
rect 19613 18717 19625 18720
rect 19659 18717 19671 18751
rect 19613 18711 19671 18717
rect 10321 18615 10379 18621
rect 10321 18581 10333 18615
rect 10367 18612 10379 18615
rect 10686 18612 10692 18624
rect 10367 18584 10692 18612
rect 10367 18581 10379 18584
rect 10321 18575 10379 18581
rect 10686 18572 10692 18584
rect 10744 18572 10750 18624
rect 11882 18612 11888 18624
rect 11795 18584 11888 18612
rect 11882 18572 11888 18584
rect 11940 18612 11946 18624
rect 12342 18612 12348 18624
rect 11940 18584 12348 18612
rect 11940 18572 11946 18584
rect 12342 18572 12348 18584
rect 12400 18572 12406 18624
rect 12434 18572 12440 18624
rect 12492 18612 12498 18624
rect 12894 18612 12900 18624
rect 12492 18584 12537 18612
rect 12855 18584 12900 18612
rect 12492 18572 12498 18584
rect 12894 18572 12900 18584
rect 12952 18572 12958 18624
rect 14734 18612 14740 18624
rect 14695 18584 14740 18612
rect 14734 18572 14740 18584
rect 14792 18572 14798 18624
rect 15470 18612 15476 18624
rect 15431 18584 15476 18612
rect 15470 18572 15476 18584
rect 15528 18572 15534 18624
rect 20070 18612 20076 18624
rect 20031 18584 20076 18612
rect 20070 18572 20076 18584
rect 20128 18572 20134 18624
rect 20806 18572 20812 18624
rect 20864 18612 20870 18624
rect 21039 18615 21097 18621
rect 21039 18612 21051 18615
rect 20864 18584 21051 18612
rect 20864 18572 20870 18584
rect 21039 18581 21051 18584
rect 21085 18581 21097 18615
rect 21450 18612 21456 18624
rect 21411 18584 21456 18612
rect 21039 18575 21097 18581
rect 21450 18572 21456 18584
rect 21508 18572 21514 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 5629 18411 5687 18417
rect 5629 18377 5641 18411
rect 5675 18408 5687 18411
rect 6178 18408 6184 18420
rect 5675 18380 6184 18408
rect 5675 18377 5687 18380
rect 5629 18371 5687 18377
rect 5442 18164 5448 18216
rect 5500 18204 5506 18216
rect 5828 18213 5856 18380
rect 6178 18368 6184 18380
rect 6236 18368 6242 18420
rect 6454 18408 6460 18420
rect 6415 18380 6460 18408
rect 6454 18368 6460 18380
rect 6512 18368 6518 18420
rect 7558 18368 7564 18420
rect 7616 18408 7622 18420
rect 8389 18411 8447 18417
rect 8389 18408 8401 18411
rect 7616 18380 8401 18408
rect 7616 18368 7622 18380
rect 8389 18377 8401 18380
rect 8435 18377 8447 18411
rect 8389 18371 8447 18377
rect 9769 18411 9827 18417
rect 9769 18377 9781 18411
rect 9815 18408 9827 18411
rect 9861 18411 9919 18417
rect 9861 18408 9873 18411
rect 9815 18380 9873 18408
rect 9815 18377 9827 18380
rect 9769 18371 9827 18377
rect 9861 18377 9873 18380
rect 9907 18408 9919 18411
rect 11238 18408 11244 18420
rect 9907 18380 11244 18408
rect 9907 18377 9919 18380
rect 9861 18371 9919 18377
rect 11238 18368 11244 18380
rect 11296 18368 11302 18420
rect 13906 18368 13912 18420
rect 13964 18408 13970 18420
rect 14553 18411 14611 18417
rect 14553 18408 14565 18411
rect 13964 18380 14565 18408
rect 13964 18368 13970 18380
rect 14553 18377 14565 18380
rect 14599 18377 14611 18411
rect 14553 18371 14611 18377
rect 7282 18232 7288 18284
rect 7340 18272 7346 18284
rect 7469 18275 7527 18281
rect 7469 18272 7481 18275
rect 7340 18244 7481 18272
rect 7340 18232 7346 18244
rect 7469 18241 7481 18244
rect 7515 18272 7527 18275
rect 8757 18275 8815 18281
rect 8757 18272 8769 18275
rect 7515 18244 8769 18272
rect 7515 18241 7527 18244
rect 7469 18235 7527 18241
rect 8757 18241 8769 18244
rect 8803 18241 8815 18275
rect 10318 18272 10324 18284
rect 10279 18244 10324 18272
rect 8757 18235 8815 18241
rect 10318 18232 10324 18244
rect 10376 18272 10382 18284
rect 11054 18272 11060 18284
rect 10376 18244 11060 18272
rect 10376 18232 10382 18244
rect 11054 18232 11060 18244
rect 11112 18232 11118 18284
rect 11885 18275 11943 18281
rect 11885 18241 11897 18275
rect 11931 18272 11943 18275
rect 13170 18272 13176 18284
rect 11931 18244 13176 18272
rect 11931 18241 11943 18244
rect 11885 18235 11943 18241
rect 13170 18232 13176 18244
rect 13228 18272 13234 18284
rect 14568 18272 14596 18371
rect 16022 18368 16028 18420
rect 16080 18408 16086 18420
rect 16117 18411 16175 18417
rect 16117 18408 16129 18411
rect 16080 18380 16129 18408
rect 16080 18368 16086 18380
rect 16117 18377 16129 18380
rect 16163 18377 16175 18411
rect 16482 18408 16488 18420
rect 16443 18380 16488 18408
rect 16117 18371 16175 18377
rect 16482 18368 16488 18380
rect 16540 18368 16546 18420
rect 19153 18411 19211 18417
rect 19153 18377 19165 18411
rect 19199 18408 19211 18411
rect 19518 18408 19524 18420
rect 19199 18380 19524 18408
rect 19199 18377 19211 18380
rect 19153 18371 19211 18377
rect 19518 18368 19524 18380
rect 19576 18368 19582 18420
rect 24670 18408 24676 18420
rect 24631 18380 24676 18408
rect 24670 18368 24676 18380
rect 24728 18368 24734 18420
rect 15470 18340 15476 18352
rect 15431 18312 15476 18340
rect 15470 18300 15476 18312
rect 15528 18300 15534 18352
rect 21818 18340 21824 18352
rect 21468 18312 21824 18340
rect 13228 18244 13676 18272
rect 14568 18244 15240 18272
rect 13228 18232 13234 18244
rect 5788 18207 5856 18213
rect 5788 18204 5800 18207
rect 5500 18176 5800 18204
rect 5500 18164 5506 18176
rect 5788 18173 5800 18176
rect 5834 18176 5856 18207
rect 9217 18207 9275 18213
rect 5834 18173 5846 18176
rect 5788 18167 5846 18173
rect 9217 18173 9229 18207
rect 9263 18204 9275 18207
rect 9861 18207 9919 18213
rect 9861 18204 9873 18207
rect 9263 18176 9873 18204
rect 9263 18173 9275 18176
rect 9217 18167 9275 18173
rect 9861 18173 9873 18176
rect 9907 18173 9919 18207
rect 9861 18167 9919 18173
rect 10962 18164 10968 18216
rect 11020 18204 11026 18216
rect 12158 18204 12164 18216
rect 11020 18176 12164 18204
rect 11020 18164 11026 18176
rect 12158 18164 12164 18176
rect 12216 18164 12222 18216
rect 12437 18207 12495 18213
rect 12437 18204 12449 18207
rect 12268 18176 12449 18204
rect 6822 18136 6828 18148
rect 6288 18108 6828 18136
rect 5859 18071 5917 18077
rect 5859 18037 5871 18071
rect 5905 18068 5917 18071
rect 6288 18068 6316 18108
rect 6822 18096 6828 18108
rect 6880 18096 6886 18148
rect 7006 18096 7012 18148
rect 7064 18136 7070 18148
rect 7285 18139 7343 18145
rect 7285 18136 7297 18139
rect 7064 18108 7297 18136
rect 7064 18096 7070 18108
rect 7285 18105 7297 18108
rect 7331 18136 7343 18139
rect 7561 18139 7619 18145
rect 7561 18136 7573 18139
rect 7331 18108 7573 18136
rect 7331 18105 7343 18108
rect 7285 18099 7343 18105
rect 7561 18105 7573 18108
rect 7607 18105 7619 18139
rect 7561 18099 7619 18105
rect 7834 18096 7840 18148
rect 7892 18136 7898 18148
rect 8113 18139 8171 18145
rect 8113 18136 8125 18139
rect 7892 18108 8125 18136
rect 7892 18096 7898 18108
rect 8113 18105 8125 18108
rect 8159 18105 8171 18139
rect 8113 18099 8171 18105
rect 10413 18139 10471 18145
rect 10413 18105 10425 18139
rect 10459 18136 10471 18139
rect 10686 18136 10692 18148
rect 10459 18108 10692 18136
rect 10459 18105 10471 18108
rect 10413 18099 10471 18105
rect 10686 18096 10692 18108
rect 10744 18096 10750 18148
rect 12268 18080 12296 18176
rect 12437 18173 12449 18176
rect 12483 18173 12495 18207
rect 12894 18204 12900 18216
rect 12855 18176 12900 18204
rect 12437 18167 12495 18173
rect 12894 18164 12900 18176
rect 12952 18164 12958 18216
rect 13648 18213 13676 18244
rect 13449 18207 13507 18213
rect 13449 18173 13461 18207
rect 13495 18173 13507 18207
rect 13449 18167 13507 18173
rect 13633 18207 13691 18213
rect 13633 18173 13645 18207
rect 13679 18173 13691 18207
rect 13633 18167 13691 18173
rect 13464 18136 13492 18167
rect 14182 18164 14188 18216
rect 14240 18204 14246 18216
rect 14734 18204 14740 18216
rect 14240 18176 14740 18204
rect 14240 18164 14246 18176
rect 14734 18164 14740 18176
rect 14792 18164 14798 18216
rect 15212 18213 15240 18244
rect 20714 18232 20720 18284
rect 20772 18272 20778 18284
rect 20901 18275 20959 18281
rect 20901 18272 20913 18275
rect 20772 18244 20913 18272
rect 20772 18232 20778 18244
rect 20901 18241 20913 18244
rect 20947 18272 20959 18275
rect 21266 18272 21272 18284
rect 20947 18244 21272 18272
rect 20947 18241 20959 18244
rect 20901 18235 20959 18241
rect 21266 18232 21272 18244
rect 21324 18232 21330 18284
rect 21468 18281 21496 18312
rect 21818 18300 21824 18312
rect 21876 18300 21882 18352
rect 21453 18275 21511 18281
rect 21453 18241 21465 18275
rect 21499 18241 21511 18275
rect 21453 18235 21511 18241
rect 21634 18232 21640 18284
rect 21692 18272 21698 18284
rect 21729 18275 21787 18281
rect 21729 18272 21741 18275
rect 21692 18244 21741 18272
rect 21692 18232 21698 18244
rect 21729 18241 21741 18244
rect 21775 18241 21787 18275
rect 21729 18235 21787 18241
rect 15197 18207 15255 18213
rect 15197 18173 15209 18207
rect 15243 18173 15255 18207
rect 15562 18204 15568 18216
rect 15523 18176 15568 18204
rect 15197 18167 15255 18173
rect 15562 18164 15568 18176
rect 15620 18164 15626 18216
rect 16574 18164 16580 18216
rect 16632 18204 16638 18216
rect 16669 18207 16727 18213
rect 16669 18204 16681 18207
rect 16632 18176 16681 18204
rect 16632 18164 16638 18176
rect 16669 18173 16681 18176
rect 16715 18204 16727 18207
rect 17129 18207 17187 18213
rect 17129 18204 17141 18207
rect 16715 18176 17141 18204
rect 16715 18173 16727 18176
rect 16669 18167 16727 18173
rect 17129 18173 17141 18176
rect 17175 18173 17187 18207
rect 17129 18167 17187 18173
rect 18325 18207 18383 18213
rect 18325 18173 18337 18207
rect 18371 18204 18383 18207
rect 18414 18204 18420 18216
rect 18371 18176 18420 18204
rect 18371 18173 18383 18176
rect 18325 18167 18383 18173
rect 18414 18164 18420 18176
rect 18472 18164 18478 18216
rect 18509 18207 18567 18213
rect 18509 18173 18521 18207
rect 18555 18173 18567 18207
rect 18509 18167 18567 18173
rect 18785 18207 18843 18213
rect 18785 18173 18797 18207
rect 18831 18204 18843 18207
rect 19058 18204 19064 18216
rect 18831 18176 19064 18204
rect 18831 18173 18843 18176
rect 18785 18167 18843 18173
rect 13906 18136 13912 18148
rect 13464 18108 13912 18136
rect 13906 18096 13912 18108
rect 13964 18096 13970 18148
rect 18524 18136 18552 18167
rect 19058 18164 19064 18176
rect 19116 18164 19122 18216
rect 19242 18164 19248 18216
rect 19300 18204 19306 18216
rect 19613 18207 19671 18213
rect 19613 18204 19625 18207
rect 19300 18176 19625 18204
rect 19300 18164 19306 18176
rect 19613 18173 19625 18176
rect 19659 18204 19671 18207
rect 20070 18204 20076 18216
rect 19659 18176 20076 18204
rect 19659 18173 19671 18176
rect 19613 18167 19671 18173
rect 20070 18164 20076 18176
rect 20128 18164 20134 18216
rect 18064 18108 18552 18136
rect 19934 18139 19992 18145
rect 18064 18080 18092 18108
rect 19934 18105 19946 18139
rect 19980 18105 19992 18139
rect 19934 18099 19992 18105
rect 9398 18068 9404 18080
rect 5905 18040 6316 18068
rect 9359 18040 9404 18068
rect 5905 18037 5917 18040
rect 5859 18031 5917 18037
rect 9398 18028 9404 18040
rect 9456 18028 9462 18080
rect 10137 18071 10195 18077
rect 10137 18037 10149 18071
rect 10183 18068 10195 18071
rect 10778 18068 10784 18080
rect 10183 18040 10784 18068
rect 10183 18037 10195 18040
rect 10137 18031 10195 18037
rect 10778 18028 10784 18040
rect 10836 18028 10842 18080
rect 11514 18068 11520 18080
rect 11475 18040 11520 18068
rect 11514 18028 11520 18040
rect 11572 18028 11578 18080
rect 12250 18068 12256 18080
rect 12211 18040 12256 18068
rect 12250 18028 12256 18040
rect 12308 18028 12314 18080
rect 12710 18068 12716 18080
rect 12671 18040 12716 18068
rect 12710 18028 12716 18040
rect 12768 18028 12774 18080
rect 13538 18028 13544 18080
rect 13596 18068 13602 18080
rect 14277 18071 14335 18077
rect 14277 18068 14289 18071
rect 13596 18040 14289 18068
rect 13596 18028 13602 18040
rect 14277 18037 14289 18040
rect 14323 18068 14335 18071
rect 14458 18068 14464 18080
rect 14323 18040 14464 18068
rect 14323 18037 14335 18040
rect 14277 18031 14335 18037
rect 14458 18028 14464 18040
rect 14516 18028 14522 18080
rect 16850 18068 16856 18080
rect 16811 18040 16856 18068
rect 16850 18028 16856 18040
rect 16908 18028 16914 18080
rect 17865 18071 17923 18077
rect 17865 18037 17877 18071
rect 17911 18068 17923 18071
rect 18046 18068 18052 18080
rect 17911 18040 18052 18068
rect 17911 18037 17923 18040
rect 17865 18031 17923 18037
rect 18046 18028 18052 18040
rect 18104 18028 18110 18080
rect 18966 18028 18972 18080
rect 19024 18068 19030 18080
rect 19521 18071 19579 18077
rect 19521 18068 19533 18071
rect 19024 18040 19533 18068
rect 19024 18028 19030 18040
rect 19521 18037 19533 18040
rect 19567 18068 19579 18071
rect 19949 18068 19977 18099
rect 20714 18096 20720 18148
rect 20772 18136 20778 18148
rect 21450 18136 21456 18148
rect 20772 18108 21456 18136
rect 20772 18096 20778 18108
rect 21450 18096 21456 18108
rect 21508 18136 21514 18148
rect 21545 18139 21603 18145
rect 21545 18136 21557 18139
rect 21508 18108 21557 18136
rect 21508 18096 21514 18108
rect 21545 18105 21557 18108
rect 21591 18105 21603 18139
rect 21545 18099 21603 18105
rect 19567 18040 19977 18068
rect 20533 18071 20591 18077
rect 19567 18037 19579 18040
rect 19521 18031 19579 18037
rect 20533 18037 20545 18071
rect 20579 18068 20591 18071
rect 20622 18068 20628 18080
rect 20579 18040 20628 18068
rect 20579 18037 20591 18040
rect 20533 18031 20591 18037
rect 20622 18028 20628 18040
rect 20680 18028 20686 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 5534 17824 5540 17876
rect 5592 17864 5598 17876
rect 5592 17836 5672 17864
rect 5592 17824 5598 17836
rect 5644 17805 5672 17836
rect 7466 17824 7472 17876
rect 7524 17864 7530 17876
rect 8113 17867 8171 17873
rect 8113 17864 8125 17867
rect 7524 17836 8125 17864
rect 7524 17824 7530 17836
rect 8113 17833 8125 17836
rect 8159 17833 8171 17867
rect 8113 17827 8171 17833
rect 10781 17867 10839 17873
rect 10781 17833 10793 17867
rect 10827 17864 10839 17867
rect 10870 17864 10876 17876
rect 10827 17836 10876 17864
rect 10827 17833 10839 17836
rect 10781 17827 10839 17833
rect 10870 17824 10876 17836
rect 10928 17824 10934 17876
rect 11054 17864 11060 17876
rect 11015 17836 11060 17864
rect 11054 17824 11060 17836
rect 11112 17824 11118 17876
rect 12342 17824 12348 17876
rect 12400 17864 12406 17876
rect 12437 17867 12495 17873
rect 12437 17864 12449 17867
rect 12400 17836 12449 17864
rect 12400 17824 12406 17836
rect 12437 17833 12449 17836
rect 12483 17833 12495 17867
rect 13906 17864 13912 17876
rect 13867 17836 13912 17864
rect 12437 17827 12495 17833
rect 13906 17824 13912 17836
rect 13964 17824 13970 17876
rect 16942 17864 16948 17876
rect 16903 17836 16948 17864
rect 16942 17824 16948 17836
rect 17000 17824 17006 17876
rect 17494 17864 17500 17876
rect 17455 17836 17500 17864
rect 17494 17824 17500 17836
rect 17552 17824 17558 17876
rect 18874 17864 18880 17876
rect 18835 17836 18880 17864
rect 18874 17824 18880 17836
rect 18932 17824 18938 17876
rect 19981 17867 20039 17873
rect 19981 17833 19993 17867
rect 20027 17864 20039 17867
rect 20530 17864 20536 17876
rect 20027 17836 20536 17864
rect 20027 17833 20039 17836
rect 19981 17827 20039 17833
rect 20530 17824 20536 17836
rect 20588 17824 20594 17876
rect 5629 17799 5687 17805
rect 5629 17765 5641 17799
rect 5675 17765 5687 17799
rect 5629 17759 5687 17765
rect 5721 17799 5779 17805
rect 5721 17765 5733 17799
rect 5767 17796 5779 17799
rect 7006 17796 7012 17808
rect 5767 17768 7012 17796
rect 5767 17765 5779 17768
rect 5721 17759 5779 17765
rect 7006 17756 7012 17768
rect 7064 17756 7070 17808
rect 7190 17796 7196 17808
rect 7151 17768 7196 17796
rect 7190 17756 7196 17768
rect 7248 17756 7254 17808
rect 7285 17799 7343 17805
rect 7285 17765 7297 17799
rect 7331 17796 7343 17799
rect 7558 17796 7564 17808
rect 7331 17768 7564 17796
rect 7331 17765 7343 17768
rect 7285 17759 7343 17765
rect 7558 17756 7564 17768
rect 7616 17756 7622 17808
rect 7834 17796 7840 17808
rect 7795 17768 7840 17796
rect 7834 17756 7840 17768
rect 7892 17796 7898 17808
rect 9398 17796 9404 17808
rect 7892 17768 9404 17796
rect 7892 17756 7898 17768
rect 9398 17756 9404 17768
rect 9456 17796 9462 17808
rect 9769 17799 9827 17805
rect 9769 17796 9781 17799
rect 9456 17768 9781 17796
rect 9456 17756 9462 17768
rect 9769 17765 9781 17768
rect 9815 17765 9827 17799
rect 9769 17759 9827 17765
rect 9858 17756 9864 17808
rect 9916 17796 9922 17808
rect 10413 17799 10471 17805
rect 9916 17768 9961 17796
rect 9916 17756 9922 17768
rect 10413 17765 10425 17799
rect 10459 17796 10471 17799
rect 10962 17796 10968 17808
rect 10459 17768 10968 17796
rect 10459 17765 10471 17768
rect 10413 17759 10471 17765
rect 10962 17756 10968 17768
rect 11020 17756 11026 17808
rect 11790 17756 11796 17808
rect 11848 17796 11854 17808
rect 13924 17796 13952 17824
rect 11848 17768 13952 17796
rect 11848 17756 11854 17768
rect 2130 17737 2136 17740
rect 2108 17731 2136 17737
rect 2108 17697 2120 17731
rect 2108 17691 2136 17697
rect 2130 17688 2136 17691
rect 2188 17688 2194 17740
rect 4614 17737 4620 17740
rect 4592 17731 4620 17737
rect 4592 17728 4604 17731
rect 4527 17700 4604 17728
rect 4592 17697 4604 17700
rect 4672 17728 4678 17740
rect 5442 17728 5448 17740
rect 4672 17700 5448 17728
rect 4592 17691 4620 17697
rect 4614 17688 4620 17691
rect 4672 17688 4678 17700
rect 5442 17688 5448 17700
rect 5500 17688 5506 17740
rect 12250 17728 12256 17740
rect 12211 17700 12256 17728
rect 12250 17688 12256 17700
rect 12308 17688 12314 17740
rect 12894 17728 12900 17740
rect 12855 17700 12900 17728
rect 12894 17688 12900 17700
rect 12952 17688 12958 17740
rect 13188 17737 13216 17768
rect 16022 17756 16028 17808
rect 16080 17796 16086 17808
rect 16346 17799 16404 17805
rect 16346 17796 16358 17799
rect 16080 17768 16358 17796
rect 16080 17756 16086 17768
rect 16346 17765 16358 17768
rect 16392 17765 16404 17799
rect 16346 17759 16404 17765
rect 18966 17756 18972 17808
rect 19024 17796 19030 17808
rect 19382 17799 19440 17805
rect 19382 17796 19394 17799
rect 19024 17768 19394 17796
rect 19024 17756 19030 17768
rect 19382 17765 19394 17768
rect 19428 17765 19440 17799
rect 19382 17759 19440 17765
rect 20714 17756 20720 17808
rect 20772 17796 20778 17808
rect 21085 17799 21143 17805
rect 21085 17796 21097 17799
rect 20772 17768 21097 17796
rect 20772 17756 20778 17768
rect 21085 17765 21097 17768
rect 21131 17796 21143 17799
rect 22278 17796 22284 17808
rect 21131 17768 22284 17796
rect 21131 17765 21143 17768
rect 21085 17759 21143 17765
rect 22278 17756 22284 17768
rect 22336 17756 22342 17808
rect 13173 17731 13231 17737
rect 13173 17697 13185 17731
rect 13219 17697 13231 17731
rect 13538 17728 13544 17740
rect 13451 17700 13544 17728
rect 13173 17691 13231 17697
rect 13538 17688 13544 17700
rect 13596 17728 13602 17740
rect 13814 17728 13820 17740
rect 13596 17700 13820 17728
rect 13596 17688 13602 17700
rect 13814 17688 13820 17700
rect 13872 17688 13878 17740
rect 17770 17728 17776 17740
rect 17731 17700 17776 17728
rect 17770 17688 17776 17700
rect 17828 17688 17834 17740
rect 15654 17620 15660 17672
rect 15712 17660 15718 17672
rect 16025 17663 16083 17669
rect 16025 17660 16037 17663
rect 15712 17632 16037 17660
rect 15712 17620 15718 17632
rect 16025 17629 16037 17632
rect 16071 17629 16083 17663
rect 19058 17660 19064 17672
rect 19019 17632 19064 17660
rect 16025 17623 16083 17629
rect 19058 17620 19064 17632
rect 19116 17620 19122 17672
rect 20717 17663 20775 17669
rect 20717 17629 20729 17663
rect 20763 17660 20775 17663
rect 20806 17660 20812 17672
rect 20763 17632 20812 17660
rect 20763 17629 20775 17632
rect 20717 17623 20775 17629
rect 20806 17620 20812 17632
rect 20864 17620 20870 17672
rect 20993 17663 21051 17669
rect 20993 17629 21005 17663
rect 21039 17660 21051 17663
rect 21634 17660 21640 17672
rect 21039 17632 21640 17660
rect 21039 17629 21051 17632
rect 20993 17623 21051 17629
rect 1394 17552 1400 17604
rect 1452 17592 1458 17604
rect 1673 17595 1731 17601
rect 1673 17592 1685 17595
rect 1452 17564 1685 17592
rect 1452 17552 1458 17564
rect 1673 17561 1685 17564
rect 1719 17592 1731 17595
rect 4062 17592 4068 17604
rect 1719 17564 4068 17592
rect 1719 17561 1731 17564
rect 1673 17555 1731 17561
rect 4062 17552 4068 17564
rect 4120 17552 4126 17604
rect 6181 17595 6239 17601
rect 6181 17561 6193 17595
rect 6227 17592 6239 17595
rect 7742 17592 7748 17604
rect 6227 17564 7748 17592
rect 6227 17561 6239 17564
rect 6181 17555 6239 17561
rect 7742 17552 7748 17564
rect 7800 17552 7806 17604
rect 20349 17595 20407 17601
rect 20349 17561 20361 17595
rect 20395 17592 20407 17595
rect 21008 17592 21036 17623
rect 21634 17620 21640 17632
rect 21692 17620 21698 17672
rect 22462 17660 22468 17672
rect 22423 17632 22468 17660
rect 22462 17620 22468 17632
rect 22520 17620 22526 17672
rect 21542 17592 21548 17604
rect 20395 17564 21036 17592
rect 21503 17564 21548 17592
rect 20395 17561 20407 17564
rect 20349 17555 20407 17561
rect 21542 17552 21548 17564
rect 21600 17552 21606 17604
rect 2179 17527 2237 17533
rect 2179 17493 2191 17527
rect 2225 17524 2237 17527
rect 2406 17524 2412 17536
rect 2225 17496 2412 17524
rect 2225 17493 2237 17496
rect 2179 17487 2237 17493
rect 2406 17484 2412 17496
rect 2464 17484 2470 17536
rect 4663 17527 4721 17533
rect 4663 17493 4675 17527
rect 4709 17524 4721 17527
rect 5074 17524 5080 17536
rect 4709 17496 5080 17524
rect 4709 17493 4721 17496
rect 4663 17487 4721 17493
rect 5074 17484 5080 17496
rect 5132 17484 5138 17536
rect 5258 17524 5264 17536
rect 5219 17496 5264 17524
rect 5258 17484 5264 17496
rect 5316 17484 5322 17536
rect 6914 17524 6920 17536
rect 6875 17496 6920 17524
rect 6914 17484 6920 17496
rect 6972 17484 6978 17536
rect 12069 17527 12127 17533
rect 12069 17493 12081 17527
rect 12115 17524 12127 17527
rect 12158 17524 12164 17536
rect 12115 17496 12164 17524
rect 12115 17493 12127 17496
rect 12069 17487 12127 17493
rect 12158 17484 12164 17496
rect 12216 17484 12222 17536
rect 14274 17524 14280 17536
rect 14235 17496 14280 17524
rect 14274 17484 14280 17496
rect 14332 17524 14338 17536
rect 14737 17527 14795 17533
rect 14737 17524 14749 17527
rect 14332 17496 14749 17524
rect 14332 17484 14338 17496
rect 14737 17493 14749 17496
rect 14783 17524 14795 17527
rect 15562 17524 15568 17536
rect 14783 17496 15568 17524
rect 14783 17493 14795 17496
rect 14737 17487 14795 17493
rect 15562 17484 15568 17496
rect 15620 17484 15626 17536
rect 15838 17524 15844 17536
rect 15799 17496 15844 17524
rect 15838 17484 15844 17496
rect 15896 17484 15902 17536
rect 17954 17524 17960 17536
rect 17915 17496 17960 17524
rect 17954 17484 17960 17496
rect 18012 17484 18018 17536
rect 18325 17527 18383 17533
rect 18325 17493 18337 17527
rect 18371 17524 18383 17527
rect 18414 17524 18420 17536
rect 18371 17496 18420 17524
rect 18371 17493 18383 17496
rect 18325 17487 18383 17493
rect 18414 17484 18420 17496
rect 18472 17484 18478 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 4062 17320 4068 17332
rect 4023 17292 4068 17320
rect 4062 17280 4068 17292
rect 4120 17280 4126 17332
rect 4614 17320 4620 17332
rect 4575 17292 4620 17320
rect 4614 17280 4620 17292
rect 4672 17280 4678 17332
rect 6273 17323 6331 17329
rect 6273 17289 6285 17323
rect 6319 17320 6331 17323
rect 7006 17320 7012 17332
rect 6319 17292 7012 17320
rect 6319 17289 6331 17292
rect 6273 17283 6331 17289
rect 7006 17280 7012 17292
rect 7064 17280 7070 17332
rect 7558 17280 7564 17332
rect 7616 17320 7622 17332
rect 7745 17323 7803 17329
rect 7745 17320 7757 17323
rect 7616 17292 7757 17320
rect 7616 17280 7622 17292
rect 7745 17289 7757 17292
rect 7791 17320 7803 17323
rect 8021 17323 8079 17329
rect 8021 17320 8033 17323
rect 7791 17292 8033 17320
rect 7791 17289 7803 17292
rect 7745 17283 7803 17289
rect 8021 17289 8033 17292
rect 8067 17289 8079 17323
rect 10778 17320 10784 17332
rect 10739 17292 10784 17320
rect 8021 17283 8079 17289
rect 10778 17280 10784 17292
rect 10836 17280 10842 17332
rect 11514 17320 11520 17332
rect 11475 17292 11520 17320
rect 11514 17280 11520 17292
rect 11572 17280 11578 17332
rect 11790 17320 11796 17332
rect 11751 17292 11796 17320
rect 11790 17280 11796 17292
rect 11848 17280 11854 17332
rect 13633 17323 13691 17329
rect 13633 17289 13645 17323
rect 13679 17320 13691 17323
rect 13906 17320 13912 17332
rect 13679 17292 13912 17320
rect 13679 17289 13691 17292
rect 13633 17283 13691 17289
rect 13906 17280 13912 17292
rect 13964 17280 13970 17332
rect 15197 17323 15255 17329
rect 15197 17289 15209 17323
rect 15243 17320 15255 17323
rect 15746 17320 15752 17332
rect 15243 17292 15752 17320
rect 15243 17289 15255 17292
rect 15197 17283 15255 17289
rect 15746 17280 15752 17292
rect 15804 17280 15810 17332
rect 15933 17323 15991 17329
rect 15933 17289 15945 17323
rect 15979 17320 15991 17323
rect 16022 17320 16028 17332
rect 15979 17292 16028 17320
rect 15979 17289 15991 17292
rect 15933 17283 15991 17289
rect 16022 17280 16028 17292
rect 16080 17320 16086 17332
rect 18601 17323 18659 17329
rect 18601 17320 18613 17323
rect 16080 17292 18613 17320
rect 16080 17280 16086 17292
rect 18601 17289 18613 17292
rect 18647 17320 18659 17323
rect 18966 17320 18972 17332
rect 18647 17292 18972 17320
rect 18647 17289 18659 17292
rect 18601 17283 18659 17289
rect 18966 17280 18972 17292
rect 19024 17280 19030 17332
rect 20714 17320 20720 17332
rect 20675 17292 20720 17320
rect 20714 17280 20720 17292
rect 20772 17280 20778 17332
rect 22278 17320 22284 17332
rect 22239 17292 22284 17320
rect 22278 17280 22284 17292
rect 22336 17280 22342 17332
rect 23017 17323 23075 17329
rect 23017 17289 23029 17323
rect 23063 17320 23075 17323
rect 23382 17320 23388 17332
rect 23063 17292 23388 17320
rect 23063 17289 23075 17292
rect 23017 17283 23075 17289
rect 11532 17252 11560 17280
rect 12342 17252 12348 17264
rect 11532 17224 12348 17252
rect 12342 17212 12348 17224
rect 12400 17212 12406 17264
rect 12158 17144 12164 17196
rect 12216 17184 12222 17196
rect 12805 17187 12863 17193
rect 12805 17184 12817 17187
rect 12216 17156 12817 17184
rect 12216 17144 12222 17156
rect 12805 17153 12817 17156
rect 12851 17153 12863 17187
rect 13924 17184 13952 17280
rect 20073 17255 20131 17261
rect 20073 17221 20085 17255
rect 20119 17252 20131 17255
rect 21082 17252 21088 17264
rect 20119 17224 21088 17252
rect 20119 17221 20131 17224
rect 20073 17215 20131 17221
rect 21082 17212 21088 17224
rect 21140 17212 21146 17264
rect 13924 17156 14596 17184
rect 12805 17147 12863 17153
rect 1394 17116 1400 17128
rect 1355 17088 1400 17116
rect 1394 17076 1400 17088
rect 1452 17076 1458 17128
rect 3580 17119 3638 17125
rect 3580 17085 3592 17119
rect 3626 17116 3638 17119
rect 4062 17116 4068 17128
rect 3626 17088 4068 17116
rect 3626 17085 3638 17088
rect 3580 17079 3638 17085
rect 4062 17076 4068 17088
rect 4120 17076 4126 17128
rect 5169 17119 5227 17125
rect 5169 17085 5181 17119
rect 5215 17085 5227 17119
rect 5169 17079 5227 17085
rect 1486 16940 1492 16992
rect 1544 16980 1550 16992
rect 1581 16983 1639 16989
rect 1581 16980 1593 16983
rect 1544 16952 1593 16980
rect 1544 16940 1550 16952
rect 1581 16949 1593 16952
rect 1627 16949 1639 16983
rect 2130 16980 2136 16992
rect 2091 16952 2136 16980
rect 1581 16943 1639 16949
rect 2130 16940 2136 16952
rect 2188 16940 2194 16992
rect 2501 16983 2559 16989
rect 2501 16949 2513 16983
rect 2547 16980 2559 16983
rect 2590 16980 2596 16992
rect 2547 16952 2596 16980
rect 2547 16949 2559 16952
rect 2501 16943 2559 16949
rect 2590 16940 2596 16952
rect 2648 16940 2654 16992
rect 2866 16940 2872 16992
rect 2924 16980 2930 16992
rect 3651 16983 3709 16989
rect 3651 16980 3663 16983
rect 2924 16952 3663 16980
rect 2924 16940 2930 16952
rect 3651 16949 3663 16952
rect 3697 16949 3709 16983
rect 3651 16943 3709 16949
rect 5077 16983 5135 16989
rect 5077 16949 5089 16983
rect 5123 16980 5135 16983
rect 5184 16980 5212 17079
rect 5258 17076 5264 17128
rect 5316 17116 5322 17128
rect 5629 17119 5687 17125
rect 5629 17116 5641 17119
rect 5316 17088 5641 17116
rect 5316 17076 5322 17088
rect 5629 17085 5641 17088
rect 5675 17085 5687 17119
rect 5629 17079 5687 17085
rect 6825 17119 6883 17125
rect 6825 17085 6837 17119
rect 6871 17116 6883 17119
rect 6914 17116 6920 17128
rect 6871 17088 6920 17116
rect 6871 17085 6883 17088
rect 6825 17079 6883 17085
rect 6914 17076 6920 17088
rect 6972 17076 6978 17128
rect 8849 17119 8907 17125
rect 8849 17085 8861 17119
rect 8895 17116 8907 17119
rect 9861 17119 9919 17125
rect 8895 17088 9444 17116
rect 8895 17085 8907 17088
rect 8849 17079 8907 17085
rect 5905 17051 5963 17057
rect 5905 17017 5917 17051
rect 5951 17048 5963 17051
rect 6270 17048 6276 17060
rect 5951 17020 6276 17048
rect 5951 17017 5963 17020
rect 5905 17011 5963 17017
rect 6270 17008 6276 17020
rect 6328 17008 6334 17060
rect 6638 17048 6644 17060
rect 6551 17020 6644 17048
rect 6638 17008 6644 17020
rect 6696 17048 6702 17060
rect 7187 17051 7245 17057
rect 7187 17048 7199 17051
rect 6696 17020 7199 17048
rect 6696 17008 6702 17020
rect 7187 17017 7199 17020
rect 7233 17048 7245 17051
rect 8202 17048 8208 17060
rect 7233 17020 8208 17048
rect 7233 17017 7245 17020
rect 7187 17011 7245 17017
rect 8202 17008 8208 17020
rect 8260 17008 8266 17060
rect 6546 16980 6552 16992
rect 5123 16952 6552 16980
rect 5123 16949 5135 16952
rect 5077 16943 5135 16949
rect 6546 16940 6552 16952
rect 6604 16940 6610 16992
rect 9030 16980 9036 16992
rect 8991 16952 9036 16980
rect 9030 16940 9036 16952
rect 9088 16940 9094 16992
rect 9416 16989 9444 17088
rect 9861 17085 9873 17119
rect 9907 17116 9919 17119
rect 9950 17116 9956 17128
rect 9907 17088 9956 17116
rect 9907 17085 9919 17088
rect 9861 17079 9919 17085
rect 9950 17076 9956 17088
rect 10008 17076 10014 17128
rect 14001 17119 14059 17125
rect 14001 17085 14013 17119
rect 14047 17116 14059 17119
rect 14369 17119 14427 17125
rect 14369 17116 14381 17119
rect 14047 17088 14381 17116
rect 14047 17085 14059 17088
rect 14001 17079 14059 17085
rect 14369 17085 14381 17088
rect 14415 17116 14427 17119
rect 14458 17116 14464 17128
rect 14415 17088 14464 17116
rect 14415 17085 14427 17088
rect 14369 17079 14427 17085
rect 14458 17076 14464 17088
rect 14516 17076 14522 17128
rect 14568 17125 14596 17156
rect 18966 17144 18972 17196
rect 19024 17184 19030 17196
rect 19024 17156 19288 17184
rect 19024 17144 19030 17156
rect 14553 17119 14611 17125
rect 14553 17085 14565 17119
rect 14599 17085 14611 17119
rect 14553 17079 14611 17085
rect 14921 17119 14979 17125
rect 14921 17085 14933 17119
rect 14967 17085 14979 17119
rect 14921 17079 14979 17085
rect 10182 17051 10240 17057
rect 10182 17048 10194 17051
rect 9784 17020 10194 17048
rect 9784 16992 9812 17020
rect 10182 17017 10194 17020
rect 10228 17017 10240 17051
rect 12526 17048 12532 17060
rect 12487 17020 12532 17048
rect 10182 17011 10240 17017
rect 12526 17008 12532 17020
rect 12584 17008 12590 17060
rect 12618 17008 12624 17060
rect 12676 17048 12682 17060
rect 12676 17020 12721 17048
rect 12676 17008 12682 17020
rect 13814 17008 13820 17060
rect 13872 17048 13878 17060
rect 14274 17048 14280 17060
rect 13872 17020 14280 17048
rect 13872 17008 13878 17020
rect 14274 17008 14280 17020
rect 14332 17048 14338 17060
rect 14936 17048 14964 17079
rect 15194 17076 15200 17128
rect 15252 17116 15258 17128
rect 15838 17116 15844 17128
rect 15252 17088 15844 17116
rect 15252 17076 15258 17088
rect 15838 17076 15844 17088
rect 15896 17116 15902 17128
rect 16025 17119 16083 17125
rect 16025 17116 16037 17119
rect 15896 17088 16037 17116
rect 15896 17076 15902 17088
rect 16025 17085 16037 17088
rect 16071 17085 16083 17119
rect 16025 17079 16083 17085
rect 18049 17119 18107 17125
rect 18049 17085 18061 17119
rect 18095 17116 18107 17119
rect 19153 17119 19211 17125
rect 18095 17088 18129 17116
rect 18095 17085 18107 17088
rect 18049 17079 18107 17085
rect 19153 17085 19165 17119
rect 19199 17085 19211 17119
rect 19153 17079 19211 17085
rect 14332 17020 14964 17048
rect 14332 17008 14338 17020
rect 16114 17008 16120 17060
rect 16172 17048 16178 17060
rect 16346 17051 16404 17057
rect 16346 17048 16358 17051
rect 16172 17020 16358 17048
rect 16172 17008 16178 17020
rect 16346 17017 16358 17020
rect 16392 17017 16404 17051
rect 16346 17011 16404 17017
rect 17497 17051 17555 17057
rect 17497 17017 17509 17051
rect 17543 17048 17555 17051
rect 17954 17048 17960 17060
rect 17543 17020 17960 17048
rect 17543 17017 17555 17020
rect 17497 17011 17555 17017
rect 17954 17008 17960 17020
rect 18012 17048 18018 17060
rect 18064 17048 18092 17079
rect 18322 17048 18328 17060
rect 18012 17020 18328 17048
rect 18012 17008 18018 17020
rect 18322 17008 18328 17020
rect 18380 17008 18386 17060
rect 9401 16983 9459 16989
rect 9401 16949 9413 16983
rect 9447 16980 9459 16983
rect 9490 16980 9496 16992
rect 9447 16952 9496 16980
rect 9447 16949 9459 16952
rect 9401 16943 9459 16949
rect 9490 16940 9496 16952
rect 9548 16940 9554 16992
rect 9766 16980 9772 16992
rect 9727 16952 9772 16980
rect 9766 16940 9772 16952
rect 9824 16940 9830 16992
rect 9858 16940 9864 16992
rect 9916 16980 9922 16992
rect 11057 16983 11115 16989
rect 11057 16980 11069 16983
rect 9916 16952 11069 16980
rect 9916 16940 9922 16952
rect 11057 16949 11069 16952
rect 11103 16949 11115 16983
rect 11057 16943 11115 16949
rect 11606 16940 11612 16992
rect 11664 16980 11670 16992
rect 12161 16983 12219 16989
rect 12161 16980 12173 16983
rect 11664 16952 12173 16980
rect 11664 16940 11670 16952
rect 12161 16949 12173 16952
rect 12207 16980 12219 16983
rect 12250 16980 12256 16992
rect 12207 16952 12256 16980
rect 12207 16949 12219 16952
rect 12161 16943 12219 16949
rect 12250 16940 12256 16952
rect 12308 16940 12314 16992
rect 12342 16940 12348 16992
rect 12400 16980 12406 16992
rect 13262 16980 13268 16992
rect 12400 16952 13268 16980
rect 12400 16940 12406 16952
rect 13262 16940 13268 16952
rect 13320 16980 13326 16992
rect 13538 16980 13544 16992
rect 13320 16952 13544 16980
rect 13320 16940 13326 16952
rect 13538 16940 13544 16952
rect 13596 16940 13602 16992
rect 15565 16983 15623 16989
rect 15565 16949 15577 16983
rect 15611 16980 15623 16983
rect 15654 16980 15660 16992
rect 15611 16952 15660 16980
rect 15611 16949 15623 16952
rect 15565 16943 15623 16949
rect 15654 16940 15660 16952
rect 15712 16940 15718 16992
rect 16942 16980 16948 16992
rect 16903 16952 16948 16980
rect 16942 16940 16948 16952
rect 17000 16940 17006 16992
rect 17770 16980 17776 16992
rect 17731 16952 17776 16980
rect 17770 16940 17776 16952
rect 17828 16940 17834 16992
rect 18230 16980 18236 16992
rect 18191 16952 18236 16980
rect 18230 16940 18236 16952
rect 18288 16940 18294 16992
rect 19168 16980 19196 17079
rect 19260 17048 19288 17156
rect 20806 17144 20812 17196
rect 20864 17184 20870 17196
rect 20993 17187 21051 17193
rect 20993 17184 21005 17187
rect 20864 17156 21005 17184
rect 20864 17144 20870 17156
rect 20993 17153 21005 17156
rect 21039 17153 21051 17187
rect 21634 17184 21640 17196
rect 21595 17156 21640 17184
rect 20993 17147 21051 17153
rect 21634 17144 21640 17156
rect 21692 17144 21698 17196
rect 22554 17125 22560 17128
rect 22532 17119 22560 17125
rect 22532 17085 22544 17119
rect 22612 17116 22618 17128
rect 23032 17116 23060 17283
rect 23382 17280 23388 17292
rect 23440 17280 23446 17332
rect 22612 17088 23060 17116
rect 22532 17079 22560 17085
rect 22554 17076 22560 17079
rect 22612 17076 22618 17088
rect 23658 17076 23664 17128
rect 23716 17125 23722 17128
rect 23716 17119 23754 17125
rect 23742 17116 23754 17119
rect 23742 17088 23888 17116
rect 23742 17085 23754 17088
rect 23716 17079 23754 17085
rect 23716 17076 23722 17079
rect 19474 17051 19532 17057
rect 19474 17048 19486 17051
rect 19260 17020 19486 17048
rect 19474 17017 19486 17020
rect 19520 17017 19532 17051
rect 19474 17011 19532 17017
rect 21085 17051 21143 17057
rect 21085 17017 21097 17051
rect 21131 17017 21143 17051
rect 23860 17048 23888 17088
rect 23934 17076 23940 17128
rect 23992 17116 23998 17128
rect 24708 17119 24766 17125
rect 24708 17116 24720 17119
rect 23992 17088 24720 17116
rect 23992 17076 23998 17088
rect 24708 17085 24720 17088
rect 24754 17116 24766 17119
rect 25133 17119 25191 17125
rect 25133 17116 25145 17119
rect 24754 17088 25145 17116
rect 24754 17085 24766 17088
rect 24708 17079 24766 17085
rect 25133 17085 25145 17088
rect 25179 17085 25191 17119
rect 25133 17079 25191 17085
rect 24121 17051 24179 17057
rect 24121 17048 24133 17051
rect 23860 17020 24133 17048
rect 21085 17011 21143 17017
rect 24121 17017 24133 17020
rect 24167 17048 24179 17051
rect 24946 17048 24952 17060
rect 24167 17020 24952 17048
rect 24167 17017 24179 17020
rect 24121 17011 24179 17017
rect 20441 16983 20499 16989
rect 20441 16980 20453 16983
rect 19168 16952 20453 16980
rect 20441 16949 20453 16952
rect 20487 16980 20499 16983
rect 20622 16980 20628 16992
rect 20487 16952 20628 16980
rect 20487 16949 20499 16952
rect 20441 16943 20499 16949
rect 20622 16940 20628 16952
rect 20680 16940 20686 16992
rect 20806 16940 20812 16992
rect 20864 16980 20870 16992
rect 21100 16980 21128 17011
rect 24946 17008 24952 17020
rect 25004 17008 25010 17060
rect 21913 16983 21971 16989
rect 21913 16980 21925 16983
rect 20864 16952 21925 16980
rect 20864 16940 20870 16952
rect 21913 16949 21925 16952
rect 21959 16949 21971 16983
rect 21913 16943 21971 16949
rect 22370 16940 22376 16992
rect 22428 16980 22434 16992
rect 23842 16989 23848 16992
rect 22603 16983 22661 16989
rect 22603 16980 22615 16983
rect 22428 16952 22615 16980
rect 22428 16940 22434 16952
rect 22603 16949 22615 16952
rect 22649 16949 22661 16983
rect 22603 16943 22661 16949
rect 23799 16983 23848 16989
rect 23799 16949 23811 16983
rect 23845 16949 23848 16983
rect 23799 16943 23848 16949
rect 23842 16940 23848 16943
rect 23900 16940 23906 16992
rect 24670 16940 24676 16992
rect 24728 16980 24734 16992
rect 24811 16983 24869 16989
rect 24811 16980 24823 16983
rect 24728 16952 24823 16980
rect 24728 16940 24734 16952
rect 24811 16949 24823 16952
rect 24857 16949 24869 16983
rect 24811 16943 24869 16949
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 1394 16736 1400 16788
rect 1452 16776 1458 16788
rect 1581 16779 1639 16785
rect 1581 16776 1593 16779
rect 1452 16748 1593 16776
rect 1452 16736 1458 16748
rect 1581 16745 1593 16748
rect 1627 16745 1639 16779
rect 1581 16739 1639 16745
rect 2406 16736 2412 16788
rect 2464 16776 2470 16788
rect 3329 16779 3387 16785
rect 3329 16776 3341 16779
rect 2464 16748 3341 16776
rect 2464 16736 2470 16748
rect 3329 16745 3341 16748
rect 3375 16745 3387 16779
rect 3329 16739 3387 16745
rect 5534 16736 5540 16788
rect 5592 16776 5598 16788
rect 5905 16779 5963 16785
rect 5905 16776 5917 16779
rect 5592 16748 5917 16776
rect 5592 16736 5598 16748
rect 5905 16745 5917 16748
rect 5951 16745 5963 16779
rect 7006 16776 7012 16788
rect 6967 16748 7012 16776
rect 5905 16739 5963 16745
rect 7006 16736 7012 16748
rect 7064 16736 7070 16788
rect 7190 16736 7196 16788
rect 7248 16776 7254 16788
rect 7653 16779 7711 16785
rect 7653 16776 7665 16779
rect 7248 16748 7665 16776
rect 7248 16736 7254 16748
rect 7653 16745 7665 16748
rect 7699 16745 7711 16779
rect 9398 16776 9404 16788
rect 9359 16748 9404 16776
rect 7653 16739 7711 16745
rect 9398 16736 9404 16748
rect 9456 16736 9462 16788
rect 10321 16779 10379 16785
rect 10321 16745 10333 16779
rect 10367 16776 10379 16779
rect 10962 16776 10968 16788
rect 10367 16748 10968 16776
rect 10367 16745 10379 16748
rect 10321 16739 10379 16745
rect 10962 16736 10968 16748
rect 11020 16736 11026 16788
rect 12069 16779 12127 16785
rect 12069 16745 12081 16779
rect 12115 16776 12127 16779
rect 12618 16776 12624 16788
rect 12115 16748 12624 16776
rect 12115 16745 12127 16748
rect 12069 16739 12127 16745
rect 12618 16736 12624 16748
rect 12676 16776 12682 16788
rect 13081 16779 13139 16785
rect 13081 16776 13093 16779
rect 12676 16748 13093 16776
rect 12676 16736 12682 16748
rect 13081 16745 13093 16748
rect 13127 16745 13139 16779
rect 13081 16739 13139 16745
rect 15378 16736 15384 16788
rect 15436 16776 15442 16788
rect 16022 16776 16028 16788
rect 15436 16748 16028 16776
rect 15436 16736 15442 16748
rect 16022 16736 16028 16748
rect 16080 16736 16086 16788
rect 19889 16779 19947 16785
rect 19889 16745 19901 16779
rect 19935 16776 19947 16779
rect 20806 16776 20812 16788
rect 19935 16748 20812 16776
rect 19935 16745 19947 16748
rect 19889 16739 19947 16745
rect 20806 16736 20812 16748
rect 20864 16736 20870 16788
rect 22370 16776 22376 16788
rect 21008 16748 22376 16776
rect 2314 16668 2320 16720
rect 2372 16708 2378 16720
rect 2639 16711 2697 16717
rect 2639 16708 2651 16711
rect 2372 16680 2651 16708
rect 2372 16668 2378 16680
rect 2639 16677 2651 16680
rect 2685 16677 2697 16711
rect 2639 16671 2697 16677
rect 6451 16711 6509 16717
rect 6451 16677 6463 16711
rect 6497 16708 6509 16711
rect 6638 16708 6644 16720
rect 6497 16680 6644 16708
rect 6497 16677 6509 16680
rect 6451 16671 6509 16677
rect 6638 16668 6644 16680
rect 6696 16668 6702 16720
rect 8202 16717 8208 16720
rect 8199 16708 8208 16717
rect 8163 16680 8208 16708
rect 8199 16671 8208 16680
rect 8202 16668 8208 16671
rect 8260 16668 8266 16720
rect 9766 16668 9772 16720
rect 9824 16708 9830 16720
rect 11470 16711 11528 16717
rect 11470 16708 11482 16711
rect 9824 16680 11482 16708
rect 9824 16668 9830 16680
rect 11470 16677 11482 16680
rect 11516 16677 11528 16711
rect 11470 16671 11528 16677
rect 12526 16668 12532 16720
rect 12584 16708 12590 16720
rect 12713 16711 12771 16717
rect 12713 16708 12725 16711
rect 12584 16680 12725 16708
rect 12584 16668 12590 16680
rect 12713 16677 12725 16680
rect 12759 16677 12771 16711
rect 14366 16708 14372 16720
rect 14327 16680 14372 16708
rect 12713 16671 12771 16677
rect 14366 16668 14372 16680
rect 14424 16668 14430 16720
rect 16669 16711 16727 16717
rect 16669 16677 16681 16711
rect 16715 16708 16727 16711
rect 16942 16708 16948 16720
rect 16715 16680 16948 16708
rect 16715 16677 16727 16680
rect 16669 16671 16727 16677
rect 16942 16668 16948 16680
rect 17000 16668 17006 16720
rect 18966 16668 18972 16720
rect 19024 16708 19030 16720
rect 19290 16711 19348 16717
rect 19290 16708 19302 16711
rect 19024 16680 19302 16708
rect 19024 16668 19030 16680
rect 19290 16677 19302 16680
rect 19336 16708 19348 16711
rect 19426 16708 19432 16720
rect 19336 16680 19432 16708
rect 19336 16677 19348 16680
rect 19290 16671 19348 16677
rect 19426 16668 19432 16680
rect 19484 16668 19490 16720
rect 20162 16708 20168 16720
rect 20123 16680 20168 16708
rect 20162 16668 20168 16680
rect 20220 16668 20226 16720
rect 21008 16717 21036 16748
rect 22370 16736 22376 16748
rect 22428 16736 22434 16788
rect 22646 16776 22652 16788
rect 22607 16748 22652 16776
rect 22646 16736 22652 16748
rect 22704 16736 22710 16788
rect 23750 16736 23756 16788
rect 23808 16776 23814 16788
rect 24673 16779 24731 16785
rect 24673 16776 24685 16779
rect 23808 16748 24685 16776
rect 23808 16736 23814 16748
rect 24673 16745 24685 16748
rect 24719 16745 24731 16779
rect 24673 16739 24731 16745
rect 20717 16711 20775 16717
rect 20717 16677 20729 16711
rect 20763 16708 20775 16711
rect 20993 16711 21051 16717
rect 20993 16708 21005 16711
rect 20763 16680 21005 16708
rect 20763 16677 20775 16680
rect 20717 16671 20775 16677
rect 20993 16677 21005 16680
rect 21039 16677 21051 16711
rect 20993 16671 21051 16677
rect 21082 16668 21088 16720
rect 21140 16708 21146 16720
rect 21634 16708 21640 16720
rect 21140 16680 21185 16708
rect 21595 16680 21640 16708
rect 21140 16668 21146 16680
rect 21634 16668 21640 16680
rect 21692 16668 21698 16720
rect 22664 16708 22692 16736
rect 22664 16680 24532 16708
rect 1397 16643 1455 16649
rect 1397 16609 1409 16643
rect 1443 16640 1455 16643
rect 2038 16640 2044 16652
rect 1443 16612 2044 16640
rect 1443 16609 1455 16612
rect 1397 16603 1455 16609
rect 2038 16600 2044 16612
rect 2096 16600 2102 16652
rect 2498 16600 2504 16652
rect 2556 16649 2562 16652
rect 2556 16643 2594 16649
rect 2582 16609 2594 16643
rect 2556 16603 2594 16609
rect 2556 16600 2562 16603
rect 2774 16600 2780 16652
rect 2832 16640 2838 16652
rect 2961 16643 3019 16649
rect 2961 16640 2973 16643
rect 2832 16612 2973 16640
rect 2832 16600 2838 16612
rect 2961 16609 2973 16612
rect 3007 16609 3019 16643
rect 4522 16640 4528 16652
rect 4483 16612 4528 16640
rect 2961 16603 3019 16609
rect 4522 16600 4528 16612
rect 4580 16600 4586 16652
rect 5077 16643 5135 16649
rect 5077 16609 5089 16643
rect 5123 16609 5135 16643
rect 5077 16603 5135 16609
rect 5261 16643 5319 16649
rect 5261 16609 5273 16643
rect 5307 16640 5319 16643
rect 5442 16640 5448 16652
rect 5307 16612 5448 16640
rect 5307 16609 5319 16612
rect 5261 16603 5319 16609
rect 5092 16572 5120 16603
rect 5442 16600 5448 16612
rect 5500 16600 5506 16652
rect 7837 16643 7895 16649
rect 7837 16609 7849 16643
rect 7883 16640 7895 16643
rect 8294 16640 8300 16652
rect 7883 16612 8300 16640
rect 7883 16609 7895 16612
rect 7837 16603 7895 16609
rect 8294 16600 8300 16612
rect 8352 16600 8358 16652
rect 8757 16643 8815 16649
rect 8757 16609 8769 16643
rect 8803 16640 8815 16643
rect 9858 16640 9864 16652
rect 8803 16612 9864 16640
rect 8803 16609 8815 16612
rect 8757 16603 8815 16609
rect 9858 16600 9864 16612
rect 9916 16600 9922 16652
rect 10134 16640 10140 16652
rect 10095 16612 10140 16640
rect 10134 16600 10140 16612
rect 10192 16600 10198 16652
rect 12437 16643 12495 16649
rect 12437 16609 12449 16643
rect 12483 16640 12495 16643
rect 12894 16640 12900 16652
rect 12483 16612 12900 16640
rect 12483 16609 12495 16612
rect 12437 16603 12495 16609
rect 12894 16600 12900 16612
rect 12952 16600 12958 16652
rect 13170 16600 13176 16652
rect 13228 16640 13234 16652
rect 13633 16643 13691 16649
rect 13633 16640 13645 16643
rect 13228 16612 13645 16640
rect 13228 16600 13234 16612
rect 13633 16609 13645 16612
rect 13679 16640 13691 16643
rect 13814 16640 13820 16652
rect 13679 16612 13820 16640
rect 13679 16609 13691 16612
rect 13633 16603 13691 16609
rect 13814 16600 13820 16612
rect 13872 16600 13878 16652
rect 13909 16643 13967 16649
rect 13909 16609 13921 16643
rect 13955 16640 13967 16643
rect 14458 16640 14464 16652
rect 13955 16612 14464 16640
rect 13955 16609 13967 16612
rect 13909 16603 13967 16609
rect 14458 16600 14464 16612
rect 14516 16640 14522 16652
rect 15286 16640 15292 16652
rect 14516 16612 15148 16640
rect 15247 16612 15292 16640
rect 14516 16600 14522 16612
rect 6086 16572 6092 16584
rect 5092 16544 5304 16572
rect 6047 16544 6092 16572
rect 5276 16448 5304 16544
rect 6086 16532 6092 16544
rect 6144 16532 6150 16584
rect 11149 16575 11207 16581
rect 11149 16541 11161 16575
rect 11195 16572 11207 16575
rect 11514 16572 11520 16584
rect 11195 16544 11520 16572
rect 11195 16541 11207 16544
rect 11149 16535 11207 16541
rect 11514 16532 11520 16544
rect 11572 16532 11578 16584
rect 15120 16572 15148 16612
rect 15286 16600 15292 16612
rect 15344 16640 15350 16652
rect 16390 16640 16396 16652
rect 15344 16612 16396 16640
rect 15344 16600 15350 16612
rect 16390 16600 16396 16612
rect 16448 16600 16454 16652
rect 19886 16600 19892 16652
rect 19944 16640 19950 16652
rect 20180 16640 20208 16668
rect 22462 16640 22468 16652
rect 19944 16612 20208 16640
rect 22423 16612 22468 16640
rect 19944 16600 19950 16612
rect 22462 16600 22468 16612
rect 22520 16600 22526 16652
rect 24504 16649 24532 16680
rect 23477 16643 23535 16649
rect 23477 16640 23489 16643
rect 23400 16612 23489 16640
rect 16577 16575 16635 16581
rect 15120 16544 15332 16572
rect 15304 16516 15332 16544
rect 16577 16541 16589 16575
rect 16623 16572 16635 16575
rect 17218 16572 17224 16584
rect 16623 16544 17224 16572
rect 16623 16541 16635 16544
rect 16577 16535 16635 16541
rect 17218 16532 17224 16544
rect 17276 16532 17282 16584
rect 18966 16572 18972 16584
rect 18927 16544 18972 16572
rect 18966 16532 18972 16544
rect 19024 16532 19030 16584
rect 23106 16532 23112 16584
rect 23164 16572 23170 16584
rect 23400 16572 23428 16612
rect 23477 16609 23489 16612
rect 23523 16609 23535 16643
rect 23477 16603 23535 16609
rect 24489 16643 24547 16649
rect 24489 16609 24501 16643
rect 24535 16640 24547 16643
rect 24762 16640 24768 16652
rect 24535 16612 24768 16640
rect 24535 16609 24547 16612
rect 24489 16603 24547 16609
rect 24762 16600 24768 16612
rect 24820 16600 24826 16652
rect 23164 16544 23428 16572
rect 23164 16532 23170 16544
rect 13722 16504 13728 16516
rect 13683 16476 13728 16504
rect 13722 16464 13728 16476
rect 13780 16464 13786 16516
rect 15286 16464 15292 16516
rect 15344 16464 15350 16516
rect 17126 16504 17132 16516
rect 17087 16476 17132 16504
rect 17126 16464 17132 16476
rect 17184 16464 17190 16516
rect 5258 16396 5264 16448
rect 5316 16436 5322 16448
rect 5537 16439 5595 16445
rect 5537 16436 5549 16439
rect 5316 16408 5549 16436
rect 5316 16396 5322 16408
rect 5537 16405 5549 16408
rect 5583 16405 5595 16439
rect 7282 16436 7288 16448
rect 7243 16408 7288 16436
rect 5537 16399 5595 16405
rect 7282 16396 7288 16408
rect 7340 16396 7346 16448
rect 9950 16436 9956 16448
rect 9911 16408 9956 16436
rect 9950 16396 9956 16408
rect 10008 16396 10014 16448
rect 10689 16439 10747 16445
rect 10689 16405 10701 16439
rect 10735 16436 10747 16439
rect 10962 16436 10968 16448
rect 10735 16408 10968 16436
rect 10735 16405 10747 16408
rect 10689 16399 10747 16405
rect 10962 16396 10968 16408
rect 11020 16396 11026 16448
rect 15470 16436 15476 16448
rect 15431 16408 15476 16436
rect 15470 16396 15476 16408
rect 15528 16396 15534 16448
rect 18322 16436 18328 16448
rect 18283 16408 18328 16436
rect 18322 16396 18328 16408
rect 18380 16396 18386 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 1578 16232 1584 16244
rect 1539 16204 1584 16232
rect 1578 16192 1584 16204
rect 1636 16192 1642 16244
rect 2409 16235 2467 16241
rect 2409 16201 2421 16235
rect 2455 16232 2467 16235
rect 2498 16232 2504 16244
rect 2455 16204 2504 16232
rect 2455 16201 2467 16204
rect 2409 16195 2467 16201
rect 2498 16192 2504 16204
rect 2556 16192 2562 16244
rect 4065 16235 4123 16241
rect 4065 16201 4077 16235
rect 4111 16232 4123 16235
rect 4522 16232 4528 16244
rect 4111 16204 4528 16232
rect 4111 16201 4123 16204
rect 4065 16195 4123 16201
rect 4522 16192 4528 16204
rect 4580 16192 4586 16244
rect 6273 16235 6331 16241
rect 6273 16201 6285 16235
rect 6319 16232 6331 16235
rect 6638 16232 6644 16244
rect 6319 16204 6644 16232
rect 6319 16201 6331 16204
rect 6273 16195 6331 16201
rect 6638 16192 6644 16204
rect 6696 16192 6702 16244
rect 8294 16232 8300 16244
rect 8255 16204 8300 16232
rect 8294 16192 8300 16204
rect 8352 16192 8358 16244
rect 10686 16232 10692 16244
rect 10647 16204 10692 16232
rect 10686 16192 10692 16204
rect 10744 16192 10750 16244
rect 11514 16232 11520 16244
rect 11475 16204 11520 16232
rect 11514 16192 11520 16204
rect 11572 16192 11578 16244
rect 15286 16232 15292 16244
rect 15247 16204 15292 16232
rect 15286 16192 15292 16204
rect 15344 16192 15350 16244
rect 16574 16192 16580 16244
rect 16632 16232 16638 16244
rect 16761 16235 16819 16241
rect 16761 16232 16773 16235
rect 16632 16204 16773 16232
rect 16632 16192 16638 16204
rect 16761 16201 16773 16204
rect 16807 16201 16819 16235
rect 17218 16232 17224 16244
rect 17179 16204 17224 16232
rect 16761 16195 16819 16201
rect 17218 16192 17224 16204
rect 17276 16192 17282 16244
rect 19337 16235 19395 16241
rect 19337 16201 19349 16235
rect 19383 16232 19395 16235
rect 19426 16232 19432 16244
rect 19383 16204 19432 16232
rect 19383 16201 19395 16204
rect 19337 16195 19395 16201
rect 19426 16192 19432 16204
rect 19484 16192 19490 16244
rect 21174 16232 21180 16244
rect 21135 16204 21180 16232
rect 21174 16192 21180 16204
rect 21232 16192 21238 16244
rect 24762 16232 24768 16244
rect 24723 16204 24768 16232
rect 24762 16192 24768 16204
rect 24820 16192 24826 16244
rect 4540 16164 4568 16192
rect 6178 16164 6184 16176
rect 4540 16136 6184 16164
rect 6178 16124 6184 16136
rect 6236 16164 6242 16176
rect 6549 16167 6607 16173
rect 6549 16164 6561 16167
rect 6236 16136 6561 16164
rect 6236 16124 6242 16136
rect 6549 16133 6561 16136
rect 6595 16133 6607 16167
rect 6549 16127 6607 16133
rect 9309 16167 9367 16173
rect 9309 16133 9321 16167
rect 9355 16164 9367 16167
rect 10134 16164 10140 16176
rect 9355 16136 10140 16164
rect 9355 16133 9367 16136
rect 9309 16127 9367 16133
rect 2406 16056 2412 16108
rect 2464 16096 2470 16108
rect 2593 16099 2651 16105
rect 2593 16096 2605 16099
rect 2464 16068 2605 16096
rect 2464 16056 2470 16068
rect 2593 16065 2605 16068
rect 2639 16065 2651 16099
rect 2593 16059 2651 16065
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 16028 1455 16031
rect 1670 16028 1676 16040
rect 1443 16000 1676 16028
rect 1443 15997 1455 16000
rect 1397 15991 1455 15997
rect 1670 15988 1676 16000
rect 1728 15988 1734 16040
rect 4246 16037 4252 16040
rect 4224 16031 4252 16037
rect 4224 15997 4236 16031
rect 4304 16028 4310 16040
rect 4617 16031 4675 16037
rect 4617 16028 4629 16031
rect 4304 16000 4629 16028
rect 4224 15991 4252 15997
rect 4246 15988 4252 15991
rect 4304 15988 4310 16000
rect 4617 15997 4629 16000
rect 4663 16028 4675 16031
rect 4982 16028 4988 16040
rect 4663 16000 4988 16028
rect 4663 15997 4675 16000
rect 4617 15991 4675 15997
rect 4982 15988 4988 16000
rect 5040 15988 5046 16040
rect 5077 16031 5135 16037
rect 5077 15997 5089 16031
rect 5123 16028 5135 16031
rect 5166 16028 5172 16040
rect 5123 16000 5172 16028
rect 5123 15997 5135 16000
rect 5077 15991 5135 15997
rect 5166 15988 5172 16000
rect 5224 15988 5230 16040
rect 5258 15988 5264 16040
rect 5316 16028 5322 16040
rect 5629 16031 5687 16037
rect 5629 16028 5641 16031
rect 5316 16000 5641 16028
rect 5316 15988 5322 16000
rect 5629 15997 5641 16000
rect 5675 15997 5687 16031
rect 6564 16028 6592 16127
rect 10134 16124 10140 16136
rect 10192 16124 10198 16176
rect 15378 16164 15384 16176
rect 11164 16136 15384 16164
rect 7929 16099 7987 16105
rect 7929 16065 7941 16099
rect 7975 16096 7987 16099
rect 8202 16096 8208 16108
rect 7975 16068 8208 16096
rect 7975 16065 7987 16068
rect 7929 16059 7987 16065
rect 8202 16056 8208 16068
rect 8260 16096 8266 16108
rect 9677 16099 9735 16105
rect 9677 16096 9689 16099
rect 8260 16068 9689 16096
rect 8260 16056 8266 16068
rect 9677 16065 9689 16068
rect 9723 16065 9735 16099
rect 9677 16059 9735 16065
rect 9769 16099 9827 16105
rect 9769 16065 9781 16099
rect 9815 16096 9827 16099
rect 10962 16096 10968 16108
rect 9815 16068 10968 16096
rect 9815 16065 9827 16068
rect 9769 16059 9827 16065
rect 6825 16031 6883 16037
rect 6825 16028 6837 16031
rect 6564 16000 6837 16028
rect 5629 15991 5687 15997
rect 6825 15997 6837 16000
rect 6871 15997 6883 16031
rect 6825 15991 6883 15997
rect 7282 15988 7288 16040
rect 7340 16028 7346 16040
rect 7377 16031 7435 16037
rect 7377 16028 7389 16031
rect 7340 16000 7389 16028
rect 7340 15988 7346 16000
rect 7377 15997 7389 16000
rect 7423 16028 7435 16031
rect 8110 16028 8116 16040
rect 7423 16000 8116 16028
rect 7423 15997 7435 16000
rect 7377 15991 7435 15997
rect 8110 15988 8116 16000
rect 8168 15988 8174 16040
rect 8757 16031 8815 16037
rect 8757 16028 8769 16031
rect 8680 16000 8769 16028
rect 2222 15920 2228 15972
rect 2280 15960 2286 15972
rect 2685 15963 2743 15969
rect 2685 15960 2697 15963
rect 2280 15932 2697 15960
rect 2280 15920 2286 15932
rect 2685 15929 2697 15932
rect 2731 15960 2743 15963
rect 2774 15960 2780 15972
rect 2731 15932 2780 15960
rect 2731 15929 2743 15932
rect 2685 15923 2743 15929
rect 2774 15920 2780 15932
rect 2832 15920 2838 15972
rect 3234 15960 3240 15972
rect 3195 15932 3240 15960
rect 3234 15920 3240 15932
rect 3292 15920 3298 15972
rect 3697 15963 3755 15969
rect 3697 15929 3709 15963
rect 3743 15960 3755 15963
rect 5276 15960 5304 15988
rect 3743 15932 5304 15960
rect 5905 15963 5963 15969
rect 3743 15929 3755 15932
rect 3697 15923 3755 15929
rect 5905 15929 5917 15963
rect 5951 15960 5963 15963
rect 6730 15960 6736 15972
rect 5951 15932 6736 15960
rect 5951 15929 5963 15932
rect 5905 15923 5963 15929
rect 6730 15920 6736 15932
rect 6788 15920 6794 15972
rect 8680 15904 8708 16000
rect 8757 15997 8769 16000
rect 8803 15997 8815 16031
rect 8757 15991 8815 15997
rect 9692 15960 9720 16059
rect 10962 16056 10968 16068
rect 11020 16056 11026 16108
rect 9766 15960 9772 15972
rect 9692 15932 9772 15960
rect 9766 15920 9772 15932
rect 9824 15960 9830 15972
rect 11164 15969 11192 16136
rect 15378 16124 15384 16136
rect 15436 16124 15442 16176
rect 20809 16167 20867 16173
rect 20809 16164 20821 16167
rect 18708 16136 20821 16164
rect 14826 16096 14832 16108
rect 14787 16068 14832 16096
rect 14826 16056 14832 16068
rect 14884 16056 14890 16108
rect 12529 16031 12587 16037
rect 12529 16028 12541 16031
rect 12176 16000 12541 16028
rect 10090 15963 10148 15969
rect 10090 15960 10102 15963
rect 9824 15932 10102 15960
rect 9824 15920 9830 15932
rect 10090 15929 10102 15932
rect 10136 15960 10148 15963
rect 11149 15963 11207 15969
rect 11149 15960 11161 15963
rect 10136 15932 11161 15960
rect 10136 15929 10148 15932
rect 10090 15923 10148 15929
rect 11149 15929 11161 15932
rect 11195 15929 11207 15963
rect 11149 15923 11207 15929
rect 12176 15904 12204 16000
rect 12529 15997 12541 16000
rect 12575 16028 12587 16031
rect 13633 16031 13691 16037
rect 13633 16028 13645 16031
rect 12575 16000 13645 16028
rect 12575 15997 12587 16000
rect 12529 15991 12587 15997
rect 13633 15997 13645 16000
rect 13679 16028 13691 16031
rect 13722 16028 13728 16040
rect 13679 16000 13728 16028
rect 13679 15997 13691 16000
rect 13633 15991 13691 15997
rect 13722 15988 13728 16000
rect 13780 15988 13786 16040
rect 14182 16028 14188 16040
rect 14143 16000 14188 16028
rect 14182 15988 14188 16000
rect 14240 15988 14246 16040
rect 14645 16031 14703 16037
rect 14645 15997 14657 16031
rect 14691 15997 14703 16031
rect 15746 16028 15752 16040
rect 15707 16000 15752 16028
rect 14645 15991 14703 15997
rect 13173 15963 13231 15969
rect 13173 15929 13185 15963
rect 13219 15960 13231 15963
rect 13354 15960 13360 15972
rect 13219 15932 13360 15960
rect 13219 15929 13231 15932
rect 13173 15923 13231 15929
rect 13354 15920 13360 15932
rect 13412 15920 13418 15972
rect 14660 15960 14688 15991
rect 15746 15988 15752 16000
rect 15804 15988 15810 16040
rect 16209 16031 16267 16037
rect 16209 15997 16221 16031
rect 16255 15997 16267 16031
rect 16209 15991 16267 15997
rect 15565 15963 15623 15969
rect 15565 15960 15577 15963
rect 14108 15932 15577 15960
rect 14108 15904 14136 15932
rect 15565 15929 15577 15932
rect 15611 15960 15623 15963
rect 16224 15960 16252 15991
rect 16390 15988 16396 16040
rect 16448 16028 16454 16040
rect 18233 16031 18291 16037
rect 18233 16028 18245 16031
rect 16448 16000 18245 16028
rect 16448 15988 16454 16000
rect 18233 15997 18245 16000
rect 18279 16028 18291 16031
rect 18322 16028 18328 16040
rect 18279 16000 18328 16028
rect 18279 15997 18291 16000
rect 18233 15991 18291 15997
rect 18322 15988 18328 16000
rect 18380 15988 18386 16040
rect 18708 16037 18736 16136
rect 20809 16133 20821 16136
rect 20855 16133 20867 16167
rect 20809 16127 20867 16133
rect 18969 16099 19027 16105
rect 18969 16065 18981 16099
rect 19015 16096 19027 16099
rect 19242 16096 19248 16108
rect 19015 16068 19248 16096
rect 19015 16065 19027 16068
rect 18969 16059 19027 16065
rect 19242 16056 19248 16068
rect 19300 16056 19306 16108
rect 19426 16056 19432 16108
rect 19484 16096 19490 16108
rect 20165 16099 20223 16105
rect 20165 16096 20177 16099
rect 19484 16068 20177 16096
rect 19484 16056 19490 16068
rect 20165 16065 20177 16068
rect 20211 16065 20223 16099
rect 20824 16096 20852 16127
rect 23109 16099 23167 16105
rect 20824 16068 21864 16096
rect 20165 16059 20223 16065
rect 18693 16031 18751 16037
rect 18693 15997 18705 16031
rect 18739 15997 18751 16031
rect 18693 15991 18751 15997
rect 17494 15960 17500 15972
rect 15611 15932 17500 15960
rect 15611 15929 15623 15932
rect 15565 15923 15623 15929
rect 17494 15920 17500 15932
rect 17552 15960 17558 15972
rect 17773 15963 17831 15969
rect 17773 15960 17785 15963
rect 17552 15932 17785 15960
rect 17552 15920 17558 15932
rect 17773 15929 17785 15932
rect 17819 15960 17831 15963
rect 18046 15960 18052 15972
rect 17819 15932 18052 15960
rect 17819 15929 17831 15932
rect 17773 15923 17831 15929
rect 18046 15920 18052 15932
rect 18104 15960 18110 15972
rect 18708 15960 18736 15991
rect 21174 15988 21180 16040
rect 21232 16028 21238 16040
rect 21836 16037 21864 16068
rect 23109 16065 23121 16099
rect 23155 16096 23167 16099
rect 23753 16099 23811 16105
rect 23753 16096 23765 16099
rect 23155 16068 23765 16096
rect 23155 16065 23167 16068
rect 23109 16059 23167 16065
rect 23753 16065 23765 16068
rect 23799 16096 23811 16099
rect 25363 16099 25421 16105
rect 25363 16096 25375 16099
rect 23799 16068 25375 16096
rect 23799 16065 23811 16068
rect 23753 16059 23811 16065
rect 25363 16065 25375 16068
rect 25409 16065 25421 16099
rect 25363 16059 25421 16065
rect 21361 16031 21419 16037
rect 21361 16028 21373 16031
rect 21232 16000 21373 16028
rect 21232 15988 21238 16000
rect 21361 15997 21373 16000
rect 21407 15997 21419 16031
rect 21361 15991 21419 15997
rect 21821 16031 21879 16037
rect 21821 15997 21833 16031
rect 21867 15997 21879 16031
rect 22462 16028 22468 16040
rect 22423 16000 22468 16028
rect 21821 15991 21879 15997
rect 22462 15988 22468 16000
rect 22520 15988 22526 16040
rect 25222 15988 25228 16040
rect 25280 16037 25286 16040
rect 25280 16031 25318 16037
rect 25306 16028 25318 16031
rect 25685 16031 25743 16037
rect 25685 16028 25697 16031
rect 25306 16000 25697 16028
rect 25306 15997 25318 16000
rect 25280 15991 25318 15997
rect 25685 15997 25697 16000
rect 25731 15997 25743 16031
rect 25685 15991 25743 15997
rect 25280 15988 25286 15991
rect 19886 15960 19892 15972
rect 18104 15932 18736 15960
rect 19847 15932 19892 15960
rect 18104 15920 18110 15932
rect 19886 15920 19892 15932
rect 19944 15920 19950 15972
rect 19978 15920 19984 15972
rect 20036 15960 20042 15972
rect 20036 15932 20081 15960
rect 20036 15920 20042 15932
rect 20714 15920 20720 15972
rect 20772 15960 20778 15972
rect 23845 15963 23903 15969
rect 23845 15960 23857 15963
rect 20772 15932 21496 15960
rect 20772 15920 20778 15932
rect 2038 15892 2044 15904
rect 1999 15864 2044 15892
rect 2038 15852 2044 15864
rect 2096 15852 2102 15904
rect 4295 15895 4353 15901
rect 4295 15861 4307 15895
rect 4341 15892 4353 15895
rect 4890 15892 4896 15904
rect 4341 15864 4896 15892
rect 4341 15861 4353 15864
rect 4295 15855 4353 15861
rect 4890 15852 4896 15864
rect 4948 15852 4954 15904
rect 6914 15892 6920 15904
rect 6875 15864 6920 15892
rect 6914 15852 6920 15864
rect 6972 15852 6978 15904
rect 8662 15892 8668 15904
rect 8623 15864 8668 15892
rect 8662 15852 8668 15864
rect 8720 15852 8726 15904
rect 8938 15892 8944 15904
rect 8899 15864 8944 15892
rect 8938 15852 8944 15864
rect 8996 15852 9002 15904
rect 12158 15892 12164 15904
rect 12119 15864 12164 15892
rect 12158 15852 12164 15864
rect 12216 15852 12222 15904
rect 14090 15892 14096 15904
rect 14051 15864 14096 15892
rect 14090 15852 14096 15864
rect 14148 15852 14154 15904
rect 15654 15852 15660 15904
rect 15712 15892 15718 15904
rect 15841 15895 15899 15901
rect 15841 15892 15853 15895
rect 15712 15864 15853 15892
rect 15712 15852 15718 15864
rect 15841 15861 15853 15864
rect 15887 15861 15899 15895
rect 15841 15855 15899 15861
rect 19705 15895 19763 15901
rect 19705 15861 19717 15895
rect 19751 15892 19763 15895
rect 19996 15892 20024 15920
rect 21468 15901 21496 15932
rect 23492 15932 23857 15960
rect 23492 15904 23520 15932
rect 23845 15929 23857 15932
rect 23891 15929 23903 15963
rect 24394 15960 24400 15972
rect 24355 15932 24400 15960
rect 23845 15923 23903 15929
rect 24394 15920 24400 15932
rect 24452 15920 24458 15972
rect 19751 15864 20024 15892
rect 21453 15895 21511 15901
rect 19751 15861 19763 15864
rect 19705 15855 19763 15861
rect 21453 15861 21465 15895
rect 21499 15861 21511 15895
rect 23474 15892 23480 15904
rect 23435 15864 23480 15892
rect 21453 15855 21511 15861
rect 23474 15852 23480 15864
rect 23532 15852 23538 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 4430 15648 4436 15700
rect 4488 15688 4494 15700
rect 4709 15691 4767 15697
rect 4709 15688 4721 15691
rect 4488 15660 4721 15688
rect 4488 15648 4494 15660
rect 4709 15657 4721 15660
rect 4755 15657 4767 15691
rect 4709 15651 4767 15657
rect 5997 15691 6055 15697
rect 5997 15657 6009 15691
rect 6043 15688 6055 15691
rect 6086 15688 6092 15700
rect 6043 15660 6092 15688
rect 6043 15657 6055 15660
rect 5997 15651 6055 15657
rect 6086 15648 6092 15660
rect 6144 15688 6150 15700
rect 6549 15691 6607 15697
rect 6549 15688 6561 15691
rect 6144 15660 6561 15688
rect 6144 15648 6150 15660
rect 6549 15657 6561 15660
rect 6595 15657 6607 15691
rect 6549 15651 6607 15657
rect 6914 15648 6920 15700
rect 6972 15688 6978 15700
rect 7469 15691 7527 15697
rect 7469 15688 7481 15691
rect 6972 15660 7481 15688
rect 6972 15648 6978 15660
rect 7469 15657 7481 15660
rect 7515 15657 7527 15691
rect 8294 15688 8300 15700
rect 8255 15660 8300 15688
rect 7469 15651 7527 15657
rect 8294 15648 8300 15660
rect 8352 15648 8358 15700
rect 9122 15688 9128 15700
rect 9083 15660 9128 15688
rect 9122 15648 9128 15660
rect 9180 15648 9186 15700
rect 9950 15688 9956 15700
rect 9911 15660 9956 15688
rect 9950 15648 9956 15660
rect 10008 15648 10014 15700
rect 10781 15691 10839 15697
rect 10781 15657 10793 15691
rect 10827 15688 10839 15691
rect 11330 15688 11336 15700
rect 10827 15660 11336 15688
rect 10827 15657 10839 15660
rect 10781 15651 10839 15657
rect 2498 15580 2504 15632
rect 2556 15620 2562 15632
rect 2593 15623 2651 15629
rect 2593 15620 2605 15623
rect 2556 15592 2605 15620
rect 2556 15580 2562 15592
rect 2593 15589 2605 15592
rect 2639 15589 2651 15623
rect 2593 15583 2651 15589
rect 3145 15623 3203 15629
rect 3145 15589 3157 15623
rect 3191 15620 3203 15623
rect 3234 15620 3240 15632
rect 3191 15592 3240 15620
rect 3191 15589 3203 15592
rect 3145 15583 3203 15589
rect 3234 15580 3240 15592
rect 3292 15580 3298 15632
rect 6365 15623 6423 15629
rect 6365 15589 6377 15623
rect 6411 15620 6423 15623
rect 6411 15592 7052 15620
rect 6411 15589 6423 15592
rect 6365 15583 6423 15589
rect 1464 15555 1522 15561
rect 1464 15521 1476 15555
rect 1510 15552 1522 15555
rect 1854 15552 1860 15564
rect 1510 15524 1860 15552
rect 1510 15521 1522 15524
rect 1464 15515 1522 15521
rect 1854 15512 1860 15524
rect 1912 15512 1918 15564
rect 4798 15552 4804 15564
rect 4759 15524 4804 15552
rect 4798 15512 4804 15524
rect 4856 15512 4862 15564
rect 5077 15555 5135 15561
rect 5077 15521 5089 15555
rect 5123 15552 5135 15555
rect 6546 15552 6552 15564
rect 5123 15524 5212 15552
rect 6507 15524 6552 15552
rect 5123 15521 5135 15524
rect 5077 15515 5135 15521
rect 5184 15496 5212 15524
rect 6546 15512 6552 15524
rect 6604 15512 6610 15564
rect 7024 15561 7052 15592
rect 7009 15555 7067 15561
rect 7009 15521 7021 15555
rect 7055 15552 7067 15555
rect 7282 15552 7288 15564
rect 7055 15524 7288 15552
rect 7055 15521 7067 15524
rect 7009 15515 7067 15521
rect 7282 15512 7288 15524
rect 7340 15512 7346 15564
rect 8018 15552 8024 15564
rect 7979 15524 8024 15552
rect 8018 15512 8024 15524
rect 8076 15512 8082 15564
rect 8110 15512 8116 15564
rect 8168 15552 8174 15564
rect 8573 15555 8631 15561
rect 8573 15552 8585 15555
rect 8168 15524 8585 15552
rect 8168 15512 8174 15524
rect 8573 15521 8585 15524
rect 8619 15521 8631 15555
rect 9766 15552 9772 15564
rect 9727 15524 9772 15552
rect 8573 15515 8631 15521
rect 2498 15484 2504 15496
rect 2459 15456 2504 15484
rect 2498 15444 2504 15456
rect 2556 15484 2562 15496
rect 2866 15484 2872 15496
rect 2556 15456 2872 15484
rect 2556 15444 2562 15456
rect 2866 15444 2872 15456
rect 2924 15444 2930 15496
rect 5166 15444 5172 15496
rect 5224 15444 5230 15496
rect 8588 15484 8616 15515
rect 9766 15512 9772 15524
rect 9824 15512 9830 15564
rect 10229 15555 10287 15561
rect 10229 15521 10241 15555
rect 10275 15552 10287 15555
rect 10796 15552 10824 15651
rect 11330 15648 11336 15660
rect 11388 15648 11394 15700
rect 11514 15688 11520 15700
rect 11475 15660 11520 15688
rect 11514 15648 11520 15660
rect 11572 15648 11578 15700
rect 14182 15648 14188 15700
rect 14240 15688 14246 15700
rect 14645 15691 14703 15697
rect 14645 15688 14657 15691
rect 14240 15660 14657 15688
rect 14240 15648 14246 15660
rect 14645 15657 14657 15660
rect 14691 15657 14703 15691
rect 15746 15688 15752 15700
rect 15707 15660 15752 15688
rect 14645 15651 14703 15657
rect 15746 15648 15752 15660
rect 15804 15648 15810 15700
rect 16942 15688 16948 15700
rect 16903 15660 16948 15688
rect 16942 15648 16948 15660
rect 17000 15648 17006 15700
rect 17494 15648 17500 15700
rect 17552 15648 17558 15700
rect 20717 15691 20775 15697
rect 20717 15657 20729 15691
rect 20763 15688 20775 15691
rect 21082 15688 21088 15700
rect 20763 15660 21088 15688
rect 20763 15657 20775 15660
rect 20717 15651 20775 15657
rect 21082 15648 21088 15660
rect 21140 15648 21146 15700
rect 24118 15688 24124 15700
rect 24079 15660 24124 15688
rect 24118 15648 24124 15660
rect 24176 15648 24182 15700
rect 24762 15688 24768 15700
rect 24723 15660 24768 15688
rect 24762 15648 24768 15660
rect 24820 15648 24826 15700
rect 10275 15524 10824 15552
rect 11241 15555 11299 15561
rect 10275 15521 10287 15524
rect 10229 15515 10287 15521
rect 11241 15521 11253 15555
rect 11287 15521 11299 15555
rect 11348 15552 11376 15648
rect 17512 15620 17540 15648
rect 18233 15623 18291 15629
rect 17512 15592 18000 15620
rect 11698 15552 11704 15564
rect 11348 15524 11704 15552
rect 11241 15515 11299 15521
rect 9030 15484 9036 15496
rect 8588 15456 9036 15484
rect 9030 15444 9036 15456
rect 9088 15484 9094 15496
rect 10244 15484 10272 15515
rect 9088 15456 10272 15484
rect 11256 15484 11284 15515
rect 11698 15512 11704 15524
rect 11756 15512 11762 15564
rect 13262 15552 13268 15564
rect 13223 15524 13268 15552
rect 13262 15512 13268 15524
rect 13320 15512 13326 15564
rect 13354 15512 13360 15564
rect 13412 15552 13418 15564
rect 13538 15552 13544 15564
rect 13412 15524 13457 15552
rect 13499 15524 13544 15552
rect 13412 15512 13418 15524
rect 13538 15512 13544 15524
rect 13596 15512 13602 15564
rect 16022 15552 16028 15564
rect 15983 15524 16028 15552
rect 16022 15512 16028 15524
rect 16080 15512 16086 15564
rect 16114 15512 16120 15564
rect 16172 15552 16178 15564
rect 16390 15552 16396 15564
rect 16172 15524 16396 15552
rect 16172 15512 16178 15524
rect 16390 15512 16396 15524
rect 16448 15512 16454 15564
rect 16574 15512 16580 15564
rect 16632 15552 16638 15564
rect 17497 15555 17555 15561
rect 17497 15552 17509 15555
rect 16632 15524 17509 15552
rect 16632 15512 16638 15524
rect 17497 15521 17509 15524
rect 17543 15552 17555 15555
rect 17862 15552 17868 15564
rect 17543 15524 17868 15552
rect 17543 15521 17555 15524
rect 17497 15515 17555 15521
rect 17862 15512 17868 15524
rect 17920 15512 17926 15564
rect 17972 15561 18000 15592
rect 18233 15589 18245 15623
rect 18279 15620 18291 15623
rect 18877 15623 18935 15629
rect 18877 15620 18889 15623
rect 18279 15592 18889 15620
rect 18279 15589 18291 15592
rect 18233 15583 18291 15589
rect 18877 15589 18889 15592
rect 18923 15620 18935 15623
rect 18966 15620 18972 15632
rect 18923 15592 18972 15620
rect 18923 15589 18935 15592
rect 18877 15583 18935 15589
rect 18966 15580 18972 15592
rect 19024 15580 19030 15632
rect 19423 15623 19481 15629
rect 19423 15589 19435 15623
rect 19469 15620 19481 15623
rect 19518 15620 19524 15632
rect 19469 15592 19524 15620
rect 19469 15589 19481 15592
rect 19423 15583 19481 15589
rect 19518 15580 19524 15592
rect 19576 15580 19582 15632
rect 21266 15620 21272 15632
rect 21227 15592 21272 15620
rect 21266 15580 21272 15592
rect 21324 15580 21330 15632
rect 23106 15620 23112 15632
rect 23067 15592 23112 15620
rect 23106 15580 23112 15592
rect 23164 15580 23170 15632
rect 23198 15580 23204 15632
rect 23256 15620 23262 15632
rect 23256 15592 23301 15620
rect 23256 15580 23262 15592
rect 23566 15580 23572 15632
rect 23624 15620 23630 15632
rect 23753 15623 23811 15629
rect 23753 15620 23765 15623
rect 23624 15592 23765 15620
rect 23624 15580 23630 15592
rect 23753 15589 23765 15592
rect 23799 15620 23811 15623
rect 24394 15620 24400 15632
rect 23799 15592 24400 15620
rect 23799 15589 23811 15592
rect 23753 15583 23811 15589
rect 24394 15580 24400 15592
rect 24452 15580 24458 15632
rect 17957 15555 18015 15561
rect 17957 15521 17969 15555
rect 18003 15521 18015 15555
rect 17957 15515 18015 15521
rect 19061 15555 19119 15561
rect 19061 15521 19073 15555
rect 19107 15552 19119 15555
rect 19242 15552 19248 15564
rect 19107 15524 19248 15552
rect 19107 15521 19119 15524
rect 19061 15515 19119 15521
rect 19242 15512 19248 15524
rect 19300 15512 19306 15564
rect 24578 15552 24584 15564
rect 24539 15524 24584 15552
rect 24578 15512 24584 15524
rect 24636 15552 24642 15564
rect 24854 15552 24860 15564
rect 24636 15524 24860 15552
rect 24636 15512 24642 15524
rect 24854 15512 24860 15524
rect 24912 15512 24918 15564
rect 11422 15484 11428 15496
rect 11256 15456 11428 15484
rect 9088 15444 9094 15456
rect 11422 15444 11428 15456
rect 11480 15444 11486 15496
rect 13814 15484 13820 15496
rect 13775 15456 13820 15484
rect 13814 15444 13820 15456
rect 13872 15444 13878 15496
rect 16482 15484 16488 15496
rect 16443 15456 16488 15484
rect 16482 15444 16488 15456
rect 16540 15444 16546 15496
rect 19426 15444 19432 15496
rect 19484 15484 19490 15496
rect 21174 15484 21180 15496
rect 19484 15456 21180 15484
rect 19484 15444 19490 15456
rect 21174 15444 21180 15456
rect 21232 15444 21238 15496
rect 21818 15484 21824 15496
rect 21779 15456 21824 15484
rect 21818 15444 21824 15456
rect 21876 15444 21882 15496
rect 1535 15419 1593 15425
rect 1535 15385 1547 15419
rect 1581 15416 1593 15419
rect 1946 15416 1952 15428
rect 1581 15388 1952 15416
rect 1581 15385 1593 15388
rect 1535 15379 1593 15385
rect 1946 15376 1952 15388
rect 2004 15376 2010 15428
rect 1670 15308 1676 15360
rect 1728 15348 1734 15360
rect 1857 15351 1915 15357
rect 1857 15348 1869 15351
rect 1728 15320 1869 15348
rect 1728 15308 1734 15320
rect 1857 15317 1869 15320
rect 1903 15317 1915 15351
rect 1857 15311 1915 15317
rect 13170 15308 13176 15360
rect 13228 15348 13234 15360
rect 14369 15351 14427 15357
rect 14369 15348 14381 15351
rect 13228 15320 14381 15348
rect 13228 15308 13234 15320
rect 14369 15317 14381 15320
rect 14415 15348 14427 15351
rect 15286 15348 15292 15360
rect 14415 15320 15292 15348
rect 14415 15317 14427 15320
rect 14369 15311 14427 15317
rect 15286 15308 15292 15320
rect 15344 15308 15350 15360
rect 18601 15351 18659 15357
rect 18601 15317 18613 15351
rect 18647 15348 18659 15351
rect 18690 15348 18696 15360
rect 18647 15320 18696 15348
rect 18647 15317 18659 15320
rect 18601 15311 18659 15317
rect 18690 15308 18696 15320
rect 18748 15348 18754 15360
rect 19978 15348 19984 15360
rect 18748 15320 19984 15348
rect 18748 15308 18754 15320
rect 19978 15308 19984 15320
rect 20036 15308 20042 15360
rect 21910 15308 21916 15360
rect 21968 15348 21974 15360
rect 22097 15351 22155 15357
rect 22097 15348 22109 15351
rect 21968 15320 22109 15348
rect 21968 15308 21974 15320
rect 22097 15317 22109 15320
rect 22143 15317 22155 15351
rect 22097 15311 22155 15317
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 1765 15147 1823 15153
rect 1765 15113 1777 15147
rect 1811 15144 1823 15147
rect 2498 15144 2504 15156
rect 1811 15116 2504 15144
rect 1811 15113 1823 15116
rect 1765 15107 1823 15113
rect 2498 15104 2504 15116
rect 2556 15104 2562 15156
rect 8481 15147 8539 15153
rect 8481 15113 8493 15147
rect 8527 15144 8539 15147
rect 8941 15147 8999 15153
rect 8941 15144 8953 15147
rect 8527 15116 8953 15144
rect 8527 15113 8539 15116
rect 8481 15107 8539 15113
rect 8941 15113 8953 15116
rect 8987 15144 8999 15147
rect 9030 15144 9036 15156
rect 8987 15116 9036 15144
rect 8987 15113 8999 15116
rect 8941 15107 8999 15113
rect 9030 15104 9036 15116
rect 9088 15104 9094 15156
rect 9766 15104 9772 15156
rect 9824 15144 9830 15156
rect 10045 15147 10103 15153
rect 10045 15144 10057 15147
rect 9824 15116 10057 15144
rect 9824 15104 9830 15116
rect 10045 15113 10057 15116
rect 10091 15113 10103 15147
rect 11698 15144 11704 15156
rect 11659 15116 11704 15144
rect 10045 15107 10103 15113
rect 11698 15104 11704 15116
rect 11756 15104 11762 15156
rect 14458 15144 14464 15156
rect 14419 15116 14464 15144
rect 14458 15104 14464 15116
rect 14516 15104 14522 15156
rect 15657 15147 15715 15153
rect 15657 15113 15669 15147
rect 15703 15144 15715 15147
rect 15746 15144 15752 15156
rect 15703 15116 15752 15144
rect 15703 15113 15715 15116
rect 15657 15107 15715 15113
rect 15746 15104 15752 15116
rect 15804 15104 15810 15156
rect 17494 15144 17500 15156
rect 17455 15116 17500 15144
rect 17494 15104 17500 15116
rect 17552 15104 17558 15156
rect 17954 15104 17960 15156
rect 18012 15144 18018 15156
rect 18233 15147 18291 15153
rect 18233 15144 18245 15147
rect 18012 15116 18245 15144
rect 18012 15104 18018 15116
rect 18233 15113 18245 15116
rect 18279 15113 18291 15147
rect 18233 15107 18291 15113
rect 18966 15104 18972 15156
rect 19024 15144 19030 15156
rect 19518 15144 19524 15156
rect 19024 15116 19524 15144
rect 19024 15104 19030 15116
rect 19518 15104 19524 15116
rect 19576 15144 19582 15156
rect 19889 15147 19947 15153
rect 19889 15144 19901 15147
rect 19576 15116 19901 15144
rect 19576 15104 19582 15116
rect 19889 15113 19901 15116
rect 19935 15113 19947 15147
rect 19889 15107 19947 15113
rect 20993 15147 21051 15153
rect 20993 15113 21005 15147
rect 21039 15144 21051 15147
rect 21266 15144 21272 15156
rect 21039 15116 21272 15144
rect 21039 15113 21051 15116
rect 20993 15107 21051 15113
rect 4798 15036 4804 15088
rect 4856 15076 4862 15088
rect 8018 15076 8024 15088
rect 4856 15048 8024 15076
rect 4856 15036 4862 15048
rect 8018 15036 8024 15048
rect 8076 15076 8082 15088
rect 8294 15076 8300 15088
rect 8076 15048 8300 15076
rect 8076 15036 8082 15048
rect 8294 15036 8300 15048
rect 8352 15036 8358 15088
rect 9677 15079 9735 15085
rect 9677 15045 9689 15079
rect 9723 15045 9735 15079
rect 9677 15039 9735 15045
rect 2314 15008 2320 15020
rect 2275 14980 2320 15008
rect 2314 14968 2320 14980
rect 2372 14968 2378 15020
rect 2961 15011 3019 15017
rect 2961 14977 2973 15011
rect 3007 15008 3019 15011
rect 3234 15008 3240 15020
rect 3007 14980 3240 15008
rect 3007 14977 3019 14980
rect 2961 14971 3019 14977
rect 3234 14968 3240 14980
rect 3292 15008 3298 15020
rect 3878 15008 3884 15020
rect 3292 14980 3884 15008
rect 3292 14968 3298 14980
rect 3878 14968 3884 14980
rect 3936 14968 3942 15020
rect 4154 15008 4160 15020
rect 4115 14980 4160 15008
rect 4154 14968 4160 14980
rect 4212 14968 4218 15020
rect 6914 15008 6920 15020
rect 6875 14980 6920 15008
rect 6914 14968 6920 14980
rect 6972 14968 6978 15020
rect 9122 15008 9128 15020
rect 9083 14980 9128 15008
rect 9122 14968 9128 14980
rect 9180 14968 9186 15020
rect 9692 15008 9720 15039
rect 11054 15036 11060 15088
rect 11112 15076 11118 15088
rect 11112 15048 11192 15076
rect 11112 15036 11118 15048
rect 11164 15017 11192 15048
rect 13262 15036 13268 15088
rect 13320 15076 13326 15088
rect 14642 15076 14648 15088
rect 13320 15048 14648 15076
rect 13320 15036 13326 15048
rect 14642 15036 14648 15048
rect 14700 15076 14706 15088
rect 15013 15079 15071 15085
rect 15013 15076 15025 15079
rect 14700 15048 15025 15076
rect 14700 15036 14706 15048
rect 15013 15045 15025 15048
rect 15059 15045 15071 15079
rect 15013 15039 15071 15045
rect 11149 15011 11207 15017
rect 9692 14980 9904 15008
rect 4522 14900 4528 14952
rect 4580 14940 4586 14952
rect 5420 14943 5478 14949
rect 5420 14940 5432 14943
rect 4580 14912 5432 14940
rect 4580 14900 4586 14912
rect 5420 14909 5432 14912
rect 5466 14940 5478 14943
rect 5466 14912 5948 14940
rect 5466 14909 5478 14912
rect 5420 14903 5478 14909
rect 2409 14875 2467 14881
rect 2409 14841 2421 14875
rect 2455 14872 2467 14875
rect 2682 14872 2688 14884
rect 2455 14844 2688 14872
rect 2455 14841 2467 14844
rect 2409 14835 2467 14841
rect 2133 14807 2191 14813
rect 2133 14773 2145 14807
rect 2179 14804 2191 14807
rect 2424 14804 2452 14835
rect 2682 14832 2688 14844
rect 2740 14832 2746 14884
rect 3697 14875 3755 14881
rect 3697 14841 3709 14875
rect 3743 14872 3755 14875
rect 3970 14872 3976 14884
rect 3743 14844 3976 14872
rect 3743 14841 3755 14844
rect 3697 14835 3755 14841
rect 3970 14832 3976 14844
rect 4028 14832 4034 14884
rect 5920 14881 5948 14912
rect 5905 14875 5963 14881
rect 5905 14841 5917 14875
rect 5951 14872 5963 14875
rect 7006 14872 7012 14884
rect 5951 14844 6684 14872
rect 6967 14844 7012 14872
rect 5951 14841 5963 14844
rect 5905 14835 5963 14841
rect 3234 14804 3240 14816
rect 2179 14776 2452 14804
rect 3195 14776 3240 14804
rect 2179 14773 2191 14776
rect 2133 14767 2191 14773
rect 3234 14764 3240 14776
rect 3292 14764 3298 14816
rect 4798 14804 4804 14816
rect 4759 14776 4804 14804
rect 4798 14764 4804 14776
rect 4856 14764 4862 14816
rect 5166 14804 5172 14816
rect 5127 14776 5172 14804
rect 5166 14764 5172 14776
rect 5224 14764 5230 14816
rect 5258 14764 5264 14816
rect 5316 14804 5322 14816
rect 5491 14807 5549 14813
rect 5491 14804 5503 14807
rect 5316 14776 5503 14804
rect 5316 14764 5322 14776
rect 5491 14773 5503 14776
rect 5537 14773 5549 14807
rect 6546 14804 6552 14816
rect 6507 14776 6552 14804
rect 5491 14767 5549 14773
rect 6546 14764 6552 14776
rect 6604 14764 6610 14816
rect 6656 14804 6684 14844
rect 7006 14832 7012 14844
rect 7064 14832 7070 14884
rect 7561 14875 7619 14881
rect 7561 14841 7573 14875
rect 7607 14872 7619 14875
rect 7650 14872 7656 14884
rect 7607 14844 7656 14872
rect 7607 14841 7619 14844
rect 7561 14835 7619 14841
rect 7650 14832 7656 14844
rect 7708 14872 7714 14884
rect 7708 14844 8248 14872
rect 7708 14832 7714 14844
rect 7190 14804 7196 14816
rect 6656 14776 7196 14804
rect 7190 14764 7196 14776
rect 7248 14764 7254 14816
rect 8220 14804 8248 14844
rect 9122 14832 9128 14884
rect 9180 14872 9186 14884
rect 9217 14875 9275 14881
rect 9217 14872 9229 14875
rect 9180 14844 9229 14872
rect 9180 14832 9186 14844
rect 9217 14841 9229 14844
rect 9263 14841 9275 14875
rect 9217 14835 9275 14841
rect 9766 14804 9772 14816
rect 8220 14776 9772 14804
rect 9766 14764 9772 14776
rect 9824 14804 9830 14816
rect 9876 14804 9904 14980
rect 11149 14977 11161 15011
rect 11195 14977 11207 15011
rect 11149 14971 11207 14977
rect 12176 14980 12618 15008
rect 10505 14943 10563 14949
rect 10505 14909 10517 14943
rect 10551 14940 10563 14943
rect 10778 14940 10784 14952
rect 10551 14912 10784 14940
rect 10551 14909 10563 14912
rect 10505 14903 10563 14909
rect 10778 14900 10784 14912
rect 10836 14900 10842 14952
rect 11057 14943 11115 14949
rect 11057 14909 11069 14943
rect 11103 14940 11115 14943
rect 11698 14940 11704 14952
rect 11103 14912 11704 14940
rect 11103 14909 11115 14912
rect 11057 14903 11115 14909
rect 11698 14900 11704 14912
rect 11756 14900 11762 14952
rect 9824 14776 9904 14804
rect 9824 14764 9830 14776
rect 11698 14764 11704 14816
rect 11756 14804 11762 14816
rect 12176 14813 12204 14980
rect 12590 14940 12618 14980
rect 12802 14968 12808 15020
rect 12860 15008 12866 15020
rect 13170 15008 13176 15020
rect 12860 14980 13176 15008
rect 12860 14968 12866 14980
rect 13170 14968 13176 14980
rect 13228 14968 13234 15020
rect 15764 15008 15792 15104
rect 19153 15079 19211 15085
rect 19153 15045 19165 15079
rect 19199 15076 19211 15079
rect 19426 15076 19432 15088
rect 19199 15048 19432 15076
rect 19199 15045 19211 15048
rect 19153 15039 19211 15045
rect 19426 15036 19432 15048
rect 19484 15036 19490 15088
rect 18598 15008 18604 15020
rect 15764 14980 16896 15008
rect 18559 14980 18604 15008
rect 12713 14943 12771 14949
rect 12713 14940 12725 14943
rect 12590 14912 12725 14940
rect 12713 14909 12725 14912
rect 12759 14909 12771 14943
rect 14093 14943 14151 14949
rect 14093 14940 14105 14943
rect 12713 14903 12771 14909
rect 13924 14912 14105 14940
rect 13924 14816 13952 14912
rect 14093 14909 14105 14912
rect 14139 14909 14151 14943
rect 16022 14940 16028 14952
rect 15935 14912 16028 14940
rect 14093 14903 14151 14909
rect 16022 14900 16028 14912
rect 16080 14940 16086 14952
rect 16666 14940 16672 14952
rect 16080 14912 16672 14940
rect 16080 14900 16086 14912
rect 16666 14900 16672 14912
rect 16724 14900 16730 14952
rect 16868 14949 16896 14980
rect 18598 14968 18604 14980
rect 18656 14968 18662 15020
rect 16853 14943 16911 14949
rect 16853 14909 16865 14943
rect 16899 14909 16911 14943
rect 16853 14903 16911 14909
rect 17126 14872 17132 14884
rect 17087 14844 17132 14872
rect 17126 14832 17132 14844
rect 17184 14832 17190 14884
rect 18690 14832 18696 14884
rect 18748 14872 18754 14884
rect 19904 14872 19932 15107
rect 21266 15104 21272 15116
rect 21324 15104 21330 15156
rect 23106 15144 23112 15156
rect 23067 15116 23112 15144
rect 23106 15104 23112 15116
rect 23164 15104 23170 15156
rect 23474 15144 23480 15156
rect 23435 15116 23480 15144
rect 23474 15104 23480 15116
rect 23532 15104 23538 15156
rect 24854 15104 24860 15156
rect 24912 15144 24918 15156
rect 24949 15147 25007 15153
rect 24949 15144 24961 15147
rect 24912 15116 24961 15144
rect 24912 15104 24918 15116
rect 24949 15113 24961 15116
rect 24995 15113 25007 15147
rect 24949 15107 25007 15113
rect 20070 15008 20076 15020
rect 20031 14980 20076 15008
rect 20070 14968 20076 14980
rect 20128 14968 20134 15020
rect 24029 15011 24087 15017
rect 24029 14977 24041 15011
rect 24075 15008 24087 15011
rect 24118 15008 24124 15020
rect 24075 14980 24124 15008
rect 24075 14977 24087 14980
rect 24029 14971 24087 14977
rect 24118 14968 24124 14980
rect 24176 14968 24182 15020
rect 21818 14940 21824 14952
rect 21779 14912 21824 14940
rect 21818 14900 21824 14912
rect 21876 14900 21882 14952
rect 24946 14900 24952 14952
rect 25004 14940 25010 14952
rect 25501 14943 25559 14949
rect 25501 14940 25513 14943
rect 25004 14912 25513 14940
rect 25004 14900 25010 14912
rect 25501 14909 25513 14912
rect 25547 14940 25559 14943
rect 26053 14943 26111 14949
rect 26053 14940 26065 14943
rect 25547 14912 26065 14940
rect 25547 14909 25559 14912
rect 25501 14903 25559 14909
rect 26053 14909 26065 14912
rect 26099 14909 26111 14943
rect 26053 14903 26111 14909
rect 20394 14875 20452 14881
rect 20394 14872 20406 14875
rect 18748 14844 18793 14872
rect 19904 14844 20406 14872
rect 18748 14832 18754 14844
rect 20394 14841 20406 14844
rect 20440 14841 20452 14875
rect 22142 14875 22200 14881
rect 22142 14872 22154 14875
rect 20394 14835 20452 14841
rect 21744 14844 22154 14872
rect 21744 14816 21772 14844
rect 22142 14841 22154 14844
rect 22188 14841 22200 14875
rect 22142 14835 22200 14841
rect 23474 14832 23480 14884
rect 23532 14872 23538 14884
rect 24121 14875 24179 14881
rect 24121 14872 24133 14875
rect 23532 14844 24133 14872
rect 23532 14832 23538 14844
rect 24121 14841 24133 14844
rect 24167 14841 24179 14875
rect 24670 14872 24676 14884
rect 24631 14844 24676 14872
rect 24121 14835 24179 14841
rect 24670 14832 24676 14844
rect 24728 14832 24734 14884
rect 12161 14807 12219 14813
rect 12161 14804 12173 14807
rect 11756 14776 12173 14804
rect 11756 14764 11762 14776
rect 12161 14773 12173 14776
rect 12207 14773 12219 14807
rect 13538 14804 13544 14816
rect 13451 14776 13544 14804
rect 12161 14767 12219 14773
rect 13538 14764 13544 14776
rect 13596 14804 13602 14816
rect 13906 14804 13912 14816
rect 13596 14776 13912 14804
rect 13596 14764 13602 14776
rect 13906 14764 13912 14776
rect 13964 14764 13970 14816
rect 21726 14804 21732 14816
rect 21687 14776 21732 14804
rect 21726 14764 21732 14776
rect 21784 14764 21790 14816
rect 22738 14804 22744 14816
rect 22699 14776 22744 14804
rect 22738 14764 22744 14776
rect 22796 14764 22802 14816
rect 25682 14804 25688 14816
rect 25643 14776 25688 14804
rect 25682 14764 25688 14776
rect 25740 14764 25746 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1854 14600 1860 14612
rect 1815 14572 1860 14600
rect 1854 14560 1860 14572
rect 1912 14560 1918 14612
rect 2130 14560 2136 14612
rect 2188 14560 2194 14612
rect 2314 14600 2320 14612
rect 2275 14572 2320 14600
rect 2314 14560 2320 14572
rect 2372 14560 2378 14612
rect 3878 14600 3884 14612
rect 3839 14572 3884 14600
rect 3878 14560 3884 14572
rect 3936 14560 3942 14612
rect 3970 14560 3976 14612
rect 4028 14600 4034 14612
rect 5353 14603 5411 14609
rect 5353 14600 5365 14603
rect 4028 14572 5365 14600
rect 4028 14560 4034 14572
rect 5353 14569 5365 14572
rect 5399 14569 5411 14603
rect 5353 14563 5411 14569
rect 7006 14560 7012 14612
rect 7064 14600 7070 14612
rect 7469 14603 7527 14609
rect 7469 14600 7481 14603
rect 7064 14572 7481 14600
rect 7064 14560 7070 14572
rect 7469 14569 7481 14572
rect 7515 14600 7527 14603
rect 7742 14600 7748 14612
rect 7515 14572 7748 14600
rect 7515 14569 7527 14572
rect 7469 14563 7527 14569
rect 7742 14560 7748 14572
rect 7800 14560 7806 14612
rect 9030 14600 9036 14612
rect 8991 14572 9036 14600
rect 9030 14560 9036 14572
rect 9088 14600 9094 14612
rect 10597 14603 10655 14609
rect 10597 14600 10609 14603
rect 9088 14572 10609 14600
rect 9088 14560 9094 14572
rect 10597 14569 10609 14572
rect 10643 14569 10655 14603
rect 10597 14563 10655 14569
rect 11333 14603 11391 14609
rect 11333 14569 11345 14603
rect 11379 14600 11391 14603
rect 11422 14600 11428 14612
rect 11379 14572 11428 14600
rect 11379 14569 11391 14572
rect 11333 14563 11391 14569
rect 11422 14560 11428 14572
rect 11480 14560 11486 14612
rect 12526 14600 12532 14612
rect 12487 14572 12532 14600
rect 12526 14560 12532 14572
rect 12584 14560 12590 14612
rect 13354 14600 13360 14612
rect 13315 14572 13360 14600
rect 13354 14560 13360 14572
rect 13412 14560 13418 14612
rect 14458 14560 14464 14612
rect 14516 14600 14522 14612
rect 15013 14603 15071 14609
rect 15013 14600 15025 14603
rect 14516 14572 15025 14600
rect 14516 14560 14522 14572
rect 15013 14569 15025 14572
rect 15059 14569 15071 14603
rect 15013 14563 15071 14569
rect 18509 14603 18567 14609
rect 18509 14569 18521 14603
rect 18555 14600 18567 14603
rect 18598 14600 18604 14612
rect 18555 14572 18604 14600
rect 18555 14569 18567 14572
rect 18509 14563 18567 14569
rect 18598 14560 18604 14572
rect 18656 14560 18662 14612
rect 19334 14560 19340 14612
rect 19392 14600 19398 14612
rect 19797 14603 19855 14609
rect 19797 14600 19809 14603
rect 19392 14572 19809 14600
rect 19392 14560 19398 14572
rect 19797 14569 19809 14572
rect 19843 14569 19855 14603
rect 19797 14563 19855 14569
rect 20070 14560 20076 14612
rect 20128 14600 20134 14612
rect 20165 14603 20223 14609
rect 20165 14600 20177 14603
rect 20128 14572 20177 14600
rect 20128 14560 20134 14572
rect 20165 14569 20177 14572
rect 20211 14569 20223 14603
rect 21174 14600 21180 14612
rect 21135 14572 21180 14600
rect 20165 14563 20223 14569
rect 21174 14560 21180 14572
rect 21232 14560 21238 14612
rect 22373 14603 22431 14609
rect 22373 14569 22385 14603
rect 22419 14600 22431 14603
rect 23198 14600 23204 14612
rect 22419 14572 23204 14600
rect 22419 14569 22431 14572
rect 22373 14563 22431 14569
rect 23198 14560 23204 14572
rect 23256 14600 23262 14612
rect 23256 14572 23428 14600
rect 23256 14560 23262 14572
rect 2148 14532 2176 14560
rect 2593 14535 2651 14541
rect 2148 14504 2360 14532
rect 2332 14476 2360 14504
rect 2593 14501 2605 14535
rect 2639 14532 2651 14535
rect 2682 14532 2688 14544
rect 2639 14504 2688 14532
rect 2639 14501 2651 14504
rect 2593 14495 2651 14501
rect 2682 14492 2688 14504
rect 2740 14492 2746 14544
rect 4774 14535 4832 14541
rect 4774 14501 4786 14535
rect 4820 14532 4832 14535
rect 4890 14532 4896 14544
rect 4820 14504 4896 14532
rect 4820 14501 4832 14504
rect 4774 14495 4832 14501
rect 4890 14492 4896 14504
rect 4948 14532 4954 14544
rect 6638 14541 6644 14544
rect 6635 14532 6644 14541
rect 4948 14504 6644 14532
rect 4948 14492 4954 14504
rect 6635 14495 6644 14504
rect 6638 14492 6644 14495
rect 6696 14492 6702 14544
rect 10042 14541 10048 14544
rect 10039 14532 10048 14541
rect 10003 14504 10048 14532
rect 10039 14495 10048 14504
rect 10042 14492 10048 14495
rect 10100 14492 10106 14544
rect 11977 14535 12035 14541
rect 11977 14501 11989 14535
rect 12023 14532 12035 14535
rect 12802 14532 12808 14544
rect 12023 14504 12808 14532
rect 12023 14501 12035 14504
rect 11977 14495 12035 14501
rect 1448 14467 1506 14473
rect 1448 14433 1460 14467
rect 1494 14464 1506 14467
rect 2130 14464 2136 14476
rect 1494 14436 2136 14464
rect 1494 14433 1506 14436
rect 1448 14427 1506 14433
rect 2130 14424 2136 14436
rect 2188 14424 2194 14476
rect 2314 14424 2320 14476
rect 2372 14424 2378 14476
rect 4430 14464 4436 14476
rect 4391 14436 4436 14464
rect 4430 14424 4436 14436
rect 4488 14424 4494 14476
rect 6270 14464 6276 14476
rect 6231 14436 6276 14464
rect 6270 14424 6276 14436
rect 6328 14424 6334 14476
rect 8202 14464 8208 14476
rect 8163 14436 8208 14464
rect 8202 14424 8208 14436
rect 8260 14424 8266 14476
rect 8478 14464 8484 14476
rect 8439 14436 8484 14464
rect 8478 14424 8484 14436
rect 8536 14424 8542 14476
rect 8662 14424 8668 14476
rect 8720 14464 8726 14476
rect 12084 14473 12112 14504
rect 12802 14492 12808 14504
rect 12860 14492 12866 14544
rect 14366 14532 14372 14544
rect 14327 14504 14372 14532
rect 14366 14492 14372 14504
rect 14424 14492 14430 14544
rect 14642 14532 14648 14544
rect 14603 14504 14648 14532
rect 14642 14492 14648 14504
rect 14700 14492 14706 14544
rect 15930 14532 15936 14544
rect 15672 14504 15936 14532
rect 9677 14467 9735 14473
rect 9677 14464 9689 14467
rect 8720 14436 9689 14464
rect 8720 14424 8726 14436
rect 9677 14433 9689 14436
rect 9723 14433 9735 14467
rect 9677 14427 9735 14433
rect 12069 14467 12127 14473
rect 12069 14433 12081 14467
rect 12115 14433 12127 14467
rect 12342 14464 12348 14476
rect 12303 14436 12348 14464
rect 12069 14427 12127 14433
rect 12342 14424 12348 14436
rect 12400 14424 12406 14476
rect 13262 14424 13268 14476
rect 13320 14464 13326 14476
rect 13633 14467 13691 14473
rect 13633 14464 13645 14467
rect 13320 14436 13645 14464
rect 13320 14424 13326 14436
rect 13633 14433 13645 14436
rect 13679 14433 13691 14467
rect 13906 14464 13912 14476
rect 13867 14436 13912 14464
rect 13633 14427 13691 14433
rect 13906 14424 13912 14436
rect 13964 14424 13970 14476
rect 15672 14473 15700 14504
rect 15930 14492 15936 14504
rect 15988 14492 15994 14544
rect 18966 14541 18972 14544
rect 16209 14535 16267 14541
rect 16209 14501 16221 14535
rect 16255 14532 16267 14535
rect 18963 14532 18972 14541
rect 16255 14504 18644 14532
rect 18927 14504 18972 14532
rect 16255 14501 16267 14504
rect 16209 14495 16267 14501
rect 15657 14467 15715 14473
rect 15657 14433 15669 14467
rect 15703 14433 15715 14467
rect 15657 14427 15715 14433
rect 15838 14424 15844 14476
rect 15896 14464 15902 14476
rect 16025 14467 16083 14473
rect 16025 14464 16037 14467
rect 15896 14436 16037 14464
rect 15896 14424 15902 14436
rect 16025 14433 16037 14436
rect 16071 14464 16083 14467
rect 16482 14464 16488 14476
rect 16071 14436 16488 14464
rect 16071 14433 16083 14436
rect 16025 14427 16083 14433
rect 16482 14424 16488 14436
rect 16540 14424 16546 14476
rect 17313 14467 17371 14473
rect 17313 14433 17325 14467
rect 17359 14464 17371 14467
rect 17402 14464 17408 14476
rect 17359 14436 17408 14464
rect 17359 14433 17371 14436
rect 17313 14427 17371 14433
rect 17402 14424 17408 14436
rect 17460 14424 17466 14476
rect 17586 14464 17592 14476
rect 17547 14436 17592 14464
rect 17586 14424 17592 14436
rect 17644 14424 17650 14476
rect 18616 14473 18644 14504
rect 18963 14495 18972 14504
rect 18966 14492 18972 14495
rect 19024 14492 19030 14544
rect 21726 14492 21732 14544
rect 21784 14541 21790 14544
rect 23400 14541 23428 14572
rect 21784 14535 21832 14541
rect 21784 14501 21786 14535
rect 21820 14501 21832 14535
rect 21784 14495 21832 14501
rect 23385 14535 23443 14541
rect 23385 14501 23397 14535
rect 23431 14501 23443 14535
rect 23385 14495 23443 14501
rect 21784 14492 21790 14495
rect 24670 14492 24676 14544
rect 24728 14532 24734 14544
rect 24857 14535 24915 14541
rect 24857 14532 24869 14535
rect 24728 14504 24869 14532
rect 24728 14492 24734 14504
rect 24857 14501 24869 14504
rect 24903 14501 24915 14535
rect 24857 14495 24915 14501
rect 24946 14492 24952 14544
rect 25004 14532 25010 14544
rect 25004 14504 25049 14532
rect 25004 14492 25010 14504
rect 18601 14467 18659 14473
rect 18601 14433 18613 14467
rect 18647 14464 18659 14467
rect 20162 14464 20168 14476
rect 18647 14436 20168 14464
rect 18647 14433 18659 14436
rect 18601 14427 18659 14433
rect 20162 14424 20168 14436
rect 20220 14424 20226 14476
rect 2501 14399 2559 14405
rect 2501 14365 2513 14399
rect 2547 14396 2559 14399
rect 2590 14396 2596 14408
rect 2547 14368 2596 14396
rect 2547 14365 2559 14368
rect 2501 14359 2559 14365
rect 2590 14356 2596 14368
rect 2648 14356 2654 14408
rect 2866 14356 2872 14408
rect 2924 14396 2930 14408
rect 3145 14399 3203 14405
rect 3145 14396 3157 14399
rect 2924 14368 3157 14396
rect 2924 14356 2930 14368
rect 3145 14365 3157 14368
rect 3191 14396 3203 14399
rect 3421 14399 3479 14405
rect 3421 14396 3433 14399
rect 3191 14368 3433 14396
rect 3191 14365 3203 14368
rect 3145 14359 3203 14365
rect 3421 14365 3433 14368
rect 3467 14365 3479 14399
rect 8754 14396 8760 14408
rect 8715 14368 8760 14396
rect 3421 14359 3479 14365
rect 8754 14356 8760 14368
rect 8812 14356 8818 14408
rect 13280 14396 13308 14424
rect 11992 14368 13308 14396
rect 16577 14399 16635 14405
rect 11992 14340 12020 14368
rect 16577 14365 16589 14399
rect 16623 14396 16635 14399
rect 16666 14396 16672 14408
rect 16623 14368 16672 14396
rect 16623 14365 16635 14368
rect 16577 14359 16635 14365
rect 16666 14356 16672 14368
rect 16724 14396 16730 14408
rect 17604 14396 17632 14424
rect 17770 14396 17776 14408
rect 16724 14368 17632 14396
rect 17731 14368 17776 14396
rect 16724 14356 16730 14368
rect 17770 14356 17776 14368
rect 17828 14356 17834 14408
rect 21450 14396 21456 14408
rect 21411 14368 21456 14396
rect 21450 14356 21456 14368
rect 21508 14356 21514 14408
rect 23293 14399 23351 14405
rect 23293 14365 23305 14399
rect 23339 14396 23351 14399
rect 23382 14396 23388 14408
rect 23339 14368 23388 14396
rect 23339 14365 23351 14368
rect 23293 14359 23351 14365
rect 23382 14356 23388 14368
rect 23440 14356 23446 14408
rect 23658 14396 23664 14408
rect 23619 14368 23664 14396
rect 23658 14356 23664 14368
rect 23716 14396 23722 14408
rect 25133 14399 25191 14405
rect 25133 14396 25145 14399
rect 23716 14368 25145 14396
rect 23716 14356 23722 14368
rect 25133 14365 25145 14368
rect 25179 14396 25191 14399
rect 25590 14396 25596 14408
rect 25179 14368 25596 14396
rect 25179 14365 25191 14368
rect 25133 14359 25191 14365
rect 25590 14356 25596 14368
rect 25648 14356 25654 14408
rect 1854 14288 1860 14340
rect 1912 14328 1918 14340
rect 4154 14328 4160 14340
rect 1912 14300 4160 14328
rect 1912 14288 1918 14300
rect 4154 14288 4160 14300
rect 4212 14288 4218 14340
rect 11974 14288 11980 14340
rect 12032 14288 12038 14340
rect 12158 14328 12164 14340
rect 12119 14300 12164 14328
rect 12158 14288 12164 14300
rect 12216 14328 12222 14340
rect 13725 14331 13783 14337
rect 13725 14328 13737 14331
rect 12216 14300 13737 14328
rect 12216 14288 12222 14300
rect 13725 14297 13737 14300
rect 13771 14328 13783 14331
rect 13998 14328 14004 14340
rect 13771 14300 14004 14328
rect 13771 14297 13783 14300
rect 13725 14291 13783 14297
rect 13998 14288 14004 14300
rect 14056 14288 14062 14340
rect 16758 14288 16764 14340
rect 16816 14328 16822 14340
rect 16853 14331 16911 14337
rect 16853 14328 16865 14331
rect 16816 14300 16865 14328
rect 16816 14288 16822 14300
rect 16853 14297 16865 14300
rect 16899 14297 16911 14331
rect 16853 14291 16911 14297
rect 1535 14263 1593 14269
rect 1535 14229 1547 14263
rect 1581 14260 1593 14263
rect 1762 14260 1768 14272
rect 1581 14232 1768 14260
rect 1581 14229 1593 14232
rect 1535 14223 1593 14229
rect 1762 14220 1768 14232
rect 1820 14220 1826 14272
rect 4338 14260 4344 14272
rect 4299 14232 4344 14260
rect 4338 14220 4344 14232
rect 4396 14220 4402 14272
rect 5074 14220 5080 14272
rect 5132 14260 5138 14272
rect 5350 14260 5356 14272
rect 5132 14232 5356 14260
rect 5132 14220 5138 14232
rect 5350 14220 5356 14232
rect 5408 14220 5414 14272
rect 7190 14260 7196 14272
rect 7151 14232 7196 14260
rect 7190 14220 7196 14232
rect 7248 14220 7254 14272
rect 19518 14260 19524 14272
rect 19479 14232 19524 14260
rect 19518 14220 19524 14232
rect 19576 14220 19582 14272
rect 23106 14260 23112 14272
rect 23067 14232 23112 14260
rect 23106 14220 23112 14232
rect 23164 14220 23170 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 1578 14056 1584 14068
rect 1539 14028 1584 14056
rect 1578 14016 1584 14028
rect 1636 14016 1642 14068
rect 2501 14059 2559 14065
rect 2501 14025 2513 14059
rect 2547 14056 2559 14059
rect 2590 14056 2596 14068
rect 2547 14028 2596 14056
rect 2547 14025 2559 14028
rect 2501 14019 2559 14025
rect 2590 14016 2596 14028
rect 2648 14016 2654 14068
rect 3881 14059 3939 14065
rect 3881 14025 3893 14059
rect 3927 14056 3939 14059
rect 4430 14056 4436 14068
rect 3927 14028 4436 14056
rect 3927 14025 3939 14028
rect 3881 14019 3939 14025
rect 4430 14016 4436 14028
rect 4488 14016 4494 14068
rect 5905 14059 5963 14065
rect 5905 14025 5917 14059
rect 5951 14056 5963 14059
rect 6270 14056 6276 14068
rect 5951 14028 6276 14056
rect 5951 14025 5963 14028
rect 5905 14019 5963 14025
rect 6270 14016 6276 14028
rect 6328 14016 6334 14068
rect 6638 14056 6644 14068
rect 6599 14028 6644 14056
rect 6638 14016 6644 14028
rect 6696 14016 6702 14068
rect 7742 14056 7748 14068
rect 7703 14028 7748 14056
rect 7742 14016 7748 14028
rect 7800 14016 7806 14068
rect 8113 14059 8171 14065
rect 8113 14025 8125 14059
rect 8159 14056 8171 14059
rect 8202 14056 8208 14068
rect 8159 14028 8208 14056
rect 8159 14025 8171 14028
rect 8113 14019 8171 14025
rect 8202 14016 8208 14028
rect 8260 14016 8266 14068
rect 8662 14016 8668 14068
rect 8720 14056 8726 14068
rect 8757 14059 8815 14065
rect 8757 14056 8769 14059
rect 8720 14028 8769 14056
rect 8720 14016 8726 14028
rect 8757 14025 8769 14028
rect 8803 14025 8815 14059
rect 13998 14056 14004 14068
rect 13959 14028 14004 14056
rect 8757 14019 8815 14025
rect 13998 14016 14004 14028
rect 14056 14056 14062 14068
rect 15286 14056 15292 14068
rect 14056 14028 14412 14056
rect 15247 14028 15292 14056
rect 14056 14016 14062 14028
rect 1394 13948 1400 14000
rect 1452 13988 1458 14000
rect 2041 13991 2099 13997
rect 2041 13988 2053 13991
rect 1452 13960 2053 13988
rect 1452 13948 1458 13960
rect 2041 13957 2053 13960
rect 2087 13988 2099 13991
rect 2130 13988 2136 14000
rect 2087 13960 2136 13988
rect 2087 13957 2099 13960
rect 2041 13951 2099 13957
rect 2130 13948 2136 13960
rect 2188 13948 2194 14000
rect 3510 13948 3516 14000
rect 3568 13988 3574 14000
rect 5261 13991 5319 13997
rect 5261 13988 5273 13991
rect 3568 13960 5273 13988
rect 3568 13948 3574 13960
rect 5261 13957 5273 13960
rect 5307 13957 5319 13991
rect 5261 13951 5319 13957
rect 6181 13991 6239 13997
rect 6181 13957 6193 13991
rect 6227 13988 6239 13991
rect 6656 13988 6684 14016
rect 9125 13991 9183 13997
rect 9125 13988 9137 13991
rect 6227 13960 9137 13988
rect 6227 13957 6239 13960
rect 6181 13951 6239 13957
rect 2866 13920 2872 13932
rect 2827 13892 2872 13920
rect 2866 13880 2872 13892
rect 2924 13880 2930 13932
rect 5534 13880 5540 13932
rect 5592 13920 5598 13932
rect 6730 13920 6736 13932
rect 5592 13892 6736 13920
rect 5592 13880 5598 13892
rect 6730 13880 6736 13892
rect 6788 13920 6794 13932
rect 6825 13923 6883 13929
rect 6825 13920 6837 13923
rect 6788 13892 6837 13920
rect 6788 13880 6794 13892
rect 6825 13889 6837 13892
rect 6871 13889 6883 13923
rect 6825 13883 6883 13889
rect 1397 13855 1455 13861
rect 1397 13821 1409 13855
rect 1443 13852 1455 13855
rect 3513 13855 3571 13861
rect 1443 13824 1716 13852
rect 1443 13821 1455 13824
rect 1397 13815 1455 13821
rect 1578 13676 1584 13728
rect 1636 13716 1642 13728
rect 1688 13716 1716 13824
rect 3513 13821 3525 13855
rect 3559 13852 3571 13855
rect 4154 13852 4160 13864
rect 3559 13824 4160 13852
rect 3559 13821 3571 13824
rect 3513 13815 3571 13821
rect 4154 13812 4160 13824
rect 4212 13812 4218 13864
rect 4338 13852 4344 13864
rect 4299 13824 4344 13852
rect 4338 13812 4344 13824
rect 4396 13812 4402 13864
rect 2961 13787 3019 13793
rect 2961 13753 2973 13787
rect 3007 13784 3019 13787
rect 3326 13784 3332 13796
rect 3007 13756 3332 13784
rect 3007 13753 3019 13756
rect 2961 13747 3019 13753
rect 3326 13744 3332 13756
rect 3384 13744 3390 13796
rect 4249 13787 4307 13793
rect 4249 13753 4261 13787
rect 4295 13784 4307 13787
rect 4430 13784 4436 13796
rect 4295 13756 4436 13784
rect 4295 13753 4307 13756
rect 4249 13747 4307 13753
rect 4430 13744 4436 13756
rect 4488 13784 4494 13796
rect 4703 13787 4761 13793
rect 4703 13784 4715 13787
rect 4488 13756 4715 13784
rect 4488 13744 4494 13756
rect 4703 13753 4715 13756
rect 4749 13784 4761 13787
rect 4890 13784 4896 13796
rect 4749 13756 4896 13784
rect 4749 13753 4761 13756
rect 4703 13747 4761 13753
rect 4890 13744 4896 13756
rect 4948 13744 4954 13796
rect 7161 13793 7189 13960
rect 9125 13957 9137 13960
rect 9171 13988 9183 13991
rect 11514 13988 11520 14000
rect 9171 13960 9628 13988
rect 11475 13960 11520 13988
rect 9171 13957 9183 13960
rect 9125 13951 9183 13957
rect 8754 13880 8760 13932
rect 8812 13920 8818 13932
rect 9306 13920 9312 13932
rect 8812 13892 9312 13920
rect 8812 13880 8818 13892
rect 9306 13880 9312 13892
rect 9364 13880 9370 13932
rect 8478 13852 8484 13864
rect 8439 13824 8484 13852
rect 8478 13812 8484 13824
rect 8536 13812 8542 13864
rect 9600 13852 9628 13960
rect 11514 13948 11520 13960
rect 11572 13948 11578 14000
rect 12713 13991 12771 13997
rect 12713 13957 12725 13991
rect 12759 13988 12771 13991
rect 13354 13988 13360 14000
rect 12759 13960 13360 13988
rect 12759 13957 12771 13960
rect 12713 13951 12771 13957
rect 13354 13948 13360 13960
rect 13412 13948 13418 14000
rect 14384 13997 14412 14028
rect 15286 14016 15292 14028
rect 15344 14016 15350 14068
rect 16114 14056 16120 14068
rect 16075 14028 16120 14056
rect 16114 14016 16120 14028
rect 16172 14016 16178 14068
rect 18693 14059 18751 14065
rect 18693 14025 18705 14059
rect 18739 14056 18751 14059
rect 18966 14056 18972 14068
rect 18739 14028 18972 14056
rect 18739 14025 18751 14028
rect 18693 14019 18751 14025
rect 18966 14016 18972 14028
rect 19024 14016 19030 14068
rect 19518 14016 19524 14068
rect 19576 14056 19582 14068
rect 20533 14059 20591 14065
rect 20533 14056 20545 14059
rect 19576 14028 20545 14056
rect 19576 14016 19582 14028
rect 20533 14025 20545 14028
rect 20579 14056 20591 14059
rect 20898 14056 20904 14068
rect 20579 14028 20904 14056
rect 20579 14025 20591 14028
rect 20533 14019 20591 14025
rect 20898 14016 20904 14028
rect 20956 14016 20962 14068
rect 21450 14016 21456 14068
rect 21508 14056 21514 14068
rect 22097 14059 22155 14065
rect 22097 14056 22109 14059
rect 21508 14028 22109 14056
rect 21508 14016 21514 14028
rect 22097 14025 22109 14028
rect 22143 14025 22155 14059
rect 22462 14056 22468 14068
rect 22423 14028 22468 14056
rect 22097 14019 22155 14025
rect 22462 14016 22468 14028
rect 22520 14016 22526 14068
rect 23198 14056 23204 14068
rect 23159 14028 23204 14056
rect 23198 14016 23204 14028
rect 23256 14016 23262 14068
rect 24946 14016 24952 14068
rect 25004 14056 25010 14068
rect 25041 14059 25099 14065
rect 25041 14056 25053 14059
rect 25004 14028 25053 14056
rect 25004 14016 25010 14028
rect 25041 14025 25053 14028
rect 25087 14025 25099 14059
rect 25041 14019 25099 14025
rect 14369 13991 14427 13997
rect 14369 13957 14381 13991
rect 14415 13957 14427 13991
rect 14369 13951 14427 13957
rect 15749 13991 15807 13997
rect 15749 13957 15761 13991
rect 15795 13988 15807 13991
rect 16022 13988 16028 14000
rect 15795 13960 16028 13988
rect 15795 13957 15807 13960
rect 15749 13951 15807 13957
rect 16022 13948 16028 13960
rect 16080 13948 16086 14000
rect 17586 13948 17592 14000
rect 17644 13988 17650 14000
rect 17865 13991 17923 13997
rect 17865 13988 17877 13991
rect 17644 13960 17877 13988
rect 17644 13948 17650 13960
rect 17865 13957 17877 13960
rect 17911 13988 17923 13991
rect 18874 13988 18880 14000
rect 17911 13960 18880 13988
rect 17911 13957 17923 13960
rect 17865 13951 17923 13957
rect 18874 13948 18880 13960
rect 18932 13948 18938 14000
rect 19886 13988 19892 14000
rect 19847 13960 19892 13988
rect 19886 13948 19892 13960
rect 19944 13948 19950 14000
rect 20162 13988 20168 14000
rect 20123 13960 20168 13988
rect 20162 13948 20168 13960
rect 20220 13948 20226 14000
rect 20916 13988 20944 14016
rect 23106 13988 23112 14000
rect 20916 13960 23112 13988
rect 23106 13948 23112 13960
rect 23164 13948 23170 14000
rect 24670 13988 24676 14000
rect 24631 13960 24676 13988
rect 24670 13948 24676 13960
rect 24728 13988 24734 14000
rect 25406 13988 25412 14000
rect 24728 13960 25412 13988
rect 24728 13948 24734 13960
rect 25406 13948 25412 13960
rect 25464 13948 25470 14000
rect 12434 13880 12440 13932
rect 12492 13920 12498 13932
rect 13081 13923 13139 13929
rect 13081 13920 13093 13923
rect 12492 13892 13093 13920
rect 12492 13880 12498 13892
rect 13081 13889 13093 13892
rect 13127 13889 13139 13923
rect 14734 13920 14740 13932
rect 14695 13892 14740 13920
rect 13081 13883 13139 13889
rect 14734 13880 14740 13892
rect 14792 13880 14798 13932
rect 16485 13923 16543 13929
rect 16485 13889 16497 13923
rect 16531 13920 16543 13923
rect 16758 13920 16764 13932
rect 16531 13892 16764 13920
rect 16531 13889 16543 13892
rect 16485 13883 16543 13889
rect 16758 13880 16764 13892
rect 16816 13880 16822 13932
rect 20809 13923 20867 13929
rect 20809 13889 20821 13923
rect 20855 13920 20867 13923
rect 20990 13920 20996 13932
rect 20855 13892 20996 13920
rect 20855 13889 20867 13892
rect 20809 13883 20867 13889
rect 20990 13880 20996 13892
rect 21048 13880 21054 13932
rect 21174 13920 21180 13932
rect 21135 13892 21180 13920
rect 21174 13880 21180 13892
rect 21232 13880 21238 13932
rect 25498 13880 25504 13932
rect 25556 13920 25562 13932
rect 25731 13923 25789 13929
rect 25731 13920 25743 13923
rect 25556 13892 25743 13920
rect 25556 13880 25562 13892
rect 25731 13889 25743 13892
rect 25777 13889 25789 13923
rect 25731 13883 25789 13889
rect 10042 13852 10048 13864
rect 9600 13824 10048 13852
rect 9692 13793 9720 13824
rect 10042 13812 10048 13824
rect 10100 13852 10106 13864
rect 10505 13855 10563 13861
rect 10505 13852 10517 13855
rect 10100 13824 10517 13852
rect 10100 13812 10106 13824
rect 10505 13821 10517 13824
rect 10551 13821 10563 13855
rect 11330 13852 11336 13864
rect 11291 13824 11336 13852
rect 10505 13815 10563 13821
rect 11330 13812 11336 13824
rect 11388 13812 11394 13864
rect 12621 13855 12679 13861
rect 12621 13821 12633 13855
rect 12667 13852 12679 13855
rect 12802 13852 12808 13864
rect 12667 13824 12808 13852
rect 12667 13821 12679 13824
rect 12621 13815 12679 13821
rect 12802 13812 12808 13824
rect 12860 13812 12866 13864
rect 12897 13855 12955 13861
rect 12897 13821 12909 13855
rect 12943 13852 12955 13855
rect 13633 13855 13691 13861
rect 13633 13852 13645 13855
rect 12943 13824 13645 13852
rect 12943 13821 12955 13824
rect 12897 13815 12955 13821
rect 13633 13821 13645 13824
rect 13679 13852 13691 13855
rect 13906 13852 13912 13864
rect 13679 13824 13912 13852
rect 13679 13821 13691 13824
rect 13633 13815 13691 13821
rect 7146 13787 7204 13793
rect 7146 13753 7158 13787
rect 7192 13753 7204 13787
rect 7146 13747 7204 13753
rect 9671 13787 9729 13793
rect 9671 13753 9683 13787
rect 9717 13753 9729 13787
rect 12158 13784 12164 13796
rect 9671 13747 9729 13753
rect 11164 13756 12164 13784
rect 4522 13716 4528 13728
rect 1636 13688 4528 13716
rect 1636 13676 1642 13688
rect 4522 13676 4528 13688
rect 4580 13676 4586 13728
rect 9858 13676 9864 13728
rect 9916 13716 9922 13728
rect 10229 13719 10287 13725
rect 10229 13716 10241 13719
rect 9916 13688 10241 13716
rect 9916 13676 9922 13688
rect 10229 13685 10241 13688
rect 10275 13685 10287 13719
rect 10229 13679 10287 13685
rect 10686 13676 10692 13728
rect 10744 13716 10750 13728
rect 11164 13725 11192 13756
rect 12158 13744 12164 13756
rect 12216 13744 12222 13796
rect 11149 13719 11207 13725
rect 11149 13716 11161 13719
rect 10744 13688 11161 13716
rect 10744 13676 10750 13688
rect 11149 13685 11161 13688
rect 11195 13685 11207 13719
rect 11149 13679 11207 13685
rect 11422 13676 11428 13728
rect 11480 13716 11486 13728
rect 11698 13716 11704 13728
rect 11480 13688 11704 13716
rect 11480 13676 11486 13688
rect 11698 13676 11704 13688
rect 11756 13676 11762 13728
rect 11790 13676 11796 13728
rect 11848 13716 11854 13728
rect 12069 13719 12127 13725
rect 12069 13716 12081 13719
rect 11848 13688 12081 13716
rect 11848 13676 11854 13688
rect 12069 13685 12081 13688
rect 12115 13716 12127 13719
rect 12342 13716 12348 13728
rect 12115 13688 12348 13716
rect 12115 13685 12127 13688
rect 12069 13679 12127 13685
rect 12342 13676 12348 13688
rect 12400 13716 12406 13728
rect 12912 13716 12940 13815
rect 13906 13812 13912 13824
rect 13964 13812 13970 13864
rect 14277 13855 14335 13861
rect 14277 13821 14289 13855
rect 14323 13821 14335 13855
rect 14277 13815 14335 13821
rect 14292 13784 14320 13815
rect 14458 13812 14464 13864
rect 14516 13852 14522 13864
rect 14553 13855 14611 13861
rect 14553 13852 14565 13855
rect 14516 13824 14565 13852
rect 14516 13812 14522 13824
rect 14553 13821 14565 13824
rect 14599 13821 14611 13855
rect 18322 13852 18328 13864
rect 18283 13824 18328 13852
rect 14553 13815 14611 13821
rect 18322 13812 18328 13824
rect 18380 13852 18386 13864
rect 18969 13855 19027 13861
rect 18969 13852 18981 13855
rect 18380 13824 18981 13852
rect 18380 13812 18386 13824
rect 18969 13821 18981 13824
rect 19015 13821 19027 13855
rect 22278 13852 22284 13864
rect 22191 13824 22284 13852
rect 18969 13815 19027 13821
rect 22278 13812 22284 13824
rect 22336 13852 22342 13864
rect 22741 13855 22799 13861
rect 22741 13852 22753 13855
rect 22336 13824 22753 13852
rect 22336 13812 22342 13824
rect 22741 13821 22753 13824
rect 22787 13821 22799 13855
rect 23845 13855 23903 13861
rect 23845 13852 23857 13855
rect 22741 13815 22799 13821
rect 23400 13824 23857 13852
rect 14642 13784 14648 13796
rect 14292 13756 14648 13784
rect 14642 13744 14648 13756
rect 14700 13744 14706 13796
rect 16574 13784 16580 13796
rect 16535 13756 16580 13784
rect 16574 13744 16580 13756
rect 16632 13744 16638 13796
rect 17129 13787 17187 13793
rect 17129 13753 17141 13787
rect 17175 13784 17187 13787
rect 17310 13784 17316 13796
rect 17175 13756 17316 13784
rect 17175 13753 17187 13756
rect 17129 13747 17187 13753
rect 17310 13744 17316 13756
rect 17368 13744 17374 13796
rect 19290 13787 19348 13793
rect 19290 13784 19302 13787
rect 18984 13756 19302 13784
rect 18984 13728 19012 13756
rect 19290 13753 19302 13756
rect 19336 13753 19348 13787
rect 19290 13747 19348 13753
rect 20898 13744 20904 13796
rect 20956 13784 20962 13796
rect 20956 13756 21001 13784
rect 20956 13744 20962 13756
rect 23290 13744 23296 13796
rect 23348 13784 23354 13796
rect 23400 13784 23428 13824
rect 23845 13821 23857 13824
rect 23891 13852 23903 13855
rect 23891 13824 23980 13852
rect 23891 13821 23903 13824
rect 23845 13815 23903 13821
rect 23348 13756 23428 13784
rect 23348 13744 23354 13756
rect 12400 13688 12940 13716
rect 12400 13676 12406 13688
rect 17402 13676 17408 13728
rect 17460 13716 17466 13728
rect 17497 13719 17555 13725
rect 17497 13716 17509 13719
rect 17460 13688 17509 13716
rect 17460 13676 17466 13688
rect 17497 13685 17509 13688
rect 17543 13716 17555 13719
rect 17586 13716 17592 13728
rect 17543 13688 17592 13716
rect 17543 13685 17555 13688
rect 17497 13679 17555 13685
rect 17586 13676 17592 13688
rect 17644 13676 17650 13728
rect 18506 13676 18512 13728
rect 18564 13716 18570 13728
rect 18966 13716 18972 13728
rect 18564 13688 18972 13716
rect 18564 13676 18570 13688
rect 18966 13676 18972 13688
rect 19024 13676 19030 13728
rect 21726 13716 21732 13728
rect 21687 13688 21732 13716
rect 21726 13676 21732 13688
rect 21784 13676 21790 13728
rect 23952 13716 23980 13824
rect 25590 13812 25596 13864
rect 25648 13861 25654 13864
rect 25648 13855 25686 13861
rect 25674 13852 25686 13855
rect 26053 13855 26111 13861
rect 26053 13852 26065 13855
rect 25674 13824 26065 13852
rect 25674 13821 25686 13824
rect 25648 13815 25686 13821
rect 26053 13821 26065 13824
rect 26099 13821 26111 13855
rect 26053 13815 26111 13821
rect 25648 13812 25654 13815
rect 24118 13784 24124 13796
rect 24079 13756 24124 13784
rect 24118 13744 24124 13756
rect 24176 13744 24182 13796
rect 24213 13787 24271 13793
rect 24213 13753 24225 13787
rect 24259 13753 24271 13787
rect 24213 13747 24271 13753
rect 24228 13716 24256 13747
rect 23952 13688 24256 13716
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1578 13512 1584 13524
rect 1539 13484 1584 13512
rect 1578 13472 1584 13484
rect 1636 13472 1642 13524
rect 3050 13512 3056 13524
rect 3011 13484 3056 13512
rect 3050 13472 3056 13484
rect 3108 13472 3114 13524
rect 3510 13512 3516 13524
rect 3471 13484 3516 13512
rect 3510 13472 3516 13484
rect 3568 13472 3574 13524
rect 4338 13472 4344 13524
rect 4396 13512 4402 13524
rect 4709 13515 4767 13521
rect 4709 13512 4721 13515
rect 4396 13484 4721 13512
rect 4396 13472 4402 13484
rect 4709 13481 4721 13484
rect 4755 13481 4767 13515
rect 6730 13512 6736 13524
rect 6691 13484 6736 13512
rect 4709 13475 4767 13481
rect 6730 13472 6736 13484
rect 6788 13472 6794 13524
rect 8757 13515 8815 13521
rect 8757 13481 8769 13515
rect 8803 13481 8815 13515
rect 9306 13512 9312 13524
rect 9267 13484 9312 13512
rect 8757 13475 8815 13481
rect 2130 13404 2136 13456
rect 2188 13444 2194 13456
rect 2225 13447 2283 13453
rect 2225 13444 2237 13447
rect 2188 13416 2237 13444
rect 2188 13404 2194 13416
rect 2225 13413 2237 13416
rect 2271 13444 2283 13447
rect 2406 13444 2412 13456
rect 2271 13416 2412 13444
rect 2271 13413 2283 13416
rect 2225 13407 2283 13413
rect 2406 13404 2412 13416
rect 2464 13404 2470 13456
rect 4430 13444 4436 13456
rect 4391 13416 4436 13444
rect 4430 13404 4436 13416
rect 4488 13404 4494 13456
rect 6178 13404 6184 13456
rect 6236 13444 6242 13456
rect 7101 13447 7159 13453
rect 7101 13444 7113 13447
rect 6236 13416 7113 13444
rect 6236 13404 6242 13416
rect 7101 13413 7113 13416
rect 7147 13444 7159 13447
rect 7190 13444 7196 13456
rect 7147 13416 7196 13444
rect 7147 13413 7159 13416
rect 7101 13407 7159 13413
rect 7190 13404 7196 13416
rect 7248 13404 7254 13456
rect 7650 13444 7656 13456
rect 7611 13416 7656 13444
rect 7650 13404 7656 13416
rect 7708 13404 7714 13456
rect 8481 13447 8539 13453
rect 8481 13413 8493 13447
rect 8527 13444 8539 13447
rect 8772 13444 8800 13475
rect 9306 13472 9312 13484
rect 9364 13472 9370 13524
rect 9692 13484 11100 13512
rect 9692 13444 9720 13484
rect 9858 13444 9864 13456
rect 8527 13416 9720 13444
rect 9819 13416 9864 13444
rect 8527 13413 8539 13416
rect 8481 13407 8539 13413
rect 9858 13404 9864 13416
rect 9916 13404 9922 13456
rect 11072 13444 11100 13484
rect 11146 13472 11152 13524
rect 11204 13512 11210 13524
rect 12069 13515 12127 13521
rect 12069 13512 12081 13515
rect 11204 13484 12081 13512
rect 11204 13472 11210 13484
rect 12069 13481 12081 13484
rect 12115 13481 12127 13515
rect 12069 13475 12127 13481
rect 13081 13515 13139 13521
rect 13081 13481 13093 13515
rect 13127 13512 13139 13515
rect 13354 13512 13360 13524
rect 13127 13484 13360 13512
rect 13127 13481 13139 13484
rect 13081 13475 13139 13481
rect 13354 13472 13360 13484
rect 13412 13472 13418 13524
rect 13998 13472 14004 13524
rect 14056 13512 14062 13524
rect 14277 13515 14335 13521
rect 14277 13512 14289 13515
rect 14056 13484 14289 13512
rect 14056 13472 14062 13484
rect 14277 13481 14289 13484
rect 14323 13481 14335 13515
rect 14277 13475 14335 13481
rect 14642 13472 14648 13524
rect 14700 13512 14706 13524
rect 15013 13515 15071 13521
rect 15013 13512 15025 13515
rect 14700 13484 15025 13512
rect 14700 13472 14706 13484
rect 15013 13481 15025 13484
rect 15059 13481 15071 13515
rect 15838 13512 15844 13524
rect 15799 13484 15844 13512
rect 15013 13475 15071 13481
rect 15838 13472 15844 13484
rect 15896 13472 15902 13524
rect 18598 13512 18604 13524
rect 17328 13484 18604 13512
rect 17328 13456 17356 13484
rect 18598 13472 18604 13484
rect 18656 13512 18662 13524
rect 18656 13484 18920 13512
rect 18656 13472 18662 13484
rect 11072 13416 11744 13444
rect 4890 13376 4896 13388
rect 4851 13348 4896 13376
rect 4890 13336 4896 13348
rect 4948 13336 4954 13388
rect 5166 13376 5172 13388
rect 5127 13348 5172 13376
rect 5166 13336 5172 13348
rect 5224 13336 5230 13388
rect 8570 13376 8576 13388
rect 8531 13348 8576 13376
rect 8570 13336 8576 13348
rect 8628 13336 8634 13388
rect 11146 13376 11152 13388
rect 11059 13348 11152 13376
rect 11146 13336 11152 13348
rect 11204 13376 11210 13388
rect 11330 13376 11336 13388
rect 11204 13348 11336 13376
rect 11204 13336 11210 13348
rect 11330 13336 11336 13348
rect 11388 13336 11394 13388
rect 11609 13379 11667 13385
rect 11609 13345 11621 13379
rect 11655 13345 11667 13379
rect 11609 13339 11667 13345
rect 2133 13311 2191 13317
rect 2133 13308 2145 13311
rect 2056 13280 2145 13308
rect 2056 13252 2084 13280
rect 2133 13277 2145 13280
rect 2179 13277 2191 13311
rect 2133 13271 2191 13277
rect 7009 13311 7067 13317
rect 7009 13277 7021 13311
rect 7055 13308 7067 13311
rect 7098 13308 7104 13320
rect 7055 13280 7104 13308
rect 7055 13277 7067 13280
rect 7009 13271 7067 13277
rect 7098 13268 7104 13280
rect 7156 13268 7162 13320
rect 9490 13268 9496 13320
rect 9548 13308 9554 13320
rect 9766 13308 9772 13320
rect 9548 13280 9772 13308
rect 9548 13268 9554 13280
rect 9766 13268 9772 13280
rect 9824 13268 9830 13320
rect 10042 13308 10048 13320
rect 10003 13280 10048 13308
rect 10042 13268 10048 13280
rect 10100 13268 10106 13320
rect 11238 13268 11244 13320
rect 11296 13308 11302 13320
rect 11624 13308 11652 13339
rect 11296 13280 11652 13308
rect 11716 13308 11744 13416
rect 11790 13404 11796 13456
rect 11848 13444 11854 13456
rect 12621 13447 12679 13453
rect 12621 13444 12633 13447
rect 11848 13416 12633 13444
rect 11848 13404 11854 13416
rect 12621 13413 12633 13416
rect 12667 13413 12679 13447
rect 12621 13407 12679 13413
rect 16761 13447 16819 13453
rect 16761 13413 16773 13447
rect 16807 13444 16819 13447
rect 17126 13444 17132 13456
rect 16807 13416 17132 13444
rect 16807 13413 16819 13416
rect 16761 13407 16819 13413
rect 17126 13404 17132 13416
rect 17184 13404 17190 13456
rect 17310 13444 17316 13456
rect 17271 13416 17316 13444
rect 17310 13404 17316 13416
rect 17368 13404 17374 13456
rect 18046 13404 18052 13456
rect 18104 13444 18110 13456
rect 18892 13453 18920 13484
rect 18966 13472 18972 13524
rect 19024 13512 19030 13524
rect 19153 13515 19211 13521
rect 19153 13512 19165 13515
rect 19024 13484 19165 13512
rect 19024 13472 19030 13484
rect 19153 13481 19165 13484
rect 19199 13481 19211 13515
rect 19153 13475 19211 13481
rect 20990 13472 20996 13524
rect 21048 13512 21054 13524
rect 21085 13515 21143 13521
rect 21085 13512 21097 13515
rect 21048 13484 21097 13512
rect 21048 13472 21054 13484
rect 21085 13481 21097 13484
rect 21131 13481 21143 13515
rect 21085 13475 21143 13481
rect 23017 13515 23075 13521
rect 23017 13481 23029 13515
rect 23063 13512 23075 13515
rect 23063 13484 23428 13512
rect 23063 13481 23075 13484
rect 23017 13475 23075 13481
rect 23400 13456 23428 13484
rect 18325 13447 18383 13453
rect 18325 13444 18337 13447
rect 18104 13416 18337 13444
rect 18104 13404 18110 13416
rect 18325 13413 18337 13416
rect 18371 13413 18383 13447
rect 18325 13407 18383 13413
rect 18877 13447 18935 13453
rect 18877 13413 18889 13447
rect 18923 13413 18935 13447
rect 21634 13444 21640 13456
rect 21595 13416 21640 13444
rect 18877 13407 18935 13413
rect 21634 13404 21640 13416
rect 21692 13404 21698 13456
rect 23290 13444 23296 13456
rect 23251 13416 23296 13444
rect 23290 13404 23296 13416
rect 23348 13404 23354 13456
rect 23382 13404 23388 13456
rect 23440 13444 23446 13456
rect 23845 13447 23903 13453
rect 23845 13444 23857 13447
rect 23440 13416 23857 13444
rect 23440 13404 23446 13416
rect 23845 13413 23857 13416
rect 23891 13413 23903 13447
rect 24762 13444 24768 13456
rect 24723 13416 24768 13444
rect 23845 13407 23903 13413
rect 24762 13404 24768 13416
rect 24820 13404 24826 13456
rect 24854 13404 24860 13456
rect 24912 13444 24918 13456
rect 25406 13444 25412 13456
rect 24912 13416 24957 13444
rect 25367 13416 25412 13444
rect 24912 13404 24918 13416
rect 25406 13404 25412 13416
rect 25464 13404 25470 13456
rect 11882 13376 11888 13388
rect 11843 13348 11888 13376
rect 11882 13336 11888 13348
rect 11940 13336 11946 13388
rect 13170 13376 13176 13388
rect 13131 13348 13176 13376
rect 13170 13336 13176 13348
rect 13228 13336 13234 13388
rect 13446 13376 13452 13388
rect 13407 13348 13452 13376
rect 13446 13336 13452 13348
rect 13504 13336 13510 13388
rect 15286 13376 15292 13388
rect 15247 13348 15292 13376
rect 15286 13336 15292 13348
rect 15344 13336 15350 13388
rect 19794 13376 19800 13388
rect 19758 13348 19800 13376
rect 19794 13336 19800 13348
rect 19852 13385 19858 13388
rect 19852 13379 19906 13385
rect 19852 13345 19860 13379
rect 19894 13376 19906 13379
rect 20806 13376 20812 13388
rect 19894 13348 20812 13376
rect 19894 13345 19906 13348
rect 19852 13339 19906 13345
rect 19852 13336 19858 13339
rect 20806 13336 20812 13348
rect 20864 13336 20870 13388
rect 13909 13311 13967 13317
rect 11716 13280 13860 13308
rect 11296 13268 11302 13280
rect 2038 13200 2044 13252
rect 2096 13200 2102 13252
rect 2682 13240 2688 13252
rect 2643 13212 2688 13240
rect 2682 13200 2688 13212
rect 2740 13200 2746 13252
rect 5994 13132 6000 13184
rect 6052 13172 6058 13184
rect 8481 13175 8539 13181
rect 8481 13172 8493 13175
rect 6052 13144 8493 13172
rect 6052 13132 6058 13144
rect 8481 13141 8493 13144
rect 8527 13141 8539 13175
rect 8481 13135 8539 13141
rect 11517 13175 11575 13181
rect 11517 13141 11529 13175
rect 11563 13172 11575 13175
rect 11624 13172 11652 13280
rect 11701 13243 11759 13249
rect 11701 13209 11713 13243
rect 11747 13240 11759 13243
rect 11790 13240 11796 13252
rect 11747 13212 11796 13240
rect 11747 13209 11759 13212
rect 11701 13203 11759 13209
rect 11790 13200 11796 13212
rect 11848 13200 11854 13252
rect 13262 13240 13268 13252
rect 13223 13212 13268 13240
rect 13262 13200 13268 13212
rect 13320 13200 13326 13252
rect 13832 13240 13860 13280
rect 13909 13277 13921 13311
rect 13955 13308 13967 13311
rect 13998 13308 14004 13320
rect 13955 13280 14004 13308
rect 13955 13277 13967 13280
rect 13909 13271 13967 13277
rect 13998 13268 14004 13280
rect 14056 13268 14062 13320
rect 16669 13311 16727 13317
rect 16669 13277 16681 13311
rect 16715 13308 16727 13311
rect 16758 13308 16764 13320
rect 16715 13280 16764 13308
rect 16715 13277 16727 13280
rect 16669 13271 16727 13277
rect 16758 13268 16764 13280
rect 16816 13268 16822 13320
rect 18233 13311 18291 13317
rect 18233 13308 18245 13311
rect 17972 13280 18245 13308
rect 17586 13240 17592 13252
rect 13832 13212 17592 13240
rect 17586 13200 17592 13212
rect 17644 13200 17650 13252
rect 17972 13184 18000 13280
rect 18233 13277 18245 13280
rect 18279 13277 18291 13311
rect 18233 13271 18291 13277
rect 19935 13311 19993 13317
rect 19935 13277 19947 13311
rect 19981 13308 19993 13311
rect 20714 13308 20720 13320
rect 19981 13280 20720 13308
rect 19981 13277 19993 13280
rect 19935 13271 19993 13277
rect 20714 13268 20720 13280
rect 20772 13308 20778 13320
rect 21545 13311 21603 13317
rect 21545 13308 21557 13311
rect 20772 13280 21557 13308
rect 20772 13268 20778 13280
rect 21545 13277 21557 13280
rect 21591 13277 21603 13311
rect 22186 13308 22192 13320
rect 22147 13280 22192 13308
rect 21545 13271 21603 13277
rect 22186 13268 22192 13280
rect 22244 13268 22250 13320
rect 23201 13311 23259 13317
rect 23201 13277 23213 13311
rect 23247 13308 23259 13311
rect 23842 13308 23848 13320
rect 23247 13280 23848 13308
rect 23247 13277 23259 13280
rect 23201 13271 23259 13277
rect 23842 13268 23848 13280
rect 23900 13268 23906 13320
rect 12618 13172 12624 13184
rect 11563 13144 12624 13172
rect 11563 13141 11575 13144
rect 11517 13135 11575 13141
rect 12618 13132 12624 13144
rect 12676 13132 12682 13184
rect 14274 13132 14280 13184
rect 14332 13172 14338 13184
rect 14645 13175 14703 13181
rect 14645 13172 14657 13175
rect 14332 13144 14657 13172
rect 14332 13132 14338 13144
rect 14645 13141 14657 13144
rect 14691 13141 14703 13175
rect 14645 13135 14703 13141
rect 14734 13132 14740 13184
rect 14792 13172 14798 13184
rect 15473 13175 15531 13181
rect 15473 13172 15485 13175
rect 14792 13144 15485 13172
rect 14792 13132 14798 13144
rect 15473 13141 15485 13144
rect 15519 13141 15531 13175
rect 15473 13135 15531 13141
rect 16485 13175 16543 13181
rect 16485 13141 16497 13175
rect 16531 13172 16543 13175
rect 16574 13172 16580 13184
rect 16531 13144 16580 13172
rect 16531 13141 16543 13144
rect 16485 13135 16543 13141
rect 16574 13132 16580 13144
rect 16632 13132 16638 13184
rect 17954 13172 17960 13184
rect 17915 13144 17960 13172
rect 17954 13132 17960 13144
rect 18012 13132 18018 13184
rect 24118 13172 24124 13184
rect 24079 13144 24124 13172
rect 24118 13132 24124 13144
rect 24176 13132 24182 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1949 12971 2007 12977
rect 1949 12937 1961 12971
rect 1995 12968 2007 12971
rect 2222 12968 2228 12980
rect 1995 12940 2228 12968
rect 1995 12937 2007 12940
rect 1949 12931 2007 12937
rect 1964 12696 1992 12931
rect 2222 12928 2228 12940
rect 2280 12928 2286 12980
rect 7098 12928 7104 12980
rect 7156 12968 7162 12980
rect 7837 12971 7895 12977
rect 7837 12968 7849 12971
rect 7156 12940 7849 12968
rect 7156 12928 7162 12940
rect 7837 12937 7849 12940
rect 7883 12937 7895 12971
rect 8570 12968 8576 12980
rect 8531 12940 8576 12968
rect 7837 12931 7895 12937
rect 8570 12928 8576 12940
rect 8628 12928 8634 12980
rect 9858 12928 9864 12980
rect 9916 12968 9922 12980
rect 10229 12971 10287 12977
rect 10229 12968 10241 12971
rect 9916 12940 10241 12968
rect 9916 12928 9922 12940
rect 10229 12937 10241 12940
rect 10275 12937 10287 12971
rect 10229 12931 10287 12937
rect 15197 12971 15255 12977
rect 15197 12937 15209 12971
rect 15243 12968 15255 12971
rect 15286 12968 15292 12980
rect 15243 12940 15292 12968
rect 15243 12937 15255 12940
rect 15197 12931 15255 12937
rect 15286 12928 15292 12940
rect 15344 12928 15350 12980
rect 16574 12968 16580 12980
rect 16535 12940 16580 12968
rect 16574 12928 16580 12940
rect 16632 12928 16638 12980
rect 17126 12928 17132 12980
rect 17184 12968 17190 12980
rect 17221 12971 17279 12977
rect 17221 12968 17233 12971
rect 17184 12940 17233 12968
rect 17184 12928 17190 12940
rect 17221 12937 17233 12940
rect 17267 12968 17279 12971
rect 17310 12968 17316 12980
rect 17267 12940 17316 12968
rect 17267 12937 17279 12940
rect 17221 12931 17279 12937
rect 17310 12928 17316 12940
rect 17368 12928 17374 12980
rect 19794 12968 19800 12980
rect 19755 12940 19800 12968
rect 19794 12928 19800 12940
rect 19852 12928 19858 12980
rect 21634 12928 21640 12980
rect 21692 12968 21698 12980
rect 23201 12971 23259 12977
rect 21692 12940 22600 12968
rect 21692 12928 21698 12940
rect 2682 12900 2688 12912
rect 2643 12872 2688 12900
rect 2682 12860 2688 12872
rect 2740 12860 2746 12912
rect 4430 12900 4436 12912
rect 4343 12872 4436 12900
rect 4430 12860 4436 12872
rect 4488 12900 4494 12912
rect 5534 12900 5540 12912
rect 4488 12872 5463 12900
rect 5495 12872 5540 12900
rect 4488 12860 4494 12872
rect 2133 12835 2191 12841
rect 2133 12801 2145 12835
rect 2179 12832 2191 12835
rect 2406 12832 2412 12844
rect 2179 12804 2412 12832
rect 2179 12801 2191 12804
rect 2133 12795 2191 12801
rect 2406 12792 2412 12804
rect 2464 12832 2470 12844
rect 3053 12835 3111 12841
rect 3053 12832 3065 12835
rect 2464 12804 3065 12832
rect 2464 12792 2470 12804
rect 3053 12801 3065 12804
rect 3099 12801 3111 12835
rect 3053 12795 3111 12801
rect 4893 12835 4951 12841
rect 4893 12801 4905 12835
rect 4939 12832 4951 12835
rect 5166 12832 5172 12844
rect 4939 12804 5172 12832
rect 4939 12801 4951 12804
rect 4893 12795 4951 12801
rect 5166 12792 5172 12804
rect 5224 12792 5230 12844
rect 5435 12832 5463 12872
rect 5534 12860 5540 12872
rect 5592 12860 5598 12912
rect 12894 12900 12900 12912
rect 12855 12872 12900 12900
rect 12894 12860 12900 12872
rect 12952 12860 12958 12912
rect 15565 12903 15623 12909
rect 15565 12869 15577 12903
rect 15611 12900 15623 12903
rect 15746 12900 15752 12912
rect 15611 12872 15752 12900
rect 15611 12869 15623 12872
rect 15565 12863 15623 12869
rect 15746 12860 15752 12872
rect 15804 12900 15810 12912
rect 18506 12900 18512 12912
rect 15804 12872 18512 12900
rect 15804 12860 15810 12872
rect 18506 12860 18512 12872
rect 18564 12860 18570 12912
rect 9585 12835 9643 12841
rect 9585 12832 9597 12835
rect 5435 12804 9597 12832
rect 9585 12801 9597 12804
rect 9631 12801 9643 12835
rect 9585 12795 9643 12801
rect 11514 12792 11520 12844
rect 11572 12832 11578 12844
rect 14274 12832 14280 12844
rect 11572 12804 14280 12832
rect 11572 12792 11578 12804
rect 5350 12764 5356 12776
rect 5311 12736 5356 12764
rect 5350 12724 5356 12736
rect 5408 12724 5414 12776
rect 6546 12724 6552 12776
rect 6604 12764 6610 12776
rect 6641 12767 6699 12773
rect 6641 12764 6653 12767
rect 6604 12736 6653 12764
rect 6604 12724 6610 12736
rect 6641 12733 6653 12736
rect 6687 12764 6699 12767
rect 7101 12767 7159 12773
rect 7101 12764 7113 12767
rect 6687 12736 7113 12764
rect 6687 12733 6699 12736
rect 6641 12727 6699 12733
rect 7101 12733 7113 12736
rect 7147 12733 7159 12767
rect 7101 12727 7159 12733
rect 7377 12767 7435 12773
rect 7377 12733 7389 12767
rect 7423 12764 7435 12767
rect 7558 12764 7564 12776
rect 7423 12736 7564 12764
rect 7423 12733 7435 12736
rect 7377 12727 7435 12733
rect 2225 12699 2283 12705
rect 2225 12696 2237 12699
rect 1964 12668 2237 12696
rect 2225 12665 2237 12668
rect 2271 12696 2283 12699
rect 2498 12696 2504 12708
rect 2271 12668 2504 12696
rect 2271 12665 2283 12668
rect 2225 12659 2283 12665
rect 2498 12656 2504 12668
rect 2556 12656 2562 12708
rect 3878 12696 3884 12708
rect 3839 12668 3884 12696
rect 3878 12656 3884 12668
rect 3936 12656 3942 12708
rect 3973 12699 4031 12705
rect 3973 12665 3985 12699
rect 4019 12665 4031 12699
rect 7116 12696 7144 12727
rect 7558 12724 7564 12736
rect 7616 12724 7622 12776
rect 10689 12767 10747 12773
rect 10689 12733 10701 12767
rect 10735 12764 10747 12767
rect 11422 12764 11428 12776
rect 10735 12736 11428 12764
rect 10735 12733 10747 12736
rect 10689 12727 10747 12733
rect 11422 12724 11428 12736
rect 11480 12764 11486 12776
rect 11882 12764 11888 12776
rect 11480 12736 11888 12764
rect 11480 12724 11486 12736
rect 11882 12724 11888 12736
rect 11940 12724 11946 12776
rect 12802 12724 12808 12776
rect 12860 12764 12866 12776
rect 14108 12773 14136 12804
rect 14274 12792 14280 12804
rect 14332 12792 14338 12844
rect 18598 12832 18604 12844
rect 18559 12804 18604 12832
rect 18598 12792 18604 12804
rect 18656 12792 18662 12844
rect 20622 12832 20628 12844
rect 20583 12804 20628 12832
rect 20622 12792 20628 12804
rect 20680 12792 20686 12844
rect 21361 12835 21419 12841
rect 21361 12801 21373 12835
rect 21407 12832 21419 12835
rect 21545 12835 21603 12841
rect 21545 12832 21557 12835
rect 21407 12804 21557 12832
rect 21407 12801 21419 12804
rect 21361 12795 21419 12801
rect 21545 12801 21557 12804
rect 21591 12832 21603 12835
rect 22002 12832 22008 12844
rect 21591 12804 22008 12832
rect 21591 12801 21603 12804
rect 21545 12795 21603 12801
rect 22002 12792 22008 12804
rect 22060 12792 22066 12844
rect 22186 12832 22192 12844
rect 22147 12804 22192 12832
rect 22186 12792 22192 12804
rect 22244 12792 22250 12844
rect 14093 12767 14151 12773
rect 12860 12736 12905 12764
rect 12860 12724 12866 12736
rect 14093 12733 14105 12767
rect 14139 12733 14151 12767
rect 14093 12727 14151 12733
rect 14645 12767 14703 12773
rect 14645 12733 14657 12767
rect 14691 12764 14703 12767
rect 14734 12764 14740 12776
rect 14691 12736 14740 12764
rect 14691 12733 14703 12736
rect 14645 12727 14703 12733
rect 14734 12724 14740 12736
rect 14792 12724 14798 12776
rect 14829 12767 14887 12773
rect 14829 12733 14841 12767
rect 14875 12764 14887 12767
rect 15657 12767 15715 12773
rect 15657 12764 15669 12767
rect 14875 12736 15669 12764
rect 14875 12733 14887 12736
rect 14829 12727 14887 12733
rect 15657 12733 15669 12736
rect 15703 12764 15715 12767
rect 16853 12767 16911 12773
rect 16853 12764 16865 12767
rect 15703 12736 16865 12764
rect 15703 12733 15715 12736
rect 15657 12727 15715 12733
rect 16853 12733 16865 12736
rect 16899 12733 16911 12767
rect 16853 12727 16911 12733
rect 19334 12724 19340 12776
rect 19392 12764 19398 12776
rect 20257 12767 20315 12773
rect 20257 12764 20269 12767
rect 19392 12736 20269 12764
rect 19392 12724 19398 12736
rect 20257 12733 20269 12736
rect 20303 12764 20315 12767
rect 20901 12767 20959 12773
rect 20901 12764 20913 12767
rect 20303 12736 20913 12764
rect 20303 12733 20315 12736
rect 20257 12727 20315 12733
rect 20901 12733 20913 12736
rect 20947 12733 20959 12767
rect 20901 12727 20959 12733
rect 7466 12696 7472 12708
rect 7116 12668 7472 12696
rect 3973 12659 4031 12665
rect 3697 12631 3755 12637
rect 3697 12597 3709 12631
rect 3743 12628 3755 12631
rect 3988 12628 4016 12659
rect 7466 12656 7472 12668
rect 7524 12656 7530 12708
rect 9030 12696 9036 12708
rect 8220 12668 9036 12696
rect 4338 12628 4344 12640
rect 3743 12600 4344 12628
rect 3743 12597 3755 12600
rect 3697 12591 3755 12597
rect 4338 12588 4344 12600
rect 4396 12588 4402 12640
rect 4890 12588 4896 12640
rect 4948 12628 4954 12640
rect 5261 12631 5319 12637
rect 5261 12628 5273 12631
rect 4948 12600 5273 12628
rect 4948 12588 4954 12600
rect 5261 12597 5273 12600
rect 5307 12628 5319 12631
rect 5994 12628 6000 12640
rect 5307 12600 6000 12628
rect 5307 12597 5319 12600
rect 5261 12591 5319 12597
rect 5994 12588 6000 12600
rect 6052 12588 6058 12640
rect 6178 12628 6184 12640
rect 6139 12600 6184 12628
rect 6178 12588 6184 12600
rect 6236 12588 6242 12640
rect 7098 12628 7104 12640
rect 7059 12600 7104 12628
rect 7098 12588 7104 12600
rect 7156 12588 7162 12640
rect 8018 12588 8024 12640
rect 8076 12628 8082 12640
rect 8220 12637 8248 12668
rect 9030 12656 9036 12668
rect 9088 12696 9094 12708
rect 9309 12699 9367 12705
rect 9309 12696 9321 12699
rect 9088 12668 9321 12696
rect 9088 12656 9094 12668
rect 9309 12665 9321 12668
rect 9355 12665 9367 12699
rect 9309 12659 9367 12665
rect 9401 12699 9459 12705
rect 9401 12665 9413 12699
rect 9447 12665 9459 12699
rect 9401 12659 9459 12665
rect 11517 12699 11575 12705
rect 11517 12665 11529 12699
rect 11563 12696 11575 12699
rect 11606 12696 11612 12708
rect 11563 12668 11612 12696
rect 11563 12665 11575 12668
rect 11517 12659 11575 12665
rect 8205 12631 8263 12637
rect 8205 12628 8217 12631
rect 8076 12600 8217 12628
rect 8076 12588 8082 12600
rect 8205 12597 8217 12600
rect 8251 12597 8263 12631
rect 8205 12591 8263 12597
rect 9125 12631 9183 12637
rect 9125 12597 9137 12631
rect 9171 12628 9183 12631
rect 9416 12628 9444 12659
rect 11606 12656 11612 12668
rect 11664 12656 11670 12708
rect 12710 12696 12716 12708
rect 12176 12668 12716 12696
rect 9674 12628 9680 12640
rect 9171 12600 9680 12628
rect 9171 12597 9183 12600
rect 9125 12591 9183 12597
rect 9674 12588 9680 12600
rect 9732 12588 9738 12640
rect 11790 12628 11796 12640
rect 11751 12600 11796 12628
rect 11790 12588 11796 12600
rect 11848 12628 11854 12640
rect 12176 12637 12204 12668
rect 12710 12656 12716 12668
rect 12768 12696 12774 12708
rect 13262 12696 13268 12708
rect 12768 12668 13268 12696
rect 12768 12656 12774 12668
rect 13262 12656 13268 12668
rect 13320 12696 13326 12708
rect 13541 12699 13599 12705
rect 13541 12696 13553 12699
rect 13320 12668 13553 12696
rect 13320 12656 13326 12668
rect 13541 12665 13553 12668
rect 13587 12665 13599 12699
rect 13541 12659 13599 12665
rect 15746 12656 15752 12708
rect 15804 12696 15810 12708
rect 15978 12699 16036 12705
rect 15978 12696 15990 12699
rect 15804 12668 15990 12696
rect 15804 12656 15810 12668
rect 15978 12665 15990 12668
rect 16024 12665 16036 12699
rect 15978 12659 16036 12665
rect 17865 12699 17923 12705
rect 17865 12665 17877 12699
rect 17911 12696 17923 12699
rect 18693 12699 18751 12705
rect 17911 12668 18552 12696
rect 17911 12665 17923 12668
rect 17865 12659 17923 12665
rect 12161 12631 12219 12637
rect 12161 12628 12173 12631
rect 11848 12600 12173 12628
rect 11848 12588 11854 12600
rect 12161 12597 12173 12600
rect 12207 12597 12219 12631
rect 12161 12591 12219 12597
rect 12802 12588 12808 12640
rect 12860 12628 12866 12640
rect 13446 12628 13452 12640
rect 12860 12600 13452 12628
rect 12860 12588 12866 12600
rect 13446 12588 13452 12600
rect 13504 12628 13510 12640
rect 13817 12631 13875 12637
rect 13817 12628 13829 12631
rect 13504 12600 13829 12628
rect 13504 12588 13510 12600
rect 13817 12597 13829 12600
rect 13863 12597 13875 12631
rect 13817 12591 13875 12597
rect 18046 12588 18052 12640
rect 18104 12628 18110 12640
rect 18233 12631 18291 12637
rect 18233 12628 18245 12631
rect 18104 12600 18245 12628
rect 18104 12588 18110 12600
rect 18233 12597 18245 12600
rect 18279 12597 18291 12631
rect 18524 12628 18552 12668
rect 18693 12665 18705 12699
rect 18739 12665 18751 12699
rect 19242 12696 19248 12708
rect 19203 12668 19248 12696
rect 18693 12659 18751 12665
rect 18708 12628 18736 12659
rect 19242 12656 19248 12668
rect 19300 12656 19306 12708
rect 20073 12699 20131 12705
rect 20073 12665 20085 12699
rect 20119 12696 20131 12699
rect 21637 12699 21695 12705
rect 20119 12668 20300 12696
rect 20119 12665 20131 12668
rect 20073 12659 20131 12665
rect 20272 12640 20300 12668
rect 21637 12665 21649 12699
rect 21683 12696 21695 12699
rect 21910 12696 21916 12708
rect 21683 12668 21916 12696
rect 21683 12665 21695 12668
rect 21637 12659 21695 12665
rect 21910 12656 21916 12668
rect 21968 12656 21974 12708
rect 22572 12705 22600 12940
rect 23201 12937 23213 12971
rect 23247 12968 23259 12971
rect 23290 12968 23296 12980
rect 23247 12940 23296 12968
rect 23247 12937 23259 12940
rect 23201 12931 23259 12937
rect 23290 12928 23296 12940
rect 23348 12928 23354 12980
rect 23842 12968 23848 12980
rect 23803 12940 23848 12968
rect 23842 12928 23848 12940
rect 23900 12928 23906 12980
rect 24489 12971 24547 12977
rect 24489 12937 24501 12971
rect 24535 12968 24547 12971
rect 24762 12968 24768 12980
rect 24535 12940 24768 12968
rect 24535 12937 24547 12940
rect 24489 12931 24547 12937
rect 24762 12928 24768 12940
rect 24820 12928 24826 12980
rect 24854 12928 24860 12980
rect 24912 12968 24918 12980
rect 25501 12971 25559 12977
rect 25501 12968 25513 12971
rect 24912 12940 25513 12968
rect 24912 12928 24918 12940
rect 25501 12937 25513 12940
rect 25547 12937 25559 12971
rect 25501 12931 25559 12937
rect 24578 12764 24584 12776
rect 24539 12736 24584 12764
rect 24578 12724 24584 12736
rect 24636 12764 24642 12776
rect 25133 12767 25191 12773
rect 25133 12764 25145 12767
rect 24636 12736 25145 12764
rect 24636 12724 24642 12736
rect 25133 12733 25145 12736
rect 25179 12733 25191 12767
rect 25133 12727 25191 12733
rect 22557 12699 22615 12705
rect 22557 12665 22569 12699
rect 22603 12696 22615 12699
rect 23382 12696 23388 12708
rect 22603 12668 23388 12696
rect 22603 12665 22615 12668
rect 22557 12659 22615 12665
rect 23382 12656 23388 12668
rect 23440 12656 23446 12708
rect 18782 12628 18788 12640
rect 18524 12600 18788 12628
rect 18233 12591 18291 12597
rect 18782 12588 18788 12600
rect 18840 12588 18846 12640
rect 20254 12588 20260 12640
rect 20312 12588 20318 12640
rect 24210 12588 24216 12640
rect 24268 12628 24274 12640
rect 24765 12631 24823 12637
rect 24765 12628 24777 12631
rect 24268 12600 24777 12628
rect 24268 12588 24274 12600
rect 24765 12597 24777 12600
rect 24811 12597 24823 12631
rect 24765 12591 24823 12597
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 2130 12424 2136 12436
rect 2091 12396 2136 12424
rect 2130 12384 2136 12396
rect 2188 12384 2194 12436
rect 3878 12424 3884 12436
rect 3068 12396 3884 12424
rect 3068 12368 3096 12396
rect 3878 12384 3884 12396
rect 3936 12384 3942 12436
rect 4522 12384 4528 12436
rect 4580 12424 4586 12436
rect 5721 12427 5779 12433
rect 5721 12424 5733 12427
rect 4580 12396 5733 12424
rect 4580 12384 4586 12396
rect 5721 12393 5733 12396
rect 5767 12393 5779 12427
rect 5721 12387 5779 12393
rect 9033 12427 9091 12433
rect 9033 12393 9045 12427
rect 9079 12424 9091 12427
rect 9490 12424 9496 12436
rect 9079 12396 9496 12424
rect 9079 12393 9091 12396
rect 9033 12387 9091 12393
rect 9490 12384 9496 12396
rect 9548 12384 9554 12436
rect 18414 12424 18420 12436
rect 18156 12396 18420 12424
rect 2038 12356 2044 12368
rect 1688 12328 2044 12356
rect 1394 12044 1400 12096
rect 1452 12084 1458 12096
rect 1688 12093 1716 12328
rect 2038 12316 2044 12328
rect 2096 12316 2102 12368
rect 2225 12359 2283 12365
rect 2225 12325 2237 12359
rect 2271 12356 2283 12359
rect 2501 12359 2559 12365
rect 2501 12356 2513 12359
rect 2271 12328 2513 12356
rect 2271 12325 2283 12328
rect 2225 12319 2283 12325
rect 2501 12325 2513 12328
rect 2547 12325 2559 12359
rect 3050 12356 3056 12368
rect 2963 12328 3056 12356
rect 2501 12319 2559 12325
rect 3050 12316 3056 12328
rect 3108 12316 3114 12368
rect 4246 12356 4252 12368
rect 4207 12328 4252 12356
rect 4246 12316 4252 12328
rect 4304 12316 4310 12368
rect 7190 12316 7196 12368
rect 7248 12356 7254 12368
rect 7469 12359 7527 12365
rect 7469 12356 7481 12359
rect 7248 12328 7481 12356
rect 7248 12316 7254 12328
rect 7469 12325 7481 12328
rect 7515 12325 7527 12359
rect 8018 12356 8024 12368
rect 7979 12328 8024 12356
rect 7469 12319 7527 12325
rect 8018 12316 8024 12328
rect 8076 12316 8082 12368
rect 8846 12316 8852 12368
rect 8904 12356 8910 12368
rect 9861 12359 9919 12365
rect 9861 12356 9873 12359
rect 8904 12328 9873 12356
rect 8904 12316 8910 12328
rect 9861 12325 9873 12328
rect 9907 12356 9919 12359
rect 10134 12356 10140 12368
rect 9907 12328 10140 12356
rect 9907 12325 9919 12328
rect 9861 12319 9919 12325
rect 10134 12316 10140 12328
rect 10192 12316 10198 12368
rect 12805 12359 12863 12365
rect 12805 12325 12817 12359
rect 12851 12356 12863 12359
rect 15473 12359 15531 12365
rect 15473 12356 15485 12359
rect 12851 12328 15485 12356
rect 12851 12325 12863 12328
rect 12805 12319 12863 12325
rect 15473 12325 15485 12328
rect 15519 12356 15531 12359
rect 15519 12328 15700 12356
rect 15519 12325 15531 12328
rect 15473 12319 15531 12325
rect 5905 12291 5963 12297
rect 5905 12257 5917 12291
rect 5951 12288 5963 12291
rect 5994 12288 6000 12300
rect 5951 12260 6000 12288
rect 5951 12257 5963 12260
rect 5905 12251 5963 12257
rect 5994 12248 6000 12260
rect 6052 12248 6058 12300
rect 6181 12291 6239 12297
rect 6181 12257 6193 12291
rect 6227 12288 6239 12291
rect 6546 12288 6552 12300
rect 6227 12260 6552 12288
rect 6227 12257 6239 12260
rect 6181 12251 6239 12257
rect 6546 12248 6552 12260
rect 6604 12248 6610 12300
rect 10594 12248 10600 12300
rect 10652 12288 10658 12300
rect 12069 12291 12127 12297
rect 12069 12288 12081 12291
rect 10652 12260 12081 12288
rect 10652 12248 10658 12260
rect 12069 12257 12081 12260
rect 12115 12257 12127 12291
rect 12069 12251 12127 12257
rect 1854 12180 1860 12232
rect 1912 12220 1918 12232
rect 2406 12220 2412 12232
rect 1912 12192 2412 12220
rect 1912 12180 1918 12192
rect 2406 12180 2412 12192
rect 2464 12180 2470 12232
rect 4154 12220 4160 12232
rect 4115 12192 4160 12220
rect 4154 12180 4160 12192
rect 4212 12180 4218 12232
rect 4430 12220 4436 12232
rect 4391 12192 4436 12220
rect 4430 12180 4436 12192
rect 4488 12180 4494 12232
rect 7377 12223 7435 12229
rect 7377 12189 7389 12223
rect 7423 12189 7435 12223
rect 7377 12183 7435 12189
rect 9769 12223 9827 12229
rect 9769 12189 9781 12223
rect 9815 12220 9827 12223
rect 9950 12220 9956 12232
rect 9815 12192 9956 12220
rect 9815 12189 9827 12192
rect 9769 12183 9827 12189
rect 2038 12112 2044 12164
rect 2096 12152 2102 12164
rect 2225 12155 2283 12161
rect 2225 12152 2237 12155
rect 2096 12124 2237 12152
rect 2096 12112 2102 12124
rect 2225 12121 2237 12124
rect 2271 12121 2283 12155
rect 7392 12152 7420 12183
rect 9950 12180 9956 12192
rect 10008 12180 10014 12232
rect 10045 12223 10103 12229
rect 10045 12189 10057 12223
rect 10091 12189 10103 12223
rect 12084 12220 12112 12251
rect 12158 12248 12164 12300
rect 12216 12288 12222 12300
rect 12621 12291 12679 12297
rect 12621 12288 12633 12291
rect 12216 12260 12633 12288
rect 12216 12248 12222 12260
rect 12621 12257 12633 12260
rect 12667 12257 12679 12291
rect 13906 12288 13912 12300
rect 13867 12260 13912 12288
rect 12621 12251 12679 12257
rect 12250 12220 12256 12232
rect 12084 12192 12256 12220
rect 10045 12183 10103 12189
rect 8478 12152 8484 12164
rect 7392 12124 8484 12152
rect 2225 12115 2283 12121
rect 8478 12112 8484 12124
rect 8536 12112 8542 12164
rect 9030 12112 9036 12164
rect 9088 12152 9094 12164
rect 10060 12152 10088 12183
rect 12250 12180 12256 12192
rect 12308 12180 12314 12232
rect 12636 12220 12664 12251
rect 13906 12248 13912 12260
rect 13964 12248 13970 12300
rect 14185 12291 14243 12297
rect 14185 12257 14197 12291
rect 14231 12288 14243 12291
rect 14734 12288 14740 12300
rect 14231 12260 14740 12288
rect 14231 12257 14243 12260
rect 14185 12251 14243 12257
rect 14200 12220 14228 12251
rect 14734 12248 14740 12260
rect 14792 12248 14798 12300
rect 15672 12297 15700 12328
rect 15746 12316 15752 12368
rect 15804 12356 15810 12368
rect 15978 12359 16036 12365
rect 15978 12356 15990 12359
rect 15804 12328 15990 12356
rect 15804 12316 15810 12328
rect 15978 12325 15990 12328
rect 16024 12325 16036 12359
rect 15978 12319 16036 12325
rect 17402 12316 17408 12368
rect 17460 12356 17466 12368
rect 18156 12356 18184 12396
rect 18414 12384 18420 12396
rect 18472 12384 18478 12436
rect 18782 12424 18788 12436
rect 18743 12396 18788 12424
rect 18782 12384 18788 12396
rect 18840 12384 18846 12436
rect 20254 12424 20260 12436
rect 20215 12396 20260 12424
rect 20254 12384 20260 12396
rect 20312 12384 20318 12436
rect 20714 12424 20720 12436
rect 20675 12396 20720 12424
rect 20714 12384 20720 12396
rect 20772 12384 20778 12436
rect 21266 12384 21272 12436
rect 21324 12424 21330 12436
rect 22186 12424 22192 12436
rect 21324 12396 22192 12424
rect 21324 12384 21330 12396
rect 22186 12384 22192 12396
rect 22244 12424 22250 12436
rect 22244 12396 23428 12424
rect 22244 12384 22250 12396
rect 17460 12328 18184 12356
rect 18227 12359 18285 12365
rect 17460 12316 17466 12328
rect 18227 12325 18239 12359
rect 18273 12356 18285 12359
rect 18506 12356 18512 12368
rect 18273 12328 18512 12356
rect 18273 12325 18285 12328
rect 18227 12319 18285 12325
rect 18506 12316 18512 12328
rect 18564 12316 18570 12368
rect 18598 12316 18604 12368
rect 18656 12356 18662 12368
rect 19061 12359 19119 12365
rect 19061 12356 19073 12359
rect 18656 12328 19073 12356
rect 18656 12316 18662 12328
rect 19061 12325 19073 12328
rect 19107 12325 19119 12359
rect 19061 12319 19119 12325
rect 20806 12316 20812 12368
rect 20864 12356 20870 12368
rect 21361 12359 21419 12365
rect 21361 12356 21373 12359
rect 20864 12328 21373 12356
rect 20864 12316 20870 12328
rect 21361 12325 21373 12328
rect 21407 12325 21419 12359
rect 21361 12319 21419 12325
rect 22830 12316 22836 12368
rect 22888 12356 22894 12368
rect 22925 12359 22983 12365
rect 22925 12356 22937 12359
rect 22888 12328 22937 12356
rect 22888 12316 22894 12328
rect 22925 12325 22937 12328
rect 22971 12325 22983 12359
rect 23400 12356 23428 12396
rect 23477 12359 23535 12365
rect 23477 12356 23489 12359
rect 23400 12328 23489 12356
rect 22925 12319 22983 12325
rect 23477 12325 23489 12328
rect 23523 12325 23535 12359
rect 23477 12319 23535 12325
rect 23566 12316 23572 12368
rect 23624 12356 23630 12368
rect 24489 12359 24547 12365
rect 24489 12356 24501 12359
rect 23624 12328 24501 12356
rect 23624 12316 23630 12328
rect 24489 12325 24501 12328
rect 24535 12356 24547 12359
rect 24670 12356 24676 12368
rect 24535 12328 24676 12356
rect 24535 12325 24547 12328
rect 24489 12319 24547 12325
rect 24670 12316 24676 12328
rect 24728 12316 24734 12368
rect 15657 12291 15715 12297
rect 15657 12257 15669 12291
rect 15703 12257 15715 12291
rect 15657 12251 15715 12257
rect 16577 12291 16635 12297
rect 16577 12257 16589 12291
rect 16623 12288 16635 12291
rect 18046 12288 18052 12300
rect 16623 12260 18052 12288
rect 16623 12257 16635 12260
rect 16577 12251 16635 12257
rect 18046 12248 18052 12260
rect 18104 12248 18110 12300
rect 19886 12297 19892 12300
rect 19864 12291 19892 12297
rect 19864 12257 19876 12291
rect 19864 12251 19892 12257
rect 19886 12248 19892 12251
rect 19944 12248 19950 12300
rect 12636 12192 14228 12220
rect 14369 12223 14427 12229
rect 14369 12189 14381 12223
rect 14415 12220 14427 12223
rect 17865 12223 17923 12229
rect 17865 12220 17877 12223
rect 14415 12192 17877 12220
rect 14415 12189 14427 12192
rect 14369 12183 14427 12189
rect 17865 12189 17877 12192
rect 17911 12220 17923 12223
rect 18414 12220 18420 12232
rect 17911 12192 18420 12220
rect 17911 12189 17923 12192
rect 17865 12183 17923 12189
rect 18414 12180 18420 12192
rect 18472 12180 18478 12232
rect 20714 12180 20720 12232
rect 20772 12220 20778 12232
rect 21266 12220 21272 12232
rect 20772 12192 21272 12220
rect 20772 12180 20778 12192
rect 21266 12180 21272 12192
rect 21324 12180 21330 12232
rect 21542 12220 21548 12232
rect 21503 12192 21548 12220
rect 21542 12180 21548 12192
rect 21600 12180 21606 12232
rect 22833 12223 22891 12229
rect 22833 12220 22845 12223
rect 21744 12192 22845 12220
rect 9088 12124 10088 12152
rect 9088 12112 9094 12124
rect 11422 12112 11428 12164
rect 11480 12152 11486 12164
rect 11701 12155 11759 12161
rect 11701 12152 11713 12155
rect 11480 12124 11713 12152
rect 11480 12112 11486 12124
rect 11701 12121 11713 12124
rect 11747 12152 11759 12155
rect 12802 12152 12808 12164
rect 11747 12124 12808 12152
rect 11747 12121 11759 12124
rect 11701 12115 11759 12121
rect 12802 12112 12808 12124
rect 12860 12112 12866 12164
rect 19935 12155 19993 12161
rect 19935 12121 19947 12155
rect 19981 12152 19993 12155
rect 21744 12152 21772 12192
rect 22833 12189 22845 12192
rect 22879 12220 22891 12223
rect 22922 12220 22928 12232
rect 22879 12192 22928 12220
rect 22879 12189 22891 12192
rect 22833 12183 22891 12189
rect 22922 12180 22928 12192
rect 22980 12180 22986 12232
rect 24210 12180 24216 12232
rect 24268 12220 24274 12232
rect 24397 12223 24455 12229
rect 24397 12220 24409 12223
rect 24268 12192 24409 12220
rect 24268 12180 24274 12192
rect 24397 12189 24409 12192
rect 24443 12189 24455 12223
rect 24397 12183 24455 12189
rect 24673 12223 24731 12229
rect 24673 12189 24685 12223
rect 24719 12189 24731 12223
rect 24673 12183 24731 12189
rect 19981 12124 21772 12152
rect 19981 12121 19993 12124
rect 19935 12115 19993 12121
rect 23750 12112 23756 12164
rect 23808 12152 23814 12164
rect 23845 12155 23903 12161
rect 23845 12152 23857 12155
rect 23808 12124 23857 12152
rect 23808 12112 23814 12124
rect 23845 12121 23857 12124
rect 23891 12152 23903 12155
rect 24688 12152 24716 12183
rect 23891 12124 24716 12152
rect 23891 12121 23903 12124
rect 23845 12115 23903 12121
rect 1673 12087 1731 12093
rect 1673 12084 1685 12087
rect 1452 12056 1685 12084
rect 1452 12044 1458 12056
rect 1673 12053 1685 12056
rect 1719 12053 1731 12087
rect 5350 12084 5356 12096
rect 5311 12056 5356 12084
rect 1673 12047 1731 12053
rect 5350 12044 5356 12056
rect 5408 12044 5414 12096
rect 6546 12044 6552 12096
rect 6604 12084 6610 12096
rect 6825 12087 6883 12093
rect 6825 12084 6837 12087
rect 6604 12056 6837 12084
rect 6604 12044 6610 12056
rect 6825 12053 6837 12056
rect 6871 12084 6883 12087
rect 7558 12084 7564 12096
rect 6871 12056 7564 12084
rect 6871 12053 6883 12056
rect 6825 12047 6883 12053
rect 7558 12044 7564 12056
rect 7616 12044 7622 12096
rect 9309 12087 9367 12093
rect 9309 12053 9321 12087
rect 9355 12084 9367 12087
rect 9582 12084 9588 12096
rect 9355 12056 9588 12084
rect 9355 12053 9367 12056
rect 9309 12047 9367 12053
rect 9582 12044 9588 12056
rect 9640 12044 9646 12096
rect 12250 12044 12256 12096
rect 12308 12084 12314 12096
rect 13081 12087 13139 12093
rect 13081 12084 13093 12087
rect 12308 12056 13093 12084
rect 12308 12044 12314 12056
rect 13081 12053 13093 12056
rect 13127 12053 13139 12087
rect 13081 12047 13139 12053
rect 13170 12044 13176 12096
rect 13228 12084 13234 12096
rect 13538 12084 13544 12096
rect 13228 12056 13544 12084
rect 13228 12044 13234 12056
rect 13538 12044 13544 12056
rect 13596 12044 13602 12096
rect 14737 12087 14795 12093
rect 14737 12053 14749 12087
rect 14783 12084 14795 12087
rect 14826 12084 14832 12096
rect 14783 12056 14832 12084
rect 14783 12053 14795 12056
rect 14737 12047 14795 12053
rect 14826 12044 14832 12056
rect 14884 12044 14890 12096
rect 16758 12044 16764 12096
rect 16816 12084 16822 12096
rect 16853 12087 16911 12093
rect 16853 12084 16865 12087
rect 16816 12056 16865 12084
rect 16816 12044 16822 12056
rect 16853 12053 16865 12056
rect 16899 12053 16911 12087
rect 16853 12047 16911 12053
rect 21910 12044 21916 12096
rect 21968 12084 21974 12096
rect 22281 12087 22339 12093
rect 22281 12084 22293 12087
rect 21968 12056 22293 12084
rect 21968 12044 21974 12056
rect 22281 12053 22293 12056
rect 22327 12084 22339 12087
rect 23658 12084 23664 12096
rect 22327 12056 23664 12084
rect 22327 12053 22339 12056
rect 22281 12047 22339 12053
rect 23658 12044 23664 12056
rect 23716 12044 23722 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 4433 11883 4491 11889
rect 4433 11849 4445 11883
rect 4479 11880 4491 11883
rect 4614 11880 4620 11892
rect 4479 11852 4620 11880
rect 4479 11849 4491 11852
rect 4433 11843 4491 11849
rect 4614 11840 4620 11852
rect 4672 11880 4678 11892
rect 6549 11883 6607 11889
rect 6549 11880 6561 11883
rect 4672 11852 6561 11880
rect 4672 11840 4678 11852
rect 6549 11849 6561 11852
rect 6595 11849 6607 11883
rect 8846 11880 8852 11892
rect 8807 11852 8852 11880
rect 6549 11843 6607 11849
rect 4065 11815 4123 11821
rect 4065 11781 4077 11815
rect 4111 11812 4123 11815
rect 4246 11812 4252 11824
rect 4111 11784 4252 11812
rect 4111 11781 4123 11784
rect 4065 11775 4123 11781
rect 4246 11772 4252 11784
rect 4304 11812 4310 11824
rect 5445 11815 5503 11821
rect 5445 11812 5457 11815
rect 4304 11784 5457 11812
rect 4304 11772 4310 11784
rect 5445 11781 5457 11784
rect 5491 11781 5503 11815
rect 6564 11812 6592 11843
rect 8846 11840 8852 11852
rect 8904 11840 8910 11892
rect 9674 11840 9680 11892
rect 9732 11880 9738 11892
rect 10229 11883 10287 11889
rect 10229 11880 10241 11883
rect 9732 11852 10241 11880
rect 9732 11840 9738 11852
rect 10229 11849 10241 11852
rect 10275 11849 10287 11883
rect 10229 11843 10287 11849
rect 10594 11840 10600 11892
rect 10652 11880 10658 11892
rect 10781 11883 10839 11889
rect 10781 11880 10793 11883
rect 10652 11852 10793 11880
rect 10652 11840 10658 11852
rect 10781 11849 10793 11852
rect 10827 11849 10839 11883
rect 10781 11843 10839 11849
rect 11517 11883 11575 11889
rect 11517 11849 11529 11883
rect 11563 11880 11575 11883
rect 11974 11880 11980 11892
rect 11563 11852 11980 11880
rect 11563 11849 11575 11852
rect 11517 11843 11575 11849
rect 11974 11840 11980 11852
rect 12032 11840 12038 11892
rect 12710 11880 12716 11892
rect 12671 11852 12716 11880
rect 12710 11840 12716 11852
rect 12768 11840 12774 11892
rect 16853 11883 16911 11889
rect 16853 11849 16865 11883
rect 16899 11880 16911 11883
rect 17310 11880 17316 11892
rect 16899 11852 17316 11880
rect 16899 11849 16911 11852
rect 16853 11843 16911 11849
rect 17310 11840 17316 11852
rect 17368 11840 17374 11892
rect 19797 11883 19855 11889
rect 19797 11849 19809 11883
rect 19843 11880 19855 11883
rect 19886 11880 19892 11892
rect 19843 11852 19892 11880
rect 19843 11849 19855 11852
rect 19797 11843 19855 11849
rect 19886 11840 19892 11852
rect 19944 11880 19950 11892
rect 21082 11880 21088 11892
rect 19944 11852 21088 11880
rect 19944 11840 19950 11852
rect 21082 11840 21088 11852
rect 21140 11840 21146 11892
rect 22830 11840 22836 11892
rect 22888 11880 22894 11892
rect 23017 11883 23075 11889
rect 23017 11880 23029 11883
rect 22888 11852 23029 11880
rect 22888 11840 22894 11852
rect 23017 11849 23029 11852
rect 23063 11880 23075 11883
rect 23566 11880 23572 11892
rect 23063 11852 23572 11880
rect 23063 11849 23075 11852
rect 23017 11843 23075 11849
rect 23566 11840 23572 11852
rect 23624 11840 23630 11892
rect 24670 11880 24676 11892
rect 24631 11852 24676 11880
rect 24670 11840 24676 11852
rect 24728 11840 24734 11892
rect 25406 11880 25412 11892
rect 25367 11852 25412 11880
rect 25406 11840 25412 11852
rect 25464 11840 25470 11892
rect 6730 11812 6736 11824
rect 6564 11784 6736 11812
rect 5445 11775 5503 11781
rect 6730 11772 6736 11784
rect 6788 11812 6794 11824
rect 9125 11815 9183 11821
rect 9125 11812 9137 11815
rect 6788 11784 9137 11812
rect 6788 11772 6794 11784
rect 1762 11704 1768 11756
rect 1820 11744 1826 11756
rect 2406 11744 2412 11756
rect 1820 11716 2412 11744
rect 1820 11704 1826 11716
rect 2406 11704 2412 11716
rect 2464 11704 2470 11756
rect 2774 11704 2780 11756
rect 2832 11744 2838 11756
rect 3050 11744 3056 11756
rect 2832 11716 3056 11744
rect 2832 11704 2838 11716
rect 3050 11704 3056 11716
rect 3108 11704 3114 11756
rect 3697 11747 3755 11753
rect 3697 11713 3709 11747
rect 3743 11744 3755 11747
rect 4522 11744 4528 11756
rect 3743 11716 4528 11744
rect 3743 11713 3755 11716
rect 3697 11707 3755 11713
rect 4522 11704 4528 11716
rect 4580 11704 4586 11756
rect 5813 11679 5871 11685
rect 5813 11645 5825 11679
rect 5859 11676 5871 11679
rect 6546 11676 6552 11688
rect 5859 11648 6552 11676
rect 5859 11645 5871 11648
rect 5813 11639 5871 11645
rect 6546 11636 6552 11648
rect 6604 11636 6610 11688
rect 6822 11676 6828 11688
rect 6783 11648 6828 11676
rect 6822 11636 6828 11648
rect 6880 11636 6886 11688
rect 7116 11676 7144 11784
rect 9125 11781 9137 11784
rect 9171 11781 9183 11815
rect 9125 11775 9183 11781
rect 11241 11815 11299 11821
rect 11241 11781 11253 11815
rect 11287 11812 11299 11815
rect 12158 11812 12164 11824
rect 11287 11784 12164 11812
rect 11287 11781 11299 11784
rect 11241 11775 11299 11781
rect 7190 11704 7196 11756
rect 7248 11744 7254 11756
rect 8021 11747 8079 11753
rect 8021 11744 8033 11747
rect 7248 11716 8033 11744
rect 7248 11704 7254 11716
rect 8021 11713 8033 11716
rect 8067 11713 8079 11747
rect 8021 11707 8079 11713
rect 7116 11648 7190 11676
rect 2225 11611 2283 11617
rect 2225 11577 2237 11611
rect 2271 11608 2283 11611
rect 2498 11608 2504 11620
rect 2271 11580 2504 11608
rect 2271 11577 2283 11580
rect 2225 11571 2283 11577
rect 2498 11568 2504 11580
rect 2556 11568 2562 11620
rect 4614 11568 4620 11620
rect 4672 11608 4678 11620
rect 7162 11617 7190 11648
rect 4846 11611 4904 11617
rect 4846 11608 4858 11611
rect 4672 11580 4858 11608
rect 4672 11568 4678 11580
rect 4846 11577 4858 11580
rect 4892 11577 4904 11611
rect 4846 11571 4904 11577
rect 7147 11611 7205 11617
rect 7147 11577 7159 11611
rect 7193 11577 7205 11611
rect 7147 11571 7205 11577
rect 1857 11543 1915 11549
rect 1857 11509 1869 11543
rect 1903 11540 1915 11543
rect 2038 11540 2044 11552
rect 1903 11512 2044 11540
rect 1903 11509 1915 11512
rect 1857 11503 1915 11509
rect 2038 11500 2044 11512
rect 2096 11500 2102 11552
rect 2774 11500 2780 11552
rect 2832 11540 2838 11552
rect 5994 11540 6000 11552
rect 2832 11512 6000 11540
rect 2832 11500 2838 11512
rect 5994 11500 6000 11512
rect 6052 11540 6058 11552
rect 6089 11543 6147 11549
rect 6089 11540 6101 11543
rect 6052 11512 6101 11540
rect 6052 11500 6058 11512
rect 6089 11509 6101 11512
rect 6135 11509 6147 11543
rect 6089 11503 6147 11509
rect 7558 11500 7564 11552
rect 7616 11540 7622 11552
rect 7745 11543 7803 11549
rect 7745 11540 7757 11543
rect 7616 11512 7757 11540
rect 7616 11500 7622 11512
rect 7745 11509 7757 11512
rect 7791 11509 7803 11543
rect 8478 11540 8484 11552
rect 8439 11512 8484 11540
rect 7745 11503 7803 11509
rect 8478 11500 8484 11512
rect 8536 11500 8542 11552
rect 9140 11540 9168 11775
rect 12158 11772 12164 11784
rect 12216 11772 12222 11824
rect 17402 11812 17408 11824
rect 17363 11784 17408 11812
rect 17402 11772 17408 11784
rect 17460 11772 17466 11824
rect 17865 11815 17923 11821
rect 17865 11781 17877 11815
rect 17911 11812 17923 11815
rect 19426 11812 19432 11824
rect 17911 11784 19432 11812
rect 17911 11781 17923 11784
rect 17865 11775 17923 11781
rect 9309 11747 9367 11753
rect 9309 11713 9321 11747
rect 9355 11744 9367 11747
rect 9582 11744 9588 11756
rect 9355 11716 9588 11744
rect 9355 11713 9367 11716
rect 9309 11707 9367 11713
rect 9582 11704 9588 11716
rect 9640 11704 9646 11756
rect 12802 11744 12808 11756
rect 12763 11716 12808 11744
rect 12802 11704 12808 11716
rect 12860 11704 12866 11756
rect 11330 11676 11336 11688
rect 11291 11648 11336 11676
rect 11330 11636 11336 11648
rect 11388 11676 11394 11688
rect 11793 11679 11851 11685
rect 11793 11676 11805 11679
rect 11388 11648 11805 11676
rect 11388 11636 11394 11648
rect 11793 11645 11805 11648
rect 11839 11645 11851 11679
rect 11793 11639 11851 11645
rect 12584 11679 12642 11685
rect 12584 11645 12596 11679
rect 12630 11676 12642 11679
rect 14642 11676 14648 11688
rect 12630 11648 13584 11676
rect 14603 11648 14648 11676
rect 12630 11645 12642 11648
rect 12584 11639 12642 11645
rect 9671 11611 9729 11617
rect 9671 11577 9683 11611
rect 9717 11577 9729 11611
rect 9671 11571 9729 11577
rect 9692 11540 9720 11571
rect 12250 11568 12256 11620
rect 12308 11608 12314 11620
rect 12437 11611 12495 11617
rect 12437 11608 12449 11611
rect 12308 11580 12449 11608
rect 12308 11568 12314 11580
rect 12437 11577 12449 11580
rect 12483 11577 12495 11611
rect 12437 11571 12495 11577
rect 10042 11540 10048 11552
rect 9140 11512 10048 11540
rect 10042 11500 10048 11512
rect 10100 11500 10106 11552
rect 11698 11500 11704 11552
rect 11756 11540 11762 11552
rect 11974 11540 11980 11552
rect 11756 11512 11980 11540
rect 11756 11500 11762 11512
rect 11974 11500 11980 11512
rect 12032 11540 12038 11552
rect 12161 11543 12219 11549
rect 12161 11540 12173 11543
rect 12032 11512 12173 11540
rect 12032 11500 12038 11512
rect 12161 11509 12173 11512
rect 12207 11509 12219 11543
rect 12161 11503 12219 11509
rect 12342 11500 12348 11552
rect 12400 11540 12406 11552
rect 13556 11549 13584 11648
rect 14642 11636 14648 11648
rect 14700 11636 14706 11688
rect 14918 11676 14924 11688
rect 14879 11648 14924 11676
rect 14918 11636 14924 11648
rect 14976 11636 14982 11688
rect 15105 11679 15163 11685
rect 15105 11645 15117 11679
rect 15151 11676 15163 11679
rect 15930 11676 15936 11688
rect 15151 11648 15936 11676
rect 15151 11645 15163 11648
rect 15105 11639 15163 11645
rect 15930 11636 15936 11648
rect 15988 11636 15994 11688
rect 17880 11676 17908 11775
rect 19426 11772 19432 11784
rect 19484 11772 19490 11824
rect 23474 11772 23480 11824
rect 23532 11812 23538 11824
rect 24210 11812 24216 11824
rect 23532 11784 24216 11812
rect 23532 11772 23538 11784
rect 24210 11772 24216 11784
rect 24268 11812 24274 11824
rect 25041 11815 25099 11821
rect 25041 11812 25053 11815
rect 24268 11784 25053 11812
rect 24268 11772 24274 11784
rect 25041 11781 25053 11784
rect 25087 11781 25099 11815
rect 25041 11775 25099 11781
rect 18874 11744 18880 11756
rect 18340 11716 18880 11744
rect 17328 11648 17908 11676
rect 13909 11611 13967 11617
rect 13909 11577 13921 11611
rect 13955 11608 13967 11611
rect 14277 11611 14335 11617
rect 14277 11608 14289 11611
rect 13955 11580 14289 11608
rect 13955 11577 13967 11580
rect 13909 11571 13967 11577
rect 14277 11577 14289 11580
rect 14323 11608 14335 11611
rect 14936 11608 14964 11636
rect 14323 11580 14964 11608
rect 15473 11611 15531 11617
rect 14323 11577 14335 11580
rect 14277 11571 14335 11577
rect 15473 11577 15485 11611
rect 15519 11608 15531 11611
rect 15746 11608 15752 11620
rect 15519 11580 15752 11608
rect 15519 11577 15531 11580
rect 15473 11571 15531 11577
rect 15746 11568 15752 11580
rect 15804 11608 15810 11620
rect 15841 11611 15899 11617
rect 15841 11608 15853 11611
rect 15804 11580 15853 11608
rect 15804 11568 15810 11580
rect 15841 11577 15853 11580
rect 15887 11608 15899 11611
rect 16295 11611 16353 11617
rect 16295 11608 16307 11611
rect 15887 11580 16307 11608
rect 15887 11577 15899 11580
rect 15841 11571 15899 11577
rect 16295 11577 16307 11580
rect 16341 11608 16353 11611
rect 17328 11608 17356 11648
rect 18138 11636 18144 11688
rect 18196 11676 18202 11688
rect 18340 11685 18368 11716
rect 18874 11704 18880 11716
rect 18932 11704 18938 11756
rect 21637 11747 21695 11753
rect 21637 11744 21649 11747
rect 20824 11716 21649 11744
rect 18325 11679 18383 11685
rect 18325 11676 18337 11679
rect 18196 11648 18337 11676
rect 18196 11636 18202 11648
rect 18325 11645 18337 11648
rect 18371 11645 18383 11679
rect 18325 11639 18383 11645
rect 18509 11679 18567 11685
rect 18509 11645 18521 11679
rect 18555 11645 18567 11679
rect 19889 11679 19947 11685
rect 19889 11676 19901 11679
rect 18509 11639 18567 11645
rect 19352 11648 19901 11676
rect 16341 11580 17356 11608
rect 16341 11577 16353 11580
rect 16295 11571 16353 11577
rect 17402 11568 17408 11620
rect 17460 11608 17466 11620
rect 18524 11608 18552 11639
rect 17460 11580 18552 11608
rect 17460 11568 17466 11580
rect 19352 11552 19380 11648
rect 19889 11645 19901 11648
rect 19935 11645 19947 11679
rect 19889 11639 19947 11645
rect 20070 11568 20076 11620
rect 20128 11608 20134 11620
rect 20210 11611 20268 11617
rect 20210 11608 20222 11611
rect 20128 11580 20222 11608
rect 20128 11568 20134 11580
rect 20210 11577 20222 11580
rect 20256 11608 20268 11611
rect 20824 11608 20852 11716
rect 21637 11713 21649 11716
rect 21683 11744 21695 11747
rect 21726 11744 21732 11756
rect 21683 11716 21732 11744
rect 21683 11713 21695 11716
rect 21637 11707 21695 11713
rect 21726 11704 21732 11716
rect 21784 11744 21790 11756
rect 23750 11744 23756 11756
rect 21784 11716 22185 11744
rect 23711 11716 23756 11744
rect 21784 11704 21790 11716
rect 21821 11679 21879 11685
rect 21821 11676 21833 11679
rect 20256 11580 20852 11608
rect 21284 11648 21833 11676
rect 20256 11577 20268 11580
rect 20210 11571 20268 11577
rect 21284 11552 21312 11648
rect 21821 11645 21833 11648
rect 21867 11645 21879 11679
rect 21821 11639 21879 11645
rect 22157 11617 22185 11716
rect 23750 11704 23756 11716
rect 23808 11704 23814 11756
rect 24026 11744 24032 11756
rect 23987 11716 24032 11744
rect 24026 11704 24032 11716
rect 24084 11704 24090 11756
rect 22741 11679 22799 11685
rect 22741 11645 22753 11679
rect 22787 11676 22799 11679
rect 23385 11679 23443 11685
rect 23385 11676 23397 11679
rect 22787 11648 23397 11676
rect 22787 11645 22799 11648
rect 22741 11639 22799 11645
rect 23385 11645 23397 11648
rect 23431 11645 23443 11679
rect 23385 11639 23443 11645
rect 22142 11611 22200 11617
rect 22142 11577 22154 11611
rect 22188 11577 22200 11611
rect 22142 11571 22200 11577
rect 13081 11543 13139 11549
rect 13081 11540 13093 11543
rect 12400 11512 13093 11540
rect 12400 11500 12406 11512
rect 13081 11509 13093 11512
rect 13127 11509 13139 11543
rect 13081 11503 13139 11509
rect 13541 11543 13599 11549
rect 13541 11509 13553 11543
rect 13587 11540 13599 11543
rect 13630 11540 13636 11552
rect 13587 11512 13636 11540
rect 13587 11509 13599 11512
rect 13541 11503 13599 11509
rect 13630 11500 13636 11512
rect 13688 11500 13694 11552
rect 18322 11540 18328 11552
rect 18283 11512 18328 11540
rect 18322 11500 18328 11512
rect 18380 11500 18386 11552
rect 19334 11540 19340 11552
rect 19295 11512 19340 11540
rect 19334 11500 19340 11512
rect 19392 11500 19398 11552
rect 20806 11540 20812 11552
rect 20767 11512 20812 11540
rect 20806 11500 20812 11512
rect 20864 11500 20870 11552
rect 21266 11540 21272 11552
rect 21227 11512 21272 11540
rect 21266 11500 21272 11512
rect 21324 11500 21330 11552
rect 23400 11540 23428 11639
rect 24854 11636 24860 11688
rect 24912 11676 24918 11688
rect 25225 11679 25283 11685
rect 25225 11676 25237 11679
rect 24912 11648 25237 11676
rect 24912 11636 24918 11648
rect 25225 11645 25237 11648
rect 25271 11676 25283 11679
rect 25777 11679 25835 11685
rect 25777 11676 25789 11679
rect 25271 11648 25789 11676
rect 25271 11645 25283 11648
rect 25225 11639 25283 11645
rect 25777 11645 25789 11648
rect 25823 11645 25835 11679
rect 25777 11639 25835 11645
rect 23845 11611 23903 11617
rect 23845 11577 23857 11611
rect 23891 11577 23903 11611
rect 23845 11571 23903 11577
rect 23860 11540 23888 11571
rect 23400 11512 23888 11540
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1854 11336 1860 11348
rect 1815 11308 1860 11336
rect 1854 11296 1860 11308
rect 1912 11296 1918 11348
rect 2406 11296 2412 11348
rect 2464 11336 2470 11348
rect 2961 11339 3019 11345
rect 2961 11336 2973 11339
rect 2464 11308 2973 11336
rect 2464 11296 2470 11308
rect 2961 11305 2973 11308
rect 3007 11305 3019 11339
rect 2961 11299 3019 11305
rect 3881 11339 3939 11345
rect 3881 11305 3893 11339
rect 3927 11336 3939 11339
rect 4154 11336 4160 11348
rect 3927 11308 4160 11336
rect 3927 11305 3939 11308
rect 3881 11299 3939 11305
rect 2038 11228 2044 11280
rect 2096 11268 2102 11280
rect 2133 11271 2191 11277
rect 2133 11268 2145 11271
rect 2096 11240 2145 11268
rect 2096 11228 2102 11240
rect 2133 11237 2145 11240
rect 2179 11237 2191 11271
rect 2133 11231 2191 11237
rect 1578 11092 1584 11144
rect 1636 11132 1642 11144
rect 2041 11135 2099 11141
rect 2041 11132 2053 11135
rect 1636 11104 2053 11132
rect 1636 11092 1642 11104
rect 2041 11101 2053 11104
rect 2087 11101 2099 11135
rect 2498 11132 2504 11144
rect 2459 11104 2504 11132
rect 2041 11095 2099 11101
rect 2056 11064 2084 11095
rect 2498 11092 2504 11104
rect 2556 11132 2562 11144
rect 3896 11132 3924 11299
rect 4154 11296 4160 11308
rect 4212 11296 4218 11348
rect 4338 11296 4344 11348
rect 4396 11336 4402 11348
rect 5445 11339 5503 11345
rect 5445 11336 5457 11339
rect 4396 11308 5457 11336
rect 4396 11296 4402 11308
rect 5445 11305 5457 11308
rect 5491 11305 5503 11339
rect 5445 11299 5503 11305
rect 7190 11296 7196 11348
rect 7248 11336 7254 11348
rect 7377 11339 7435 11345
rect 7377 11336 7389 11339
rect 7248 11308 7389 11336
rect 7248 11296 7254 11308
rect 7377 11305 7389 11308
rect 7423 11305 7435 11339
rect 7377 11299 7435 11305
rect 10134 11296 10140 11348
rect 10192 11336 10198 11348
rect 10597 11339 10655 11345
rect 10597 11336 10609 11339
rect 10192 11308 10609 11336
rect 10192 11296 10198 11308
rect 10597 11305 10609 11308
rect 10643 11305 10655 11339
rect 10597 11299 10655 11305
rect 11974 11296 11980 11348
rect 12032 11336 12038 11348
rect 12710 11336 12716 11348
rect 12032 11308 12716 11336
rect 12032 11296 12038 11308
rect 12710 11296 12716 11308
rect 12768 11296 12774 11348
rect 13906 11296 13912 11348
rect 13964 11336 13970 11348
rect 14369 11339 14427 11345
rect 14369 11336 14381 11339
rect 13964 11308 14381 11336
rect 13964 11296 13970 11308
rect 14369 11305 14381 11308
rect 14415 11305 14427 11339
rect 14369 11299 14427 11305
rect 14642 11296 14648 11348
rect 14700 11336 14706 11348
rect 14737 11339 14795 11345
rect 14737 11336 14749 11339
rect 14700 11308 14749 11336
rect 14700 11296 14706 11308
rect 14737 11305 14749 11308
rect 14783 11305 14795 11339
rect 14737 11299 14795 11305
rect 15930 11296 15936 11348
rect 15988 11336 15994 11348
rect 16669 11339 16727 11345
rect 16669 11336 16681 11339
rect 15988 11308 16681 11336
rect 15988 11296 15994 11308
rect 16669 11305 16681 11308
rect 16715 11305 16727 11339
rect 17494 11336 17500 11348
rect 17455 11308 17500 11336
rect 16669 11299 16727 11305
rect 17494 11296 17500 11308
rect 17552 11296 17558 11348
rect 18138 11336 18144 11348
rect 18099 11308 18144 11336
rect 18138 11296 18144 11308
rect 18196 11296 18202 11348
rect 18414 11336 18420 11348
rect 18375 11308 18420 11336
rect 18414 11296 18420 11308
rect 18472 11296 18478 11348
rect 20714 11336 20720 11348
rect 20675 11308 20720 11336
rect 20714 11296 20720 11308
rect 20772 11296 20778 11348
rect 20806 11296 20812 11348
rect 20864 11336 20870 11348
rect 21913 11339 21971 11345
rect 21913 11336 21925 11339
rect 20864 11308 21925 11336
rect 20864 11296 20870 11308
rect 21913 11305 21925 11308
rect 21959 11305 21971 11339
rect 21913 11299 21971 11305
rect 22603 11339 22661 11345
rect 22603 11305 22615 11339
rect 22649 11336 22661 11339
rect 25222 11336 25228 11348
rect 22649 11308 25084 11336
rect 25183 11308 25228 11336
rect 22649 11305 22661 11308
rect 22603 11299 22661 11305
rect 4614 11228 4620 11280
rect 4672 11268 4678 11280
rect 4846 11271 4904 11277
rect 4846 11268 4858 11271
rect 4672 11240 4858 11268
rect 4672 11228 4678 11240
rect 4846 11237 4858 11240
rect 4892 11237 4904 11271
rect 4846 11231 4904 11237
rect 6730 11228 6736 11280
rect 6788 11277 6794 11280
rect 6788 11271 6836 11277
rect 6788 11237 6790 11271
rect 6824 11237 6836 11271
rect 8754 11268 8760 11280
rect 8715 11240 8760 11268
rect 6788 11231 6836 11237
rect 6788 11228 6794 11231
rect 8754 11228 8760 11240
rect 8812 11228 8818 11280
rect 10042 11277 10048 11280
rect 10039 11268 10048 11277
rect 10003 11240 10048 11268
rect 10039 11231 10048 11240
rect 10042 11228 10048 11231
rect 10100 11228 10106 11280
rect 11793 11271 11851 11277
rect 11793 11237 11805 11271
rect 11839 11268 11851 11271
rect 12158 11268 12164 11280
rect 11839 11240 12164 11268
rect 11839 11237 11851 11240
rect 11793 11231 11851 11237
rect 12158 11228 12164 11240
rect 12216 11228 12222 11280
rect 12250 11228 12256 11280
rect 12308 11268 12314 11280
rect 13814 11268 13820 11280
rect 12308 11240 13820 11268
rect 12308 11228 12314 11240
rect 6546 11160 6552 11212
rect 6604 11200 6610 11212
rect 8202 11200 8208 11212
rect 6604 11172 7788 11200
rect 8163 11172 8208 11200
rect 6604 11160 6610 11172
rect 2556 11104 3924 11132
rect 4525 11135 4583 11141
rect 2556 11092 2562 11104
rect 4525 11101 4537 11135
rect 4571 11132 4583 11135
rect 6457 11135 6515 11141
rect 4571 11104 4605 11132
rect 4571 11101 4583 11104
rect 4525 11095 4583 11101
rect 6457 11101 6469 11135
rect 6503 11132 6515 11135
rect 6503 11104 6868 11132
rect 6503 11101 6515 11104
rect 6457 11095 6515 11101
rect 3329 11067 3387 11073
rect 3329 11064 3341 11067
rect 2056 11036 3341 11064
rect 3329 11033 3341 11036
rect 3375 11033 3387 11067
rect 3329 11027 3387 11033
rect 4433 11067 4491 11073
rect 4433 11033 4445 11067
rect 4479 11064 4491 11067
rect 4540 11064 4568 11095
rect 4479 11036 5580 11064
rect 4479 11033 4491 11036
rect 4433 11027 4491 11033
rect 5552 11008 5580 11036
rect 5534 10956 5540 11008
rect 5592 10956 5598 11008
rect 6840 10996 6868 11104
rect 6914 11092 6920 11144
rect 6972 11132 6978 11144
rect 7653 11135 7711 11141
rect 7653 11132 7665 11135
rect 6972 11104 7665 11132
rect 6972 11092 6978 11104
rect 7653 11101 7665 11104
rect 7699 11101 7711 11135
rect 7760 11132 7788 11172
rect 8202 11160 8208 11172
rect 8260 11160 8266 11212
rect 8389 11203 8447 11209
rect 8389 11169 8401 11203
rect 8435 11200 8447 11203
rect 8570 11200 8576 11212
rect 8435 11172 8576 11200
rect 8435 11169 8447 11172
rect 8389 11163 8447 11169
rect 8570 11160 8576 11172
rect 8628 11200 8634 11212
rect 11606 11200 11612 11212
rect 8628 11172 11612 11200
rect 8628 11160 8634 11172
rect 11606 11160 11612 11172
rect 11664 11160 11670 11212
rect 11974 11160 11980 11212
rect 12032 11209 12038 11212
rect 12032 11203 12081 11209
rect 12032 11169 12035 11203
rect 12069 11169 12081 11203
rect 12176 11200 12204 11228
rect 13173 11203 13231 11209
rect 13173 11200 13185 11203
rect 12176 11172 13185 11200
rect 12032 11163 12081 11169
rect 13173 11169 13185 11172
rect 13219 11169 13231 11203
rect 13173 11163 13231 11169
rect 13357 11203 13415 11209
rect 13357 11169 13369 11203
rect 13403 11200 13415 11203
rect 13538 11200 13544 11212
rect 13403 11172 13544 11200
rect 13403 11169 13415 11172
rect 13357 11163 13415 11169
rect 12032 11160 12038 11163
rect 13538 11160 13544 11172
rect 13596 11160 13602 11212
rect 13648 11209 13676 11240
rect 13814 11228 13820 11240
rect 13872 11228 13878 11280
rect 15565 11271 15623 11277
rect 15565 11237 15577 11271
rect 15611 11268 15623 11271
rect 15841 11271 15899 11277
rect 15841 11268 15853 11271
rect 15611 11240 15853 11268
rect 15611 11237 15623 11240
rect 15565 11231 15623 11237
rect 15841 11237 15853 11240
rect 15887 11268 15899 11271
rect 16022 11268 16028 11280
rect 15887 11240 16028 11268
rect 15887 11237 15899 11240
rect 15841 11231 15899 11237
rect 16022 11228 16028 11240
rect 16080 11228 16086 11280
rect 19334 11268 19340 11280
rect 19295 11240 19340 11268
rect 19334 11228 19340 11240
rect 19392 11228 19398 11280
rect 21085 11271 21143 11277
rect 21085 11237 21097 11271
rect 21131 11268 21143 11271
rect 21450 11268 21456 11280
rect 21131 11240 21456 11268
rect 21131 11237 21143 11240
rect 21085 11231 21143 11237
rect 21450 11228 21456 11240
rect 21508 11228 21514 11280
rect 22922 11268 22928 11280
rect 22883 11240 22928 11268
rect 22922 11228 22928 11240
rect 22980 11228 22986 11280
rect 23658 11268 23664 11280
rect 23619 11240 23664 11268
rect 23658 11228 23664 11240
rect 23716 11228 23722 11280
rect 13633 11203 13691 11209
rect 13633 11169 13645 11203
rect 13679 11169 13691 11203
rect 13633 11163 13691 11169
rect 16850 11160 16856 11212
rect 16908 11200 16914 11212
rect 17221 11203 17279 11209
rect 17221 11200 17233 11203
rect 16908 11172 17233 11200
rect 16908 11160 16914 11172
rect 17221 11169 17233 11172
rect 17267 11169 17279 11203
rect 17402 11200 17408 11212
rect 17363 11172 17408 11200
rect 17221 11163 17279 11169
rect 17402 11160 17408 11172
rect 17460 11160 17466 11212
rect 17586 11160 17592 11212
rect 17644 11200 17650 11212
rect 18601 11203 18659 11209
rect 18601 11200 18613 11203
rect 17644 11172 18613 11200
rect 17644 11160 17650 11172
rect 18601 11169 18613 11172
rect 18647 11169 18659 11203
rect 19058 11200 19064 11212
rect 19019 11172 19064 11200
rect 18601 11163 18659 11169
rect 9674 11132 9680 11144
rect 7760 11104 9168 11132
rect 9635 11104 9680 11132
rect 7653 11095 7711 11101
rect 7098 10996 7104 11008
rect 6840 10968 7104 10996
rect 7098 10956 7104 10968
rect 7156 10956 7162 11008
rect 7466 10956 7472 11008
rect 7524 10996 7530 11008
rect 9140 11005 9168 11104
rect 9674 11092 9680 11104
rect 9732 11092 9738 11144
rect 11624 11132 11652 11160
rect 12161 11135 12219 11141
rect 12161 11132 12173 11135
rect 11624 11104 12173 11132
rect 12161 11101 12173 11104
rect 12207 11132 12219 11135
rect 12250 11132 12256 11144
rect 12207 11104 12256 11132
rect 12207 11101 12219 11104
rect 12161 11095 12219 11101
rect 12250 11092 12256 11104
rect 12308 11092 12314 11144
rect 12526 11132 12532 11144
rect 12487 11104 12532 11132
rect 12526 11092 12532 11104
rect 12584 11092 12590 11144
rect 12894 11092 12900 11144
rect 12952 11132 12958 11144
rect 13449 11135 13507 11141
rect 13449 11132 13461 11135
rect 12952 11104 13461 11132
rect 12952 11092 12958 11104
rect 13449 11101 13461 11104
rect 13495 11101 13507 11135
rect 13906 11132 13912 11144
rect 13867 11104 13912 11132
rect 13449 11095 13507 11101
rect 13906 11092 13912 11104
rect 13964 11092 13970 11144
rect 15749 11135 15807 11141
rect 15749 11101 15761 11135
rect 15795 11101 15807 11135
rect 16206 11132 16212 11144
rect 16167 11104 16212 11132
rect 15749 11095 15807 11101
rect 9493 11067 9551 11073
rect 9493 11033 9505 11067
rect 9539 11064 9551 11067
rect 9950 11064 9956 11076
rect 9539 11036 9956 11064
rect 9539 11033 9551 11036
rect 9493 11027 9551 11033
rect 9950 11024 9956 11036
rect 10008 11024 10014 11076
rect 10965 11067 11023 11073
rect 10965 11064 10977 11067
rect 10060 11036 10977 11064
rect 8021 10999 8079 11005
rect 8021 10996 8033 10999
rect 7524 10968 8033 10996
rect 7524 10956 7530 10968
rect 8021 10965 8033 10968
rect 8067 10965 8079 10999
rect 8021 10959 8079 10965
rect 9125 10999 9183 11005
rect 9125 10965 9137 10999
rect 9171 10996 9183 10999
rect 9398 10996 9404 11008
rect 9171 10968 9404 10996
rect 9171 10965 9183 10968
rect 9125 10959 9183 10965
rect 9398 10956 9404 10968
rect 9456 10996 9462 11008
rect 10060 10996 10088 11036
rect 10965 11033 10977 11036
rect 11011 11033 11023 11067
rect 15764 11064 15792 11095
rect 16206 11092 16212 11104
rect 16264 11092 16270 11144
rect 18616 11132 18644 11163
rect 19058 11160 19064 11172
rect 19116 11160 19122 11212
rect 21634 11160 21640 11212
rect 21692 11200 21698 11212
rect 22370 11200 22376 11212
rect 21692 11172 22376 11200
rect 21692 11160 21698 11172
rect 22370 11160 22376 11172
rect 22428 11200 22434 11212
rect 25056 11209 25084 11308
rect 25222 11296 25228 11308
rect 25280 11296 25286 11348
rect 22500 11203 22558 11209
rect 22500 11200 22512 11203
rect 22428 11172 22512 11200
rect 22428 11160 22434 11172
rect 22500 11169 22512 11172
rect 22546 11200 22558 11203
rect 25041 11203 25099 11209
rect 22546 11172 23152 11200
rect 22546 11169 22558 11172
rect 22500 11163 22558 11169
rect 19334 11132 19340 11144
rect 18616 11104 19340 11132
rect 19334 11092 19340 11104
rect 19392 11092 19398 11144
rect 20714 11092 20720 11144
rect 20772 11132 20778 11144
rect 20993 11135 21051 11141
rect 20993 11132 21005 11135
rect 20772 11104 21005 11132
rect 20772 11092 20778 11104
rect 20993 11101 21005 11104
rect 21039 11101 21051 11135
rect 20993 11095 21051 11101
rect 21174 11092 21180 11144
rect 21232 11132 21238 11144
rect 21269 11135 21327 11141
rect 21269 11132 21281 11135
rect 21232 11104 21281 11132
rect 21232 11092 21238 11104
rect 21269 11101 21281 11104
rect 21315 11101 21327 11135
rect 21269 11095 21327 11101
rect 16390 11064 16396 11076
rect 15764 11036 16396 11064
rect 10965 11027 11023 11033
rect 9456 10968 10088 10996
rect 10980 10996 11008 11027
rect 16390 11024 16396 11036
rect 16448 11024 16454 11076
rect 17037 11067 17095 11073
rect 17037 11064 17049 11067
rect 16500 11036 17049 11064
rect 11146 10996 11152 11008
rect 10980 10968 11152 10996
rect 9456 10956 9462 10968
rect 11146 10956 11152 10968
rect 11204 10956 11210 11008
rect 11882 10956 11888 11008
rect 11940 11005 11946 11008
rect 11940 10999 11989 11005
rect 11940 10965 11943 10999
rect 11977 10965 11989 10999
rect 11940 10959 11989 10965
rect 11940 10956 11946 10959
rect 12802 10956 12808 11008
rect 12860 10996 12866 11008
rect 12897 10999 12955 11005
rect 12897 10996 12909 10999
rect 12860 10968 12909 10996
rect 12860 10956 12866 10968
rect 12897 10965 12909 10968
rect 12943 10996 12955 10999
rect 15286 10996 15292 11008
rect 12943 10968 15292 10996
rect 12943 10965 12955 10968
rect 12897 10959 12955 10965
rect 15286 10956 15292 10968
rect 15344 10956 15350 11008
rect 15838 10956 15844 11008
rect 15896 10996 15902 11008
rect 16500 10996 16528 11036
rect 17037 11033 17049 11036
rect 17083 11033 17095 11067
rect 23124 11064 23152 11172
rect 25041 11169 25053 11203
rect 25087 11200 25099 11203
rect 25130 11200 25136 11212
rect 25087 11172 25136 11200
rect 25087 11169 25099 11172
rect 25041 11163 25099 11169
rect 25130 11160 25136 11172
rect 25188 11160 25194 11212
rect 23566 11132 23572 11144
rect 23527 11104 23572 11132
rect 23566 11092 23572 11104
rect 23624 11092 23630 11144
rect 23750 11092 23756 11144
rect 23808 11132 23814 11144
rect 23845 11135 23903 11141
rect 23845 11132 23857 11135
rect 23808 11104 23857 11132
rect 23808 11092 23814 11104
rect 23845 11101 23857 11104
rect 23891 11101 23903 11135
rect 23845 11095 23903 11101
rect 24026 11064 24032 11076
rect 23124 11036 24032 11064
rect 17037 11027 17095 11033
rect 24026 11024 24032 11036
rect 24084 11024 24090 11076
rect 15896 10968 16528 10996
rect 15896 10956 15902 10968
rect 19426 10956 19432 11008
rect 19484 10996 19490 11008
rect 19889 10999 19947 11005
rect 19889 10996 19901 10999
rect 19484 10968 19901 10996
rect 19484 10956 19490 10968
rect 19889 10965 19901 10968
rect 19935 10996 19947 10999
rect 20070 10996 20076 11008
rect 19935 10968 20076 10996
rect 19935 10965 19947 10968
rect 19889 10959 19947 10965
rect 20070 10956 20076 10968
rect 20128 10956 20134 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 4614 10792 4620 10804
rect 4575 10764 4620 10792
rect 4614 10752 4620 10764
rect 4672 10752 4678 10804
rect 6549 10795 6607 10801
rect 6549 10761 6561 10795
rect 6595 10792 6607 10795
rect 6730 10792 6736 10804
rect 6595 10764 6736 10792
rect 6595 10761 6607 10764
rect 6549 10755 6607 10761
rect 6730 10752 6736 10764
rect 6788 10752 6794 10804
rect 7098 10792 7104 10804
rect 7059 10764 7104 10792
rect 7098 10752 7104 10764
rect 7156 10752 7162 10804
rect 8294 10752 8300 10804
rect 8352 10792 8358 10804
rect 8389 10795 8447 10801
rect 8389 10792 8401 10795
rect 8352 10764 8401 10792
rect 8352 10752 8358 10764
rect 8389 10761 8401 10764
rect 8435 10761 8447 10795
rect 8389 10755 8447 10761
rect 1949 10727 2007 10733
rect 1949 10693 1961 10727
rect 1995 10724 2007 10727
rect 2038 10724 2044 10736
rect 1995 10696 2044 10724
rect 1995 10693 2007 10696
rect 1949 10687 2007 10693
rect 2038 10684 2044 10696
rect 2096 10684 2102 10736
rect 2682 10724 2688 10736
rect 2643 10696 2688 10724
rect 2682 10684 2688 10696
rect 2740 10684 2746 10736
rect 8018 10724 8024 10736
rect 7979 10696 8024 10724
rect 8018 10684 8024 10696
rect 8076 10684 8082 10736
rect 8404 10724 8432 10755
rect 8570 10752 8576 10804
rect 8628 10792 8634 10804
rect 8757 10795 8815 10801
rect 8757 10792 8769 10795
rect 8628 10764 8769 10792
rect 8628 10752 8634 10764
rect 8757 10761 8769 10764
rect 8803 10761 8815 10795
rect 8757 10755 8815 10761
rect 12713 10795 12771 10801
rect 12713 10761 12725 10795
rect 12759 10792 12771 10795
rect 12894 10792 12900 10804
rect 12759 10764 12900 10792
rect 12759 10761 12771 10764
rect 12713 10755 12771 10761
rect 12894 10752 12900 10764
rect 12952 10752 12958 10804
rect 13814 10792 13820 10804
rect 13775 10764 13820 10792
rect 13814 10752 13820 10764
rect 13872 10752 13878 10804
rect 15654 10792 15660 10804
rect 15615 10764 15660 10792
rect 15654 10752 15660 10764
rect 15712 10752 15718 10804
rect 16942 10752 16948 10804
rect 17000 10792 17006 10804
rect 17773 10795 17831 10801
rect 17773 10792 17785 10795
rect 17000 10764 17785 10792
rect 17000 10752 17006 10764
rect 17773 10761 17785 10764
rect 17819 10761 17831 10795
rect 17773 10755 17831 10761
rect 11974 10724 11980 10736
rect 8404 10696 11980 10724
rect 11974 10684 11980 10696
rect 12032 10684 12038 10736
rect 3145 10659 3203 10665
rect 3145 10625 3157 10659
rect 3191 10656 3203 10659
rect 3786 10656 3792 10668
rect 3191 10628 3792 10656
rect 3191 10625 3203 10628
rect 3145 10619 3203 10625
rect 2130 10520 2136 10532
rect 2091 10492 2136 10520
rect 2130 10480 2136 10492
rect 2188 10480 2194 10532
rect 2225 10523 2283 10529
rect 2225 10489 2237 10523
rect 2271 10520 2283 10523
rect 3160 10520 3188 10619
rect 3786 10616 3792 10628
rect 3844 10616 3850 10668
rect 4154 10656 4160 10668
rect 4115 10628 4160 10656
rect 4154 10616 4160 10628
rect 4212 10616 4218 10668
rect 5534 10616 5540 10668
rect 5592 10656 5598 10668
rect 5721 10659 5779 10665
rect 5721 10656 5733 10659
rect 5592 10628 5733 10656
rect 5592 10616 5598 10628
rect 5721 10625 5733 10628
rect 5767 10625 5779 10659
rect 9582 10656 9588 10668
rect 9543 10628 9588 10656
rect 5721 10619 5779 10625
rect 9582 10616 9588 10628
rect 9640 10616 9646 10668
rect 12253 10659 12311 10665
rect 12253 10625 12265 10659
rect 12299 10656 12311 10659
rect 12802 10656 12808 10668
rect 12299 10628 12808 10656
rect 12299 10625 12311 10628
rect 12253 10619 12311 10625
rect 12802 10616 12808 10628
rect 12860 10616 12866 10668
rect 15838 10656 15844 10668
rect 15799 10628 15844 10656
rect 15838 10616 15844 10628
rect 15896 10616 15902 10668
rect 16206 10656 16212 10668
rect 16167 10628 16212 10656
rect 16206 10616 16212 10628
rect 16264 10616 16270 10668
rect 5169 10591 5227 10597
rect 5169 10588 5181 10591
rect 5000 10560 5181 10588
rect 3697 10523 3755 10529
rect 3697 10520 3709 10523
rect 2271 10492 3188 10520
rect 3436 10492 3709 10520
rect 2271 10489 2283 10492
rect 2225 10483 2283 10489
rect 3436 10464 3464 10492
rect 3697 10489 3709 10492
rect 3743 10489 3755 10523
rect 3697 10483 3755 10489
rect 3786 10480 3792 10532
rect 3844 10520 3850 10532
rect 3844 10492 3889 10520
rect 3844 10480 3850 10492
rect 3418 10452 3424 10464
rect 3379 10424 3424 10452
rect 3418 10412 3424 10424
rect 3476 10412 3482 10464
rect 4798 10412 4804 10464
rect 4856 10452 4862 10464
rect 5000 10461 5028 10560
rect 5169 10557 5181 10560
rect 5215 10557 5227 10591
rect 5169 10551 5227 10557
rect 5258 10548 5264 10600
rect 5316 10588 5322 10600
rect 5629 10591 5687 10597
rect 5629 10588 5641 10591
rect 5316 10560 5641 10588
rect 5316 10548 5322 10560
rect 5629 10557 5641 10560
rect 5675 10588 5687 10591
rect 6546 10588 6552 10600
rect 5675 10560 6552 10588
rect 5675 10557 5687 10560
rect 5629 10551 5687 10557
rect 6546 10548 6552 10560
rect 6604 10548 6610 10600
rect 9214 10588 9220 10600
rect 9175 10560 9220 10588
rect 9214 10548 9220 10560
rect 9272 10548 9278 10600
rect 9398 10588 9404 10600
rect 9359 10560 9404 10588
rect 9398 10548 9404 10560
rect 9456 10548 9462 10600
rect 10413 10591 10471 10597
rect 10413 10557 10425 10591
rect 10459 10588 10471 10591
rect 10778 10588 10784 10600
rect 10459 10560 10784 10588
rect 10459 10557 10471 10560
rect 10413 10551 10471 10557
rect 10778 10548 10784 10560
rect 10836 10548 10842 10600
rect 11057 10591 11115 10597
rect 11057 10557 11069 10591
rect 11103 10588 11115 10591
rect 11146 10588 11152 10600
rect 11103 10560 11152 10588
rect 11103 10557 11115 10560
rect 11057 10551 11115 10557
rect 11146 10548 11152 10560
rect 11204 10548 11210 10600
rect 12584 10591 12642 10597
rect 12584 10557 12596 10591
rect 12630 10588 12642 10591
rect 13173 10591 13231 10597
rect 12630 10560 13124 10588
rect 12630 10557 12642 10560
rect 12584 10551 12642 10557
rect 7466 10520 7472 10532
rect 7427 10492 7472 10520
rect 7466 10480 7472 10492
rect 7524 10480 7530 10532
rect 7558 10480 7564 10532
rect 7616 10520 7622 10532
rect 7616 10492 7661 10520
rect 7616 10480 7622 10492
rect 9766 10480 9772 10532
rect 9824 10520 9830 10532
rect 9824 10492 10640 10520
rect 9824 10480 9830 10492
rect 4985 10455 5043 10461
rect 4985 10452 4997 10455
rect 4856 10424 4997 10452
rect 4856 10412 4862 10424
rect 4985 10421 4997 10424
rect 5031 10421 5043 10455
rect 10042 10452 10048 10464
rect 10003 10424 10048 10452
rect 4985 10415 5043 10421
rect 10042 10412 10048 10424
rect 10100 10412 10106 10464
rect 10612 10461 10640 10492
rect 12158 10480 12164 10532
rect 12216 10520 12222 10532
rect 12437 10523 12495 10529
rect 12437 10520 12449 10523
rect 12216 10492 12449 10520
rect 12216 10480 12222 10492
rect 12437 10489 12449 10492
rect 12483 10489 12495 10523
rect 13096 10520 13124 10560
rect 13173 10557 13185 10591
rect 13219 10588 13231 10591
rect 13814 10588 13820 10600
rect 13219 10560 13820 10588
rect 13219 10557 13231 10560
rect 13173 10551 13231 10557
rect 13814 10548 13820 10560
rect 13872 10548 13878 10600
rect 14274 10588 14280 10600
rect 14235 10560 14280 10588
rect 14274 10548 14280 10560
rect 14332 10548 14338 10600
rect 14737 10591 14795 10597
rect 14737 10557 14749 10591
rect 14783 10557 14795 10591
rect 17788 10588 17816 10755
rect 19334 10752 19340 10804
rect 19392 10792 19398 10804
rect 19521 10795 19579 10801
rect 19521 10792 19533 10795
rect 19392 10764 19533 10792
rect 19392 10752 19398 10764
rect 19521 10761 19533 10764
rect 19567 10761 19579 10795
rect 19521 10755 19579 10761
rect 20714 10752 20720 10804
rect 20772 10792 20778 10804
rect 21821 10795 21879 10801
rect 21821 10792 21833 10795
rect 20772 10764 21833 10792
rect 20772 10752 20778 10764
rect 21821 10761 21833 10764
rect 21867 10761 21879 10795
rect 22370 10792 22376 10804
rect 22331 10764 22376 10792
rect 21821 10755 21879 10761
rect 22370 10752 22376 10764
rect 22428 10752 22434 10804
rect 22695 10795 22753 10801
rect 22695 10761 22707 10795
rect 22741 10792 22753 10795
rect 23382 10792 23388 10804
rect 22741 10764 23388 10792
rect 22741 10761 22753 10764
rect 22695 10755 22753 10761
rect 23382 10752 23388 10764
rect 23440 10752 23446 10804
rect 23474 10752 23480 10804
rect 23532 10792 23538 10804
rect 23842 10792 23848 10804
rect 23532 10764 23848 10792
rect 23532 10752 23538 10764
rect 23842 10752 23848 10764
rect 23900 10752 23906 10804
rect 25406 10792 25412 10804
rect 25367 10764 25412 10792
rect 25406 10752 25412 10764
rect 25464 10752 25470 10804
rect 20438 10684 20444 10736
rect 20496 10684 20502 10736
rect 21450 10724 21456 10736
rect 21411 10696 21456 10724
rect 21450 10684 21456 10696
rect 21508 10684 21514 10736
rect 19242 10656 19248 10668
rect 19203 10628 19248 10656
rect 19242 10616 19248 10628
rect 19300 10616 19306 10668
rect 20456 10656 20484 10684
rect 20533 10659 20591 10665
rect 20533 10656 20545 10659
rect 20456 10628 20545 10656
rect 20533 10625 20545 10628
rect 20579 10625 20591 10659
rect 21174 10656 21180 10668
rect 21135 10628 21180 10656
rect 20533 10619 20591 10625
rect 21174 10616 21180 10628
rect 21232 10616 21238 10668
rect 23750 10616 23756 10668
rect 23808 10656 23814 10668
rect 24029 10659 24087 10665
rect 24029 10656 24041 10659
rect 23808 10628 24041 10656
rect 23808 10616 23814 10628
rect 24029 10625 24041 10628
rect 24075 10625 24087 10659
rect 24029 10619 24087 10625
rect 18230 10588 18236 10600
rect 17788 10560 18236 10588
rect 14737 10551 14795 10557
rect 13096 10492 13584 10520
rect 12437 10483 12495 10489
rect 10597 10455 10655 10461
rect 10597 10421 10609 10455
rect 10643 10421 10655 10455
rect 10597 10415 10655 10421
rect 11885 10455 11943 10461
rect 11885 10421 11897 10455
rect 11931 10452 11943 10455
rect 11974 10452 11980 10464
rect 11931 10424 11980 10452
rect 11931 10421 11943 10424
rect 11885 10415 11943 10421
rect 11974 10412 11980 10424
rect 12032 10412 12038 10464
rect 13556 10461 13584 10492
rect 14752 10464 14780 10551
rect 18230 10548 18236 10560
rect 18288 10588 18294 10600
rect 18509 10591 18567 10597
rect 18509 10588 18521 10591
rect 18288 10560 18521 10588
rect 18288 10548 18294 10560
rect 18509 10557 18521 10560
rect 18555 10557 18567 10591
rect 18969 10591 19027 10597
rect 18969 10588 18981 10591
rect 18509 10551 18567 10557
rect 18616 10560 18981 10588
rect 14826 10480 14832 10532
rect 14884 10520 14890 10532
rect 14921 10523 14979 10529
rect 14921 10520 14933 10523
rect 14884 10492 14933 10520
rect 14884 10480 14890 10492
rect 14921 10489 14933 10492
rect 14967 10489 14979 10523
rect 14921 10483 14979 10489
rect 15933 10523 15991 10529
rect 15933 10489 15945 10523
rect 15979 10520 15991 10523
rect 16298 10520 16304 10532
rect 15979 10492 16304 10520
rect 15979 10489 15991 10492
rect 15933 10483 15991 10489
rect 16298 10480 16304 10492
rect 16356 10480 16362 10532
rect 16408 10492 16988 10520
rect 13541 10455 13599 10461
rect 13541 10421 13553 10455
rect 13587 10452 13599 10455
rect 13630 10452 13636 10464
rect 13587 10424 13636 10452
rect 13587 10421 13599 10424
rect 13541 10415 13599 10421
rect 13630 10412 13636 10424
rect 13688 10412 13694 10464
rect 14734 10412 14740 10464
rect 14792 10452 14798 10464
rect 15197 10455 15255 10461
rect 15197 10452 15209 10455
rect 14792 10424 15209 10452
rect 14792 10412 14798 10424
rect 15197 10421 15209 10424
rect 15243 10421 15255 10455
rect 15197 10415 15255 10421
rect 15286 10412 15292 10464
rect 15344 10452 15350 10464
rect 16408 10452 16436 10492
rect 16960 10464 16988 10492
rect 18616 10464 18644 10560
rect 18969 10557 18981 10560
rect 19015 10588 19027 10591
rect 19058 10588 19064 10600
rect 19015 10560 19064 10588
rect 19015 10557 19027 10560
rect 18969 10551 19027 10557
rect 19058 10548 19064 10560
rect 19116 10548 19122 10600
rect 22624 10591 22682 10597
rect 22624 10557 22636 10591
rect 22670 10588 22682 10591
rect 25222 10588 25228 10600
rect 22670 10560 23060 10588
rect 25183 10560 25228 10588
rect 22670 10557 22682 10560
rect 22624 10551 22682 10557
rect 20254 10520 20260 10532
rect 20215 10492 20260 10520
rect 20254 10480 20260 10492
rect 20312 10520 20318 10532
rect 20625 10523 20683 10529
rect 20625 10520 20637 10523
rect 20312 10492 20637 10520
rect 20312 10480 20318 10492
rect 20625 10489 20637 10492
rect 20671 10489 20683 10523
rect 20625 10483 20683 10489
rect 23032 10464 23060 10560
rect 25222 10548 25228 10560
rect 25280 10588 25286 10600
rect 25777 10591 25835 10597
rect 25777 10588 25789 10591
rect 25280 10560 25789 10588
rect 25280 10548 25286 10560
rect 25777 10557 25789 10560
rect 25823 10557 25835 10591
rect 25777 10551 25835 10557
rect 23753 10523 23811 10529
rect 23753 10489 23765 10523
rect 23799 10489 23811 10523
rect 23753 10483 23811 10489
rect 16850 10452 16856 10464
rect 15344 10424 16436 10452
rect 16811 10424 16856 10452
rect 15344 10412 15350 10424
rect 16850 10412 16856 10424
rect 16908 10412 16914 10464
rect 16942 10412 16948 10464
rect 17000 10452 17006 10464
rect 17221 10455 17279 10461
rect 17221 10452 17233 10455
rect 17000 10424 17233 10452
rect 17000 10412 17006 10424
rect 17221 10421 17233 10424
rect 17267 10452 17279 10455
rect 17402 10452 17408 10464
rect 17267 10424 17408 10452
rect 17267 10421 17279 10424
rect 17221 10415 17279 10421
rect 17402 10412 17408 10424
rect 17460 10412 17466 10464
rect 18417 10455 18475 10461
rect 18417 10421 18429 10455
rect 18463 10452 18475 10455
rect 18598 10452 18604 10464
rect 18463 10424 18604 10452
rect 18463 10421 18475 10424
rect 18417 10415 18475 10421
rect 18598 10412 18604 10424
rect 18656 10412 18662 10464
rect 23014 10452 23020 10464
rect 22975 10424 23020 10452
rect 23014 10412 23020 10424
rect 23072 10412 23078 10464
rect 23768 10452 23796 10483
rect 23842 10480 23848 10532
rect 23900 10520 23906 10532
rect 23900 10492 23945 10520
rect 23900 10480 23906 10492
rect 24210 10452 24216 10464
rect 23768 10424 24216 10452
rect 24210 10412 24216 10424
rect 24268 10452 24274 10464
rect 24673 10455 24731 10461
rect 24673 10452 24685 10455
rect 24268 10424 24685 10452
rect 24268 10412 24274 10424
rect 24673 10421 24685 10424
rect 24719 10421 24731 10455
rect 25038 10452 25044 10464
rect 24999 10424 25044 10452
rect 24673 10415 24731 10421
rect 25038 10412 25044 10424
rect 25096 10412 25102 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 3697 10251 3755 10257
rect 3697 10217 3709 10251
rect 3743 10248 3755 10251
rect 3786 10248 3792 10260
rect 3743 10220 3792 10248
rect 3743 10217 3755 10220
rect 3697 10211 3755 10217
rect 3786 10208 3792 10220
rect 3844 10208 3850 10260
rect 5258 10248 5264 10260
rect 5219 10220 5264 10248
rect 5258 10208 5264 10220
rect 5316 10208 5322 10260
rect 7469 10251 7527 10257
rect 7469 10217 7481 10251
rect 7515 10248 7527 10251
rect 7558 10248 7564 10260
rect 7515 10220 7564 10248
rect 7515 10217 7527 10220
rect 7469 10211 7527 10217
rect 7558 10208 7564 10220
rect 7616 10208 7622 10260
rect 9033 10251 9091 10257
rect 9033 10217 9045 10251
rect 9079 10248 9091 10251
rect 9214 10248 9220 10260
rect 9079 10220 9220 10248
rect 9079 10217 9091 10220
rect 9033 10211 9091 10217
rect 9214 10208 9220 10220
rect 9272 10208 9278 10260
rect 9493 10251 9551 10257
rect 9493 10217 9505 10251
rect 9539 10248 9551 10251
rect 9582 10248 9588 10260
rect 9539 10220 9588 10248
rect 9539 10217 9551 10220
rect 9493 10211 9551 10217
rect 9582 10208 9588 10220
rect 9640 10208 9646 10260
rect 11882 10248 11888 10260
rect 11843 10220 11888 10248
rect 11882 10208 11888 10220
rect 11940 10208 11946 10260
rect 12894 10208 12900 10260
rect 12952 10248 12958 10260
rect 13541 10251 13599 10257
rect 13541 10248 13553 10251
rect 12952 10220 13553 10248
rect 12952 10208 12958 10220
rect 13541 10217 13553 10220
rect 13587 10248 13599 10251
rect 13722 10248 13728 10260
rect 13587 10220 13728 10248
rect 13587 10217 13599 10220
rect 13541 10211 13599 10217
rect 13722 10208 13728 10220
rect 13780 10248 13786 10260
rect 13909 10251 13967 10257
rect 13909 10248 13921 10251
rect 13780 10220 13921 10248
rect 13780 10208 13786 10220
rect 13909 10217 13921 10220
rect 13955 10217 13967 10251
rect 13909 10211 13967 10217
rect 14090 10208 14096 10260
rect 14148 10248 14154 10260
rect 14277 10251 14335 10257
rect 14277 10248 14289 10251
rect 14148 10220 14289 10248
rect 14148 10208 14154 10220
rect 14277 10217 14289 10220
rect 14323 10217 14335 10251
rect 16298 10248 16304 10260
rect 16259 10220 16304 10248
rect 14277 10211 14335 10217
rect 16298 10208 16304 10220
rect 16356 10248 16362 10260
rect 16577 10251 16635 10257
rect 16577 10248 16589 10251
rect 16356 10220 16589 10248
rect 16356 10208 16362 10220
rect 16577 10217 16589 10220
rect 16623 10217 16635 10251
rect 18598 10248 18604 10260
rect 18559 10220 18604 10248
rect 16577 10211 16635 10217
rect 18598 10208 18604 10220
rect 18656 10208 18662 10260
rect 19981 10251 20039 10257
rect 19981 10217 19993 10251
rect 20027 10248 20039 10251
rect 20027 10220 21128 10248
rect 20027 10217 20039 10220
rect 19981 10211 20039 10217
rect 2133 10183 2191 10189
rect 2133 10149 2145 10183
rect 2179 10180 2191 10183
rect 2406 10180 2412 10192
rect 2179 10152 2412 10180
rect 2179 10149 2191 10152
rect 2133 10143 2191 10149
rect 2406 10140 2412 10152
rect 2464 10140 2470 10192
rect 4246 10180 4252 10192
rect 4207 10152 4252 10180
rect 4246 10140 4252 10152
rect 4304 10140 4310 10192
rect 6733 10183 6791 10189
rect 6733 10149 6745 10183
rect 6779 10180 6791 10183
rect 6822 10180 6828 10192
rect 6779 10152 6828 10180
rect 6779 10149 6791 10152
rect 6733 10143 6791 10149
rect 6822 10140 6828 10152
rect 6880 10140 6886 10192
rect 7190 10140 7196 10192
rect 7248 10180 7254 10192
rect 7745 10183 7803 10189
rect 7745 10180 7757 10183
rect 7248 10152 7757 10180
rect 7248 10140 7254 10152
rect 7745 10149 7757 10152
rect 7791 10149 7803 10183
rect 7745 10143 7803 10149
rect 9861 10183 9919 10189
rect 9861 10149 9873 10183
rect 9907 10180 9919 10183
rect 10134 10180 10140 10192
rect 9907 10152 10140 10180
rect 9907 10149 9919 10152
rect 9861 10143 9919 10149
rect 10134 10140 10140 10152
rect 10192 10140 10198 10192
rect 1394 10072 1400 10124
rect 1452 10072 1458 10124
rect 6270 10112 6276 10124
rect 6231 10084 6276 10112
rect 6270 10072 6276 10084
rect 6328 10072 6334 10124
rect 6546 10112 6552 10124
rect 6507 10084 6552 10112
rect 6546 10072 6552 10084
rect 6604 10072 6610 10124
rect 11900 10112 11928 10208
rect 21100 10192 21128 10220
rect 22002 10208 22008 10260
rect 22060 10248 22066 10260
rect 22465 10251 22523 10257
rect 22465 10248 22477 10251
rect 22060 10220 22477 10248
rect 22060 10208 22066 10220
rect 22465 10217 22477 10220
rect 22511 10217 22523 10251
rect 22465 10211 22523 10217
rect 23566 10208 23572 10260
rect 23624 10208 23630 10260
rect 24762 10248 24768 10260
rect 24723 10220 24768 10248
rect 24762 10208 24768 10220
rect 24820 10208 24826 10260
rect 25130 10248 25136 10260
rect 25091 10220 25136 10248
rect 25130 10208 25136 10220
rect 25188 10208 25194 10260
rect 15746 10189 15752 10192
rect 14921 10183 14979 10189
rect 14921 10180 14933 10183
rect 14108 10152 14933 10180
rect 12069 10115 12127 10121
rect 12069 10112 12081 10115
rect 11900 10084 12081 10112
rect 12069 10081 12081 10084
rect 12115 10081 12127 10115
rect 12069 10075 12127 10081
rect 12434 10072 12440 10124
rect 12492 10112 12498 10124
rect 13081 10115 13139 10121
rect 12492 10084 12537 10112
rect 12492 10072 12498 10084
rect 13081 10081 13093 10115
rect 13127 10112 13139 10115
rect 13446 10112 13452 10124
rect 13127 10084 13452 10112
rect 13127 10081 13139 10084
rect 13081 10075 13139 10081
rect 13446 10072 13452 10084
rect 13504 10072 13510 10124
rect 13998 10072 14004 10124
rect 14056 10112 14062 10124
rect 14108 10121 14136 10152
rect 14921 10149 14933 10152
rect 14967 10149 14979 10183
rect 15743 10180 15752 10189
rect 15707 10152 15752 10180
rect 14921 10143 14979 10149
rect 15743 10143 15752 10152
rect 15746 10140 15752 10143
rect 15804 10140 15810 10192
rect 17678 10180 17684 10192
rect 17639 10152 17684 10180
rect 17678 10140 17684 10152
rect 17736 10140 17742 10192
rect 19426 10189 19432 10192
rect 19423 10180 19432 10189
rect 19387 10152 19432 10180
rect 19423 10143 19432 10152
rect 19426 10140 19432 10143
rect 19484 10140 19490 10192
rect 21082 10180 21088 10192
rect 20995 10152 21088 10180
rect 21082 10140 21088 10152
rect 21140 10140 21146 10192
rect 23584 10180 23612 10208
rect 23707 10183 23765 10189
rect 23707 10180 23719 10183
rect 23584 10152 23719 10180
rect 23707 10149 23719 10152
rect 23753 10180 23765 10183
rect 25038 10180 25044 10192
rect 23753 10152 25044 10180
rect 23753 10149 23765 10152
rect 23707 10143 23765 10149
rect 25038 10140 25044 10152
rect 25096 10140 25102 10192
rect 14093 10115 14151 10121
rect 14093 10112 14105 10115
rect 14056 10084 14105 10112
rect 14056 10072 14062 10084
rect 14093 10081 14105 10084
rect 14139 10081 14151 10115
rect 14093 10075 14151 10081
rect 14274 10072 14280 10124
rect 14332 10112 14338 10124
rect 14553 10115 14611 10121
rect 14553 10112 14565 10115
rect 14332 10084 14565 10112
rect 14332 10072 14338 10084
rect 14553 10081 14565 10084
rect 14599 10081 14611 10115
rect 14553 10075 14611 10081
rect 23566 10072 23572 10124
rect 23624 10121 23630 10124
rect 23624 10115 23662 10121
rect 23650 10081 23662 10115
rect 23624 10075 23662 10081
rect 23624 10072 23630 10075
rect 24026 10072 24032 10124
rect 24084 10112 24090 10124
rect 24302 10112 24308 10124
rect 24084 10084 24308 10112
rect 24084 10072 24090 10084
rect 24302 10072 24308 10084
rect 24360 10112 24366 10124
rect 24581 10115 24639 10121
rect 24581 10112 24593 10115
rect 24360 10084 24593 10112
rect 24360 10072 24366 10084
rect 24581 10081 24593 10084
rect 24627 10081 24639 10115
rect 24581 10075 24639 10081
rect 1412 9920 1440 10072
rect 2038 10044 2044 10056
rect 1999 10016 2044 10044
rect 2038 10004 2044 10016
rect 2096 10004 2102 10056
rect 2498 10044 2504 10056
rect 2459 10016 2504 10044
rect 2498 10004 2504 10016
rect 2556 10004 2562 10056
rect 4154 10044 4160 10056
rect 4115 10016 4160 10044
rect 4154 10004 4160 10016
rect 4212 10004 4218 10056
rect 4614 10044 4620 10056
rect 4575 10016 4620 10044
rect 4614 10004 4620 10016
rect 4672 10004 4678 10056
rect 7653 10047 7711 10053
rect 7653 10013 7665 10047
rect 7699 10044 7711 10047
rect 8018 10044 8024 10056
rect 7699 10016 8024 10044
rect 7699 10013 7711 10016
rect 7653 10007 7711 10013
rect 8018 10004 8024 10016
rect 8076 10004 8082 10056
rect 9766 10044 9772 10056
rect 9727 10016 9772 10044
rect 9766 10004 9772 10016
rect 9824 10004 9830 10056
rect 10045 10047 10103 10053
rect 10045 10013 10057 10047
rect 10091 10013 10103 10047
rect 10045 10007 10103 10013
rect 13265 10047 13323 10053
rect 13265 10013 13277 10047
rect 13311 10044 13323 10047
rect 13538 10044 13544 10056
rect 13311 10016 13544 10044
rect 13311 10013 13323 10016
rect 13265 10007 13323 10013
rect 2130 9936 2136 9988
rect 2188 9976 2194 9988
rect 2188 9948 2728 9976
rect 2188 9936 2194 9948
rect 1394 9868 1400 9920
rect 1452 9868 1458 9920
rect 1673 9911 1731 9917
rect 1673 9877 1685 9911
rect 1719 9908 1731 9911
rect 2590 9908 2596 9920
rect 1719 9880 2596 9908
rect 1719 9877 1731 9880
rect 1673 9871 1731 9877
rect 2590 9868 2596 9880
rect 2648 9868 2654 9920
rect 2700 9908 2728 9948
rect 4522 9936 4528 9988
rect 4580 9976 4586 9988
rect 5074 9976 5080 9988
rect 4580 9948 5080 9976
rect 4580 9936 4586 9948
rect 5074 9936 5080 9948
rect 5132 9936 5138 9988
rect 8205 9979 8263 9985
rect 8205 9945 8217 9979
rect 8251 9976 8263 9979
rect 8665 9979 8723 9985
rect 8665 9976 8677 9979
rect 8251 9948 8677 9976
rect 8251 9945 8263 9948
rect 8205 9939 8263 9945
rect 8665 9945 8677 9948
rect 8711 9976 8723 9979
rect 9214 9976 9220 9988
rect 8711 9948 9220 9976
rect 8711 9945 8723 9948
rect 8665 9939 8723 9945
rect 9214 9936 9220 9948
rect 9272 9976 9278 9988
rect 10060 9976 10088 10007
rect 13538 10004 13544 10016
rect 13596 10004 13602 10056
rect 15286 10004 15292 10056
rect 15344 10044 15350 10056
rect 15381 10047 15439 10053
rect 15381 10044 15393 10047
rect 15344 10016 15393 10044
rect 15344 10004 15350 10016
rect 15381 10013 15393 10016
rect 15427 10013 15439 10047
rect 15381 10007 15439 10013
rect 16206 10004 16212 10056
rect 16264 10044 16270 10056
rect 17589 10047 17647 10053
rect 17589 10044 17601 10047
rect 16264 10016 17601 10044
rect 16264 10004 16270 10016
rect 17589 10013 17601 10016
rect 17635 10044 17647 10047
rect 17954 10044 17960 10056
rect 17635 10016 17960 10044
rect 17635 10013 17647 10016
rect 17589 10007 17647 10013
rect 17954 10004 17960 10016
rect 18012 10004 18018 10056
rect 19058 10044 19064 10056
rect 19019 10016 19064 10044
rect 19058 10004 19064 10016
rect 19116 10004 19122 10056
rect 20993 10047 21051 10053
rect 20993 10013 21005 10047
rect 21039 10044 21051 10047
rect 21174 10044 21180 10056
rect 21039 10016 21180 10044
rect 21039 10013 21051 10016
rect 20993 10007 21051 10013
rect 21174 10004 21180 10016
rect 21232 10004 21238 10056
rect 21269 10047 21327 10053
rect 21269 10013 21281 10047
rect 21315 10013 21327 10047
rect 21269 10007 21327 10013
rect 9272 9948 10088 9976
rect 9272 9936 9278 9948
rect 11974 9936 11980 9988
rect 12032 9976 12038 9988
rect 13998 9976 14004 9988
rect 12032 9948 14004 9976
rect 12032 9936 12038 9948
rect 13998 9936 14004 9948
rect 14056 9936 14062 9988
rect 18141 9979 18199 9985
rect 18141 9945 18153 9979
rect 18187 9976 18199 9979
rect 21284 9976 21312 10007
rect 21634 9976 21640 9988
rect 18187 9948 21640 9976
rect 18187 9945 18199 9948
rect 18141 9939 18199 9945
rect 21634 9936 21640 9948
rect 21692 9936 21698 9988
rect 23658 9936 23664 9988
rect 23716 9976 23722 9988
rect 24029 9979 24087 9985
rect 24029 9976 24041 9979
rect 23716 9948 24041 9976
rect 23716 9936 23722 9948
rect 24029 9945 24041 9948
rect 24075 9945 24087 9979
rect 24029 9939 24087 9945
rect 2961 9911 3019 9917
rect 2961 9908 2973 9911
rect 2700 9880 2973 9908
rect 2961 9877 2973 9880
rect 3007 9877 3019 9911
rect 2961 9871 3019 9877
rect 10781 9911 10839 9917
rect 10781 9877 10793 9911
rect 10827 9908 10839 9911
rect 10962 9908 10968 9920
rect 10827 9880 10968 9908
rect 10827 9877 10839 9880
rect 10781 9871 10839 9877
rect 10962 9868 10968 9880
rect 11020 9868 11026 9920
rect 11517 9911 11575 9917
rect 11517 9877 11529 9911
rect 11563 9908 11575 9911
rect 12158 9908 12164 9920
rect 11563 9880 12164 9908
rect 11563 9877 11575 9880
rect 11517 9871 11575 9877
rect 12158 9868 12164 9880
rect 12216 9868 12222 9920
rect 16574 9868 16580 9920
rect 16632 9908 16638 9920
rect 16945 9911 17003 9917
rect 16945 9908 16957 9911
rect 16632 9880 16957 9908
rect 16632 9868 16638 9880
rect 16945 9877 16957 9880
rect 16991 9877 17003 9911
rect 20438 9908 20444 9920
rect 20399 9880 20444 9908
rect 16945 9871 17003 9877
rect 20438 9868 20444 9880
rect 20496 9868 20502 9920
rect 21358 9868 21364 9920
rect 21416 9908 21422 9920
rect 21913 9911 21971 9917
rect 21913 9908 21925 9911
rect 21416 9880 21925 9908
rect 21416 9868 21422 9880
rect 21913 9877 21925 9880
rect 21959 9877 21971 9911
rect 21913 9871 21971 9877
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 2406 9704 2412 9716
rect 2367 9676 2412 9704
rect 2406 9664 2412 9676
rect 2464 9664 2470 9716
rect 4154 9664 4160 9716
rect 4212 9704 4218 9716
rect 5258 9704 5264 9716
rect 4212 9676 5264 9704
rect 4212 9664 4218 9676
rect 5258 9664 5264 9676
rect 5316 9704 5322 9716
rect 6086 9704 6092 9716
rect 5316 9676 5488 9704
rect 5999 9676 6092 9704
rect 5316 9664 5322 9676
rect 1854 9596 1860 9648
rect 1912 9596 1918 9648
rect 5460 9636 5488 9676
rect 6086 9664 6092 9676
rect 6144 9704 6150 9716
rect 6270 9704 6276 9716
rect 6144 9676 6276 9704
rect 6144 9664 6150 9676
rect 6270 9664 6276 9676
rect 6328 9664 6334 9716
rect 6457 9707 6515 9713
rect 6457 9673 6469 9707
rect 6503 9704 6515 9707
rect 6546 9704 6552 9716
rect 6503 9676 6552 9704
rect 6503 9673 6515 9676
rect 6457 9667 6515 9673
rect 6546 9664 6552 9676
rect 6604 9664 6610 9716
rect 10134 9704 10140 9716
rect 10095 9676 10140 9704
rect 10134 9664 10140 9676
rect 10192 9664 10198 9716
rect 10597 9707 10655 9713
rect 10597 9673 10609 9707
rect 10643 9704 10655 9707
rect 10778 9704 10784 9716
rect 10643 9676 10784 9704
rect 10643 9673 10655 9676
rect 10597 9667 10655 9673
rect 10778 9664 10784 9676
rect 10836 9664 10842 9716
rect 13630 9704 13636 9716
rect 12452 9676 13636 9704
rect 5537 9639 5595 9645
rect 5537 9636 5549 9639
rect 5460 9608 5549 9636
rect 5537 9605 5549 9608
rect 5583 9605 5595 9639
rect 11882 9636 11888 9648
rect 11843 9608 11888 9636
rect 5537 9599 5595 9605
rect 11882 9596 11888 9608
rect 11940 9636 11946 9648
rect 12161 9639 12219 9645
rect 12161 9636 12173 9639
rect 11940 9608 12173 9636
rect 11940 9596 11946 9608
rect 12161 9605 12173 9608
rect 12207 9636 12219 9639
rect 12452 9636 12480 9676
rect 13630 9664 13636 9676
rect 13688 9664 13694 9716
rect 15286 9664 15292 9716
rect 15344 9704 15350 9716
rect 15344 9676 16528 9704
rect 15344 9664 15350 9676
rect 12207 9608 12480 9636
rect 12207 9605 12219 9608
rect 12161 9599 12219 9605
rect 1872 9568 1900 9596
rect 2682 9568 2688 9580
rect 1688 9540 2688 9568
rect 1688 9509 1716 9540
rect 2682 9528 2688 9540
rect 2740 9528 2746 9580
rect 3142 9528 3148 9580
rect 3200 9568 3206 9580
rect 3697 9571 3755 9577
rect 3697 9568 3709 9571
rect 3200 9540 3709 9568
rect 3200 9528 3206 9540
rect 3697 9537 3709 9540
rect 3743 9568 3755 9571
rect 4614 9568 4620 9580
rect 3743 9540 4620 9568
rect 3743 9537 3755 9540
rect 3697 9531 3755 9537
rect 4614 9528 4620 9540
rect 4672 9528 4678 9580
rect 4890 9568 4896 9580
rect 4851 9540 4896 9568
rect 4890 9528 4896 9540
rect 4948 9528 4954 9580
rect 8297 9571 8355 9577
rect 8297 9537 8309 9571
rect 8343 9568 8355 9571
rect 9214 9568 9220 9580
rect 8343 9540 9220 9568
rect 8343 9537 8355 9540
rect 8297 9531 8355 9537
rect 9214 9528 9220 9540
rect 9272 9528 9278 9580
rect 9674 9568 9680 9580
rect 9635 9540 9680 9568
rect 9674 9528 9680 9540
rect 9732 9528 9738 9580
rect 1673 9503 1731 9509
rect 1673 9469 1685 9503
rect 1719 9469 1731 9503
rect 1673 9463 1731 9469
rect 1949 9503 2007 9509
rect 1949 9469 1961 9503
rect 1995 9500 2007 9503
rect 2590 9500 2596 9512
rect 1995 9472 2596 9500
rect 1995 9469 2007 9472
rect 1949 9463 2007 9469
rect 2590 9460 2596 9472
rect 2648 9460 2654 9512
rect 10778 9500 10784 9512
rect 10739 9472 10784 9500
rect 10778 9460 10784 9472
rect 10836 9460 10842 9512
rect 10962 9460 10968 9512
rect 11020 9500 11026 9512
rect 11238 9500 11244 9512
rect 11020 9472 11244 9500
rect 11020 9460 11026 9472
rect 11238 9460 11244 9472
rect 11296 9460 11302 9512
rect 12452 9509 12480 9608
rect 12529 9639 12587 9645
rect 12529 9605 12541 9639
rect 12575 9636 12587 9639
rect 13078 9636 13084 9648
rect 12575 9608 13084 9636
rect 12575 9605 12587 9608
rect 12529 9599 12587 9605
rect 13078 9596 13084 9608
rect 13136 9596 13142 9648
rect 13446 9636 13452 9648
rect 13407 9608 13452 9636
rect 13446 9596 13452 9608
rect 13504 9596 13510 9648
rect 13814 9636 13820 9648
rect 13775 9608 13820 9636
rect 13814 9596 13820 9608
rect 13872 9596 13878 9648
rect 16500 9636 16528 9676
rect 21082 9664 21088 9716
rect 21140 9704 21146 9716
rect 21140 9676 22140 9704
rect 21140 9664 21146 9676
rect 16669 9639 16727 9645
rect 16669 9636 16681 9639
rect 16500 9608 16681 9636
rect 16669 9605 16681 9608
rect 16715 9605 16727 9639
rect 16669 9599 16727 9605
rect 17954 9596 17960 9648
rect 18012 9636 18018 9648
rect 18233 9639 18291 9645
rect 18233 9636 18245 9639
rect 18012 9608 18245 9636
rect 18012 9596 18018 9608
rect 18233 9605 18245 9608
rect 18279 9605 18291 9639
rect 18233 9599 18291 9605
rect 21174 9596 21180 9648
rect 21232 9636 21238 9648
rect 22112 9636 22140 9676
rect 24026 9664 24032 9716
rect 24084 9704 24090 9716
rect 24397 9707 24455 9713
rect 24397 9704 24409 9707
rect 24084 9676 24409 9704
rect 24084 9664 24090 9676
rect 24397 9673 24409 9676
rect 24443 9673 24455 9707
rect 24397 9667 24455 9673
rect 22281 9639 22339 9645
rect 22281 9636 22293 9639
rect 21232 9608 22048 9636
rect 22112 9608 22293 9636
rect 21232 9596 21238 9608
rect 12618 9528 12624 9580
rect 12676 9568 12682 9580
rect 12897 9571 12955 9577
rect 12897 9568 12909 9571
rect 12676 9540 12909 9568
rect 12676 9528 12682 9540
rect 12897 9537 12909 9540
rect 12943 9537 12955 9571
rect 12897 9531 12955 9537
rect 12437 9503 12495 9509
rect 12437 9469 12449 9503
rect 12483 9469 12495 9503
rect 12710 9500 12716 9512
rect 12671 9472 12716 9500
rect 12437 9463 12495 9469
rect 12710 9460 12716 9472
rect 12768 9460 12774 9512
rect 13832 9500 13860 9596
rect 21358 9568 21364 9580
rect 21319 9540 21364 9568
rect 21358 9528 21364 9540
rect 21416 9528 21422 9580
rect 21634 9568 21640 9580
rect 21595 9540 21640 9568
rect 21634 9528 21640 9540
rect 21692 9528 21698 9580
rect 14001 9503 14059 9509
rect 14001 9500 14013 9503
rect 13832 9472 14013 9500
rect 14001 9469 14013 9472
rect 14047 9469 14059 9503
rect 15102 9500 15108 9512
rect 15063 9472 15108 9500
rect 14001 9463 14059 9469
rect 15102 9460 15108 9472
rect 15160 9500 15166 9512
rect 16301 9503 16359 9509
rect 16301 9500 16313 9503
rect 15160 9472 16313 9500
rect 15160 9460 15166 9472
rect 16301 9469 16313 9472
rect 16347 9469 16359 9503
rect 16301 9463 16359 9469
rect 16758 9460 16764 9512
rect 16816 9500 16822 9512
rect 16888 9503 16946 9509
rect 16888 9500 16900 9503
rect 16816 9472 16900 9500
rect 16816 9460 16822 9472
rect 16888 9469 16900 9472
rect 16934 9500 16946 9503
rect 17313 9503 17371 9509
rect 17313 9500 17325 9503
rect 16934 9472 17325 9500
rect 16934 9469 16946 9472
rect 16888 9463 16946 9469
rect 17313 9469 17325 9472
rect 17359 9469 17371 9503
rect 19518 9500 19524 9512
rect 19479 9472 19524 9500
rect 17313 9463 17371 9469
rect 19518 9460 19524 9472
rect 19576 9460 19582 9512
rect 20441 9503 20499 9509
rect 20441 9469 20453 9503
rect 20487 9500 20499 9503
rect 21085 9503 21143 9509
rect 21085 9500 21097 9503
rect 20487 9472 21097 9500
rect 20487 9469 20499 9472
rect 20441 9463 20499 9469
rect 21085 9469 21097 9472
rect 21131 9469 21143 9503
rect 21085 9463 21143 9469
rect 2130 9432 2136 9444
rect 2091 9404 2136 9432
rect 2130 9392 2136 9404
rect 2188 9392 2194 9444
rect 3050 9432 3056 9444
rect 3011 9404 3056 9432
rect 3050 9392 3056 9404
rect 3108 9392 3114 9444
rect 3145 9435 3203 9441
rect 3145 9401 3157 9435
rect 3191 9432 3203 9435
rect 3234 9432 3240 9444
rect 3191 9404 3240 9432
rect 3191 9401 3203 9404
rect 3145 9395 3203 9401
rect 1670 9364 1676 9376
rect 1044 9336 1676 9364
rect 1044 9160 1072 9336
rect 1670 9324 1676 9336
rect 1728 9324 1734 9376
rect 2869 9367 2927 9373
rect 2869 9333 2881 9367
rect 2915 9364 2927 9367
rect 3160 9364 3188 9395
rect 3234 9392 3240 9404
rect 3292 9392 3298 9444
rect 3878 9392 3884 9444
rect 3936 9432 3942 9444
rect 4617 9435 4675 9441
rect 4617 9432 4629 9435
rect 3936 9404 4629 9432
rect 3936 9392 3942 9404
rect 4617 9401 4629 9404
rect 4663 9401 4675 9435
rect 4617 9395 4675 9401
rect 4706 9392 4712 9444
rect 4764 9432 4770 9444
rect 4764 9404 4809 9432
rect 4764 9392 4770 9404
rect 7282 9392 7288 9444
rect 7340 9432 7346 9444
rect 7377 9435 7435 9441
rect 7377 9432 7389 9435
rect 7340 9404 7389 9432
rect 7340 9392 7346 9404
rect 7377 9401 7389 9404
rect 7423 9401 7435 9435
rect 7377 9395 7435 9401
rect 7653 9435 7711 9441
rect 7653 9401 7665 9435
rect 7699 9401 7711 9435
rect 7653 9395 7711 9401
rect 4062 9364 4068 9376
rect 2915 9336 3188 9364
rect 4023 9336 4068 9364
rect 2915 9333 2927 9336
rect 2869 9327 2927 9333
rect 4062 9324 4068 9336
rect 4120 9364 4126 9376
rect 4246 9364 4252 9376
rect 4120 9336 4252 9364
rect 4120 9324 4126 9336
rect 4246 9324 4252 9336
rect 4304 9324 4310 9376
rect 7006 9364 7012 9376
rect 6967 9336 7012 9364
rect 7006 9324 7012 9336
rect 7064 9324 7070 9376
rect 7668 9364 7696 9395
rect 7742 9392 7748 9444
rect 7800 9432 7806 9444
rect 9033 9435 9091 9441
rect 7800 9404 7845 9432
rect 7800 9392 7806 9404
rect 9033 9401 9045 9435
rect 9079 9432 9091 9435
rect 9306 9432 9312 9444
rect 9079 9404 9312 9432
rect 9079 9401 9091 9404
rect 9033 9395 9091 9401
rect 9306 9392 9312 9404
rect 9364 9392 9370 9444
rect 10042 9392 10048 9444
rect 10100 9432 10106 9444
rect 14553 9435 14611 9441
rect 14553 9432 14565 9435
rect 10100 9404 14565 9432
rect 10100 9392 10106 9404
rect 14553 9401 14565 9404
rect 14599 9401 14611 9435
rect 14553 9395 14611 9401
rect 15013 9435 15071 9441
rect 15013 9401 15025 9435
rect 15059 9432 15071 9435
rect 15467 9435 15525 9441
rect 15467 9432 15479 9435
rect 15059 9404 15479 9432
rect 15059 9401 15071 9404
rect 15013 9395 15071 9401
rect 15467 9401 15479 9404
rect 15513 9432 15525 9435
rect 15746 9432 15752 9444
rect 15513 9404 15752 9432
rect 15513 9401 15525 9404
rect 15467 9395 15525 9401
rect 15746 9392 15752 9404
rect 15804 9392 15810 9444
rect 16390 9392 16396 9444
rect 16448 9432 16454 9444
rect 16991 9435 17049 9441
rect 16991 9432 17003 9435
rect 16448 9404 17003 9432
rect 16448 9392 16454 9404
rect 16991 9401 17003 9404
rect 17037 9401 17049 9435
rect 16991 9395 17049 9401
rect 19153 9435 19211 9441
rect 19153 9401 19165 9435
rect 19199 9432 19211 9435
rect 19426 9432 19432 9444
rect 19199 9404 19432 9432
rect 19199 9401 19211 9404
rect 19153 9395 19211 9401
rect 19426 9392 19432 9404
rect 19484 9432 19490 9444
rect 19883 9435 19941 9441
rect 19883 9432 19895 9435
rect 19484 9404 19895 9432
rect 19484 9392 19490 9404
rect 19883 9401 19895 9404
rect 19929 9432 19941 9435
rect 19929 9404 20852 9432
rect 19929 9401 19941 9404
rect 19883 9395 19941 9401
rect 20824 9376 20852 9404
rect 8570 9364 8576 9376
rect 7668 9336 8576 9364
rect 8570 9324 8576 9336
rect 8628 9324 8634 9376
rect 10778 9364 10784 9376
rect 10739 9336 10784 9364
rect 10778 9324 10784 9336
rect 10836 9324 10842 9376
rect 14182 9364 14188 9376
rect 14143 9336 14188 9364
rect 14182 9324 14188 9336
rect 14240 9324 14246 9376
rect 16025 9367 16083 9373
rect 16025 9333 16037 9367
rect 16071 9364 16083 9367
rect 16114 9364 16120 9376
rect 16071 9336 16120 9364
rect 16071 9333 16083 9336
rect 16025 9327 16083 9333
rect 16114 9324 16120 9336
rect 16172 9324 16178 9376
rect 17678 9324 17684 9376
rect 17736 9364 17742 9376
rect 17773 9367 17831 9373
rect 17773 9364 17785 9367
rect 17736 9336 17785 9364
rect 17736 9324 17742 9336
rect 17773 9333 17785 9336
rect 17819 9364 17831 9367
rect 17954 9364 17960 9376
rect 17819 9336 17960 9364
rect 17819 9333 17831 9336
rect 17773 9327 17831 9333
rect 17954 9324 17960 9336
rect 18012 9324 18018 9376
rect 18506 9364 18512 9376
rect 18467 9336 18512 9364
rect 18506 9324 18512 9336
rect 18564 9324 18570 9376
rect 20806 9364 20812 9376
rect 20767 9336 20812 9364
rect 20806 9324 20812 9336
rect 20864 9324 20870 9376
rect 21100 9364 21128 9463
rect 21453 9435 21511 9441
rect 21453 9401 21465 9435
rect 21499 9401 21511 9435
rect 21453 9395 21511 9401
rect 21468 9364 21496 9395
rect 21100 9336 21496 9364
rect 22020 9364 22048 9608
rect 22281 9605 22293 9608
rect 22327 9605 22339 9639
rect 24762 9636 24768 9648
rect 24723 9608 24768 9636
rect 22281 9599 22339 9605
rect 24762 9596 24768 9608
rect 24820 9596 24826 9648
rect 25225 9639 25283 9645
rect 25225 9605 25237 9639
rect 25271 9636 25283 9639
rect 25314 9636 25320 9648
rect 25271 9608 25320 9636
rect 25271 9605 25283 9608
rect 25225 9599 25283 9605
rect 24581 9503 24639 9509
rect 24581 9469 24593 9503
rect 24627 9500 24639 9503
rect 25240 9500 25268 9599
rect 25314 9596 25320 9608
rect 25372 9596 25378 9648
rect 24627 9472 25268 9500
rect 24627 9469 24639 9472
rect 24581 9463 24639 9469
rect 22649 9367 22707 9373
rect 22649 9364 22661 9367
rect 22020 9336 22661 9364
rect 22649 9333 22661 9336
rect 22695 9333 22707 9367
rect 22649 9327 22707 9333
rect 23566 9324 23572 9376
rect 23624 9364 23630 9376
rect 23845 9367 23903 9373
rect 23845 9364 23857 9367
rect 23624 9336 23857 9364
rect 23624 9324 23630 9336
rect 23845 9333 23857 9336
rect 23891 9333 23903 9367
rect 23845 9327 23903 9333
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 1535 9163 1593 9169
rect 1535 9160 1547 9163
rect 1044 9132 1547 9160
rect 1535 9129 1547 9132
rect 1581 9129 1593 9163
rect 1854 9160 1860 9172
rect 1815 9132 1860 9160
rect 1535 9123 1593 9129
rect 1854 9120 1860 9132
rect 1912 9120 1918 9172
rect 3878 9160 3884 9172
rect 3839 9132 3884 9160
rect 3878 9120 3884 9132
rect 3936 9120 3942 9172
rect 7006 9120 7012 9172
rect 7064 9160 7070 9172
rect 7742 9160 7748 9172
rect 7064 9132 7748 9160
rect 7064 9120 7070 9132
rect 7742 9120 7748 9132
rect 7800 9120 7806 9172
rect 8478 9120 8484 9172
rect 8536 9160 8542 9172
rect 8711 9163 8769 9169
rect 8711 9160 8723 9163
rect 8536 9132 8723 9160
rect 8536 9120 8542 9132
rect 8711 9129 8723 9132
rect 8757 9129 8769 9163
rect 8711 9123 8769 9129
rect 9306 9120 9312 9172
rect 9364 9160 9370 9172
rect 10597 9163 10655 9169
rect 10597 9160 10609 9163
rect 9364 9132 10609 9160
rect 9364 9120 9370 9132
rect 10597 9129 10609 9132
rect 10643 9129 10655 9163
rect 10597 9123 10655 9129
rect 11974 9120 11980 9172
rect 12032 9160 12038 9172
rect 12710 9160 12716 9172
rect 12032 9132 12716 9160
rect 12032 9120 12038 9132
rect 12710 9120 12716 9132
rect 12768 9160 12774 9172
rect 13265 9163 13323 9169
rect 13265 9160 13277 9163
rect 12768 9132 13277 9160
rect 12768 9120 12774 9132
rect 13265 9129 13277 9132
rect 13311 9129 13323 9163
rect 13265 9123 13323 9129
rect 16022 9120 16028 9172
rect 16080 9160 16086 9172
rect 16209 9163 16267 9169
rect 16209 9160 16221 9163
rect 16080 9132 16221 9160
rect 16080 9120 16086 9132
rect 16209 9129 16221 9132
rect 16255 9129 16267 9163
rect 16209 9123 16267 9129
rect 17954 9120 17960 9172
rect 18012 9160 18018 9172
rect 18417 9163 18475 9169
rect 18417 9160 18429 9163
rect 18012 9132 18429 9160
rect 18012 9120 18018 9132
rect 18417 9129 18429 9132
rect 18463 9129 18475 9163
rect 19058 9160 19064 9172
rect 19019 9132 19064 9160
rect 18417 9123 18475 9129
rect 19058 9120 19064 9132
rect 19116 9160 19122 9172
rect 19337 9163 19395 9169
rect 19337 9160 19349 9163
rect 19116 9132 19349 9160
rect 19116 9120 19122 9132
rect 19337 9129 19349 9132
rect 19383 9129 19395 9163
rect 19337 9123 19395 9129
rect 20898 9120 20904 9172
rect 20956 9160 20962 9172
rect 21266 9160 21272 9172
rect 20956 9132 21272 9160
rect 20956 9120 20962 9132
rect 2593 9095 2651 9101
rect 2593 9061 2605 9095
rect 2639 9092 2651 9095
rect 2774 9092 2780 9104
rect 2639 9064 2780 9092
rect 2639 9061 2651 9064
rect 2593 9055 2651 9061
rect 2774 9052 2780 9064
rect 2832 9052 2838 9104
rect 3142 9092 3148 9104
rect 3103 9064 3148 9092
rect 3142 9052 3148 9064
rect 3200 9052 3206 9104
rect 5163 9095 5221 9101
rect 5163 9061 5175 9095
rect 5209 9092 5221 9095
rect 5442 9092 5448 9104
rect 5209 9064 5448 9092
rect 5209 9061 5221 9064
rect 5163 9055 5221 9061
rect 5442 9052 5448 9064
rect 5500 9052 5506 9104
rect 7190 9101 7196 9104
rect 7187 9092 7196 9101
rect 7151 9064 7196 9092
rect 7187 9055 7196 9064
rect 7190 9052 7196 9055
rect 7248 9052 7254 9104
rect 10042 9101 10048 9104
rect 10039 9092 10048 9101
rect 10003 9064 10048 9092
rect 10039 9055 10048 9064
rect 10042 9052 10048 9055
rect 10100 9052 10106 9104
rect 14369 9095 14427 9101
rect 14369 9061 14381 9095
rect 14415 9092 14427 9095
rect 15102 9092 15108 9104
rect 14415 9064 15108 9092
rect 14415 9061 14427 9064
rect 14369 9055 14427 9061
rect 15102 9052 15108 9064
rect 15160 9052 15166 9104
rect 15651 9095 15709 9101
rect 15651 9061 15663 9095
rect 15697 9092 15709 9095
rect 15746 9092 15752 9104
rect 15697 9064 15752 9092
rect 15697 9061 15709 9064
rect 15651 9055 15709 9061
rect 15746 9052 15752 9064
rect 15804 9092 15810 9104
rect 17586 9092 17592 9104
rect 15804 9064 17592 9092
rect 15804 9052 15810 9064
rect 17586 9052 17592 9064
rect 17644 9092 17650 9104
rect 17859 9095 17917 9101
rect 17859 9092 17871 9095
rect 17644 9064 17871 9092
rect 17644 9052 17650 9064
rect 17859 9061 17871 9064
rect 17905 9092 17917 9095
rect 19426 9092 19432 9104
rect 17905 9064 19432 9092
rect 17905 9061 17917 9064
rect 17859 9055 17917 9061
rect 19426 9052 19432 9064
rect 19484 9052 19490 9104
rect 20990 9092 20996 9104
rect 20951 9064 20996 9092
rect 20990 9052 20996 9064
rect 21048 9052 21054 9104
rect 21100 9101 21128 9132
rect 21266 9120 21272 9132
rect 21324 9160 21330 9172
rect 21913 9163 21971 9169
rect 21913 9160 21925 9163
rect 21324 9132 21925 9160
rect 21324 9120 21330 9132
rect 21913 9129 21925 9132
rect 21959 9160 21971 9163
rect 22094 9160 22100 9172
rect 21959 9132 22100 9160
rect 21959 9129 21971 9132
rect 21913 9123 21971 9129
rect 22094 9120 22100 9132
rect 22152 9120 22158 9172
rect 21085 9095 21143 9101
rect 21085 9061 21097 9095
rect 21131 9061 21143 9095
rect 22646 9092 22652 9104
rect 22607 9064 22652 9092
rect 21085 9055 21143 9061
rect 22646 9052 22652 9064
rect 22704 9052 22710 9104
rect 1464 9027 1522 9033
rect 1464 8993 1476 9027
rect 1510 9024 1522 9027
rect 2314 9024 2320 9036
rect 1510 8996 2320 9024
rect 1510 8993 1522 8996
rect 1464 8987 1522 8993
rect 2314 8984 2320 8996
rect 2372 8984 2378 9036
rect 4617 9027 4675 9033
rect 4617 8993 4629 9027
rect 4663 9024 4675 9027
rect 4706 9024 4712 9036
rect 4663 8996 4712 9024
rect 4663 8993 4675 8996
rect 4617 8987 4675 8993
rect 4706 8984 4712 8996
rect 4764 9024 4770 9036
rect 5721 9027 5779 9033
rect 5721 9024 5733 9027
rect 4764 8996 5733 9024
rect 4764 8984 4770 8996
rect 5721 8993 5733 8996
rect 5767 8993 5779 9027
rect 5721 8987 5779 8993
rect 8478 8984 8484 9036
rect 8536 9024 8542 9036
rect 8608 9027 8666 9033
rect 8608 9024 8620 9027
rect 8536 8996 8620 9024
rect 8536 8984 8542 8996
rect 8608 8993 8620 8996
rect 8654 8993 8666 9027
rect 8608 8987 8666 8993
rect 12529 9027 12587 9033
rect 12529 8993 12541 9027
rect 12575 8993 12587 9027
rect 12529 8987 12587 8993
rect 2130 8916 2136 8968
rect 2188 8956 2194 8968
rect 2225 8959 2283 8965
rect 2225 8956 2237 8959
rect 2188 8928 2237 8956
rect 2188 8916 2194 8928
rect 2225 8925 2237 8928
rect 2271 8925 2283 8959
rect 2225 8919 2283 8925
rect 2501 8959 2559 8965
rect 2501 8925 2513 8959
rect 2547 8956 2559 8959
rect 2682 8956 2688 8968
rect 2547 8928 2688 8956
rect 2547 8925 2559 8928
rect 2501 8919 2559 8925
rect 2682 8916 2688 8928
rect 2740 8916 2746 8968
rect 4430 8916 4436 8968
rect 4488 8956 4494 8968
rect 4801 8959 4859 8965
rect 4801 8956 4813 8959
rect 4488 8928 4813 8956
rect 4488 8916 4494 8928
rect 4801 8925 4813 8928
rect 4847 8956 4859 8959
rect 5534 8956 5540 8968
rect 4847 8928 5540 8956
rect 4847 8925 4859 8928
rect 4801 8919 4859 8925
rect 5534 8916 5540 8928
rect 5592 8916 5598 8968
rect 6825 8959 6883 8965
rect 6825 8925 6837 8959
rect 6871 8956 6883 8959
rect 7926 8956 7932 8968
rect 6871 8928 7932 8956
rect 6871 8925 6883 8928
rect 6825 8919 6883 8925
rect 7926 8916 7932 8928
rect 7984 8916 7990 8968
rect 9677 8959 9735 8965
rect 9677 8925 9689 8959
rect 9723 8956 9735 8959
rect 10778 8956 10784 8968
rect 9723 8928 10784 8956
rect 9723 8925 9735 8928
rect 9677 8919 9735 8925
rect 10778 8916 10784 8928
rect 10836 8916 10842 8968
rect 12434 8956 12440 8968
rect 11900 8928 12440 8956
rect 11900 8832 11928 8928
rect 12434 8916 12440 8928
rect 12492 8916 12498 8968
rect 12544 8956 12572 8987
rect 13354 8984 13360 9036
rect 13412 9024 13418 9036
rect 13633 9027 13691 9033
rect 13633 9024 13645 9027
rect 13412 8996 13645 9024
rect 13412 8984 13418 8996
rect 13633 8993 13645 8996
rect 13679 8993 13691 9027
rect 13633 8987 13691 8993
rect 14185 9027 14243 9033
rect 14185 8993 14197 9027
rect 14231 9024 14243 9027
rect 14734 9024 14740 9036
rect 14231 8996 14740 9024
rect 14231 8993 14243 8996
rect 14185 8987 14243 8993
rect 14734 8984 14740 8996
rect 14792 8984 14798 9036
rect 14826 8984 14832 9036
rect 14884 9024 14890 9036
rect 15289 9027 15347 9033
rect 15289 9024 15301 9027
rect 14884 8996 15301 9024
rect 14884 8984 14890 8996
rect 15289 8993 15301 8996
rect 15335 9024 15347 9027
rect 16574 9024 16580 9036
rect 15335 8996 16580 9024
rect 15335 8993 15347 8996
rect 15289 8987 15347 8993
rect 16574 8984 16580 8996
rect 16632 8984 16638 9036
rect 19334 9024 19340 9036
rect 19295 8996 19340 9024
rect 19334 8984 19340 8996
rect 19392 8984 19398 9036
rect 19702 9024 19708 9036
rect 19663 8996 19708 9024
rect 19702 8984 19708 8996
rect 19760 8984 19766 9036
rect 24581 9027 24639 9033
rect 24581 8993 24593 9027
rect 24627 9024 24639 9027
rect 25498 9024 25504 9036
rect 24627 8996 25504 9024
rect 24627 8993 24639 8996
rect 24581 8987 24639 8993
rect 25498 8984 25504 8996
rect 25556 8984 25562 9036
rect 12618 8956 12624 8968
rect 12531 8928 12624 8956
rect 12618 8916 12624 8928
rect 12676 8956 12682 8968
rect 13446 8956 13452 8968
rect 12676 8928 13452 8956
rect 12676 8916 12682 8928
rect 13446 8916 13452 8928
rect 13504 8916 13510 8968
rect 17126 8916 17132 8968
rect 17184 8956 17190 8968
rect 17497 8959 17555 8965
rect 17497 8956 17509 8959
rect 17184 8928 17509 8956
rect 17184 8916 17190 8928
rect 17497 8925 17509 8928
rect 17543 8925 17555 8959
rect 17497 8919 17555 8925
rect 21174 8916 21180 8968
rect 21232 8956 21238 8968
rect 21269 8959 21327 8965
rect 21269 8956 21281 8959
rect 21232 8928 21281 8956
rect 21232 8916 21238 8928
rect 21269 8925 21281 8928
rect 21315 8925 21327 8959
rect 22554 8956 22560 8968
rect 22515 8928 22560 8956
rect 21269 8919 21327 8925
rect 22554 8916 22560 8928
rect 22612 8916 22618 8968
rect 22833 8959 22891 8965
rect 22833 8925 22845 8959
rect 22879 8925 22891 8959
rect 22833 8919 22891 8925
rect 11974 8848 11980 8900
rect 12032 8888 12038 8900
rect 12161 8891 12219 8897
rect 12161 8888 12173 8891
rect 12032 8860 12173 8888
rect 12032 8848 12038 8860
rect 12161 8857 12173 8860
rect 12207 8857 12219 8891
rect 12161 8851 12219 8857
rect 19518 8848 19524 8900
rect 19576 8888 19582 8900
rect 20257 8891 20315 8897
rect 20257 8888 20269 8891
rect 19576 8860 20269 8888
rect 19576 8848 19582 8860
rect 20257 8857 20269 8860
rect 20303 8857 20315 8891
rect 20257 8851 20315 8857
rect 21358 8848 21364 8900
rect 21416 8888 21422 8900
rect 22848 8888 22876 8919
rect 21416 8860 22876 8888
rect 21416 8848 21422 8860
rect 2038 8780 2044 8832
rect 2096 8820 2102 8832
rect 2222 8820 2228 8832
rect 2096 8792 2228 8820
rect 2096 8780 2102 8792
rect 2222 8780 2228 8792
rect 2280 8780 2286 8832
rect 3142 8780 3148 8832
rect 3200 8820 3206 8832
rect 3421 8823 3479 8829
rect 3421 8820 3433 8823
rect 3200 8792 3433 8820
rect 3200 8780 3206 8792
rect 3421 8789 3433 8792
rect 3467 8789 3479 8823
rect 8018 8820 8024 8832
rect 7979 8792 8024 8820
rect 3421 8783 3479 8789
rect 8018 8780 8024 8792
rect 8076 8780 8082 8832
rect 9122 8820 9128 8832
rect 9083 8792 9128 8820
rect 9122 8780 9128 8792
rect 9180 8780 9186 8832
rect 9493 8823 9551 8829
rect 9493 8789 9505 8823
rect 9539 8820 9551 8823
rect 9582 8820 9588 8832
rect 9539 8792 9588 8820
rect 9539 8789 9551 8792
rect 9493 8783 9551 8789
rect 9582 8780 9588 8792
rect 9640 8780 9646 8832
rect 11793 8823 11851 8829
rect 11793 8789 11805 8823
rect 11839 8820 11851 8823
rect 11882 8820 11888 8832
rect 11839 8792 11888 8820
rect 11839 8789 11851 8792
rect 11793 8783 11851 8789
rect 11882 8780 11888 8792
rect 11940 8780 11946 8832
rect 12989 8823 13047 8829
rect 12989 8789 13001 8823
rect 13035 8820 13047 8823
rect 13078 8820 13084 8832
rect 13035 8792 13084 8820
rect 13035 8789 13047 8792
rect 12989 8783 13047 8789
rect 13078 8780 13084 8792
rect 13136 8780 13142 8832
rect 14734 8820 14740 8832
rect 14695 8792 14740 8820
rect 14734 8780 14740 8792
rect 14792 8780 14798 8832
rect 24762 8820 24768 8832
rect 24723 8792 24768 8820
rect 24762 8780 24768 8792
rect 24820 8780 24826 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 1578 8616 1584 8628
rect 1539 8588 1584 8616
rect 1578 8576 1584 8588
rect 1636 8576 1642 8628
rect 2222 8576 2228 8628
rect 2280 8616 2286 8628
rect 2774 8616 2780 8628
rect 2280 8588 2780 8616
rect 2280 8576 2286 8588
rect 2774 8576 2780 8588
rect 2832 8576 2838 8628
rect 7282 8576 7288 8628
rect 7340 8616 7346 8628
rect 7745 8619 7803 8625
rect 7745 8616 7757 8619
rect 7340 8588 7757 8616
rect 7340 8576 7346 8588
rect 7745 8585 7757 8588
rect 7791 8585 7803 8619
rect 7745 8579 7803 8585
rect 8478 8576 8484 8628
rect 8536 8616 8542 8628
rect 8573 8619 8631 8625
rect 8573 8616 8585 8619
rect 8536 8588 8585 8616
rect 8536 8576 8542 8588
rect 8573 8585 8585 8588
rect 8619 8585 8631 8619
rect 8573 8579 8631 8585
rect 10042 8576 10048 8628
rect 10100 8616 10106 8628
rect 10229 8619 10287 8625
rect 10229 8616 10241 8619
rect 10100 8588 10241 8616
rect 10100 8576 10106 8588
rect 10229 8585 10241 8588
rect 10275 8585 10287 8619
rect 10229 8579 10287 8585
rect 10689 8619 10747 8625
rect 10689 8585 10701 8619
rect 10735 8616 10747 8619
rect 10778 8616 10784 8628
rect 10735 8588 10784 8616
rect 10735 8585 10747 8588
rect 10689 8579 10747 8585
rect 10778 8576 10784 8588
rect 10836 8576 10842 8628
rect 11333 8619 11391 8625
rect 11333 8585 11345 8619
rect 11379 8616 11391 8619
rect 12066 8616 12072 8628
rect 11379 8588 12072 8616
rect 11379 8585 11391 8588
rect 11333 8579 11391 8585
rect 9950 8508 9956 8560
rect 10008 8548 10014 8560
rect 10919 8551 10977 8557
rect 10919 8548 10931 8551
rect 10008 8520 10931 8548
rect 10008 8508 10014 8520
rect 10919 8517 10931 8520
rect 10965 8517 10977 8551
rect 10919 8511 10977 8517
rect 1302 8440 1308 8492
rect 1360 8480 1366 8492
rect 1578 8480 1584 8492
rect 1360 8452 1584 8480
rect 1360 8440 1366 8452
rect 1578 8440 1584 8452
rect 1636 8440 1642 8492
rect 2774 8440 2780 8492
rect 2832 8480 2838 8492
rect 2832 8452 2877 8480
rect 2832 8440 2838 8452
rect 3142 8440 3148 8492
rect 3200 8480 3206 8492
rect 3421 8483 3479 8489
rect 3421 8480 3433 8483
rect 3200 8452 3433 8480
rect 3200 8440 3206 8452
rect 3421 8449 3433 8452
rect 3467 8480 3479 8483
rect 3878 8480 3884 8492
rect 3467 8452 3884 8480
rect 3467 8449 3479 8452
rect 3421 8443 3479 8449
rect 3878 8440 3884 8452
rect 3936 8440 3942 8492
rect 11348 8424 11376 8579
rect 12066 8576 12072 8588
rect 12124 8576 12130 8628
rect 12618 8576 12624 8628
rect 12676 8576 12682 8628
rect 13354 8576 13360 8628
rect 13412 8616 13418 8628
rect 13449 8619 13507 8625
rect 13449 8616 13461 8619
rect 13412 8588 13461 8616
rect 13412 8576 13418 8588
rect 13449 8585 13461 8588
rect 13495 8585 13507 8619
rect 13449 8579 13507 8585
rect 15381 8619 15439 8625
rect 15381 8585 15393 8619
rect 15427 8616 15439 8619
rect 15746 8616 15752 8628
rect 15427 8588 15752 8616
rect 15427 8585 15439 8588
rect 15381 8579 15439 8585
rect 15746 8576 15752 8588
rect 15804 8576 15810 8628
rect 16574 8616 16580 8628
rect 16535 8588 16580 8616
rect 16574 8576 16580 8588
rect 16632 8576 16638 8628
rect 17586 8616 17592 8628
rect 17547 8588 17592 8616
rect 17586 8576 17592 8588
rect 17644 8576 17650 8628
rect 19334 8576 19340 8628
rect 19392 8616 19398 8628
rect 19613 8619 19671 8625
rect 19613 8616 19625 8619
rect 19392 8588 19625 8616
rect 19392 8576 19398 8588
rect 19613 8585 19625 8588
rect 19659 8585 19671 8619
rect 19613 8579 19671 8585
rect 20211 8619 20269 8625
rect 20211 8585 20223 8619
rect 20257 8616 20269 8619
rect 20622 8616 20628 8628
rect 20257 8588 20628 8616
rect 20257 8585 20269 8588
rect 20211 8579 20269 8585
rect 20622 8576 20628 8588
rect 20680 8576 20686 8628
rect 20990 8616 20996 8628
rect 20951 8588 20996 8616
rect 20990 8576 20996 8588
rect 21048 8576 21054 8628
rect 22094 8616 22100 8628
rect 22055 8588 22100 8616
rect 22094 8576 22100 8588
rect 22152 8576 22158 8628
rect 22557 8619 22615 8625
rect 22557 8585 22569 8619
rect 22603 8616 22615 8619
rect 22646 8616 22652 8628
rect 22603 8588 22652 8616
rect 22603 8585 22615 8588
rect 22557 8579 22615 8585
rect 22646 8576 22652 8588
rect 22704 8576 22710 8628
rect 25498 8616 25504 8628
rect 25459 8588 25504 8616
rect 25498 8576 25504 8588
rect 25556 8576 25562 8628
rect 11790 8508 11796 8560
rect 11848 8548 11854 8560
rect 11885 8551 11943 8557
rect 11885 8548 11897 8551
rect 11848 8520 11897 8548
rect 11848 8508 11854 8520
rect 11885 8517 11897 8520
rect 11931 8548 11943 8551
rect 12636 8548 12664 8576
rect 16206 8548 16212 8560
rect 11931 8520 12664 8548
rect 16167 8520 16212 8548
rect 11931 8517 11943 8520
rect 11885 8511 11943 8517
rect 16206 8508 16212 8520
rect 16264 8508 16270 8560
rect 19245 8551 19303 8557
rect 19245 8548 19257 8551
rect 18800 8520 19257 8548
rect 12434 8440 12440 8492
rect 12492 8480 12498 8492
rect 13909 8483 13967 8489
rect 12492 8452 12537 8480
rect 12492 8440 12498 8452
rect 13909 8449 13921 8483
rect 13955 8480 13967 8483
rect 14642 8480 14648 8492
rect 13955 8452 14648 8480
rect 13955 8449 13967 8452
rect 13909 8443 13967 8449
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8412 1455 8415
rect 1946 8412 1952 8424
rect 1443 8384 1952 8412
rect 1443 8381 1455 8384
rect 1397 8375 1455 8381
rect 1946 8372 1952 8384
rect 2004 8372 2010 8424
rect 3973 8415 4031 8421
rect 3973 8381 3985 8415
rect 4019 8412 4031 8415
rect 4801 8415 4859 8421
rect 4801 8412 4813 8415
rect 4019 8384 4813 8412
rect 4019 8381 4031 8384
rect 3973 8375 4031 8381
rect 4801 8381 4813 8384
rect 4847 8412 4859 8415
rect 4982 8412 4988 8424
rect 4847 8384 4988 8412
rect 4847 8381 4859 8384
rect 4801 8375 4859 8381
rect 4982 8372 4988 8384
rect 5040 8372 5046 8424
rect 5534 8372 5540 8424
rect 5592 8412 5598 8424
rect 5721 8415 5779 8421
rect 5721 8412 5733 8415
rect 5592 8384 5733 8412
rect 5592 8372 5598 8384
rect 5721 8381 5733 8384
rect 5767 8381 5779 8415
rect 6822 8412 6828 8424
rect 6783 8384 6828 8412
rect 5721 8375 5779 8381
rect 6822 8372 6828 8384
rect 6880 8372 6886 8424
rect 9033 8415 9091 8421
rect 9033 8381 9045 8415
rect 9079 8412 9091 8415
rect 9122 8412 9128 8424
rect 9079 8384 9128 8412
rect 9079 8381 9091 8384
rect 9033 8375 9091 8381
rect 9122 8372 9128 8384
rect 9180 8412 9186 8424
rect 9582 8412 9588 8424
rect 9180 8384 9588 8412
rect 9180 8372 9186 8384
rect 9582 8372 9588 8384
rect 9640 8372 9646 8424
rect 9953 8415 10011 8421
rect 9953 8381 9965 8415
rect 9999 8412 10011 8415
rect 10134 8412 10140 8424
rect 9999 8384 10140 8412
rect 9999 8381 10011 8384
rect 9953 8375 10011 8381
rect 10134 8372 10140 8384
rect 10192 8372 10198 8424
rect 10848 8415 10906 8421
rect 10848 8381 10860 8415
rect 10894 8412 10906 8415
rect 11330 8412 11336 8424
rect 10894 8384 11336 8412
rect 10894 8381 10906 8384
rect 10848 8375 10906 8381
rect 11330 8372 11336 8384
rect 11388 8372 11394 8424
rect 12253 8415 12311 8421
rect 12253 8381 12265 8415
rect 12299 8412 12311 8415
rect 13078 8412 13084 8424
rect 12299 8384 13084 8412
rect 12299 8381 12311 8384
rect 12253 8375 12311 8381
rect 13078 8372 13084 8384
rect 13136 8372 13142 8424
rect 14292 8421 14320 8452
rect 14642 8440 14648 8452
rect 14700 8440 14706 8492
rect 14737 8483 14795 8489
rect 14737 8449 14749 8483
rect 14783 8480 14795 8483
rect 15286 8480 15292 8492
rect 14783 8452 15292 8480
rect 14783 8449 14795 8452
rect 14737 8443 14795 8449
rect 15286 8440 15292 8452
rect 15344 8440 15350 8492
rect 15657 8483 15715 8489
rect 15657 8449 15669 8483
rect 15703 8480 15715 8483
rect 16390 8480 16396 8492
rect 15703 8452 16396 8480
rect 15703 8449 15715 8452
rect 15657 8443 15715 8449
rect 16390 8440 16396 8452
rect 16448 8440 16454 8492
rect 14277 8415 14335 8421
rect 14277 8381 14289 8415
rect 14323 8381 14335 8415
rect 14277 8375 14335 8381
rect 14553 8415 14611 8421
rect 14553 8381 14565 8415
rect 14599 8412 14611 8415
rect 18230 8412 18236 8424
rect 14599 8384 14780 8412
rect 18191 8384 18236 8412
rect 14599 8381 14611 8384
rect 14553 8375 14611 8381
rect 14752 8356 14780 8384
rect 18230 8372 18236 8384
rect 18288 8372 18294 8424
rect 18690 8372 18696 8424
rect 18748 8412 18754 8424
rect 18800 8421 18828 8520
rect 19245 8517 19257 8520
rect 19291 8548 19303 8551
rect 19702 8548 19708 8560
rect 19291 8520 19708 8548
rect 19291 8517 19303 8520
rect 19245 8511 19303 8517
rect 19702 8508 19708 8520
rect 19760 8508 19766 8560
rect 20530 8548 20536 8560
rect 20491 8520 20536 8548
rect 20530 8508 20536 8520
rect 20588 8508 20594 8560
rect 18969 8483 19027 8489
rect 18969 8449 18981 8483
rect 19015 8480 19027 8483
rect 19518 8480 19524 8492
rect 19015 8452 19524 8480
rect 19015 8449 19027 8452
rect 18969 8443 19027 8449
rect 19518 8440 19524 8452
rect 19576 8440 19582 8492
rect 18785 8415 18843 8421
rect 18785 8412 18797 8415
rect 18748 8384 18797 8412
rect 18748 8372 18754 8384
rect 18785 8381 18797 8384
rect 18831 8381 18843 8415
rect 18785 8375 18843 8381
rect 20140 8415 20198 8421
rect 20140 8381 20152 8415
rect 20186 8412 20198 8415
rect 20548 8412 20576 8508
rect 21358 8440 21364 8492
rect 21416 8480 21422 8492
rect 21453 8483 21511 8489
rect 21453 8480 21465 8483
rect 21416 8452 21465 8480
rect 21416 8440 21422 8452
rect 21453 8449 21465 8452
rect 21499 8449 21511 8483
rect 21453 8443 21511 8449
rect 22554 8440 22560 8492
rect 22612 8480 22618 8492
rect 22925 8483 22983 8489
rect 22925 8480 22937 8483
rect 22612 8452 22937 8480
rect 22612 8440 22618 8452
rect 22925 8449 22937 8452
rect 22971 8480 22983 8483
rect 24719 8483 24777 8489
rect 24719 8480 24731 8483
rect 22971 8452 24731 8480
rect 22971 8449 22983 8452
rect 22925 8443 22983 8449
rect 24719 8449 24731 8452
rect 24765 8449 24777 8483
rect 24719 8443 24777 8449
rect 20186 8384 20576 8412
rect 24632 8415 24690 8421
rect 20186 8381 20198 8384
rect 20140 8375 20198 8381
rect 24632 8381 24644 8415
rect 24678 8412 24690 8415
rect 24678 8384 24808 8412
rect 24678 8381 24690 8384
rect 24632 8375 24690 8381
rect 24780 8356 24808 8384
rect 2869 8347 2927 8353
rect 2869 8313 2881 8347
rect 2915 8344 2927 8347
rect 4062 8344 4068 8356
rect 2915 8316 4068 8344
rect 2915 8313 2927 8316
rect 2869 8307 2927 8313
rect 2222 8276 2228 8288
rect 2183 8248 2228 8276
rect 2222 8236 2228 8248
rect 2280 8236 2286 8288
rect 2593 8279 2651 8285
rect 2593 8245 2605 8279
rect 2639 8276 2651 8279
rect 2884 8276 2912 8307
rect 4062 8304 4068 8316
rect 4120 8304 4126 8356
rect 4341 8347 4399 8353
rect 4341 8313 4353 8347
rect 4387 8344 4399 8347
rect 4709 8347 4767 8353
rect 4709 8344 4721 8347
rect 4387 8316 4721 8344
rect 4387 8313 4399 8316
rect 4341 8307 4399 8313
rect 4709 8313 4721 8316
rect 4755 8344 4767 8347
rect 5163 8347 5221 8353
rect 5163 8344 5175 8347
rect 4755 8316 5175 8344
rect 4755 8313 4767 8316
rect 4709 8307 4767 8313
rect 5163 8313 5175 8316
rect 5209 8344 5221 8347
rect 5442 8344 5448 8356
rect 5209 8316 5448 8344
rect 5209 8313 5221 8316
rect 5163 8307 5221 8313
rect 5442 8304 5448 8316
rect 5500 8344 5506 8356
rect 7190 8353 7196 8356
rect 6273 8347 6331 8353
rect 6273 8344 6285 8347
rect 5500 8316 6285 8344
rect 5500 8304 5506 8316
rect 6273 8313 6285 8316
rect 6319 8344 6331 8347
rect 6641 8347 6699 8353
rect 6641 8344 6653 8347
rect 6319 8316 6653 8344
rect 6319 8313 6331 8316
rect 6273 8307 6331 8313
rect 6641 8313 6653 8316
rect 6687 8344 6699 8347
rect 7187 8344 7196 8353
rect 6687 8316 7196 8344
rect 6687 8313 6699 8316
rect 6641 8307 6699 8313
rect 7187 8307 7196 8316
rect 7248 8344 7254 8356
rect 9214 8344 9220 8356
rect 7248 8316 9220 8344
rect 7190 8304 7196 8307
rect 7248 8304 7254 8316
rect 9214 8304 9220 8316
rect 9272 8344 9278 8356
rect 9395 8347 9453 8353
rect 9395 8344 9407 8347
rect 9272 8316 9407 8344
rect 9272 8304 9278 8316
rect 9395 8313 9407 8316
rect 9441 8344 9453 8347
rect 10042 8344 10048 8356
rect 9441 8316 10048 8344
rect 9441 8313 9453 8316
rect 9395 8307 9453 8313
rect 10042 8304 10048 8316
rect 10100 8304 10106 8356
rect 14734 8304 14740 8356
rect 14792 8304 14798 8356
rect 15749 8347 15807 8353
rect 15749 8313 15761 8347
rect 15795 8344 15807 8347
rect 16114 8344 16120 8356
rect 15795 8316 16120 8344
rect 15795 8313 15807 8316
rect 15749 8307 15807 8313
rect 16114 8304 16120 8316
rect 16172 8304 16178 8356
rect 21174 8344 21180 8356
rect 21135 8316 21180 8344
rect 21174 8304 21180 8316
rect 21232 8304 21238 8356
rect 21266 8304 21272 8356
rect 21324 8344 21330 8356
rect 21324 8316 21369 8344
rect 21324 8304 21330 8316
rect 24762 8304 24768 8356
rect 24820 8344 24826 8356
rect 25041 8347 25099 8353
rect 25041 8344 25053 8347
rect 24820 8316 25053 8344
rect 24820 8304 24826 8316
rect 25041 8313 25053 8316
rect 25087 8313 25099 8347
rect 25041 8307 25099 8313
rect 2639 8248 2912 8276
rect 2639 8245 2651 8248
rect 2593 8239 2651 8245
rect 7926 8236 7932 8288
rect 7984 8276 7990 8288
rect 8021 8279 8079 8285
rect 8021 8276 8033 8279
rect 7984 8248 8033 8276
rect 7984 8236 7990 8248
rect 8021 8245 8033 8248
rect 8067 8245 8079 8279
rect 17126 8276 17132 8288
rect 17087 8248 17132 8276
rect 8021 8239 8079 8245
rect 17126 8236 17132 8248
rect 17184 8236 17190 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1535 8075 1593 8081
rect 1535 8041 1547 8075
rect 1581 8072 1593 8075
rect 1670 8072 1676 8084
rect 1581 8044 1676 8072
rect 1581 8041 1593 8044
rect 1535 8035 1593 8041
rect 1670 8032 1676 8044
rect 1728 8032 1734 8084
rect 1946 8072 1952 8084
rect 1907 8044 1952 8072
rect 1946 8032 1952 8044
rect 2004 8032 2010 8084
rect 2314 8072 2320 8084
rect 2275 8044 2320 8072
rect 2314 8032 2320 8044
rect 2372 8032 2378 8084
rect 2774 8032 2780 8084
rect 2832 8072 2838 8084
rect 3694 8072 3700 8084
rect 2832 8044 3700 8072
rect 2832 8032 2838 8044
rect 3694 8032 3700 8044
rect 3752 8072 3758 8084
rect 3789 8075 3847 8081
rect 3789 8072 3801 8075
rect 3752 8044 3801 8072
rect 3752 8032 3758 8044
rect 3789 8041 3801 8044
rect 3835 8041 3847 8075
rect 5626 8072 5632 8084
rect 5587 8044 5632 8072
rect 3789 8035 3847 8041
rect 5626 8032 5632 8044
rect 5684 8032 5690 8084
rect 6730 8072 6736 8084
rect 6288 8044 6736 8072
rect 2222 7964 2228 8016
rect 2280 8004 2286 8016
rect 2593 8007 2651 8013
rect 2593 8004 2605 8007
rect 2280 7976 2605 8004
rect 2280 7964 2286 7976
rect 2593 7973 2605 7976
rect 2639 8004 2651 8007
rect 2866 8004 2872 8016
rect 2639 7976 2872 8004
rect 2639 7973 2651 7976
rect 2593 7967 2651 7973
rect 2866 7964 2872 7976
rect 2924 7964 2930 8016
rect 3142 8004 3148 8016
rect 3103 7976 3148 8004
rect 3142 7964 3148 7976
rect 3200 7964 3206 8016
rect 4430 7964 4436 8016
rect 4488 8004 4494 8016
rect 4801 8007 4859 8013
rect 4801 8004 4813 8007
rect 4488 7976 4813 8004
rect 4488 7964 4494 7976
rect 4801 7973 4813 7976
rect 4847 8004 4859 8007
rect 5534 8004 5540 8016
rect 4847 7976 5540 8004
rect 4847 7973 4859 7976
rect 4801 7967 4859 7973
rect 5534 7964 5540 7976
rect 5592 7964 5598 8016
rect 6288 7948 6316 8044
rect 6730 8032 6736 8044
rect 6788 8032 6794 8084
rect 7466 8032 7472 8084
rect 7524 8072 7530 8084
rect 7975 8075 8033 8081
rect 7975 8072 7987 8075
rect 7524 8044 7987 8072
rect 7524 8032 7530 8044
rect 7975 8041 7987 8044
rect 8021 8041 8033 8075
rect 7975 8035 8033 8041
rect 9125 8075 9183 8081
rect 9125 8041 9137 8075
rect 9171 8072 9183 8075
rect 9214 8072 9220 8084
rect 9171 8044 9220 8072
rect 9171 8041 9183 8044
rect 9125 8035 9183 8041
rect 9214 8032 9220 8044
rect 9272 8032 9278 8084
rect 9674 8032 9680 8084
rect 9732 8072 9738 8084
rect 9769 8075 9827 8081
rect 9769 8072 9781 8075
rect 9732 8044 9781 8072
rect 9732 8032 9738 8044
rect 9769 8041 9781 8044
rect 9815 8041 9827 8075
rect 12158 8072 12164 8084
rect 12119 8044 12164 8072
rect 9769 8035 9827 8041
rect 12158 8032 12164 8044
rect 12216 8032 12222 8084
rect 14553 8075 14611 8081
rect 14553 8041 14565 8075
rect 14599 8072 14611 8075
rect 14734 8072 14740 8084
rect 14599 8044 14740 8072
rect 14599 8041 14611 8044
rect 14553 8035 14611 8041
rect 14734 8032 14740 8044
rect 14792 8032 14798 8084
rect 15562 8081 15568 8084
rect 15519 8075 15568 8081
rect 15519 8041 15531 8075
rect 15565 8041 15568 8075
rect 15519 8035 15568 8041
rect 15562 8032 15568 8035
rect 15620 8032 15626 8084
rect 15933 8075 15991 8081
rect 15933 8041 15945 8075
rect 15979 8072 15991 8075
rect 16114 8072 16120 8084
rect 15979 8044 16120 8072
rect 15979 8041 15991 8044
rect 15933 8035 15991 8041
rect 16114 8032 16120 8044
rect 16172 8032 16178 8084
rect 16301 8075 16359 8081
rect 16301 8041 16313 8075
rect 16347 8072 16359 8075
rect 16390 8072 16396 8084
rect 16347 8044 16396 8072
rect 16347 8041 16359 8044
rect 16301 8035 16359 8041
rect 16390 8032 16396 8044
rect 16448 8032 16454 8084
rect 17126 8072 17132 8084
rect 17087 8044 17132 8072
rect 17126 8032 17132 8044
rect 17184 8032 17190 8084
rect 18230 8072 18236 8084
rect 18191 8044 18236 8072
rect 18230 8032 18236 8044
rect 18288 8032 18294 8084
rect 18690 8072 18696 8084
rect 18651 8044 18696 8072
rect 18690 8032 18696 8044
rect 18748 8032 18754 8084
rect 19935 8075 19993 8081
rect 19935 8041 19947 8075
rect 19981 8072 19993 8075
rect 20438 8072 20444 8084
rect 19981 8044 20444 8072
rect 19981 8041 19993 8044
rect 19935 8035 19993 8041
rect 20438 8032 20444 8044
rect 20496 8032 20502 8084
rect 20717 8075 20775 8081
rect 20717 8041 20729 8075
rect 20763 8072 20775 8075
rect 21174 8072 21180 8084
rect 20763 8044 21180 8072
rect 20763 8041 20775 8044
rect 20717 8035 20775 8041
rect 21174 8032 21180 8044
rect 21232 8032 21238 8084
rect 21450 8072 21456 8084
rect 21284 8044 21456 8072
rect 6822 7964 6828 8016
rect 6880 8004 6886 8016
rect 7009 8007 7067 8013
rect 7009 8004 7021 8007
rect 6880 7976 7021 8004
rect 6880 7964 6886 7976
rect 7009 7973 7021 7976
rect 7055 8004 7067 8007
rect 7285 8007 7343 8013
rect 7285 8004 7297 8007
rect 7055 7976 7297 8004
rect 7055 7973 7067 7976
rect 7009 7967 7067 7973
rect 7285 7973 7297 7976
rect 7331 7973 7343 8007
rect 10870 8004 10876 8016
rect 7285 7967 7343 7973
rect 9968 7976 10876 8004
rect 9968 7948 9996 7976
rect 10870 7964 10876 7976
rect 10928 7964 10934 8016
rect 13633 8007 13691 8013
rect 13633 7973 13645 8007
rect 13679 8004 13691 8007
rect 14185 8007 14243 8013
rect 13679 7976 13952 8004
rect 13679 7973 13691 7976
rect 13633 7967 13691 7973
rect 1394 7896 1400 7948
rect 1452 7945 1458 7948
rect 1452 7939 1490 7945
rect 1478 7905 1490 7939
rect 6270 7936 6276 7948
rect 6231 7908 6276 7936
rect 1452 7899 1490 7905
rect 1452 7896 1458 7899
rect 6270 7896 6276 7908
rect 6328 7896 6334 7948
rect 6730 7936 6736 7948
rect 6691 7908 6736 7936
rect 6730 7896 6736 7908
rect 6788 7896 6794 7948
rect 7904 7939 7962 7945
rect 7904 7905 7916 7939
rect 7950 7936 7962 7939
rect 8110 7936 8116 7948
rect 7950 7908 8116 7936
rect 7950 7905 7962 7908
rect 7904 7899 7962 7905
rect 8110 7896 8116 7908
rect 8168 7896 8174 7948
rect 9950 7936 9956 7948
rect 9863 7908 9956 7936
rect 9950 7896 9956 7908
rect 10008 7896 10014 7948
rect 10042 7896 10048 7948
rect 10100 7936 10106 7948
rect 10229 7939 10287 7945
rect 10229 7936 10241 7939
rect 10100 7908 10241 7936
rect 10100 7896 10106 7908
rect 10229 7905 10241 7908
rect 10275 7936 10287 7939
rect 10962 7936 10968 7948
rect 10275 7908 10968 7936
rect 10275 7905 10287 7908
rect 10229 7899 10287 7905
rect 10962 7896 10968 7908
rect 11020 7896 11026 7948
rect 11882 7936 11888 7948
rect 11843 7908 11888 7936
rect 11882 7896 11888 7908
rect 11940 7896 11946 7948
rect 11974 7896 11980 7948
rect 12032 7936 12038 7948
rect 12069 7939 12127 7945
rect 12069 7936 12081 7939
rect 12032 7908 12081 7936
rect 12032 7896 12038 7908
rect 12069 7905 12081 7908
rect 12115 7905 12127 7939
rect 12069 7899 12127 7905
rect 13538 7896 13544 7948
rect 13596 7936 13602 7948
rect 13817 7939 13875 7945
rect 13817 7936 13829 7939
rect 13596 7908 13829 7936
rect 13596 7896 13602 7908
rect 13817 7905 13829 7908
rect 13863 7905 13875 7939
rect 13924 7936 13952 7976
rect 14185 7973 14197 8007
rect 14231 8004 14243 8007
rect 14366 8004 14372 8016
rect 14231 7976 14372 8004
rect 14231 7973 14243 7976
rect 14185 7967 14243 7973
rect 14366 7964 14372 7976
rect 14424 7964 14430 8016
rect 14550 7936 14556 7948
rect 13924 7908 14556 7936
rect 13817 7899 13875 7905
rect 14550 7896 14556 7908
rect 14608 7896 14614 7948
rect 15378 7896 15384 7948
rect 15436 7945 15442 7948
rect 15436 7939 15474 7945
rect 15462 7905 15474 7939
rect 17034 7936 17040 7948
rect 16995 7908 17040 7936
rect 15436 7899 15474 7905
rect 15436 7896 15442 7899
rect 17034 7896 17040 7908
rect 17092 7896 17098 7948
rect 17494 7896 17500 7948
rect 17552 7936 17558 7948
rect 17589 7939 17647 7945
rect 17589 7936 17601 7939
rect 17552 7908 17601 7936
rect 17552 7896 17558 7908
rect 17589 7905 17601 7908
rect 17635 7936 17647 7939
rect 18708 7936 18736 8032
rect 21284 8013 21312 8044
rect 21450 8032 21456 8044
rect 21508 8032 21514 8084
rect 23474 8032 23480 8084
rect 23532 8072 23538 8084
rect 24719 8075 24777 8081
rect 24719 8072 24731 8075
rect 23532 8044 24731 8072
rect 23532 8032 23538 8044
rect 24719 8041 24731 8044
rect 24765 8041 24777 8075
rect 24719 8035 24777 8041
rect 21269 8007 21327 8013
rect 21269 7973 21281 8007
rect 21315 7973 21327 8007
rect 21269 7967 21327 7973
rect 21358 7964 21364 8016
rect 21416 8004 21422 8016
rect 21821 8007 21879 8013
rect 21821 8004 21833 8007
rect 21416 7976 21833 8004
rect 21416 7964 21422 7976
rect 21821 7973 21833 7976
rect 21867 7973 21879 8007
rect 21821 7967 21879 7973
rect 23615 8007 23673 8013
rect 23615 7973 23627 8007
rect 23661 8004 23673 8007
rect 24486 8004 24492 8016
rect 23661 7976 24492 8004
rect 23661 7973 23673 7976
rect 23615 7967 23673 7973
rect 24486 7964 24492 7976
rect 24544 7964 24550 8016
rect 19886 7945 19892 7948
rect 19864 7939 19892 7945
rect 19864 7936 19876 7939
rect 17635 7908 18736 7936
rect 19799 7908 19876 7936
rect 17635 7905 17647 7908
rect 17589 7899 17647 7905
rect 19864 7905 19876 7908
rect 19944 7936 19950 7948
rect 20346 7936 20352 7948
rect 19944 7908 20352 7936
rect 19864 7899 19892 7905
rect 19886 7896 19892 7899
rect 19944 7896 19950 7908
rect 20346 7896 20352 7908
rect 20404 7896 20410 7948
rect 23528 7939 23586 7945
rect 23528 7905 23540 7939
rect 23574 7936 23586 7939
rect 23750 7936 23756 7948
rect 23574 7908 23756 7936
rect 23574 7905 23586 7908
rect 23528 7899 23586 7905
rect 23750 7896 23756 7908
rect 23808 7896 23814 7948
rect 24670 7945 24676 7948
rect 24648 7939 24676 7945
rect 24648 7905 24660 7939
rect 24648 7899 24676 7905
rect 24670 7896 24676 7899
rect 24728 7896 24734 7948
rect 2501 7871 2559 7877
rect 2501 7868 2513 7871
rect 2424 7840 2513 7868
rect 2424 7744 2452 7840
rect 2501 7837 2513 7840
rect 2547 7837 2559 7871
rect 4706 7868 4712 7880
rect 4667 7840 4712 7868
rect 2501 7831 2559 7837
rect 4706 7828 4712 7840
rect 4764 7828 4770 7880
rect 4890 7828 4896 7880
rect 4948 7868 4954 7880
rect 4985 7871 5043 7877
rect 4985 7868 4997 7871
rect 4948 7840 4997 7868
rect 4948 7828 4954 7840
rect 4985 7837 4997 7840
rect 5031 7837 5043 7871
rect 4985 7831 5043 7837
rect 21177 7871 21235 7877
rect 21177 7837 21189 7871
rect 21223 7868 21235 7871
rect 21542 7868 21548 7880
rect 21223 7840 21548 7868
rect 21223 7837 21235 7840
rect 21177 7831 21235 7837
rect 21542 7828 21548 7840
rect 21600 7828 21606 7880
rect 2406 7692 2412 7744
rect 2464 7692 2470 7744
rect 2774 7692 2780 7744
rect 2832 7732 2838 7744
rect 3510 7732 3516 7744
rect 2832 7704 3516 7732
rect 2832 7692 2838 7704
rect 3510 7692 3516 7704
rect 3568 7692 3574 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 1394 7488 1400 7540
rect 1452 7528 1458 7540
rect 2317 7531 2375 7537
rect 2317 7528 2329 7531
rect 1452 7500 2329 7528
rect 1452 7488 1458 7500
rect 2317 7497 2329 7500
rect 2363 7497 2375 7531
rect 2317 7491 2375 7497
rect 2777 7531 2835 7537
rect 2777 7497 2789 7531
rect 2823 7528 2835 7531
rect 2866 7528 2872 7540
rect 2823 7500 2872 7528
rect 2823 7497 2835 7500
rect 2777 7491 2835 7497
rect 2866 7488 2872 7500
rect 2924 7488 2930 7540
rect 4430 7528 4436 7540
rect 4391 7500 4436 7528
rect 4430 7488 4436 7500
rect 4488 7488 4494 7540
rect 4798 7528 4804 7540
rect 4759 7500 4804 7528
rect 4798 7488 4804 7500
rect 4856 7488 4862 7540
rect 6086 7488 6092 7540
rect 6144 7528 6150 7540
rect 6549 7531 6607 7537
rect 6549 7528 6561 7531
rect 6144 7500 6561 7528
rect 6144 7488 6150 7500
rect 6549 7497 6561 7500
rect 6595 7497 6607 7531
rect 6549 7491 6607 7497
rect 7929 7531 7987 7537
rect 7929 7497 7941 7531
rect 7975 7528 7987 7531
rect 8110 7528 8116 7540
rect 7975 7500 8116 7528
rect 7975 7497 7987 7500
rect 7929 7491 7987 7497
rect 1486 7420 1492 7472
rect 1544 7460 1550 7472
rect 1581 7463 1639 7469
rect 1581 7460 1593 7463
rect 1544 7432 1593 7460
rect 1544 7420 1550 7432
rect 1581 7429 1593 7432
rect 1627 7429 1639 7463
rect 2038 7460 2044 7472
rect 1999 7432 2044 7460
rect 1581 7423 1639 7429
rect 2038 7420 2044 7432
rect 2096 7420 2102 7472
rect 6270 7460 6276 7472
rect 6231 7432 6276 7460
rect 6270 7420 6276 7432
rect 6328 7420 6334 7472
rect 1397 7327 1455 7333
rect 1397 7293 1409 7327
rect 1443 7324 1455 7327
rect 2056 7324 2084 7420
rect 3878 7392 3884 7404
rect 3839 7364 3884 7392
rect 3878 7352 3884 7364
rect 3936 7352 3942 7404
rect 1443 7296 2084 7324
rect 1443 7293 1455 7296
rect 1397 7287 1455 7293
rect 4798 7284 4804 7336
rect 4856 7324 4862 7336
rect 4893 7327 4951 7333
rect 4893 7324 4905 7327
rect 4856 7296 4905 7324
rect 4856 7284 4862 7296
rect 4893 7293 4905 7296
rect 4939 7293 4951 7327
rect 4893 7287 4951 7293
rect 5445 7327 5503 7333
rect 5445 7293 5457 7327
rect 5491 7293 5503 7327
rect 6564 7324 6592 7491
rect 8110 7488 8116 7500
rect 8168 7488 8174 7540
rect 8570 7537 8576 7540
rect 8527 7531 8576 7537
rect 8527 7497 8539 7531
rect 8573 7497 8576 7531
rect 8527 7491 8576 7497
rect 8570 7488 8576 7491
rect 8628 7488 8634 7540
rect 9769 7531 9827 7537
rect 9769 7497 9781 7531
rect 9815 7528 9827 7531
rect 9950 7528 9956 7540
rect 9815 7500 9956 7528
rect 9815 7497 9827 7500
rect 9769 7491 9827 7497
rect 9950 7488 9956 7500
rect 10008 7488 10014 7540
rect 10183 7531 10241 7537
rect 10183 7497 10195 7531
rect 10229 7528 10241 7531
rect 10318 7528 10324 7540
rect 10229 7500 10324 7528
rect 10229 7497 10241 7500
rect 10183 7491 10241 7497
rect 10318 7488 10324 7500
rect 10376 7488 10382 7540
rect 11054 7488 11060 7540
rect 11112 7528 11118 7540
rect 11241 7531 11299 7537
rect 11241 7528 11253 7531
rect 11112 7500 11253 7528
rect 11112 7488 11118 7500
rect 11241 7497 11253 7500
rect 11287 7497 11299 7531
rect 11974 7528 11980 7540
rect 11935 7500 11980 7528
rect 11241 7491 11299 7497
rect 11974 7488 11980 7500
rect 12032 7488 12038 7540
rect 12618 7528 12624 7540
rect 12579 7500 12624 7528
rect 12618 7488 12624 7500
rect 12676 7488 12682 7540
rect 13538 7528 13544 7540
rect 13499 7500 13544 7528
rect 13538 7488 13544 7500
rect 13596 7488 13602 7540
rect 13909 7531 13967 7537
rect 13909 7497 13921 7531
rect 13955 7528 13967 7531
rect 14734 7528 14740 7540
rect 13955 7500 14740 7528
rect 13955 7497 13967 7500
rect 13909 7491 13967 7497
rect 14734 7488 14740 7500
rect 14792 7488 14798 7540
rect 17034 7528 17040 7540
rect 16995 7500 17040 7528
rect 17034 7488 17040 7500
rect 17092 7488 17098 7540
rect 17494 7528 17500 7540
rect 17455 7500 17500 7528
rect 17494 7488 17500 7500
rect 17552 7488 17558 7540
rect 19886 7528 19892 7540
rect 19847 7500 19892 7528
rect 19886 7488 19892 7500
rect 19944 7488 19950 7540
rect 21177 7531 21235 7537
rect 21177 7497 21189 7531
rect 21223 7528 21235 7531
rect 21450 7528 21456 7540
rect 21223 7500 21456 7528
rect 21223 7497 21235 7500
rect 21177 7491 21235 7497
rect 21450 7488 21456 7500
rect 21508 7488 21514 7540
rect 23750 7488 23756 7540
rect 23808 7528 23814 7540
rect 23845 7531 23903 7537
rect 23845 7528 23857 7531
rect 23808 7500 23857 7528
rect 23808 7488 23814 7500
rect 23845 7497 23857 7500
rect 23891 7497 23903 7531
rect 24670 7528 24676 7540
rect 24631 7500 24676 7528
rect 23845 7491 23903 7497
rect 24670 7488 24676 7500
rect 24728 7488 24734 7540
rect 6730 7420 6736 7472
rect 6788 7460 6794 7472
rect 9401 7463 9459 7469
rect 9401 7460 9413 7463
rect 6788 7432 9413 7460
rect 6788 7420 6794 7432
rect 7392 7333 7420 7432
rect 9401 7429 9413 7432
rect 9447 7460 9459 7463
rect 10042 7460 10048 7472
rect 9447 7432 10048 7460
rect 9447 7429 9459 7432
rect 9401 7423 9459 7429
rect 10042 7420 10048 7432
rect 10100 7420 10106 7472
rect 11609 7463 11667 7469
rect 11609 7429 11621 7463
rect 11655 7460 11667 7463
rect 12342 7460 12348 7472
rect 11655 7432 12348 7460
rect 11655 7429 11667 7432
rect 11609 7423 11667 7429
rect 7561 7395 7619 7401
rect 7561 7361 7573 7395
rect 7607 7392 7619 7395
rect 7926 7392 7932 7404
rect 7607 7364 7932 7392
rect 7607 7361 7619 7364
rect 7561 7355 7619 7361
rect 7926 7352 7932 7364
rect 7984 7352 7990 7404
rect 6825 7327 6883 7333
rect 6825 7324 6837 7327
rect 6564 7296 6837 7324
rect 5445 7287 5503 7293
rect 6825 7293 6837 7296
rect 6871 7293 6883 7327
rect 6825 7287 6883 7293
rect 7377 7327 7435 7333
rect 7377 7293 7389 7327
rect 7423 7293 7435 7327
rect 7377 7287 7435 7293
rect 2958 7216 2964 7268
rect 3016 7256 3022 7268
rect 3237 7259 3295 7265
rect 3237 7256 3249 7259
rect 3016 7228 3249 7256
rect 3016 7216 3022 7228
rect 3237 7225 3249 7228
rect 3283 7256 3295 7259
rect 3421 7259 3479 7265
rect 3421 7256 3433 7259
rect 3283 7228 3433 7256
rect 3283 7225 3295 7228
rect 3237 7219 3295 7225
rect 3421 7225 3433 7228
rect 3467 7225 3479 7259
rect 3421 7219 3479 7225
rect 3513 7259 3571 7265
rect 3513 7225 3525 7259
rect 3559 7256 3571 7259
rect 3602 7256 3608 7268
rect 3559 7228 3608 7256
rect 3559 7225 3571 7228
rect 3513 7219 3571 7225
rect 3602 7216 3608 7228
rect 3660 7216 3666 7268
rect 5460 7256 5488 7287
rect 8386 7284 8392 7336
rect 8444 7333 8450 7336
rect 8444 7327 8482 7333
rect 8470 7324 8482 7327
rect 8849 7327 8907 7333
rect 8849 7324 8861 7327
rect 8470 7296 8861 7324
rect 8470 7293 8482 7296
rect 8444 7287 8482 7293
rect 8849 7293 8861 7296
rect 8895 7293 8907 7327
rect 8849 7287 8907 7293
rect 8444 7284 8450 7287
rect 9858 7284 9864 7336
rect 9916 7324 9922 7336
rect 10080 7327 10138 7333
rect 10080 7324 10092 7327
rect 9916 7296 10092 7324
rect 9916 7284 9922 7296
rect 10080 7293 10092 7296
rect 10126 7324 10138 7327
rect 10505 7327 10563 7333
rect 10505 7324 10517 7327
rect 10126 7296 10517 7324
rect 10126 7293 10138 7296
rect 10080 7287 10138 7293
rect 10505 7293 10517 7296
rect 10551 7293 10563 7327
rect 10505 7287 10563 7293
rect 11057 7327 11115 7333
rect 11057 7293 11069 7327
rect 11103 7324 11115 7327
rect 11624 7324 11652 7423
rect 12342 7420 12348 7432
rect 12400 7420 12406 7472
rect 14277 7463 14335 7469
rect 14277 7429 14289 7463
rect 14323 7460 14335 7463
rect 14550 7460 14556 7472
rect 14323 7432 14556 7460
rect 14323 7429 14335 7432
rect 14277 7423 14335 7429
rect 14550 7420 14556 7432
rect 14608 7420 14614 7472
rect 24118 7352 24124 7404
rect 24176 7392 24182 7404
rect 24670 7392 24676 7404
rect 24176 7364 24676 7392
rect 24176 7352 24182 7364
rect 24670 7352 24676 7364
rect 24728 7352 24734 7404
rect 11103 7296 11652 7324
rect 12437 7327 12495 7333
rect 11103 7293 11115 7296
rect 11057 7287 11115 7293
rect 12437 7293 12449 7327
rect 12483 7324 12495 7327
rect 12526 7324 12532 7336
rect 12483 7296 12532 7324
rect 12483 7293 12495 7296
rect 12437 7287 12495 7293
rect 12526 7284 12532 7296
rect 12584 7324 12590 7336
rect 12897 7327 12955 7333
rect 12897 7324 12909 7327
rect 12584 7296 12909 7324
rect 12584 7284 12590 7296
rect 12897 7293 12909 7296
rect 12943 7293 12955 7327
rect 12897 7287 12955 7293
rect 13725 7327 13783 7333
rect 13725 7293 13737 7327
rect 13771 7324 13783 7327
rect 13906 7324 13912 7336
rect 13771 7296 13912 7324
rect 13771 7293 13783 7296
rect 13725 7287 13783 7293
rect 13906 7284 13912 7296
rect 13964 7324 13970 7336
rect 14553 7327 14611 7333
rect 14553 7324 14565 7327
rect 13964 7296 14565 7324
rect 13964 7284 13970 7296
rect 14553 7293 14565 7296
rect 14599 7293 14611 7327
rect 15378 7324 15384 7336
rect 15339 7296 15384 7324
rect 14553 7287 14611 7293
rect 15378 7284 15384 7296
rect 15436 7284 15442 7336
rect 6730 7256 6736 7268
rect 5460 7228 6736 7256
rect 6730 7216 6736 7228
rect 6788 7216 6794 7268
rect 4982 7188 4988 7200
rect 4943 7160 4988 7188
rect 4982 7148 4988 7160
rect 5040 7148 5046 7200
rect 21542 7188 21548 7200
rect 21503 7160 21548 7188
rect 21542 7148 21548 7160
rect 21600 7148 21606 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 2958 6984 2964 6996
rect 2919 6956 2964 6984
rect 2958 6944 2964 6956
rect 3016 6944 3022 6996
rect 3510 6944 3516 6996
rect 3568 6984 3574 6996
rect 4203 6987 4261 6993
rect 4203 6984 4215 6987
rect 3568 6956 4215 6984
rect 3568 6944 3574 6956
rect 4203 6953 4215 6956
rect 4249 6953 4261 6987
rect 4203 6947 4261 6953
rect 4617 6987 4675 6993
rect 4617 6953 4629 6987
rect 4663 6984 4675 6987
rect 4706 6984 4712 6996
rect 4663 6956 4712 6984
rect 4663 6953 4675 6956
rect 4617 6947 4675 6953
rect 4706 6944 4712 6956
rect 4764 6944 4770 6996
rect 4798 6944 4804 6996
rect 4856 6984 4862 6996
rect 4985 6987 5043 6993
rect 4985 6984 4997 6987
rect 4856 6956 4997 6984
rect 4856 6944 4862 6956
rect 4985 6953 4997 6956
rect 5031 6984 5043 6987
rect 6365 6987 6423 6993
rect 6365 6984 6377 6987
rect 5031 6956 6377 6984
rect 5031 6953 5043 6956
rect 4985 6947 5043 6953
rect 6365 6953 6377 6956
rect 6411 6984 6423 6987
rect 6730 6984 6736 6996
rect 6411 6956 6736 6984
rect 6411 6953 6423 6956
rect 6365 6947 6423 6953
rect 6730 6944 6736 6956
rect 6788 6984 6794 6996
rect 6825 6987 6883 6993
rect 6825 6984 6837 6987
rect 6788 6956 6837 6984
rect 6788 6944 6794 6956
rect 6825 6953 6837 6956
rect 6871 6953 6883 6987
rect 11882 6984 11888 6996
rect 11843 6956 11888 6984
rect 6825 6947 6883 6953
rect 11882 6944 11888 6956
rect 11940 6944 11946 6996
rect 8110 6876 8116 6928
rect 8168 6916 8174 6928
rect 8168 6888 8248 6916
rect 8168 6876 8174 6888
rect 1397 6851 1455 6857
rect 1397 6817 1409 6851
rect 1443 6848 1455 6851
rect 1578 6848 1584 6860
rect 1443 6820 1584 6848
rect 1443 6817 1455 6820
rect 1397 6811 1455 6817
rect 1578 6808 1584 6820
rect 1636 6808 1642 6860
rect 3513 6851 3571 6857
rect 3513 6817 3525 6851
rect 3559 6848 3571 6851
rect 3602 6848 3608 6860
rect 3559 6820 3608 6848
rect 3559 6817 3571 6820
rect 3513 6811 3571 6817
rect 3602 6808 3608 6820
rect 3660 6808 3666 6860
rect 4154 6857 4160 6860
rect 4132 6851 4160 6857
rect 4132 6848 4144 6851
rect 4067 6820 4144 6848
rect 4132 6817 4144 6820
rect 4212 6848 4218 6860
rect 4522 6848 4528 6860
rect 4212 6820 4528 6848
rect 4132 6811 4160 6817
rect 4154 6808 4160 6811
rect 4212 6808 4218 6820
rect 4522 6808 4528 6820
rect 4580 6808 4586 6860
rect 5074 6808 5080 6860
rect 5132 6857 5138 6860
rect 5258 6857 5264 6860
rect 5132 6851 5170 6857
rect 5158 6817 5170 6851
rect 5132 6811 5170 6817
rect 5215 6851 5264 6857
rect 5215 6817 5227 6851
rect 5261 6817 5264 6851
rect 5215 6811 5264 6817
rect 5132 6808 5138 6811
rect 5258 6808 5264 6811
rect 5316 6808 5322 6860
rect 7374 6857 7380 6860
rect 7352 6851 7380 6857
rect 7352 6817 7364 6851
rect 7352 6811 7380 6817
rect 7374 6808 7380 6811
rect 7432 6808 7438 6860
rect 8220 6848 8248 6888
rect 8294 6848 8300 6860
rect 8352 6857 8358 6860
rect 10318 6857 10324 6860
rect 8352 6851 8390 6857
rect 8207 6820 8300 6848
rect 8294 6808 8300 6820
rect 8378 6817 8390 6851
rect 8352 6811 8390 6817
rect 10296 6851 10324 6857
rect 10296 6817 10308 6851
rect 10296 6811 10324 6817
rect 8352 6808 8358 6811
rect 10318 6808 10324 6811
rect 10376 6808 10382 6860
rect 11330 6808 11336 6860
rect 11388 6857 11394 6860
rect 11514 6857 11520 6860
rect 11388 6851 11426 6857
rect 11414 6817 11426 6851
rect 11388 6811 11426 6817
rect 11471 6851 11520 6857
rect 11471 6817 11483 6851
rect 11517 6817 11520 6851
rect 11471 6811 11520 6817
rect 11388 6808 11394 6811
rect 11514 6808 11520 6811
rect 11572 6808 11578 6860
rect 1581 6715 1639 6721
rect 1581 6681 1593 6715
rect 1627 6712 1639 6715
rect 2866 6712 2872 6724
rect 1627 6684 2872 6712
rect 1627 6681 1639 6684
rect 1581 6675 1639 6681
rect 2866 6672 2872 6684
rect 2924 6672 2930 6724
rect 7423 6715 7481 6721
rect 7423 6681 7435 6715
rect 7469 6712 7481 6715
rect 8018 6712 8024 6724
rect 7469 6684 8024 6712
rect 7469 6681 7481 6684
rect 7423 6675 7481 6681
rect 8018 6672 8024 6684
rect 8076 6672 8082 6724
rect 8435 6715 8493 6721
rect 8435 6681 8447 6715
rect 8481 6712 8493 6715
rect 9582 6712 9588 6724
rect 8481 6684 9588 6712
rect 8481 6681 8493 6684
rect 8435 6675 8493 6681
rect 9582 6672 9588 6684
rect 9640 6672 9646 6724
rect 9766 6672 9772 6724
rect 9824 6712 9830 6724
rect 10367 6715 10425 6721
rect 10367 6712 10379 6715
rect 9824 6684 10379 6712
rect 9824 6672 9830 6684
rect 10367 6681 10379 6684
rect 10413 6681 10425 6715
rect 10367 6675 10425 6681
rect 2406 6644 2412 6656
rect 2367 6616 2412 6644
rect 2406 6604 2412 6616
rect 2464 6604 2470 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6440 1639 6443
rect 1762 6440 1768 6452
rect 1627 6412 1768 6440
rect 1627 6409 1639 6412
rect 1581 6403 1639 6409
rect 1762 6400 1768 6412
rect 1820 6400 1826 6452
rect 2038 6440 2044 6452
rect 1999 6412 2044 6440
rect 2038 6400 2044 6412
rect 2096 6400 2102 6452
rect 3694 6449 3700 6452
rect 3651 6443 3700 6449
rect 3651 6409 3663 6443
rect 3697 6409 3700 6443
rect 3651 6403 3700 6409
rect 3694 6400 3700 6403
rect 3752 6400 3758 6452
rect 4154 6440 4160 6452
rect 4115 6412 4160 6440
rect 4154 6400 4160 6412
rect 4212 6400 4218 6452
rect 5074 6440 5080 6452
rect 5035 6412 5080 6440
rect 5074 6400 5080 6412
rect 5132 6400 5138 6452
rect 7374 6440 7380 6452
rect 7335 6412 7380 6440
rect 7374 6400 7380 6412
rect 7432 6400 7438 6452
rect 8294 6440 8300 6452
rect 8255 6412 8300 6440
rect 8294 6400 8300 6412
rect 8352 6400 8358 6452
rect 10318 6440 10324 6452
rect 10279 6412 10324 6440
rect 10318 6400 10324 6412
rect 10376 6400 10382 6452
rect 11330 6440 11336 6452
rect 11291 6412 11336 6440
rect 11330 6400 11336 6412
rect 11388 6400 11394 6452
rect 1578 6264 1584 6316
rect 1636 6304 1642 6316
rect 2317 6307 2375 6313
rect 2317 6304 2329 6307
rect 1636 6276 2329 6304
rect 1636 6264 1642 6276
rect 2317 6273 2329 6276
rect 2363 6273 2375 6307
rect 2498 6304 2504 6316
rect 2459 6276 2504 6304
rect 2317 6267 2375 6273
rect 2498 6264 2504 6276
rect 2556 6264 2562 6316
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6236 1455 6239
rect 2038 6236 2044 6248
rect 1443 6208 2044 6236
rect 1443 6205 1455 6208
rect 1397 6199 1455 6205
rect 2038 6196 2044 6208
rect 2096 6196 2102 6248
rect 3548 6239 3606 6245
rect 3548 6236 3560 6239
rect 3344 6208 3560 6236
rect 3344 6112 3372 6208
rect 3548 6205 3560 6208
rect 3594 6205 3606 6239
rect 3548 6199 3606 6205
rect 3326 6100 3332 6112
rect 3287 6072 3332 6100
rect 3326 6060 3332 6072
rect 3384 6060 3390 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 1394 5856 1400 5908
rect 1452 5896 1458 5908
rect 2590 5905 2596 5908
rect 1535 5899 1593 5905
rect 1535 5896 1547 5899
rect 1452 5868 1547 5896
rect 1452 5856 1458 5868
rect 1535 5865 1547 5868
rect 1581 5865 1593 5899
rect 1535 5859 1593 5865
rect 2547 5899 2596 5905
rect 2547 5865 2559 5899
rect 2593 5865 2596 5899
rect 2547 5859 2596 5865
rect 2590 5856 2596 5859
rect 2648 5856 2654 5908
rect 1394 5720 1400 5772
rect 1452 5769 1458 5772
rect 2498 5769 2504 5772
rect 1452 5763 1490 5769
rect 1478 5729 1490 5763
rect 1452 5723 1490 5729
rect 2476 5763 2504 5769
rect 2476 5729 2488 5763
rect 2476 5723 2504 5729
rect 1452 5720 1458 5723
rect 2498 5720 2504 5723
rect 2556 5720 2562 5772
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 1394 5312 1400 5364
rect 1452 5352 1458 5364
rect 1857 5355 1915 5361
rect 1857 5352 1869 5355
rect 1452 5324 1869 5352
rect 1452 5312 1458 5324
rect 1857 5321 1869 5324
rect 1903 5321 1915 5355
rect 1857 5315 1915 5321
rect 2498 5312 2504 5364
rect 2556 5352 2562 5364
rect 2593 5355 2651 5361
rect 2593 5352 2605 5355
rect 2556 5324 2605 5352
rect 2556 5312 2562 5324
rect 2593 5321 2605 5324
rect 2639 5321 2651 5355
rect 2593 5315 2651 5321
rect 1535 5287 1593 5293
rect 1535 5253 1547 5287
rect 1581 5284 1593 5287
rect 2406 5284 2412 5296
rect 1581 5256 2412 5284
rect 1581 5253 1593 5256
rect 1535 5247 1593 5253
rect 2406 5244 2412 5256
rect 2464 5244 2470 5296
rect 1486 5157 1492 5160
rect 1464 5151 1492 5157
rect 1464 5117 1476 5151
rect 1544 5148 1550 5160
rect 2225 5151 2283 5157
rect 2225 5148 2237 5151
rect 1544 5120 2237 5148
rect 1464 5111 1492 5117
rect 1486 5108 1492 5111
rect 1544 5108 1550 5120
rect 2225 5117 2237 5120
rect 2271 5117 2283 5151
rect 2225 5111 2283 5117
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1535 4811 1593 4817
rect 1535 4777 1547 4811
rect 1581 4808 1593 4811
rect 2130 4808 2136 4820
rect 1581 4780 2136 4808
rect 1581 4777 1593 4780
rect 1535 4771 1593 4777
rect 2130 4768 2136 4780
rect 2188 4768 2194 4820
rect 1394 4632 1400 4684
rect 1452 4681 1458 4684
rect 1452 4675 1490 4681
rect 1478 4641 1490 4675
rect 1452 4635 1490 4641
rect 1452 4632 1458 4635
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 1394 4224 1400 4276
rect 1452 4264 1458 4276
rect 1581 4267 1639 4273
rect 1581 4264 1593 4267
rect 1452 4236 1593 4264
rect 1452 4224 1458 4236
rect 1581 4233 1593 4236
rect 1627 4233 1639 4267
rect 1581 4227 1639 4233
rect 10686 4156 10692 4208
rect 10744 4196 10750 4208
rect 10870 4196 10876 4208
rect 10744 4168 10876 4196
rect 10744 4156 10750 4168
rect 10870 4156 10876 4168
rect 10928 4156 10934 4208
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1535 3179 1593 3185
rect 1535 3145 1547 3179
rect 1581 3176 1593 3179
rect 1854 3176 1860 3188
rect 1581 3148 1860 3176
rect 1581 3145 1593 3148
rect 1535 3139 1593 3145
rect 1854 3136 1860 3148
rect 1912 3136 1918 3188
rect 24670 3136 24676 3188
rect 24728 3185 24734 3188
rect 24728 3179 24777 3185
rect 24728 3145 24731 3179
rect 24765 3145 24777 3179
rect 24728 3139 24777 3145
rect 24728 3136 24734 3139
rect 1486 2981 1492 2984
rect 1464 2975 1492 2981
rect 1464 2972 1476 2975
rect 1399 2944 1476 2972
rect 1464 2941 1476 2944
rect 1544 2972 1550 2984
rect 1857 2975 1915 2981
rect 1857 2972 1869 2975
rect 1544 2944 1869 2972
rect 1464 2935 1492 2941
rect 1486 2932 1492 2935
rect 1544 2932 1550 2944
rect 1857 2941 1869 2944
rect 1903 2941 1915 2975
rect 1857 2935 1915 2941
rect 24648 2975 24706 2981
rect 24648 2941 24660 2975
rect 24694 2972 24706 2975
rect 24694 2944 25176 2972
rect 24694 2941 24706 2944
rect 24648 2935 24706 2941
rect 25148 2848 25176 2944
rect 25130 2836 25136 2848
rect 25091 2808 25136 2836
rect 25130 2796 25136 2808
rect 25188 2796 25194 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 1535 2635 1593 2641
rect 1535 2601 1547 2635
rect 1581 2632 1593 2635
rect 1946 2632 1952 2644
rect 1581 2604 1952 2632
rect 1581 2601 1593 2604
rect 1535 2595 1593 2601
rect 1946 2592 1952 2604
rect 2004 2592 2010 2644
rect 2547 2635 2605 2641
rect 2547 2601 2559 2635
rect 2593 2632 2605 2635
rect 2682 2632 2688 2644
rect 2593 2604 2688 2632
rect 2593 2601 2605 2604
rect 2547 2595 2605 2601
rect 2682 2592 2688 2604
rect 2740 2592 2746 2644
rect 24210 2641 24216 2644
rect 24167 2635 24216 2641
rect 24167 2601 24179 2635
rect 24213 2601 24216 2635
rect 24167 2595 24216 2601
rect 24210 2592 24216 2595
rect 24268 2592 24274 2644
rect 24854 2592 24860 2644
rect 24912 2632 24918 2644
rect 25179 2635 25237 2641
rect 25179 2632 25191 2635
rect 24912 2604 25191 2632
rect 24912 2592 24918 2604
rect 25179 2601 25191 2604
rect 25225 2601 25237 2635
rect 25179 2595 25237 2601
rect 1394 2456 1400 2508
rect 1452 2505 1458 2508
rect 1452 2499 1490 2505
rect 1478 2496 1490 2499
rect 1857 2499 1915 2505
rect 1857 2496 1869 2499
rect 1478 2468 1869 2496
rect 1478 2465 1490 2468
rect 1452 2459 1490 2465
rect 1857 2465 1869 2468
rect 1903 2465 1915 2499
rect 1857 2459 1915 2465
rect 2476 2499 2534 2505
rect 2476 2465 2488 2499
rect 2522 2496 2534 2499
rect 2774 2496 2780 2508
rect 2522 2468 2780 2496
rect 2522 2465 2534 2468
rect 2476 2459 2534 2465
rect 1452 2456 1458 2459
rect 2774 2456 2780 2468
rect 2832 2496 2838 2508
rect 2869 2499 2927 2505
rect 2869 2496 2881 2499
rect 2832 2468 2881 2496
rect 2832 2456 2838 2468
rect 2869 2465 2881 2468
rect 2915 2465 2927 2499
rect 2869 2459 2927 2465
rect 24096 2499 24154 2505
rect 24096 2465 24108 2499
rect 24142 2496 24154 2499
rect 25108 2499 25166 2505
rect 24142 2468 24624 2496
rect 24142 2465 24154 2468
rect 24096 2459 24154 2465
rect 24596 2301 24624 2468
rect 25108 2465 25120 2499
rect 25154 2496 25166 2499
rect 25590 2496 25596 2508
rect 25154 2468 25596 2496
rect 25154 2465 25166 2468
rect 25108 2459 25166 2465
rect 25590 2456 25596 2468
rect 25648 2456 25654 2508
rect 24581 2295 24639 2301
rect 24581 2261 24593 2295
rect 24627 2292 24639 2295
rect 24670 2292 24676 2304
rect 24627 2264 24676 2292
rect 24627 2261 24639 2264
rect 24581 2255 24639 2261
rect 24670 2252 24676 2264
rect 24728 2252 24734 2304
rect 25590 2292 25596 2304
rect 25551 2264 25596 2292
rect 25590 2252 25596 2264
rect 25648 2252 25654 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 7650 552 7656 604
rect 7708 592 7714 604
rect 7834 592 7840 604
rect 7708 564 7840 592
rect 7708 552 7714 564
rect 7834 552 7840 564
rect 7892 552 7898 604
rect 10778 552 10784 604
rect 10836 592 10842 604
rect 10870 592 10876 604
rect 10836 564 10876 592
rect 10836 552 10842 564
rect 10870 552 10876 564
rect 10928 552 10934 604
<< via1 >>
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 16396 24395 16448 24404
rect 16396 24361 16405 24395
rect 16405 24361 16439 24395
rect 16439 24361 16448 24395
rect 16396 24352 16448 24361
rect 664 24216 716 24268
rect 2228 24216 2280 24268
rect 16120 24216 16172 24268
rect 17408 24259 17460 24268
rect 17408 24225 17426 24259
rect 17426 24225 17460 24259
rect 17408 24216 17460 24225
rect 2688 24012 2740 24064
rect 16488 24012 16540 24064
rect 17500 24012 17552 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 2228 23851 2280 23860
rect 2228 23817 2237 23851
rect 2237 23817 2271 23851
rect 2271 23817 2280 23851
rect 2228 23808 2280 23817
rect 12992 23851 13044 23860
rect 12992 23817 13001 23851
rect 13001 23817 13035 23851
rect 13035 23817 13044 23851
rect 12992 23808 13044 23817
rect 16028 23808 16080 23860
rect 17408 23851 17460 23860
rect 17408 23817 17417 23851
rect 17417 23817 17451 23851
rect 17451 23817 17460 23851
rect 17408 23808 17460 23817
rect 18788 23808 18840 23860
rect 23848 23851 23900 23860
rect 23848 23817 23857 23851
rect 23857 23817 23891 23851
rect 23891 23817 23900 23851
rect 23848 23808 23900 23817
rect 25320 23851 25372 23860
rect 25320 23817 25329 23851
rect 25329 23817 25363 23851
rect 25363 23817 25372 23851
rect 25320 23808 25372 23817
rect 1400 23647 1452 23656
rect 1400 23613 1444 23647
rect 1444 23613 1452 23647
rect 1400 23604 1452 23613
rect 12440 23604 12492 23656
rect 15292 23647 15344 23656
rect 15292 23613 15301 23647
rect 15301 23613 15335 23647
rect 15335 23613 15344 23647
rect 15292 23604 15344 23613
rect 2688 23536 2740 23588
rect 16488 23579 16540 23588
rect 16120 23468 16172 23520
rect 16488 23545 16497 23579
rect 16497 23545 16531 23579
rect 16531 23545 16540 23579
rect 16488 23536 16540 23545
rect 16948 23536 17000 23588
rect 17132 23579 17184 23588
rect 17132 23545 17141 23579
rect 17141 23545 17175 23579
rect 17175 23545 17184 23579
rect 17132 23536 17184 23545
rect 22468 23647 22520 23656
rect 22468 23613 22512 23647
rect 22512 23613 22520 23647
rect 22468 23604 22520 23613
rect 25320 23604 25372 23656
rect 18696 23511 18748 23520
rect 18696 23477 18705 23511
rect 18705 23477 18739 23511
rect 18739 23477 18748 23511
rect 18696 23468 18748 23477
rect 24860 23468 24912 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 15292 23264 15344 23316
rect 21640 23264 21692 23316
rect 22652 23307 22704 23316
rect 22652 23273 22661 23307
rect 22661 23273 22695 23307
rect 22695 23273 22704 23307
rect 22652 23264 22704 23273
rect 16580 23196 16632 23248
rect 15476 23171 15528 23180
rect 15476 23137 15520 23171
rect 15520 23137 15528 23171
rect 15476 23128 15528 23137
rect 18604 23128 18656 23180
rect 20904 23171 20956 23180
rect 20904 23137 20913 23171
rect 20913 23137 20947 23171
rect 20947 23137 20956 23171
rect 20904 23128 20956 23137
rect 22468 23171 22520 23180
rect 22468 23137 22477 23171
rect 22477 23137 22511 23171
rect 22511 23137 22520 23171
rect 22468 23128 22520 23137
rect 16672 23060 16724 23112
rect 17316 22992 17368 23044
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 17500 22763 17552 22772
rect 17500 22729 17509 22763
rect 17509 22729 17543 22763
rect 17543 22729 17552 22763
rect 17500 22720 17552 22729
rect 18604 22763 18656 22772
rect 18604 22729 18613 22763
rect 18613 22729 18647 22763
rect 18647 22729 18656 22763
rect 18604 22720 18656 22729
rect 16764 22627 16816 22636
rect 16764 22593 16773 22627
rect 16773 22593 16807 22627
rect 16807 22593 16816 22627
rect 16764 22584 16816 22593
rect 15660 22516 15712 22568
rect 15568 22491 15620 22500
rect 15568 22457 15577 22491
rect 15577 22457 15611 22491
rect 15611 22457 15620 22491
rect 15568 22448 15620 22457
rect 16580 22491 16632 22500
rect 16580 22457 16589 22491
rect 16589 22457 16623 22491
rect 16623 22457 16632 22491
rect 16580 22448 16632 22457
rect 20904 22491 20956 22500
rect 20904 22457 20913 22491
rect 20913 22457 20947 22491
rect 20947 22457 20956 22491
rect 20904 22448 20956 22457
rect 15752 22380 15804 22432
rect 17868 22380 17920 22432
rect 22468 22423 22520 22432
rect 22468 22389 22477 22423
rect 22477 22389 22511 22423
rect 22511 22389 22520 22423
rect 22468 22380 22520 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 15476 22219 15528 22228
rect 15476 22185 15485 22219
rect 15485 22185 15519 22219
rect 15519 22185 15528 22219
rect 17316 22219 17368 22228
rect 15476 22176 15528 22185
rect 17316 22185 17325 22219
rect 17325 22185 17359 22219
rect 17359 22185 17368 22219
rect 17316 22176 17368 22185
rect 13268 22108 13320 22160
rect 15568 22108 15620 22160
rect 15936 22108 15988 22160
rect 16488 22108 16540 22160
rect 17960 22151 18012 22160
rect 17960 22117 17969 22151
rect 17969 22117 18003 22151
rect 18003 22117 18012 22151
rect 17960 22108 18012 22117
rect 19432 22040 19484 22092
rect 21824 22083 21876 22092
rect 21824 22049 21833 22083
rect 21833 22049 21867 22083
rect 21867 22049 21876 22083
rect 21824 22040 21876 22049
rect 13268 22015 13320 22024
rect 13268 21981 13277 22015
rect 13277 21981 13311 22015
rect 13311 21981 13320 22015
rect 13268 21972 13320 21981
rect 13912 22015 13964 22024
rect 13912 21981 13921 22015
rect 13921 21981 13955 22015
rect 13955 21981 13964 22015
rect 13912 21972 13964 21981
rect 16304 22015 16356 22024
rect 16304 21981 16313 22015
rect 16313 21981 16347 22015
rect 16347 21981 16356 22015
rect 16304 21972 16356 21981
rect 16488 21972 16540 22024
rect 17868 22015 17920 22024
rect 17868 21981 17877 22015
rect 17877 21981 17911 22015
rect 17911 21981 17920 22015
rect 17868 21972 17920 21981
rect 18144 22015 18196 22024
rect 18144 21981 18153 22015
rect 18153 21981 18187 22015
rect 18187 21981 18196 22015
rect 18144 21972 18196 21981
rect 16212 21904 16264 21956
rect 16764 21904 16816 21956
rect 20168 21904 20220 21956
rect 22008 21947 22060 21956
rect 22008 21913 22017 21947
rect 22017 21913 22051 21947
rect 22051 21913 22060 21947
rect 22008 21904 22060 21913
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 13176 21632 13228 21684
rect 15936 21675 15988 21684
rect 15936 21641 15945 21675
rect 15945 21641 15979 21675
rect 15979 21641 15988 21675
rect 15936 21632 15988 21641
rect 17868 21632 17920 21684
rect 19432 21675 19484 21684
rect 19432 21641 19441 21675
rect 19441 21641 19475 21675
rect 19475 21641 19484 21675
rect 19432 21632 19484 21641
rect 16396 21564 16448 21616
rect 13912 21539 13964 21548
rect 13912 21505 13921 21539
rect 13921 21505 13955 21539
rect 13955 21505 13964 21539
rect 13912 21496 13964 21505
rect 16212 21539 16264 21548
rect 1492 21471 1544 21480
rect 1492 21437 1510 21471
rect 1510 21437 1544 21471
rect 1492 21428 1544 21437
rect 16212 21505 16221 21539
rect 16221 21505 16255 21539
rect 16255 21505 16264 21539
rect 16212 21496 16264 21505
rect 16488 21539 16540 21548
rect 16488 21505 16497 21539
rect 16497 21505 16531 21539
rect 16531 21505 16540 21539
rect 16488 21496 16540 21505
rect 18052 21428 18104 21480
rect 21824 21471 21876 21480
rect 21824 21437 21833 21471
rect 21833 21437 21867 21471
rect 21867 21437 21876 21471
rect 21824 21428 21876 21437
rect 13636 21403 13688 21412
rect 13636 21369 13645 21403
rect 13645 21369 13679 21403
rect 13679 21369 13688 21403
rect 13636 21360 13688 21369
rect 13728 21403 13780 21412
rect 13728 21369 13737 21403
rect 13737 21369 13771 21403
rect 13771 21369 13780 21403
rect 15660 21403 15712 21412
rect 13728 21360 13780 21369
rect 15660 21369 15669 21403
rect 15669 21369 15703 21403
rect 15703 21369 15712 21403
rect 15660 21360 15712 21369
rect 16212 21360 16264 21412
rect 1768 21292 1820 21344
rect 16396 21292 16448 21344
rect 17960 21292 18012 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 13268 21131 13320 21140
rect 10784 21063 10836 21072
rect 10784 21029 10793 21063
rect 10793 21029 10827 21063
rect 10827 21029 10836 21063
rect 10784 21020 10836 21029
rect 11888 21020 11940 21072
rect 13268 21097 13277 21131
rect 13277 21097 13311 21131
rect 13311 21097 13320 21131
rect 13268 21088 13320 21097
rect 13636 21131 13688 21140
rect 13636 21097 13645 21131
rect 13645 21097 13679 21131
rect 13679 21097 13688 21131
rect 13636 21088 13688 21097
rect 19432 21088 19484 21140
rect 10692 20927 10744 20936
rect 10692 20893 10701 20927
rect 10701 20893 10735 20927
rect 10735 20893 10744 20927
rect 10692 20884 10744 20893
rect 12532 20884 12584 20936
rect 16396 21020 16448 21072
rect 17776 20995 17828 21004
rect 17776 20961 17785 20995
rect 17785 20961 17819 20995
rect 17819 20961 17828 20995
rect 17776 20952 17828 20961
rect 19340 20995 19392 21004
rect 19340 20961 19358 20995
rect 19358 20961 19392 20995
rect 19340 20952 19392 20961
rect 16580 20884 16632 20936
rect 16304 20816 16356 20868
rect 16764 20859 16816 20868
rect 16764 20825 16773 20859
rect 16773 20825 16807 20859
rect 16807 20825 16816 20859
rect 16764 20816 16816 20825
rect 14832 20748 14884 20800
rect 17960 20791 18012 20800
rect 17960 20757 17969 20791
rect 17969 20757 18003 20791
rect 18003 20757 18012 20791
rect 17960 20748 18012 20757
rect 18788 20791 18840 20800
rect 18788 20757 18797 20791
rect 18797 20757 18831 20791
rect 18831 20757 18840 20791
rect 18788 20748 18840 20757
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 11888 20587 11940 20596
rect 11888 20553 11897 20587
rect 11897 20553 11931 20587
rect 11931 20553 11940 20587
rect 11888 20544 11940 20553
rect 13176 20544 13228 20596
rect 15752 20544 15804 20596
rect 16396 20544 16448 20596
rect 16580 20587 16632 20596
rect 16580 20553 16589 20587
rect 16589 20553 16623 20587
rect 16623 20553 16632 20587
rect 16580 20544 16632 20553
rect 17960 20544 18012 20596
rect 10784 20451 10836 20460
rect 10784 20417 10793 20451
rect 10793 20417 10827 20451
rect 10827 20417 10836 20451
rect 10784 20408 10836 20417
rect 18788 20476 18840 20528
rect 18604 20451 18656 20460
rect 18604 20417 18613 20451
rect 18613 20417 18647 20451
rect 18647 20417 18656 20451
rect 18604 20408 18656 20417
rect 19340 20408 19392 20460
rect 20812 20451 20864 20460
rect 20812 20417 20821 20451
rect 20821 20417 20855 20451
rect 20855 20417 20864 20451
rect 20812 20408 20864 20417
rect 11888 20340 11940 20392
rect 12716 20383 12768 20392
rect 12716 20349 12725 20383
rect 12725 20349 12759 20383
rect 12759 20349 12768 20383
rect 12716 20340 12768 20349
rect 14832 20340 14884 20392
rect 16672 20383 16724 20392
rect 16672 20349 16716 20383
rect 16716 20349 16724 20383
rect 16672 20340 16724 20349
rect 19800 20383 19852 20392
rect 19800 20349 19844 20383
rect 19844 20349 19852 20383
rect 20260 20383 20312 20392
rect 19800 20340 19852 20349
rect 20260 20349 20269 20383
rect 20269 20349 20303 20383
rect 20303 20349 20312 20383
rect 20260 20340 20312 20349
rect 11980 20272 12032 20324
rect 15568 20272 15620 20324
rect 13452 20204 13504 20256
rect 17960 20204 18012 20256
rect 19432 20204 19484 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 10692 20043 10744 20052
rect 10692 20009 10701 20043
rect 10701 20009 10735 20043
rect 10735 20009 10744 20043
rect 10692 20000 10744 20009
rect 11888 20000 11940 20052
rect 13176 20000 13228 20052
rect 11980 19932 12032 19984
rect 9864 19907 9916 19916
rect 9864 19873 9908 19907
rect 9908 19873 9916 19907
rect 9864 19864 9916 19873
rect 10968 19864 11020 19916
rect 13820 20000 13872 20052
rect 16212 20043 16264 20052
rect 16212 20009 16221 20043
rect 16221 20009 16255 20043
rect 16255 20009 16264 20043
rect 16212 20000 16264 20009
rect 17776 20043 17828 20052
rect 17776 20009 17785 20043
rect 17785 20009 17819 20043
rect 17819 20009 17828 20043
rect 17776 20000 17828 20009
rect 15568 19932 15620 19984
rect 18604 19975 18656 19984
rect 18604 19941 18613 19975
rect 18613 19941 18647 19975
rect 18647 19941 18656 19975
rect 18604 19932 18656 19941
rect 19524 19907 19576 19916
rect 19524 19873 19542 19907
rect 19542 19873 19576 19907
rect 19524 19864 19576 19873
rect 11888 19839 11940 19848
rect 11888 19805 11897 19839
rect 11897 19805 11931 19839
rect 11931 19805 11940 19839
rect 11888 19796 11940 19805
rect 15476 19796 15528 19848
rect 18420 19796 18472 19848
rect 11336 19728 11388 19780
rect 10048 19660 10100 19712
rect 11428 19703 11480 19712
rect 11428 19669 11437 19703
rect 11437 19669 11471 19703
rect 11471 19669 11480 19703
rect 11428 19660 11480 19669
rect 12716 19660 12768 19712
rect 14740 19703 14792 19712
rect 14740 19669 14749 19703
rect 14749 19669 14783 19703
rect 14783 19669 14792 19703
rect 14740 19660 14792 19669
rect 16672 19660 16724 19712
rect 19340 19660 19392 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 9864 19499 9916 19508
rect 9864 19465 9873 19499
rect 9873 19465 9907 19499
rect 9907 19465 9916 19499
rect 9864 19456 9916 19465
rect 11980 19499 12032 19508
rect 11980 19465 11989 19499
rect 11989 19465 12023 19499
rect 12023 19465 12032 19499
rect 11980 19456 12032 19465
rect 15568 19456 15620 19508
rect 16028 19499 16080 19508
rect 16028 19465 16037 19499
rect 16037 19465 16071 19499
rect 16071 19465 16080 19499
rect 16028 19456 16080 19465
rect 17776 19456 17828 19508
rect 14832 19431 14884 19440
rect 14832 19397 14841 19431
rect 14841 19397 14875 19431
rect 14875 19397 14884 19431
rect 14832 19388 14884 19397
rect 16672 19320 16724 19372
rect 18420 19363 18472 19372
rect 18420 19329 18429 19363
rect 18429 19329 18463 19363
rect 18463 19329 18472 19363
rect 18420 19320 18472 19329
rect 1400 19295 1452 19304
rect 1400 19261 1444 19295
rect 1444 19261 1452 19295
rect 1400 19252 1452 19261
rect 1768 19116 1820 19168
rect 7288 19116 7340 19168
rect 8392 19252 8444 19304
rect 9036 19252 9088 19304
rect 9588 19252 9640 19304
rect 11428 19252 11480 19304
rect 12256 19252 12308 19304
rect 12440 19295 12492 19304
rect 12440 19261 12484 19295
rect 12484 19261 12492 19295
rect 14188 19295 14240 19304
rect 12440 19252 12492 19261
rect 14188 19261 14197 19295
rect 14197 19261 14231 19295
rect 14231 19261 14240 19295
rect 14188 19252 14240 19261
rect 13636 19184 13688 19236
rect 13912 19227 13964 19236
rect 13912 19193 13921 19227
rect 13921 19193 13955 19227
rect 13955 19193 13964 19227
rect 14740 19252 14792 19304
rect 15752 19252 15804 19304
rect 13912 19184 13964 19193
rect 16028 19184 16080 19236
rect 18144 19227 18196 19236
rect 18144 19193 18153 19227
rect 18153 19193 18187 19227
rect 18187 19193 18196 19227
rect 18144 19184 18196 19193
rect 7656 19116 7708 19168
rect 8944 19116 8996 19168
rect 9128 19116 9180 19168
rect 10140 19116 10192 19168
rect 10968 19159 11020 19168
rect 10968 19125 10977 19159
rect 10977 19125 11011 19159
rect 11011 19125 11020 19159
rect 10968 19116 11020 19125
rect 11428 19116 11480 19168
rect 12532 19116 12584 19168
rect 13452 19116 13504 19168
rect 14188 19116 14240 19168
rect 18328 19184 18380 19236
rect 21180 19295 21232 19304
rect 21180 19261 21224 19295
rect 21224 19261 21232 19295
rect 21180 19252 21232 19261
rect 24768 19252 24820 19304
rect 19524 19159 19576 19168
rect 19524 19125 19533 19159
rect 19533 19125 19567 19159
rect 19567 19125 19576 19159
rect 19524 19116 19576 19125
rect 20996 19116 21048 19168
rect 23480 19116 23532 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 12348 18912 12400 18964
rect 17500 18912 17552 18964
rect 7564 18887 7616 18896
rect 7564 18853 7573 18887
rect 7573 18853 7607 18887
rect 7607 18853 7616 18887
rect 7564 18844 7616 18853
rect 10508 18887 10560 18896
rect 10508 18853 10517 18887
rect 10517 18853 10551 18887
rect 10551 18853 10560 18887
rect 10508 18844 10560 18853
rect 10784 18844 10836 18896
rect 16028 18844 16080 18896
rect 17592 18887 17644 18896
rect 17592 18853 17601 18887
rect 17601 18853 17635 18887
rect 17635 18853 17644 18887
rect 17592 18844 17644 18853
rect 18144 18912 18196 18964
rect 19248 18912 19300 18964
rect 21824 18955 21876 18964
rect 21824 18921 21833 18955
rect 21833 18921 21867 18955
rect 21867 18921 21876 18955
rect 21824 18912 21876 18921
rect 18052 18844 18104 18896
rect 18420 18844 18472 18896
rect 23480 18844 23532 18896
rect 6368 18819 6420 18828
rect 6368 18785 6412 18819
rect 6412 18785 6420 18819
rect 6368 18776 6420 18785
rect 12164 18776 12216 18828
rect 13544 18819 13596 18828
rect 13544 18785 13553 18819
rect 13553 18785 13587 18819
rect 13587 18785 13596 18819
rect 13544 18776 13596 18785
rect 13912 18819 13964 18828
rect 13912 18785 13921 18819
rect 13921 18785 13955 18819
rect 13955 18785 13964 18819
rect 13912 18776 13964 18785
rect 7472 18751 7524 18760
rect 7472 18717 7481 18751
rect 7481 18717 7515 18751
rect 7515 18717 7524 18751
rect 7472 18708 7524 18717
rect 7748 18751 7800 18760
rect 7748 18717 7757 18751
rect 7757 18717 7791 18751
rect 7791 18717 7800 18751
rect 7748 18708 7800 18717
rect 10324 18708 10376 18760
rect 13820 18708 13872 18760
rect 14740 18776 14792 18828
rect 18880 18776 18932 18828
rect 19524 18819 19576 18828
rect 19524 18785 19533 18819
rect 19533 18785 19567 18819
rect 19567 18785 19576 18819
rect 19524 18776 19576 18785
rect 20720 18776 20772 18828
rect 24584 18819 24636 18828
rect 24584 18785 24628 18819
rect 24628 18785 24636 18819
rect 24584 18776 24636 18785
rect 16488 18708 16540 18760
rect 19340 18708 19392 18760
rect 10692 18572 10744 18624
rect 11888 18615 11940 18624
rect 11888 18581 11897 18615
rect 11897 18581 11931 18615
rect 11931 18581 11940 18615
rect 11888 18572 11940 18581
rect 12348 18572 12400 18624
rect 12440 18615 12492 18624
rect 12440 18581 12449 18615
rect 12449 18581 12483 18615
rect 12483 18581 12492 18615
rect 12900 18615 12952 18624
rect 12440 18572 12492 18581
rect 12900 18581 12909 18615
rect 12909 18581 12943 18615
rect 12943 18581 12952 18615
rect 12900 18572 12952 18581
rect 14740 18615 14792 18624
rect 14740 18581 14749 18615
rect 14749 18581 14783 18615
rect 14783 18581 14792 18615
rect 14740 18572 14792 18581
rect 15476 18615 15528 18624
rect 15476 18581 15485 18615
rect 15485 18581 15519 18615
rect 15519 18581 15528 18615
rect 15476 18572 15528 18581
rect 20076 18615 20128 18624
rect 20076 18581 20085 18615
rect 20085 18581 20119 18615
rect 20119 18581 20128 18615
rect 20076 18572 20128 18581
rect 20812 18572 20864 18624
rect 21456 18615 21508 18624
rect 21456 18581 21465 18615
rect 21465 18581 21499 18615
rect 21499 18581 21508 18615
rect 21456 18572 21508 18581
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 5448 18164 5500 18216
rect 6184 18368 6236 18420
rect 6460 18411 6512 18420
rect 6460 18377 6469 18411
rect 6469 18377 6503 18411
rect 6503 18377 6512 18411
rect 6460 18368 6512 18377
rect 7564 18368 7616 18420
rect 11244 18368 11296 18420
rect 13912 18368 13964 18420
rect 7288 18232 7340 18284
rect 10324 18275 10376 18284
rect 10324 18241 10333 18275
rect 10333 18241 10367 18275
rect 10367 18241 10376 18275
rect 10324 18232 10376 18241
rect 11060 18232 11112 18284
rect 13176 18232 13228 18284
rect 16028 18368 16080 18420
rect 16488 18411 16540 18420
rect 16488 18377 16497 18411
rect 16497 18377 16531 18411
rect 16531 18377 16540 18411
rect 16488 18368 16540 18377
rect 19524 18368 19576 18420
rect 24676 18411 24728 18420
rect 24676 18377 24685 18411
rect 24685 18377 24719 18411
rect 24719 18377 24728 18411
rect 24676 18368 24728 18377
rect 15476 18343 15528 18352
rect 15476 18309 15485 18343
rect 15485 18309 15519 18343
rect 15519 18309 15528 18343
rect 15476 18300 15528 18309
rect 10968 18207 11020 18216
rect 10968 18173 10977 18207
rect 10977 18173 11011 18207
rect 11011 18173 11020 18207
rect 10968 18164 11020 18173
rect 12164 18164 12216 18216
rect 6828 18096 6880 18148
rect 7012 18096 7064 18148
rect 7840 18096 7892 18148
rect 10692 18096 10744 18148
rect 12900 18207 12952 18216
rect 12900 18173 12909 18207
rect 12909 18173 12943 18207
rect 12943 18173 12952 18207
rect 12900 18164 12952 18173
rect 14188 18164 14240 18216
rect 14740 18207 14792 18216
rect 14740 18173 14749 18207
rect 14749 18173 14783 18207
rect 14783 18173 14792 18207
rect 14740 18164 14792 18173
rect 20720 18232 20772 18284
rect 21272 18232 21324 18284
rect 21824 18300 21876 18352
rect 21640 18232 21692 18284
rect 15568 18207 15620 18216
rect 15568 18173 15577 18207
rect 15577 18173 15611 18207
rect 15611 18173 15620 18207
rect 15568 18164 15620 18173
rect 16580 18164 16632 18216
rect 18420 18164 18472 18216
rect 13912 18096 13964 18148
rect 19064 18164 19116 18216
rect 19248 18164 19300 18216
rect 20076 18164 20128 18216
rect 9404 18071 9456 18080
rect 9404 18037 9413 18071
rect 9413 18037 9447 18071
rect 9447 18037 9456 18071
rect 9404 18028 9456 18037
rect 10784 18028 10836 18080
rect 11520 18071 11572 18080
rect 11520 18037 11529 18071
rect 11529 18037 11563 18071
rect 11563 18037 11572 18071
rect 11520 18028 11572 18037
rect 12256 18071 12308 18080
rect 12256 18037 12265 18071
rect 12265 18037 12299 18071
rect 12299 18037 12308 18071
rect 12256 18028 12308 18037
rect 12716 18071 12768 18080
rect 12716 18037 12725 18071
rect 12725 18037 12759 18071
rect 12759 18037 12768 18071
rect 12716 18028 12768 18037
rect 13544 18028 13596 18080
rect 14464 18028 14516 18080
rect 16856 18071 16908 18080
rect 16856 18037 16865 18071
rect 16865 18037 16899 18071
rect 16899 18037 16908 18071
rect 16856 18028 16908 18037
rect 18052 18028 18104 18080
rect 18972 18028 19024 18080
rect 20720 18096 20772 18148
rect 21456 18096 21508 18148
rect 20628 18028 20680 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 5540 17824 5592 17876
rect 7472 17824 7524 17876
rect 10876 17824 10928 17876
rect 11060 17867 11112 17876
rect 11060 17833 11069 17867
rect 11069 17833 11103 17867
rect 11103 17833 11112 17867
rect 11060 17824 11112 17833
rect 12348 17824 12400 17876
rect 13912 17867 13964 17876
rect 13912 17833 13921 17867
rect 13921 17833 13955 17867
rect 13955 17833 13964 17867
rect 13912 17824 13964 17833
rect 16948 17867 17000 17876
rect 16948 17833 16957 17867
rect 16957 17833 16991 17867
rect 16991 17833 17000 17867
rect 16948 17824 17000 17833
rect 17500 17867 17552 17876
rect 17500 17833 17509 17867
rect 17509 17833 17543 17867
rect 17543 17833 17552 17867
rect 17500 17824 17552 17833
rect 18880 17867 18932 17876
rect 18880 17833 18889 17867
rect 18889 17833 18923 17867
rect 18923 17833 18932 17867
rect 18880 17824 18932 17833
rect 20536 17824 20588 17876
rect 7012 17756 7064 17808
rect 7196 17799 7248 17808
rect 7196 17765 7205 17799
rect 7205 17765 7239 17799
rect 7239 17765 7248 17799
rect 7196 17756 7248 17765
rect 7564 17756 7616 17808
rect 7840 17799 7892 17808
rect 7840 17765 7849 17799
rect 7849 17765 7883 17799
rect 7883 17765 7892 17799
rect 7840 17756 7892 17765
rect 9404 17756 9456 17808
rect 9864 17799 9916 17808
rect 9864 17765 9873 17799
rect 9873 17765 9907 17799
rect 9907 17765 9916 17799
rect 9864 17756 9916 17765
rect 10968 17756 11020 17808
rect 11796 17756 11848 17808
rect 2136 17731 2188 17740
rect 2136 17697 2154 17731
rect 2154 17697 2188 17731
rect 2136 17688 2188 17697
rect 4620 17731 4672 17740
rect 4620 17697 4638 17731
rect 4638 17697 4672 17731
rect 4620 17688 4672 17697
rect 5448 17688 5500 17740
rect 12256 17731 12308 17740
rect 12256 17697 12265 17731
rect 12265 17697 12299 17731
rect 12299 17697 12308 17731
rect 12256 17688 12308 17697
rect 12900 17731 12952 17740
rect 12900 17697 12909 17731
rect 12909 17697 12943 17731
rect 12943 17697 12952 17731
rect 12900 17688 12952 17697
rect 16028 17756 16080 17808
rect 18972 17756 19024 17808
rect 20720 17756 20772 17808
rect 22284 17756 22336 17808
rect 13544 17731 13596 17740
rect 13544 17697 13553 17731
rect 13553 17697 13587 17731
rect 13587 17697 13596 17731
rect 13544 17688 13596 17697
rect 13820 17688 13872 17740
rect 17776 17731 17828 17740
rect 17776 17697 17785 17731
rect 17785 17697 17819 17731
rect 17819 17697 17828 17731
rect 17776 17688 17828 17697
rect 15660 17620 15712 17672
rect 19064 17663 19116 17672
rect 19064 17629 19073 17663
rect 19073 17629 19107 17663
rect 19107 17629 19116 17663
rect 19064 17620 19116 17629
rect 20812 17620 20864 17672
rect 1400 17552 1452 17604
rect 4068 17552 4120 17604
rect 7748 17552 7800 17604
rect 21640 17620 21692 17672
rect 22468 17663 22520 17672
rect 22468 17629 22477 17663
rect 22477 17629 22511 17663
rect 22511 17629 22520 17663
rect 22468 17620 22520 17629
rect 21548 17595 21600 17604
rect 21548 17561 21557 17595
rect 21557 17561 21591 17595
rect 21591 17561 21600 17595
rect 21548 17552 21600 17561
rect 2412 17484 2464 17536
rect 5080 17484 5132 17536
rect 5264 17527 5316 17536
rect 5264 17493 5273 17527
rect 5273 17493 5307 17527
rect 5307 17493 5316 17527
rect 5264 17484 5316 17493
rect 6920 17527 6972 17536
rect 6920 17493 6929 17527
rect 6929 17493 6963 17527
rect 6963 17493 6972 17527
rect 6920 17484 6972 17493
rect 12164 17484 12216 17536
rect 14280 17527 14332 17536
rect 14280 17493 14289 17527
rect 14289 17493 14323 17527
rect 14323 17493 14332 17527
rect 14280 17484 14332 17493
rect 15568 17484 15620 17536
rect 15844 17527 15896 17536
rect 15844 17493 15853 17527
rect 15853 17493 15887 17527
rect 15887 17493 15896 17527
rect 15844 17484 15896 17493
rect 17960 17527 18012 17536
rect 17960 17493 17969 17527
rect 17969 17493 18003 17527
rect 18003 17493 18012 17527
rect 17960 17484 18012 17493
rect 18420 17484 18472 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 4068 17323 4120 17332
rect 4068 17289 4077 17323
rect 4077 17289 4111 17323
rect 4111 17289 4120 17323
rect 4068 17280 4120 17289
rect 4620 17323 4672 17332
rect 4620 17289 4629 17323
rect 4629 17289 4663 17323
rect 4663 17289 4672 17323
rect 4620 17280 4672 17289
rect 7012 17280 7064 17332
rect 7564 17280 7616 17332
rect 10784 17323 10836 17332
rect 10784 17289 10793 17323
rect 10793 17289 10827 17323
rect 10827 17289 10836 17323
rect 10784 17280 10836 17289
rect 11520 17323 11572 17332
rect 11520 17289 11529 17323
rect 11529 17289 11563 17323
rect 11563 17289 11572 17323
rect 11520 17280 11572 17289
rect 11796 17323 11848 17332
rect 11796 17289 11805 17323
rect 11805 17289 11839 17323
rect 11839 17289 11848 17323
rect 11796 17280 11848 17289
rect 13912 17280 13964 17332
rect 15752 17280 15804 17332
rect 16028 17280 16080 17332
rect 18972 17323 19024 17332
rect 18972 17289 18981 17323
rect 18981 17289 19015 17323
rect 19015 17289 19024 17323
rect 18972 17280 19024 17289
rect 20720 17323 20772 17332
rect 20720 17289 20729 17323
rect 20729 17289 20763 17323
rect 20763 17289 20772 17323
rect 20720 17280 20772 17289
rect 22284 17323 22336 17332
rect 22284 17289 22293 17323
rect 22293 17289 22327 17323
rect 22327 17289 22336 17323
rect 22284 17280 22336 17289
rect 12348 17212 12400 17264
rect 12164 17144 12216 17196
rect 21088 17212 21140 17264
rect 1400 17119 1452 17128
rect 1400 17085 1409 17119
rect 1409 17085 1443 17119
rect 1443 17085 1452 17119
rect 1400 17076 1452 17085
rect 4068 17076 4120 17128
rect 1492 16940 1544 16992
rect 2136 16983 2188 16992
rect 2136 16949 2145 16983
rect 2145 16949 2179 16983
rect 2179 16949 2188 16983
rect 2136 16940 2188 16949
rect 2596 16940 2648 16992
rect 2872 16940 2924 16992
rect 5264 17076 5316 17128
rect 6920 17076 6972 17128
rect 6276 17008 6328 17060
rect 6644 17051 6696 17060
rect 6644 17017 6653 17051
rect 6653 17017 6687 17051
rect 6687 17017 6696 17051
rect 6644 17008 6696 17017
rect 8208 17008 8260 17060
rect 6552 16940 6604 16992
rect 9036 16983 9088 16992
rect 9036 16949 9045 16983
rect 9045 16949 9079 16983
rect 9079 16949 9088 16983
rect 9036 16940 9088 16949
rect 9956 17076 10008 17128
rect 14464 17076 14516 17128
rect 18972 17144 19024 17196
rect 12532 17051 12584 17060
rect 12532 17017 12541 17051
rect 12541 17017 12575 17051
rect 12575 17017 12584 17051
rect 12532 17008 12584 17017
rect 12624 17051 12676 17060
rect 12624 17017 12633 17051
rect 12633 17017 12667 17051
rect 12667 17017 12676 17051
rect 12624 17008 12676 17017
rect 13820 17008 13872 17060
rect 14280 17008 14332 17060
rect 15200 17076 15252 17128
rect 15844 17076 15896 17128
rect 16120 17008 16172 17060
rect 17960 17008 18012 17060
rect 18328 17008 18380 17060
rect 9496 16940 9548 16992
rect 9772 16983 9824 16992
rect 9772 16949 9781 16983
rect 9781 16949 9815 16983
rect 9815 16949 9824 16983
rect 9772 16940 9824 16949
rect 9864 16940 9916 16992
rect 11612 16940 11664 16992
rect 12256 16940 12308 16992
rect 12348 16940 12400 16992
rect 13268 16940 13320 16992
rect 13544 16940 13596 16992
rect 15660 16940 15712 16992
rect 16948 16983 17000 16992
rect 16948 16949 16957 16983
rect 16957 16949 16991 16983
rect 16991 16949 17000 16983
rect 16948 16940 17000 16949
rect 17776 16983 17828 16992
rect 17776 16949 17785 16983
rect 17785 16949 17819 16983
rect 17819 16949 17828 16983
rect 17776 16940 17828 16949
rect 18236 16983 18288 16992
rect 18236 16949 18245 16983
rect 18245 16949 18279 16983
rect 18279 16949 18288 16983
rect 18236 16940 18288 16949
rect 20812 17144 20864 17196
rect 21640 17187 21692 17196
rect 21640 17153 21649 17187
rect 21649 17153 21683 17187
rect 21683 17153 21692 17187
rect 21640 17144 21692 17153
rect 22560 17119 22612 17128
rect 22560 17085 22578 17119
rect 22578 17085 22612 17119
rect 23388 17280 23440 17332
rect 22560 17076 22612 17085
rect 23664 17119 23716 17128
rect 23664 17085 23708 17119
rect 23708 17085 23716 17119
rect 23664 17076 23716 17085
rect 23940 17076 23992 17128
rect 20628 16940 20680 16992
rect 20812 16940 20864 16992
rect 24952 17008 25004 17060
rect 22376 16940 22428 16992
rect 23848 16940 23900 16992
rect 24676 16940 24728 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 1400 16736 1452 16788
rect 2412 16736 2464 16788
rect 5540 16736 5592 16788
rect 7012 16779 7064 16788
rect 7012 16745 7021 16779
rect 7021 16745 7055 16779
rect 7055 16745 7064 16779
rect 7012 16736 7064 16745
rect 7196 16736 7248 16788
rect 9404 16779 9456 16788
rect 9404 16745 9413 16779
rect 9413 16745 9447 16779
rect 9447 16745 9456 16779
rect 9404 16736 9456 16745
rect 10968 16736 11020 16788
rect 12624 16736 12676 16788
rect 15384 16736 15436 16788
rect 16028 16779 16080 16788
rect 16028 16745 16037 16779
rect 16037 16745 16071 16779
rect 16071 16745 16080 16779
rect 16028 16736 16080 16745
rect 20812 16736 20864 16788
rect 2320 16668 2372 16720
rect 6644 16668 6696 16720
rect 8208 16711 8260 16720
rect 8208 16677 8211 16711
rect 8211 16677 8245 16711
rect 8245 16677 8260 16711
rect 8208 16668 8260 16677
rect 9772 16668 9824 16720
rect 12532 16668 12584 16720
rect 14372 16711 14424 16720
rect 14372 16677 14381 16711
rect 14381 16677 14415 16711
rect 14415 16677 14424 16711
rect 14372 16668 14424 16677
rect 16948 16668 17000 16720
rect 18972 16668 19024 16720
rect 19432 16668 19484 16720
rect 20168 16711 20220 16720
rect 20168 16677 20177 16711
rect 20177 16677 20211 16711
rect 20211 16677 20220 16711
rect 20168 16668 20220 16677
rect 22376 16736 22428 16788
rect 22652 16779 22704 16788
rect 22652 16745 22661 16779
rect 22661 16745 22695 16779
rect 22695 16745 22704 16779
rect 22652 16736 22704 16745
rect 23756 16736 23808 16788
rect 21088 16711 21140 16720
rect 21088 16677 21097 16711
rect 21097 16677 21131 16711
rect 21131 16677 21140 16711
rect 21640 16711 21692 16720
rect 21088 16668 21140 16677
rect 21640 16677 21649 16711
rect 21649 16677 21683 16711
rect 21683 16677 21692 16711
rect 21640 16668 21692 16677
rect 2044 16600 2096 16652
rect 2504 16643 2556 16652
rect 2504 16609 2548 16643
rect 2548 16609 2556 16643
rect 2504 16600 2556 16609
rect 2780 16600 2832 16652
rect 4528 16643 4580 16652
rect 4528 16609 4537 16643
rect 4537 16609 4571 16643
rect 4571 16609 4580 16643
rect 4528 16600 4580 16609
rect 5448 16600 5500 16652
rect 8300 16600 8352 16652
rect 9864 16600 9916 16652
rect 10140 16643 10192 16652
rect 10140 16609 10149 16643
rect 10149 16609 10183 16643
rect 10183 16609 10192 16643
rect 10140 16600 10192 16609
rect 12900 16600 12952 16652
rect 13176 16600 13228 16652
rect 13820 16600 13872 16652
rect 14464 16600 14516 16652
rect 15292 16643 15344 16652
rect 6092 16575 6144 16584
rect 6092 16541 6101 16575
rect 6101 16541 6135 16575
rect 6135 16541 6144 16575
rect 6092 16532 6144 16541
rect 11520 16532 11572 16584
rect 15292 16609 15301 16643
rect 15301 16609 15335 16643
rect 15335 16609 15344 16643
rect 15292 16600 15344 16609
rect 16396 16600 16448 16652
rect 19892 16600 19944 16652
rect 22468 16643 22520 16652
rect 22468 16609 22477 16643
rect 22477 16609 22511 16643
rect 22511 16609 22520 16643
rect 22468 16600 22520 16609
rect 17224 16532 17276 16584
rect 18972 16575 19024 16584
rect 18972 16541 18981 16575
rect 18981 16541 19015 16575
rect 19015 16541 19024 16575
rect 18972 16532 19024 16541
rect 23112 16532 23164 16584
rect 24768 16600 24820 16652
rect 13728 16507 13780 16516
rect 13728 16473 13737 16507
rect 13737 16473 13771 16507
rect 13771 16473 13780 16507
rect 13728 16464 13780 16473
rect 15292 16464 15344 16516
rect 17132 16507 17184 16516
rect 17132 16473 17141 16507
rect 17141 16473 17175 16507
rect 17175 16473 17184 16507
rect 17132 16464 17184 16473
rect 5264 16396 5316 16448
rect 7288 16439 7340 16448
rect 7288 16405 7297 16439
rect 7297 16405 7331 16439
rect 7331 16405 7340 16439
rect 7288 16396 7340 16405
rect 9956 16439 10008 16448
rect 9956 16405 9965 16439
rect 9965 16405 9999 16439
rect 9999 16405 10008 16439
rect 9956 16396 10008 16405
rect 10968 16396 11020 16448
rect 15476 16439 15528 16448
rect 15476 16405 15485 16439
rect 15485 16405 15519 16439
rect 15519 16405 15528 16439
rect 15476 16396 15528 16405
rect 18328 16439 18380 16448
rect 18328 16405 18337 16439
rect 18337 16405 18371 16439
rect 18371 16405 18380 16439
rect 18328 16396 18380 16405
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 1584 16235 1636 16244
rect 1584 16201 1593 16235
rect 1593 16201 1627 16235
rect 1627 16201 1636 16235
rect 1584 16192 1636 16201
rect 2504 16192 2556 16244
rect 4528 16192 4580 16244
rect 6644 16192 6696 16244
rect 8300 16235 8352 16244
rect 8300 16201 8309 16235
rect 8309 16201 8343 16235
rect 8343 16201 8352 16235
rect 8300 16192 8352 16201
rect 10692 16235 10744 16244
rect 10692 16201 10701 16235
rect 10701 16201 10735 16235
rect 10735 16201 10744 16235
rect 10692 16192 10744 16201
rect 11520 16235 11572 16244
rect 11520 16201 11529 16235
rect 11529 16201 11563 16235
rect 11563 16201 11572 16235
rect 11520 16192 11572 16201
rect 15292 16235 15344 16244
rect 15292 16201 15301 16235
rect 15301 16201 15335 16235
rect 15335 16201 15344 16235
rect 15292 16192 15344 16201
rect 16580 16192 16632 16244
rect 17224 16235 17276 16244
rect 17224 16201 17233 16235
rect 17233 16201 17267 16235
rect 17267 16201 17276 16235
rect 17224 16192 17276 16201
rect 19432 16192 19484 16244
rect 21180 16235 21232 16244
rect 21180 16201 21189 16235
rect 21189 16201 21223 16235
rect 21223 16201 21232 16235
rect 21180 16192 21232 16201
rect 24768 16235 24820 16244
rect 24768 16201 24777 16235
rect 24777 16201 24811 16235
rect 24811 16201 24820 16235
rect 24768 16192 24820 16201
rect 6184 16124 6236 16176
rect 2412 16056 2464 16108
rect 1676 15988 1728 16040
rect 4252 16031 4304 16040
rect 4252 15997 4270 16031
rect 4270 15997 4304 16031
rect 4252 15988 4304 15997
rect 4988 15988 5040 16040
rect 5172 16031 5224 16040
rect 5172 15997 5181 16031
rect 5181 15997 5215 16031
rect 5215 15997 5224 16031
rect 5172 15988 5224 15997
rect 5264 15988 5316 16040
rect 10140 16124 10192 16176
rect 8208 16056 8260 16108
rect 7288 15988 7340 16040
rect 8116 15988 8168 16040
rect 2228 15920 2280 15972
rect 2780 15920 2832 15972
rect 3240 15963 3292 15972
rect 3240 15929 3249 15963
rect 3249 15929 3283 15963
rect 3283 15929 3292 15963
rect 3240 15920 3292 15929
rect 6736 15920 6788 15972
rect 10968 16056 11020 16108
rect 9772 15920 9824 15972
rect 15384 16124 15436 16176
rect 14832 16099 14884 16108
rect 14832 16065 14841 16099
rect 14841 16065 14875 16099
rect 14875 16065 14884 16099
rect 14832 16056 14884 16065
rect 13728 15988 13780 16040
rect 14188 16031 14240 16040
rect 14188 15997 14197 16031
rect 14197 15997 14231 16031
rect 14231 15997 14240 16031
rect 14188 15988 14240 15997
rect 15752 16031 15804 16040
rect 13360 15920 13412 15972
rect 15752 15997 15761 16031
rect 15761 15997 15795 16031
rect 15795 15997 15804 16031
rect 15752 15988 15804 15997
rect 16396 15988 16448 16040
rect 18328 15988 18380 16040
rect 19248 16056 19300 16108
rect 19432 16056 19484 16108
rect 17500 15920 17552 15972
rect 18052 15920 18104 15972
rect 21180 15988 21232 16040
rect 22468 16031 22520 16040
rect 22468 15997 22477 16031
rect 22477 15997 22511 16031
rect 22511 15997 22520 16031
rect 22468 15988 22520 15997
rect 25228 16031 25280 16040
rect 25228 15997 25272 16031
rect 25272 15997 25280 16031
rect 25228 15988 25280 15997
rect 19892 15963 19944 15972
rect 19892 15929 19901 15963
rect 19901 15929 19935 15963
rect 19935 15929 19944 15963
rect 19892 15920 19944 15929
rect 19984 15963 20036 15972
rect 19984 15929 19993 15963
rect 19993 15929 20027 15963
rect 20027 15929 20036 15963
rect 19984 15920 20036 15929
rect 20720 15920 20772 15972
rect 2044 15895 2096 15904
rect 2044 15861 2053 15895
rect 2053 15861 2087 15895
rect 2087 15861 2096 15895
rect 2044 15852 2096 15861
rect 4896 15852 4948 15904
rect 6920 15895 6972 15904
rect 6920 15861 6929 15895
rect 6929 15861 6963 15895
rect 6963 15861 6972 15895
rect 6920 15852 6972 15861
rect 8668 15895 8720 15904
rect 8668 15861 8677 15895
rect 8677 15861 8711 15895
rect 8711 15861 8720 15895
rect 8668 15852 8720 15861
rect 8944 15895 8996 15904
rect 8944 15861 8953 15895
rect 8953 15861 8987 15895
rect 8987 15861 8996 15895
rect 8944 15852 8996 15861
rect 12164 15895 12216 15904
rect 12164 15861 12173 15895
rect 12173 15861 12207 15895
rect 12207 15861 12216 15895
rect 12164 15852 12216 15861
rect 14096 15895 14148 15904
rect 14096 15861 14105 15895
rect 14105 15861 14139 15895
rect 14139 15861 14148 15895
rect 14096 15852 14148 15861
rect 15660 15852 15712 15904
rect 24400 15963 24452 15972
rect 24400 15929 24409 15963
rect 24409 15929 24443 15963
rect 24443 15929 24452 15963
rect 24400 15920 24452 15929
rect 23480 15895 23532 15904
rect 23480 15861 23489 15895
rect 23489 15861 23523 15895
rect 23523 15861 23532 15895
rect 23480 15852 23532 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 4436 15648 4488 15700
rect 6092 15648 6144 15700
rect 6920 15648 6972 15700
rect 8300 15691 8352 15700
rect 8300 15657 8309 15691
rect 8309 15657 8343 15691
rect 8343 15657 8352 15691
rect 8300 15648 8352 15657
rect 9128 15691 9180 15700
rect 9128 15657 9137 15691
rect 9137 15657 9171 15691
rect 9171 15657 9180 15691
rect 9128 15648 9180 15657
rect 9956 15691 10008 15700
rect 9956 15657 9965 15691
rect 9965 15657 9999 15691
rect 9999 15657 10008 15691
rect 9956 15648 10008 15657
rect 2504 15580 2556 15632
rect 3240 15580 3292 15632
rect 1860 15512 1912 15564
rect 4804 15555 4856 15564
rect 4804 15521 4813 15555
rect 4813 15521 4847 15555
rect 4847 15521 4856 15555
rect 4804 15512 4856 15521
rect 6552 15555 6604 15564
rect 6552 15521 6561 15555
rect 6561 15521 6595 15555
rect 6595 15521 6604 15555
rect 6552 15512 6604 15521
rect 7288 15512 7340 15564
rect 8024 15555 8076 15564
rect 8024 15521 8033 15555
rect 8033 15521 8067 15555
rect 8067 15521 8076 15555
rect 8024 15512 8076 15521
rect 8116 15512 8168 15564
rect 9772 15555 9824 15564
rect 2504 15487 2556 15496
rect 2504 15453 2513 15487
rect 2513 15453 2547 15487
rect 2547 15453 2556 15487
rect 2504 15444 2556 15453
rect 2872 15444 2924 15496
rect 5172 15444 5224 15496
rect 9772 15521 9781 15555
rect 9781 15521 9815 15555
rect 9815 15521 9824 15555
rect 9772 15512 9824 15521
rect 11336 15648 11388 15700
rect 11520 15691 11572 15700
rect 11520 15657 11529 15691
rect 11529 15657 11563 15691
rect 11563 15657 11572 15691
rect 11520 15648 11572 15657
rect 14188 15648 14240 15700
rect 15752 15691 15804 15700
rect 15752 15657 15761 15691
rect 15761 15657 15795 15691
rect 15795 15657 15804 15691
rect 15752 15648 15804 15657
rect 16948 15691 17000 15700
rect 16948 15657 16957 15691
rect 16957 15657 16991 15691
rect 16991 15657 17000 15691
rect 16948 15648 17000 15657
rect 17500 15648 17552 15700
rect 21088 15648 21140 15700
rect 24124 15691 24176 15700
rect 24124 15657 24133 15691
rect 24133 15657 24167 15691
rect 24167 15657 24176 15691
rect 24124 15648 24176 15657
rect 24768 15691 24820 15700
rect 24768 15657 24777 15691
rect 24777 15657 24811 15691
rect 24811 15657 24820 15691
rect 24768 15648 24820 15657
rect 11704 15555 11756 15564
rect 9036 15444 9088 15496
rect 11704 15521 11713 15555
rect 11713 15521 11747 15555
rect 11747 15521 11756 15555
rect 11704 15512 11756 15521
rect 13268 15555 13320 15564
rect 13268 15521 13277 15555
rect 13277 15521 13311 15555
rect 13311 15521 13320 15555
rect 13268 15512 13320 15521
rect 13360 15555 13412 15564
rect 13360 15521 13369 15555
rect 13369 15521 13403 15555
rect 13403 15521 13412 15555
rect 13544 15555 13596 15564
rect 13360 15512 13412 15521
rect 13544 15521 13553 15555
rect 13553 15521 13587 15555
rect 13587 15521 13596 15555
rect 13544 15512 13596 15521
rect 16028 15555 16080 15564
rect 16028 15521 16037 15555
rect 16037 15521 16071 15555
rect 16071 15521 16080 15555
rect 16028 15512 16080 15521
rect 16120 15512 16172 15564
rect 16396 15555 16448 15564
rect 16396 15521 16405 15555
rect 16405 15521 16439 15555
rect 16439 15521 16448 15555
rect 16396 15512 16448 15521
rect 16580 15512 16632 15564
rect 17868 15512 17920 15564
rect 18972 15580 19024 15632
rect 19524 15580 19576 15632
rect 21272 15623 21324 15632
rect 21272 15589 21281 15623
rect 21281 15589 21315 15623
rect 21315 15589 21324 15623
rect 21272 15580 21324 15589
rect 23112 15623 23164 15632
rect 23112 15589 23121 15623
rect 23121 15589 23155 15623
rect 23155 15589 23164 15623
rect 23112 15580 23164 15589
rect 23204 15623 23256 15632
rect 23204 15589 23213 15623
rect 23213 15589 23247 15623
rect 23247 15589 23256 15623
rect 23204 15580 23256 15589
rect 23572 15580 23624 15632
rect 24400 15580 24452 15632
rect 19248 15512 19300 15564
rect 24584 15555 24636 15564
rect 24584 15521 24593 15555
rect 24593 15521 24627 15555
rect 24627 15521 24636 15555
rect 24584 15512 24636 15521
rect 24860 15512 24912 15564
rect 11428 15444 11480 15496
rect 13820 15487 13872 15496
rect 13820 15453 13829 15487
rect 13829 15453 13863 15487
rect 13863 15453 13872 15487
rect 13820 15444 13872 15453
rect 16488 15487 16540 15496
rect 16488 15453 16497 15487
rect 16497 15453 16531 15487
rect 16531 15453 16540 15487
rect 16488 15444 16540 15453
rect 19432 15444 19484 15496
rect 21180 15487 21232 15496
rect 21180 15453 21189 15487
rect 21189 15453 21223 15487
rect 21223 15453 21232 15487
rect 21180 15444 21232 15453
rect 21824 15487 21876 15496
rect 21824 15453 21833 15487
rect 21833 15453 21867 15487
rect 21867 15453 21876 15487
rect 21824 15444 21876 15453
rect 1952 15376 2004 15428
rect 1676 15308 1728 15360
rect 13176 15308 13228 15360
rect 15292 15308 15344 15360
rect 18696 15308 18748 15360
rect 19984 15351 20036 15360
rect 19984 15317 19993 15351
rect 19993 15317 20027 15351
rect 20027 15317 20036 15351
rect 19984 15308 20036 15317
rect 21916 15308 21968 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 2504 15104 2556 15156
rect 9036 15104 9088 15156
rect 9772 15104 9824 15156
rect 11704 15147 11756 15156
rect 11704 15113 11713 15147
rect 11713 15113 11747 15147
rect 11747 15113 11756 15147
rect 11704 15104 11756 15113
rect 14464 15147 14516 15156
rect 14464 15113 14473 15147
rect 14473 15113 14507 15147
rect 14507 15113 14516 15147
rect 14464 15104 14516 15113
rect 15752 15104 15804 15156
rect 17500 15147 17552 15156
rect 17500 15113 17509 15147
rect 17509 15113 17543 15147
rect 17543 15113 17552 15147
rect 17500 15104 17552 15113
rect 17960 15104 18012 15156
rect 18972 15104 19024 15156
rect 19524 15147 19576 15156
rect 19524 15113 19533 15147
rect 19533 15113 19567 15147
rect 19567 15113 19576 15147
rect 19524 15104 19576 15113
rect 21272 15147 21324 15156
rect 4804 15036 4856 15088
rect 8024 15079 8076 15088
rect 8024 15045 8033 15079
rect 8033 15045 8067 15079
rect 8067 15045 8076 15079
rect 8024 15036 8076 15045
rect 8300 15036 8352 15088
rect 2320 15011 2372 15020
rect 2320 14977 2329 15011
rect 2329 14977 2363 15011
rect 2363 14977 2372 15011
rect 2320 14968 2372 14977
rect 3240 14968 3292 15020
rect 3884 15011 3936 15020
rect 3884 14977 3893 15011
rect 3893 14977 3927 15011
rect 3927 14977 3936 15011
rect 3884 14968 3936 14977
rect 4160 15011 4212 15020
rect 4160 14977 4169 15011
rect 4169 14977 4203 15011
rect 4203 14977 4212 15011
rect 4160 14968 4212 14977
rect 6920 15011 6972 15020
rect 6920 14977 6929 15011
rect 6929 14977 6963 15011
rect 6963 14977 6972 15011
rect 6920 14968 6972 14977
rect 9128 15011 9180 15020
rect 9128 14977 9137 15011
rect 9137 14977 9171 15011
rect 9171 14977 9180 15011
rect 9128 14968 9180 14977
rect 11060 15036 11112 15088
rect 13268 15036 13320 15088
rect 14648 15036 14700 15088
rect 4528 14900 4580 14952
rect 2688 14832 2740 14884
rect 3976 14875 4028 14884
rect 3976 14841 3985 14875
rect 3985 14841 4019 14875
rect 4019 14841 4028 14875
rect 3976 14832 4028 14841
rect 7012 14875 7064 14884
rect 3240 14807 3292 14816
rect 3240 14773 3249 14807
rect 3249 14773 3283 14807
rect 3283 14773 3292 14807
rect 3240 14764 3292 14773
rect 4804 14807 4856 14816
rect 4804 14773 4813 14807
rect 4813 14773 4847 14807
rect 4847 14773 4856 14807
rect 4804 14764 4856 14773
rect 5172 14807 5224 14816
rect 5172 14773 5181 14807
rect 5181 14773 5215 14807
rect 5215 14773 5224 14807
rect 5172 14764 5224 14773
rect 5264 14764 5316 14816
rect 6552 14807 6604 14816
rect 6552 14773 6561 14807
rect 6561 14773 6595 14807
rect 6595 14773 6604 14807
rect 6552 14764 6604 14773
rect 7012 14841 7021 14875
rect 7021 14841 7055 14875
rect 7055 14841 7064 14875
rect 7012 14832 7064 14841
rect 7656 14832 7708 14884
rect 7196 14764 7248 14816
rect 9128 14832 9180 14884
rect 9772 14764 9824 14816
rect 10784 14943 10836 14952
rect 10784 14909 10793 14943
rect 10793 14909 10827 14943
rect 10827 14909 10836 14943
rect 10784 14900 10836 14909
rect 11704 14900 11756 14952
rect 11704 14764 11756 14816
rect 12808 14968 12860 15020
rect 13176 15011 13228 15020
rect 13176 14977 13185 15011
rect 13185 14977 13219 15011
rect 13219 14977 13228 15011
rect 13176 14968 13228 14977
rect 19432 15036 19484 15088
rect 18604 15011 18656 15020
rect 16028 14943 16080 14952
rect 16028 14909 16037 14943
rect 16037 14909 16071 14943
rect 16071 14909 16080 14943
rect 16672 14943 16724 14952
rect 16028 14900 16080 14909
rect 16672 14909 16681 14943
rect 16681 14909 16715 14943
rect 16715 14909 16724 14943
rect 16672 14900 16724 14909
rect 18604 14977 18613 15011
rect 18613 14977 18647 15011
rect 18647 14977 18656 15011
rect 18604 14968 18656 14977
rect 17132 14875 17184 14884
rect 17132 14841 17141 14875
rect 17141 14841 17175 14875
rect 17175 14841 17184 14875
rect 17132 14832 17184 14841
rect 18696 14875 18748 14884
rect 18696 14841 18705 14875
rect 18705 14841 18739 14875
rect 18739 14841 18748 14875
rect 21272 15113 21281 15147
rect 21281 15113 21315 15147
rect 21315 15113 21324 15147
rect 21272 15104 21324 15113
rect 23112 15147 23164 15156
rect 23112 15113 23121 15147
rect 23121 15113 23155 15147
rect 23155 15113 23164 15147
rect 23112 15104 23164 15113
rect 23480 15147 23532 15156
rect 23480 15113 23489 15147
rect 23489 15113 23523 15147
rect 23523 15113 23532 15147
rect 23480 15104 23532 15113
rect 24860 15104 24912 15156
rect 20076 15011 20128 15020
rect 20076 14977 20085 15011
rect 20085 14977 20119 15011
rect 20119 14977 20128 15011
rect 20076 14968 20128 14977
rect 24124 14968 24176 15020
rect 21824 14943 21876 14952
rect 21824 14909 21833 14943
rect 21833 14909 21867 14943
rect 21867 14909 21876 14943
rect 21824 14900 21876 14909
rect 24952 14900 25004 14952
rect 18696 14832 18748 14841
rect 23480 14832 23532 14884
rect 24676 14875 24728 14884
rect 24676 14841 24685 14875
rect 24685 14841 24719 14875
rect 24719 14841 24728 14875
rect 24676 14832 24728 14841
rect 13544 14807 13596 14816
rect 13544 14773 13553 14807
rect 13553 14773 13587 14807
rect 13587 14773 13596 14807
rect 13912 14807 13964 14816
rect 13544 14764 13596 14773
rect 13912 14773 13921 14807
rect 13921 14773 13955 14807
rect 13955 14773 13964 14807
rect 13912 14764 13964 14773
rect 21732 14807 21784 14816
rect 21732 14773 21741 14807
rect 21741 14773 21775 14807
rect 21775 14773 21784 14807
rect 21732 14764 21784 14773
rect 22744 14807 22796 14816
rect 22744 14773 22753 14807
rect 22753 14773 22787 14807
rect 22787 14773 22796 14807
rect 22744 14764 22796 14773
rect 25688 14807 25740 14816
rect 25688 14773 25697 14807
rect 25697 14773 25731 14807
rect 25731 14773 25740 14807
rect 25688 14764 25740 14773
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 1860 14603 1912 14612
rect 1860 14569 1869 14603
rect 1869 14569 1903 14603
rect 1903 14569 1912 14603
rect 1860 14560 1912 14569
rect 2136 14560 2188 14612
rect 2320 14603 2372 14612
rect 2320 14569 2329 14603
rect 2329 14569 2363 14603
rect 2363 14569 2372 14603
rect 2320 14560 2372 14569
rect 3884 14603 3936 14612
rect 3884 14569 3893 14603
rect 3893 14569 3927 14603
rect 3927 14569 3936 14603
rect 3884 14560 3936 14569
rect 3976 14560 4028 14612
rect 7012 14560 7064 14612
rect 7748 14560 7800 14612
rect 9036 14603 9088 14612
rect 9036 14569 9045 14603
rect 9045 14569 9079 14603
rect 9079 14569 9088 14603
rect 9036 14560 9088 14569
rect 11428 14560 11480 14612
rect 12532 14603 12584 14612
rect 12532 14569 12541 14603
rect 12541 14569 12575 14603
rect 12575 14569 12584 14603
rect 12532 14560 12584 14569
rect 13360 14603 13412 14612
rect 13360 14569 13369 14603
rect 13369 14569 13403 14603
rect 13403 14569 13412 14603
rect 13360 14560 13412 14569
rect 14464 14560 14516 14612
rect 18604 14560 18656 14612
rect 19340 14560 19392 14612
rect 20076 14560 20128 14612
rect 21180 14603 21232 14612
rect 21180 14569 21189 14603
rect 21189 14569 21223 14603
rect 21223 14569 21232 14603
rect 21180 14560 21232 14569
rect 23204 14560 23256 14612
rect 2688 14492 2740 14544
rect 4896 14492 4948 14544
rect 6644 14535 6696 14544
rect 6644 14501 6647 14535
rect 6647 14501 6681 14535
rect 6681 14501 6696 14535
rect 6644 14492 6696 14501
rect 10048 14535 10100 14544
rect 10048 14501 10051 14535
rect 10051 14501 10085 14535
rect 10085 14501 10100 14535
rect 10048 14492 10100 14501
rect 2136 14424 2188 14476
rect 2320 14424 2372 14476
rect 4436 14467 4488 14476
rect 4436 14433 4445 14467
rect 4445 14433 4479 14467
rect 4479 14433 4488 14467
rect 4436 14424 4488 14433
rect 6276 14467 6328 14476
rect 6276 14433 6285 14467
rect 6285 14433 6319 14467
rect 6319 14433 6328 14467
rect 6276 14424 6328 14433
rect 8208 14467 8260 14476
rect 8208 14433 8217 14467
rect 8217 14433 8251 14467
rect 8251 14433 8260 14467
rect 8208 14424 8260 14433
rect 8484 14467 8536 14476
rect 8484 14433 8493 14467
rect 8493 14433 8527 14467
rect 8527 14433 8536 14467
rect 8484 14424 8536 14433
rect 8668 14424 8720 14476
rect 12808 14492 12860 14544
rect 14372 14535 14424 14544
rect 14372 14501 14381 14535
rect 14381 14501 14415 14535
rect 14415 14501 14424 14535
rect 14372 14492 14424 14501
rect 14648 14535 14700 14544
rect 14648 14501 14657 14535
rect 14657 14501 14691 14535
rect 14691 14501 14700 14535
rect 14648 14492 14700 14501
rect 12348 14467 12400 14476
rect 12348 14433 12357 14467
rect 12357 14433 12391 14467
rect 12391 14433 12400 14467
rect 12348 14424 12400 14433
rect 13268 14424 13320 14476
rect 13912 14467 13964 14476
rect 13912 14433 13921 14467
rect 13921 14433 13955 14467
rect 13955 14433 13964 14467
rect 13912 14424 13964 14433
rect 15936 14492 15988 14544
rect 18972 14535 19024 14544
rect 15844 14424 15896 14476
rect 16488 14424 16540 14476
rect 17408 14424 17460 14476
rect 17592 14467 17644 14476
rect 17592 14433 17601 14467
rect 17601 14433 17635 14467
rect 17635 14433 17644 14467
rect 17592 14424 17644 14433
rect 18972 14501 18975 14535
rect 18975 14501 19009 14535
rect 19009 14501 19024 14535
rect 18972 14492 19024 14501
rect 21732 14492 21784 14544
rect 24676 14492 24728 14544
rect 24952 14535 25004 14544
rect 24952 14501 24961 14535
rect 24961 14501 24995 14535
rect 24995 14501 25004 14535
rect 24952 14492 25004 14501
rect 20168 14424 20220 14476
rect 2596 14356 2648 14408
rect 2872 14356 2924 14408
rect 8760 14399 8812 14408
rect 8760 14365 8769 14399
rect 8769 14365 8803 14399
rect 8803 14365 8812 14399
rect 8760 14356 8812 14365
rect 16672 14356 16724 14408
rect 17776 14399 17828 14408
rect 17776 14365 17785 14399
rect 17785 14365 17819 14399
rect 17819 14365 17828 14399
rect 17776 14356 17828 14365
rect 21456 14399 21508 14408
rect 21456 14365 21465 14399
rect 21465 14365 21499 14399
rect 21499 14365 21508 14399
rect 21456 14356 21508 14365
rect 23388 14356 23440 14408
rect 23664 14399 23716 14408
rect 23664 14365 23673 14399
rect 23673 14365 23707 14399
rect 23707 14365 23716 14399
rect 23664 14356 23716 14365
rect 25596 14356 25648 14408
rect 1860 14288 1912 14340
rect 4160 14288 4212 14340
rect 11980 14288 12032 14340
rect 12164 14331 12216 14340
rect 12164 14297 12173 14331
rect 12173 14297 12207 14331
rect 12207 14297 12216 14331
rect 12164 14288 12216 14297
rect 14004 14288 14056 14340
rect 16764 14288 16816 14340
rect 1768 14220 1820 14272
rect 4344 14263 4396 14272
rect 4344 14229 4353 14263
rect 4353 14229 4387 14263
rect 4387 14229 4396 14263
rect 4344 14220 4396 14229
rect 5080 14220 5132 14272
rect 5356 14220 5408 14272
rect 7196 14263 7248 14272
rect 7196 14229 7205 14263
rect 7205 14229 7239 14263
rect 7239 14229 7248 14263
rect 7196 14220 7248 14229
rect 19524 14263 19576 14272
rect 19524 14229 19533 14263
rect 19533 14229 19567 14263
rect 19567 14229 19576 14263
rect 19524 14220 19576 14229
rect 23112 14263 23164 14272
rect 23112 14229 23121 14263
rect 23121 14229 23155 14263
rect 23155 14229 23164 14263
rect 23112 14220 23164 14229
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 1584 14059 1636 14068
rect 1584 14025 1593 14059
rect 1593 14025 1627 14059
rect 1627 14025 1636 14059
rect 1584 14016 1636 14025
rect 2596 14016 2648 14068
rect 4436 14016 4488 14068
rect 6276 14016 6328 14068
rect 6644 14059 6696 14068
rect 6644 14025 6653 14059
rect 6653 14025 6687 14059
rect 6687 14025 6696 14059
rect 6644 14016 6696 14025
rect 7748 14059 7800 14068
rect 7748 14025 7757 14059
rect 7757 14025 7791 14059
rect 7791 14025 7800 14059
rect 7748 14016 7800 14025
rect 8208 14016 8260 14068
rect 8668 14016 8720 14068
rect 14004 14059 14056 14068
rect 14004 14025 14013 14059
rect 14013 14025 14047 14059
rect 14047 14025 14056 14059
rect 15292 14059 15344 14068
rect 14004 14016 14056 14025
rect 1400 13948 1452 14000
rect 2136 13948 2188 14000
rect 3516 13948 3568 14000
rect 2872 13923 2924 13932
rect 2872 13889 2881 13923
rect 2881 13889 2915 13923
rect 2915 13889 2924 13923
rect 2872 13880 2924 13889
rect 5540 13880 5592 13932
rect 6736 13880 6788 13932
rect 1584 13676 1636 13728
rect 4160 13812 4212 13864
rect 4344 13855 4396 13864
rect 4344 13821 4353 13855
rect 4353 13821 4387 13855
rect 4387 13821 4396 13855
rect 4344 13812 4396 13821
rect 3332 13744 3384 13796
rect 4436 13744 4488 13796
rect 4896 13744 4948 13796
rect 11520 13991 11572 14000
rect 8760 13880 8812 13932
rect 9312 13923 9364 13932
rect 9312 13889 9321 13923
rect 9321 13889 9355 13923
rect 9355 13889 9364 13923
rect 9312 13880 9364 13889
rect 8484 13855 8536 13864
rect 8484 13821 8493 13855
rect 8493 13821 8527 13855
rect 8527 13821 8536 13855
rect 8484 13812 8536 13821
rect 11520 13957 11529 13991
rect 11529 13957 11563 13991
rect 11563 13957 11572 13991
rect 11520 13948 11572 13957
rect 13360 13948 13412 14000
rect 15292 14025 15301 14059
rect 15301 14025 15335 14059
rect 15335 14025 15344 14059
rect 15292 14016 15344 14025
rect 16120 14059 16172 14068
rect 16120 14025 16129 14059
rect 16129 14025 16163 14059
rect 16163 14025 16172 14059
rect 16120 14016 16172 14025
rect 18972 14016 19024 14068
rect 19524 14016 19576 14068
rect 20904 14016 20956 14068
rect 21456 14016 21508 14068
rect 22468 14059 22520 14068
rect 22468 14025 22477 14059
rect 22477 14025 22511 14059
rect 22511 14025 22520 14059
rect 22468 14016 22520 14025
rect 23204 14059 23256 14068
rect 23204 14025 23213 14059
rect 23213 14025 23247 14059
rect 23247 14025 23256 14059
rect 23204 14016 23256 14025
rect 24952 14016 25004 14068
rect 16028 13948 16080 14000
rect 17592 13948 17644 14000
rect 18880 13948 18932 14000
rect 19892 13991 19944 14000
rect 19892 13957 19901 13991
rect 19901 13957 19935 13991
rect 19935 13957 19944 13991
rect 19892 13948 19944 13957
rect 20168 13991 20220 14000
rect 20168 13957 20177 13991
rect 20177 13957 20211 13991
rect 20211 13957 20220 13991
rect 20168 13948 20220 13957
rect 23112 13948 23164 14000
rect 24676 13991 24728 14000
rect 24676 13957 24685 13991
rect 24685 13957 24719 13991
rect 24719 13957 24728 13991
rect 25412 13991 25464 14000
rect 24676 13948 24728 13957
rect 25412 13957 25421 13991
rect 25421 13957 25455 13991
rect 25455 13957 25464 13991
rect 25412 13948 25464 13957
rect 12440 13880 12492 13932
rect 14740 13923 14792 13932
rect 14740 13889 14749 13923
rect 14749 13889 14783 13923
rect 14783 13889 14792 13923
rect 14740 13880 14792 13889
rect 16764 13880 16816 13932
rect 20996 13880 21048 13932
rect 21180 13923 21232 13932
rect 21180 13889 21189 13923
rect 21189 13889 21223 13923
rect 21223 13889 21232 13923
rect 21180 13880 21232 13889
rect 25504 13880 25556 13932
rect 10048 13812 10100 13864
rect 11336 13855 11388 13864
rect 11336 13821 11345 13855
rect 11345 13821 11379 13855
rect 11379 13821 11388 13855
rect 11336 13812 11388 13821
rect 12808 13812 12860 13864
rect 4528 13676 4580 13728
rect 9864 13676 9916 13728
rect 10692 13676 10744 13728
rect 12164 13744 12216 13796
rect 11428 13676 11480 13728
rect 11704 13676 11756 13728
rect 11796 13676 11848 13728
rect 12348 13676 12400 13728
rect 13912 13812 13964 13864
rect 14464 13812 14516 13864
rect 18328 13855 18380 13864
rect 18328 13821 18337 13855
rect 18337 13821 18371 13855
rect 18371 13821 18380 13855
rect 18328 13812 18380 13821
rect 22284 13855 22336 13864
rect 22284 13821 22293 13855
rect 22293 13821 22327 13855
rect 22327 13821 22336 13855
rect 22284 13812 22336 13821
rect 14648 13744 14700 13796
rect 16580 13787 16632 13796
rect 16580 13753 16589 13787
rect 16589 13753 16623 13787
rect 16623 13753 16632 13787
rect 16580 13744 16632 13753
rect 17316 13744 17368 13796
rect 20904 13787 20956 13796
rect 20904 13753 20913 13787
rect 20913 13753 20947 13787
rect 20947 13753 20956 13787
rect 20904 13744 20956 13753
rect 23296 13744 23348 13796
rect 17408 13676 17460 13728
rect 17592 13676 17644 13728
rect 18512 13676 18564 13728
rect 18972 13676 19024 13728
rect 21732 13719 21784 13728
rect 21732 13685 21741 13719
rect 21741 13685 21775 13719
rect 21775 13685 21784 13719
rect 21732 13676 21784 13685
rect 25596 13855 25648 13864
rect 25596 13821 25640 13855
rect 25640 13821 25648 13855
rect 25596 13812 25648 13821
rect 24124 13787 24176 13796
rect 24124 13753 24133 13787
rect 24133 13753 24167 13787
rect 24167 13753 24176 13787
rect 24124 13744 24176 13753
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 1584 13515 1636 13524
rect 1584 13481 1593 13515
rect 1593 13481 1627 13515
rect 1627 13481 1636 13515
rect 1584 13472 1636 13481
rect 3056 13515 3108 13524
rect 3056 13481 3065 13515
rect 3065 13481 3099 13515
rect 3099 13481 3108 13515
rect 3056 13472 3108 13481
rect 3516 13515 3568 13524
rect 3516 13481 3525 13515
rect 3525 13481 3559 13515
rect 3559 13481 3568 13515
rect 3516 13472 3568 13481
rect 4344 13472 4396 13524
rect 6736 13515 6788 13524
rect 6736 13481 6745 13515
rect 6745 13481 6779 13515
rect 6779 13481 6788 13515
rect 6736 13472 6788 13481
rect 9312 13515 9364 13524
rect 2136 13404 2188 13456
rect 2412 13404 2464 13456
rect 4436 13447 4488 13456
rect 4436 13413 4445 13447
rect 4445 13413 4479 13447
rect 4479 13413 4488 13447
rect 4436 13404 4488 13413
rect 6184 13404 6236 13456
rect 7196 13404 7248 13456
rect 7656 13447 7708 13456
rect 7656 13413 7665 13447
rect 7665 13413 7699 13447
rect 7699 13413 7708 13447
rect 7656 13404 7708 13413
rect 9312 13481 9321 13515
rect 9321 13481 9355 13515
rect 9355 13481 9364 13515
rect 9312 13472 9364 13481
rect 9864 13447 9916 13456
rect 9864 13413 9873 13447
rect 9873 13413 9907 13447
rect 9907 13413 9916 13447
rect 9864 13404 9916 13413
rect 11152 13472 11204 13524
rect 13360 13472 13412 13524
rect 14004 13472 14056 13524
rect 14648 13472 14700 13524
rect 15844 13515 15896 13524
rect 15844 13481 15853 13515
rect 15853 13481 15887 13515
rect 15887 13481 15896 13515
rect 15844 13472 15896 13481
rect 18604 13472 18656 13524
rect 4896 13379 4948 13388
rect 4896 13345 4905 13379
rect 4905 13345 4939 13379
rect 4939 13345 4948 13379
rect 4896 13336 4948 13345
rect 5172 13379 5224 13388
rect 5172 13345 5181 13379
rect 5181 13345 5215 13379
rect 5215 13345 5224 13379
rect 5172 13336 5224 13345
rect 8576 13379 8628 13388
rect 8576 13345 8585 13379
rect 8585 13345 8619 13379
rect 8619 13345 8628 13379
rect 8576 13336 8628 13345
rect 11152 13379 11204 13388
rect 11152 13345 11161 13379
rect 11161 13345 11195 13379
rect 11195 13345 11204 13379
rect 11152 13336 11204 13345
rect 11336 13336 11388 13388
rect 7104 13268 7156 13320
rect 9496 13268 9548 13320
rect 9772 13311 9824 13320
rect 9772 13277 9781 13311
rect 9781 13277 9815 13311
rect 9815 13277 9824 13311
rect 9772 13268 9824 13277
rect 10048 13311 10100 13320
rect 10048 13277 10057 13311
rect 10057 13277 10091 13311
rect 10091 13277 10100 13311
rect 10048 13268 10100 13277
rect 11244 13268 11296 13320
rect 11796 13404 11848 13456
rect 17132 13404 17184 13456
rect 17316 13447 17368 13456
rect 17316 13413 17325 13447
rect 17325 13413 17359 13447
rect 17359 13413 17368 13447
rect 17316 13404 17368 13413
rect 18052 13404 18104 13456
rect 18972 13472 19024 13524
rect 20996 13472 21048 13524
rect 21640 13447 21692 13456
rect 21640 13413 21649 13447
rect 21649 13413 21683 13447
rect 21683 13413 21692 13447
rect 21640 13404 21692 13413
rect 23296 13447 23348 13456
rect 23296 13413 23305 13447
rect 23305 13413 23339 13447
rect 23339 13413 23348 13447
rect 23296 13404 23348 13413
rect 23388 13404 23440 13456
rect 24768 13447 24820 13456
rect 24768 13413 24777 13447
rect 24777 13413 24811 13447
rect 24811 13413 24820 13447
rect 24768 13404 24820 13413
rect 24860 13447 24912 13456
rect 24860 13413 24869 13447
rect 24869 13413 24903 13447
rect 24903 13413 24912 13447
rect 25412 13447 25464 13456
rect 24860 13404 24912 13413
rect 25412 13413 25421 13447
rect 25421 13413 25455 13447
rect 25455 13413 25464 13447
rect 25412 13404 25464 13413
rect 11888 13379 11940 13388
rect 11888 13345 11897 13379
rect 11897 13345 11931 13379
rect 11931 13345 11940 13379
rect 11888 13336 11940 13345
rect 13176 13379 13228 13388
rect 13176 13345 13185 13379
rect 13185 13345 13219 13379
rect 13219 13345 13228 13379
rect 13176 13336 13228 13345
rect 13452 13379 13504 13388
rect 13452 13345 13461 13379
rect 13461 13345 13495 13379
rect 13495 13345 13504 13379
rect 13452 13336 13504 13345
rect 15292 13379 15344 13388
rect 15292 13345 15301 13379
rect 15301 13345 15335 13379
rect 15335 13345 15344 13379
rect 15292 13336 15344 13345
rect 19800 13336 19852 13388
rect 20812 13336 20864 13388
rect 2044 13200 2096 13252
rect 2688 13243 2740 13252
rect 2688 13209 2697 13243
rect 2697 13209 2731 13243
rect 2731 13209 2740 13243
rect 2688 13200 2740 13209
rect 6000 13132 6052 13184
rect 11796 13200 11848 13252
rect 13268 13243 13320 13252
rect 13268 13209 13277 13243
rect 13277 13209 13311 13243
rect 13311 13209 13320 13243
rect 13268 13200 13320 13209
rect 14004 13268 14056 13320
rect 16764 13268 16816 13320
rect 17592 13200 17644 13252
rect 20720 13268 20772 13320
rect 22192 13311 22244 13320
rect 22192 13277 22201 13311
rect 22201 13277 22235 13311
rect 22235 13277 22244 13311
rect 22192 13268 22244 13277
rect 23848 13268 23900 13320
rect 12624 13132 12676 13184
rect 14280 13132 14332 13184
rect 14740 13132 14792 13184
rect 16580 13132 16632 13184
rect 17960 13175 18012 13184
rect 17960 13141 17969 13175
rect 17969 13141 18003 13175
rect 18003 13141 18012 13175
rect 17960 13132 18012 13141
rect 24124 13175 24176 13184
rect 24124 13141 24133 13175
rect 24133 13141 24167 13175
rect 24167 13141 24176 13175
rect 24124 13132 24176 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 2228 12928 2280 12980
rect 7104 12928 7156 12980
rect 8576 12971 8628 12980
rect 8576 12937 8585 12971
rect 8585 12937 8619 12971
rect 8619 12937 8628 12971
rect 8576 12928 8628 12937
rect 9864 12928 9916 12980
rect 15292 12928 15344 12980
rect 16580 12971 16632 12980
rect 16580 12937 16589 12971
rect 16589 12937 16623 12971
rect 16623 12937 16632 12971
rect 16580 12928 16632 12937
rect 17132 12928 17184 12980
rect 17316 12928 17368 12980
rect 19800 12971 19852 12980
rect 19800 12937 19809 12971
rect 19809 12937 19843 12971
rect 19843 12937 19852 12971
rect 19800 12928 19852 12937
rect 21640 12928 21692 12980
rect 2688 12903 2740 12912
rect 2688 12869 2697 12903
rect 2697 12869 2731 12903
rect 2731 12869 2740 12903
rect 2688 12860 2740 12869
rect 4436 12903 4488 12912
rect 4436 12869 4445 12903
rect 4445 12869 4479 12903
rect 4479 12869 4488 12903
rect 5540 12903 5592 12912
rect 4436 12860 4488 12869
rect 2412 12792 2464 12844
rect 5172 12792 5224 12844
rect 5540 12869 5549 12903
rect 5549 12869 5583 12903
rect 5583 12869 5592 12903
rect 5540 12860 5592 12869
rect 12900 12903 12952 12912
rect 12900 12869 12909 12903
rect 12909 12869 12943 12903
rect 12943 12869 12952 12903
rect 12900 12860 12952 12869
rect 15752 12860 15804 12912
rect 18512 12860 18564 12912
rect 11520 12792 11572 12844
rect 5356 12767 5408 12776
rect 5356 12733 5365 12767
rect 5365 12733 5399 12767
rect 5399 12733 5408 12767
rect 5356 12724 5408 12733
rect 6552 12724 6604 12776
rect 2504 12656 2556 12708
rect 3884 12699 3936 12708
rect 3884 12665 3893 12699
rect 3893 12665 3927 12699
rect 3927 12665 3936 12699
rect 3884 12656 3936 12665
rect 7564 12724 7616 12776
rect 11428 12767 11480 12776
rect 11428 12733 11437 12767
rect 11437 12733 11471 12767
rect 11471 12733 11480 12767
rect 11428 12724 11480 12733
rect 11888 12724 11940 12776
rect 12808 12767 12860 12776
rect 12808 12733 12817 12767
rect 12817 12733 12851 12767
rect 12851 12733 12860 12767
rect 14280 12792 14332 12844
rect 18604 12835 18656 12844
rect 18604 12801 18613 12835
rect 18613 12801 18647 12835
rect 18647 12801 18656 12835
rect 18604 12792 18656 12801
rect 20628 12835 20680 12844
rect 20628 12801 20637 12835
rect 20637 12801 20671 12835
rect 20671 12801 20680 12835
rect 20628 12792 20680 12801
rect 22008 12792 22060 12844
rect 22192 12835 22244 12844
rect 22192 12801 22201 12835
rect 22201 12801 22235 12835
rect 22235 12801 22244 12835
rect 22192 12792 22244 12801
rect 12808 12724 12860 12733
rect 14740 12724 14792 12776
rect 19340 12724 19392 12776
rect 7472 12656 7524 12708
rect 4344 12588 4396 12640
rect 4896 12588 4948 12640
rect 6000 12588 6052 12640
rect 6184 12631 6236 12640
rect 6184 12597 6193 12631
rect 6193 12597 6227 12631
rect 6227 12597 6236 12631
rect 6184 12588 6236 12597
rect 7104 12631 7156 12640
rect 7104 12597 7113 12631
rect 7113 12597 7147 12631
rect 7147 12597 7156 12631
rect 7104 12588 7156 12597
rect 8024 12588 8076 12640
rect 9036 12656 9088 12708
rect 11612 12656 11664 12708
rect 9680 12588 9732 12640
rect 11796 12631 11848 12640
rect 11796 12597 11805 12631
rect 11805 12597 11839 12631
rect 11839 12597 11848 12631
rect 12716 12656 12768 12708
rect 13268 12656 13320 12708
rect 15752 12656 15804 12708
rect 11796 12588 11848 12597
rect 12808 12588 12860 12640
rect 13452 12588 13504 12640
rect 18052 12588 18104 12640
rect 19248 12699 19300 12708
rect 19248 12665 19257 12699
rect 19257 12665 19291 12699
rect 19291 12665 19300 12699
rect 19248 12656 19300 12665
rect 21916 12656 21968 12708
rect 23296 12928 23348 12980
rect 23848 12971 23900 12980
rect 23848 12937 23857 12971
rect 23857 12937 23891 12971
rect 23891 12937 23900 12971
rect 23848 12928 23900 12937
rect 24768 12928 24820 12980
rect 24860 12928 24912 12980
rect 24584 12767 24636 12776
rect 24584 12733 24593 12767
rect 24593 12733 24627 12767
rect 24627 12733 24636 12767
rect 24584 12724 24636 12733
rect 23388 12656 23440 12708
rect 18788 12588 18840 12640
rect 20260 12588 20312 12640
rect 24216 12588 24268 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 2136 12427 2188 12436
rect 2136 12393 2145 12427
rect 2145 12393 2179 12427
rect 2179 12393 2188 12427
rect 2136 12384 2188 12393
rect 3884 12427 3936 12436
rect 3884 12393 3893 12427
rect 3893 12393 3927 12427
rect 3927 12393 3936 12427
rect 3884 12384 3936 12393
rect 4528 12384 4580 12436
rect 9496 12384 9548 12436
rect 1400 12044 1452 12096
rect 2044 12316 2096 12368
rect 3056 12359 3108 12368
rect 3056 12325 3065 12359
rect 3065 12325 3099 12359
rect 3099 12325 3108 12359
rect 3056 12316 3108 12325
rect 4252 12359 4304 12368
rect 4252 12325 4261 12359
rect 4261 12325 4295 12359
rect 4295 12325 4304 12359
rect 4252 12316 4304 12325
rect 7196 12316 7248 12368
rect 8024 12359 8076 12368
rect 8024 12325 8033 12359
rect 8033 12325 8067 12359
rect 8067 12325 8076 12359
rect 8024 12316 8076 12325
rect 8852 12316 8904 12368
rect 10140 12316 10192 12368
rect 6000 12248 6052 12300
rect 6552 12248 6604 12300
rect 10600 12248 10652 12300
rect 1860 12180 1912 12232
rect 2412 12223 2464 12232
rect 2412 12189 2421 12223
rect 2421 12189 2455 12223
rect 2455 12189 2464 12223
rect 2412 12180 2464 12189
rect 4160 12223 4212 12232
rect 4160 12189 4169 12223
rect 4169 12189 4203 12223
rect 4203 12189 4212 12223
rect 4160 12180 4212 12189
rect 4436 12223 4488 12232
rect 4436 12189 4445 12223
rect 4445 12189 4479 12223
rect 4479 12189 4488 12223
rect 4436 12180 4488 12189
rect 2044 12112 2096 12164
rect 9956 12180 10008 12232
rect 12164 12248 12216 12300
rect 13912 12291 13964 12300
rect 8484 12112 8536 12164
rect 9036 12112 9088 12164
rect 12256 12180 12308 12232
rect 13912 12257 13921 12291
rect 13921 12257 13955 12291
rect 13955 12257 13964 12291
rect 13912 12248 13964 12257
rect 14740 12248 14792 12300
rect 15752 12316 15804 12368
rect 17408 12316 17460 12368
rect 18420 12384 18472 12436
rect 18788 12427 18840 12436
rect 18788 12393 18797 12427
rect 18797 12393 18831 12427
rect 18831 12393 18840 12427
rect 18788 12384 18840 12393
rect 20260 12427 20312 12436
rect 20260 12393 20269 12427
rect 20269 12393 20303 12427
rect 20303 12393 20312 12427
rect 20260 12384 20312 12393
rect 20720 12427 20772 12436
rect 20720 12393 20729 12427
rect 20729 12393 20763 12427
rect 20763 12393 20772 12427
rect 20720 12384 20772 12393
rect 21272 12384 21324 12436
rect 22192 12384 22244 12436
rect 18512 12316 18564 12368
rect 18604 12316 18656 12368
rect 20812 12316 20864 12368
rect 22836 12316 22888 12368
rect 23572 12316 23624 12368
rect 24676 12316 24728 12368
rect 18052 12248 18104 12300
rect 19892 12291 19944 12300
rect 19892 12257 19910 12291
rect 19910 12257 19944 12291
rect 19892 12248 19944 12257
rect 18420 12180 18472 12232
rect 20720 12180 20772 12232
rect 21272 12223 21324 12232
rect 21272 12189 21281 12223
rect 21281 12189 21315 12223
rect 21315 12189 21324 12223
rect 21272 12180 21324 12189
rect 21548 12223 21600 12232
rect 21548 12189 21557 12223
rect 21557 12189 21591 12223
rect 21591 12189 21600 12223
rect 21548 12180 21600 12189
rect 11428 12112 11480 12164
rect 12808 12112 12860 12164
rect 22928 12180 22980 12232
rect 24216 12180 24268 12232
rect 23756 12112 23808 12164
rect 5356 12087 5408 12096
rect 5356 12053 5365 12087
rect 5365 12053 5399 12087
rect 5399 12053 5408 12087
rect 5356 12044 5408 12053
rect 6552 12044 6604 12096
rect 7564 12044 7616 12096
rect 9588 12044 9640 12096
rect 12256 12044 12308 12096
rect 13176 12044 13228 12096
rect 13544 12087 13596 12096
rect 13544 12053 13553 12087
rect 13553 12053 13587 12087
rect 13587 12053 13596 12087
rect 13544 12044 13596 12053
rect 14832 12044 14884 12096
rect 16764 12044 16816 12096
rect 21916 12044 21968 12096
rect 23664 12044 23716 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 4620 11840 4672 11892
rect 8852 11883 8904 11892
rect 4252 11772 4304 11824
rect 8852 11849 8861 11883
rect 8861 11849 8895 11883
rect 8895 11849 8904 11883
rect 8852 11840 8904 11849
rect 9680 11840 9732 11892
rect 10600 11840 10652 11892
rect 11980 11840 12032 11892
rect 12716 11883 12768 11892
rect 12716 11849 12725 11883
rect 12725 11849 12759 11883
rect 12759 11849 12768 11883
rect 12716 11840 12768 11849
rect 17316 11840 17368 11892
rect 19892 11840 19944 11892
rect 21088 11840 21140 11892
rect 22836 11840 22888 11892
rect 23572 11840 23624 11892
rect 24676 11883 24728 11892
rect 24676 11849 24685 11883
rect 24685 11849 24719 11883
rect 24719 11849 24728 11883
rect 24676 11840 24728 11849
rect 25412 11883 25464 11892
rect 25412 11849 25421 11883
rect 25421 11849 25455 11883
rect 25455 11849 25464 11883
rect 25412 11840 25464 11849
rect 6736 11772 6788 11824
rect 1768 11704 1820 11756
rect 2412 11747 2464 11756
rect 2412 11713 2421 11747
rect 2421 11713 2455 11747
rect 2455 11713 2464 11747
rect 2412 11704 2464 11713
rect 2780 11704 2832 11756
rect 3056 11747 3108 11756
rect 3056 11713 3065 11747
rect 3065 11713 3099 11747
rect 3099 11713 3108 11747
rect 3056 11704 3108 11713
rect 4528 11747 4580 11756
rect 4528 11713 4537 11747
rect 4537 11713 4571 11747
rect 4571 11713 4580 11747
rect 4528 11704 4580 11713
rect 6552 11636 6604 11688
rect 6828 11679 6880 11688
rect 6828 11645 6837 11679
rect 6837 11645 6871 11679
rect 6871 11645 6880 11679
rect 6828 11636 6880 11645
rect 7196 11704 7248 11756
rect 2504 11611 2556 11620
rect 2504 11577 2513 11611
rect 2513 11577 2547 11611
rect 2547 11577 2556 11611
rect 2504 11568 2556 11577
rect 4620 11568 4672 11620
rect 2044 11500 2096 11552
rect 2780 11500 2832 11552
rect 6000 11500 6052 11552
rect 7564 11500 7616 11552
rect 8484 11543 8536 11552
rect 8484 11509 8493 11543
rect 8493 11509 8527 11543
rect 8527 11509 8536 11543
rect 8484 11500 8536 11509
rect 12164 11772 12216 11824
rect 17408 11815 17460 11824
rect 17408 11781 17417 11815
rect 17417 11781 17451 11815
rect 17451 11781 17460 11815
rect 17408 11772 17460 11781
rect 9588 11704 9640 11756
rect 12808 11747 12860 11756
rect 12808 11713 12817 11747
rect 12817 11713 12851 11747
rect 12851 11713 12860 11747
rect 12808 11704 12860 11713
rect 11336 11679 11388 11688
rect 11336 11645 11345 11679
rect 11345 11645 11379 11679
rect 11379 11645 11388 11679
rect 11336 11636 11388 11645
rect 14648 11679 14700 11688
rect 12256 11568 12308 11620
rect 10048 11500 10100 11552
rect 11704 11500 11756 11552
rect 11980 11500 12032 11552
rect 12348 11500 12400 11552
rect 14648 11645 14657 11679
rect 14657 11645 14691 11679
rect 14691 11645 14700 11679
rect 14648 11636 14700 11645
rect 14924 11679 14976 11688
rect 14924 11645 14933 11679
rect 14933 11645 14967 11679
rect 14967 11645 14976 11679
rect 14924 11636 14976 11645
rect 15936 11679 15988 11688
rect 15936 11645 15945 11679
rect 15945 11645 15979 11679
rect 15979 11645 15988 11679
rect 15936 11636 15988 11645
rect 19432 11772 19484 11824
rect 23480 11772 23532 11824
rect 24216 11772 24268 11824
rect 15752 11568 15804 11620
rect 18144 11636 18196 11688
rect 18880 11704 18932 11756
rect 17408 11568 17460 11620
rect 20076 11568 20128 11620
rect 21732 11704 21784 11756
rect 23756 11747 23808 11756
rect 23756 11713 23765 11747
rect 23765 11713 23799 11747
rect 23799 11713 23808 11747
rect 23756 11704 23808 11713
rect 24032 11747 24084 11756
rect 24032 11713 24041 11747
rect 24041 11713 24075 11747
rect 24075 11713 24084 11747
rect 24032 11704 24084 11713
rect 13636 11500 13688 11552
rect 18328 11543 18380 11552
rect 18328 11509 18337 11543
rect 18337 11509 18371 11543
rect 18371 11509 18380 11543
rect 18328 11500 18380 11509
rect 19340 11543 19392 11552
rect 19340 11509 19349 11543
rect 19349 11509 19383 11543
rect 19383 11509 19392 11543
rect 19340 11500 19392 11509
rect 20812 11543 20864 11552
rect 20812 11509 20821 11543
rect 20821 11509 20855 11543
rect 20855 11509 20864 11543
rect 20812 11500 20864 11509
rect 21272 11543 21324 11552
rect 21272 11509 21281 11543
rect 21281 11509 21315 11543
rect 21315 11509 21324 11543
rect 21272 11500 21324 11509
rect 24860 11636 24912 11688
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 1860 11339 1912 11348
rect 1860 11305 1869 11339
rect 1869 11305 1903 11339
rect 1903 11305 1912 11339
rect 1860 11296 1912 11305
rect 2412 11296 2464 11348
rect 2044 11228 2096 11280
rect 1584 11092 1636 11144
rect 2504 11135 2556 11144
rect 2504 11101 2513 11135
rect 2513 11101 2547 11135
rect 2547 11101 2556 11135
rect 4160 11296 4212 11348
rect 4344 11296 4396 11348
rect 7196 11296 7248 11348
rect 10140 11296 10192 11348
rect 11980 11296 12032 11348
rect 12716 11296 12768 11348
rect 13912 11296 13964 11348
rect 14648 11296 14700 11348
rect 15936 11296 15988 11348
rect 17500 11339 17552 11348
rect 17500 11305 17509 11339
rect 17509 11305 17543 11339
rect 17543 11305 17552 11339
rect 17500 11296 17552 11305
rect 18144 11339 18196 11348
rect 18144 11305 18153 11339
rect 18153 11305 18187 11339
rect 18187 11305 18196 11339
rect 18144 11296 18196 11305
rect 18420 11339 18472 11348
rect 18420 11305 18429 11339
rect 18429 11305 18463 11339
rect 18463 11305 18472 11339
rect 18420 11296 18472 11305
rect 20720 11339 20772 11348
rect 20720 11305 20729 11339
rect 20729 11305 20763 11339
rect 20763 11305 20772 11339
rect 20720 11296 20772 11305
rect 20812 11296 20864 11348
rect 25228 11339 25280 11348
rect 4620 11228 4672 11280
rect 6736 11228 6788 11280
rect 8760 11271 8812 11280
rect 8760 11237 8769 11271
rect 8769 11237 8803 11271
rect 8803 11237 8812 11271
rect 8760 11228 8812 11237
rect 10048 11271 10100 11280
rect 10048 11237 10051 11271
rect 10051 11237 10085 11271
rect 10085 11237 10100 11271
rect 10048 11228 10100 11237
rect 12164 11228 12216 11280
rect 12256 11228 12308 11280
rect 6552 11160 6604 11212
rect 8208 11203 8260 11212
rect 2504 11092 2556 11101
rect 5540 10956 5592 11008
rect 6920 11092 6972 11144
rect 8208 11169 8217 11203
rect 8217 11169 8251 11203
rect 8251 11169 8260 11203
rect 8208 11160 8260 11169
rect 8576 11160 8628 11212
rect 11612 11203 11664 11212
rect 11612 11169 11621 11203
rect 11621 11169 11655 11203
rect 11655 11169 11664 11203
rect 11612 11160 11664 11169
rect 11980 11160 12032 11212
rect 13544 11160 13596 11212
rect 13820 11228 13872 11280
rect 16028 11228 16080 11280
rect 19340 11271 19392 11280
rect 19340 11237 19349 11271
rect 19349 11237 19383 11271
rect 19383 11237 19392 11271
rect 19340 11228 19392 11237
rect 21456 11228 21508 11280
rect 22928 11271 22980 11280
rect 22928 11237 22937 11271
rect 22937 11237 22971 11271
rect 22971 11237 22980 11271
rect 22928 11228 22980 11237
rect 23664 11271 23716 11280
rect 23664 11237 23673 11271
rect 23673 11237 23707 11271
rect 23707 11237 23716 11271
rect 23664 11228 23716 11237
rect 16856 11160 16908 11212
rect 17408 11203 17460 11212
rect 17408 11169 17417 11203
rect 17417 11169 17451 11203
rect 17451 11169 17460 11203
rect 17408 11160 17460 11169
rect 17592 11160 17644 11212
rect 19064 11203 19116 11212
rect 9680 11135 9732 11144
rect 7104 10956 7156 11008
rect 7472 10956 7524 11008
rect 9680 11101 9689 11135
rect 9689 11101 9723 11135
rect 9723 11101 9732 11135
rect 9680 11092 9732 11101
rect 12256 11092 12308 11144
rect 12532 11135 12584 11144
rect 12532 11101 12541 11135
rect 12541 11101 12575 11135
rect 12575 11101 12584 11135
rect 12532 11092 12584 11101
rect 12900 11092 12952 11144
rect 13912 11135 13964 11144
rect 13912 11101 13921 11135
rect 13921 11101 13955 11135
rect 13955 11101 13964 11135
rect 13912 11092 13964 11101
rect 16212 11135 16264 11144
rect 9956 11024 10008 11076
rect 9404 10956 9456 11008
rect 16212 11101 16221 11135
rect 16221 11101 16255 11135
rect 16255 11101 16264 11135
rect 16212 11092 16264 11101
rect 19064 11169 19073 11203
rect 19073 11169 19107 11203
rect 19107 11169 19116 11203
rect 19064 11160 19116 11169
rect 21640 11160 21692 11212
rect 22376 11160 22428 11212
rect 25228 11305 25237 11339
rect 25237 11305 25271 11339
rect 25271 11305 25280 11339
rect 25228 11296 25280 11305
rect 19340 11092 19392 11144
rect 20720 11092 20772 11144
rect 21180 11092 21232 11144
rect 16396 11024 16448 11076
rect 11152 10956 11204 11008
rect 11888 10956 11940 11008
rect 12808 10956 12860 11008
rect 15292 10956 15344 11008
rect 15844 10956 15896 11008
rect 25136 11160 25188 11212
rect 23572 11135 23624 11144
rect 23572 11101 23581 11135
rect 23581 11101 23615 11135
rect 23615 11101 23624 11135
rect 23572 11092 23624 11101
rect 23756 11092 23808 11144
rect 24032 11024 24084 11076
rect 19432 10956 19484 11008
rect 20076 10956 20128 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 4620 10795 4672 10804
rect 4620 10761 4629 10795
rect 4629 10761 4663 10795
rect 4663 10761 4672 10795
rect 4620 10752 4672 10761
rect 6736 10752 6788 10804
rect 7104 10795 7156 10804
rect 7104 10761 7113 10795
rect 7113 10761 7147 10795
rect 7147 10761 7156 10795
rect 7104 10752 7156 10761
rect 8300 10752 8352 10804
rect 2044 10684 2096 10736
rect 2688 10727 2740 10736
rect 2688 10693 2697 10727
rect 2697 10693 2731 10727
rect 2731 10693 2740 10727
rect 2688 10684 2740 10693
rect 8024 10727 8076 10736
rect 8024 10693 8033 10727
rect 8033 10693 8067 10727
rect 8067 10693 8076 10727
rect 8024 10684 8076 10693
rect 8576 10752 8628 10804
rect 12900 10752 12952 10804
rect 13820 10795 13872 10804
rect 13820 10761 13829 10795
rect 13829 10761 13863 10795
rect 13863 10761 13872 10795
rect 13820 10752 13872 10761
rect 15660 10795 15712 10804
rect 15660 10761 15669 10795
rect 15669 10761 15703 10795
rect 15703 10761 15712 10795
rect 15660 10752 15712 10761
rect 16948 10752 17000 10804
rect 11980 10684 12032 10736
rect 2136 10523 2188 10532
rect 2136 10489 2145 10523
rect 2145 10489 2179 10523
rect 2179 10489 2188 10523
rect 2136 10480 2188 10489
rect 3792 10616 3844 10668
rect 4160 10659 4212 10668
rect 4160 10625 4169 10659
rect 4169 10625 4203 10659
rect 4203 10625 4212 10659
rect 4160 10616 4212 10625
rect 5540 10616 5592 10668
rect 9588 10659 9640 10668
rect 9588 10625 9597 10659
rect 9597 10625 9631 10659
rect 9631 10625 9640 10659
rect 9588 10616 9640 10625
rect 12808 10659 12860 10668
rect 12808 10625 12814 10659
rect 12814 10625 12848 10659
rect 12848 10625 12860 10659
rect 12808 10616 12860 10625
rect 15844 10659 15896 10668
rect 15844 10625 15853 10659
rect 15853 10625 15887 10659
rect 15887 10625 15896 10659
rect 15844 10616 15896 10625
rect 16212 10659 16264 10668
rect 16212 10625 16221 10659
rect 16221 10625 16255 10659
rect 16255 10625 16264 10659
rect 16212 10616 16264 10625
rect 3792 10523 3844 10532
rect 3792 10489 3801 10523
rect 3801 10489 3835 10523
rect 3835 10489 3844 10523
rect 3792 10480 3844 10489
rect 3424 10455 3476 10464
rect 3424 10421 3433 10455
rect 3433 10421 3467 10455
rect 3467 10421 3476 10455
rect 3424 10412 3476 10421
rect 4804 10412 4856 10464
rect 5264 10548 5316 10600
rect 6552 10548 6604 10600
rect 9220 10591 9272 10600
rect 9220 10557 9229 10591
rect 9229 10557 9263 10591
rect 9263 10557 9272 10591
rect 9220 10548 9272 10557
rect 9404 10591 9456 10600
rect 9404 10557 9413 10591
rect 9413 10557 9447 10591
rect 9447 10557 9456 10591
rect 9404 10548 9456 10557
rect 10784 10591 10836 10600
rect 10784 10557 10793 10591
rect 10793 10557 10827 10591
rect 10827 10557 10836 10591
rect 10784 10548 10836 10557
rect 11152 10548 11204 10600
rect 7472 10523 7524 10532
rect 7472 10489 7481 10523
rect 7481 10489 7515 10523
rect 7515 10489 7524 10523
rect 7472 10480 7524 10489
rect 7564 10523 7616 10532
rect 7564 10489 7573 10523
rect 7573 10489 7607 10523
rect 7607 10489 7616 10523
rect 7564 10480 7616 10489
rect 9772 10480 9824 10532
rect 10048 10455 10100 10464
rect 10048 10421 10057 10455
rect 10057 10421 10091 10455
rect 10091 10421 10100 10455
rect 10048 10412 10100 10421
rect 12164 10480 12216 10532
rect 13820 10548 13872 10600
rect 14280 10591 14332 10600
rect 14280 10557 14289 10591
rect 14289 10557 14323 10591
rect 14323 10557 14332 10591
rect 14280 10548 14332 10557
rect 19340 10752 19392 10804
rect 20720 10752 20772 10804
rect 22376 10795 22428 10804
rect 22376 10761 22385 10795
rect 22385 10761 22419 10795
rect 22419 10761 22428 10795
rect 22376 10752 22428 10761
rect 23388 10752 23440 10804
rect 23480 10795 23532 10804
rect 23480 10761 23489 10795
rect 23489 10761 23523 10795
rect 23523 10761 23532 10795
rect 23480 10752 23532 10761
rect 23848 10752 23900 10804
rect 25412 10795 25464 10804
rect 25412 10761 25421 10795
rect 25421 10761 25455 10795
rect 25455 10761 25464 10795
rect 25412 10752 25464 10761
rect 20444 10684 20496 10736
rect 21456 10727 21508 10736
rect 21456 10693 21465 10727
rect 21465 10693 21499 10727
rect 21499 10693 21508 10727
rect 21456 10684 21508 10693
rect 19248 10659 19300 10668
rect 19248 10625 19257 10659
rect 19257 10625 19291 10659
rect 19291 10625 19300 10659
rect 19248 10616 19300 10625
rect 21180 10659 21232 10668
rect 21180 10625 21189 10659
rect 21189 10625 21223 10659
rect 21223 10625 21232 10659
rect 21180 10616 21232 10625
rect 23756 10616 23808 10668
rect 11980 10412 12032 10464
rect 18236 10548 18288 10600
rect 14832 10480 14884 10532
rect 16304 10480 16356 10532
rect 13636 10412 13688 10464
rect 14740 10412 14792 10464
rect 15292 10412 15344 10464
rect 19064 10548 19116 10600
rect 25228 10591 25280 10600
rect 20260 10523 20312 10532
rect 20260 10489 20269 10523
rect 20269 10489 20303 10523
rect 20303 10489 20312 10523
rect 20260 10480 20312 10489
rect 25228 10557 25237 10591
rect 25237 10557 25271 10591
rect 25271 10557 25280 10591
rect 25228 10548 25280 10557
rect 16856 10455 16908 10464
rect 16856 10421 16865 10455
rect 16865 10421 16899 10455
rect 16899 10421 16908 10455
rect 16856 10412 16908 10421
rect 16948 10412 17000 10464
rect 17408 10412 17460 10464
rect 18604 10412 18656 10464
rect 23020 10455 23072 10464
rect 23020 10421 23029 10455
rect 23029 10421 23063 10455
rect 23063 10421 23072 10455
rect 23020 10412 23072 10421
rect 23848 10523 23900 10532
rect 23848 10489 23857 10523
rect 23857 10489 23891 10523
rect 23891 10489 23900 10523
rect 23848 10480 23900 10489
rect 24216 10412 24268 10464
rect 25044 10455 25096 10464
rect 25044 10421 25053 10455
rect 25053 10421 25087 10455
rect 25087 10421 25096 10455
rect 25044 10412 25096 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 3792 10208 3844 10260
rect 5264 10251 5316 10260
rect 5264 10217 5273 10251
rect 5273 10217 5307 10251
rect 5307 10217 5316 10251
rect 5264 10208 5316 10217
rect 7564 10208 7616 10260
rect 9220 10208 9272 10260
rect 9588 10208 9640 10260
rect 11888 10251 11940 10260
rect 11888 10217 11897 10251
rect 11897 10217 11931 10251
rect 11931 10217 11940 10251
rect 11888 10208 11940 10217
rect 12900 10208 12952 10260
rect 13728 10208 13780 10260
rect 14096 10208 14148 10260
rect 16304 10251 16356 10260
rect 16304 10217 16313 10251
rect 16313 10217 16347 10251
rect 16347 10217 16356 10251
rect 16304 10208 16356 10217
rect 18604 10251 18656 10260
rect 18604 10217 18613 10251
rect 18613 10217 18647 10251
rect 18647 10217 18656 10251
rect 18604 10208 18656 10217
rect 2412 10140 2464 10192
rect 4252 10183 4304 10192
rect 4252 10149 4261 10183
rect 4261 10149 4295 10183
rect 4295 10149 4304 10183
rect 4252 10140 4304 10149
rect 6828 10140 6880 10192
rect 7196 10140 7248 10192
rect 10140 10140 10192 10192
rect 1400 10072 1452 10124
rect 6276 10115 6328 10124
rect 6276 10081 6285 10115
rect 6285 10081 6319 10115
rect 6319 10081 6328 10115
rect 6276 10072 6328 10081
rect 6552 10115 6604 10124
rect 6552 10081 6561 10115
rect 6561 10081 6595 10115
rect 6595 10081 6604 10115
rect 6552 10072 6604 10081
rect 22008 10208 22060 10260
rect 23572 10208 23624 10260
rect 24768 10251 24820 10260
rect 24768 10217 24777 10251
rect 24777 10217 24811 10251
rect 24811 10217 24820 10251
rect 24768 10208 24820 10217
rect 25136 10251 25188 10260
rect 25136 10217 25145 10251
rect 25145 10217 25179 10251
rect 25179 10217 25188 10251
rect 25136 10208 25188 10217
rect 12440 10115 12492 10124
rect 12440 10081 12449 10115
rect 12449 10081 12483 10115
rect 12483 10081 12492 10115
rect 12440 10072 12492 10081
rect 13452 10072 13504 10124
rect 14004 10072 14056 10124
rect 15752 10183 15804 10192
rect 15752 10149 15755 10183
rect 15755 10149 15789 10183
rect 15789 10149 15804 10183
rect 15752 10140 15804 10149
rect 17684 10183 17736 10192
rect 17684 10149 17693 10183
rect 17693 10149 17727 10183
rect 17727 10149 17736 10183
rect 17684 10140 17736 10149
rect 19432 10183 19484 10192
rect 19432 10149 19435 10183
rect 19435 10149 19469 10183
rect 19469 10149 19484 10183
rect 19432 10140 19484 10149
rect 21088 10183 21140 10192
rect 21088 10149 21097 10183
rect 21097 10149 21131 10183
rect 21131 10149 21140 10183
rect 21088 10140 21140 10149
rect 25044 10140 25096 10192
rect 14280 10072 14332 10124
rect 23572 10115 23624 10124
rect 23572 10081 23616 10115
rect 23616 10081 23624 10115
rect 23572 10072 23624 10081
rect 24032 10072 24084 10124
rect 24308 10072 24360 10124
rect 2044 10047 2096 10056
rect 2044 10013 2053 10047
rect 2053 10013 2087 10047
rect 2087 10013 2096 10047
rect 2044 10004 2096 10013
rect 2504 10047 2556 10056
rect 2504 10013 2513 10047
rect 2513 10013 2547 10047
rect 2547 10013 2556 10047
rect 2504 10004 2556 10013
rect 4160 10047 4212 10056
rect 4160 10013 4169 10047
rect 4169 10013 4203 10047
rect 4203 10013 4212 10047
rect 4160 10004 4212 10013
rect 4620 10047 4672 10056
rect 4620 10013 4629 10047
rect 4629 10013 4663 10047
rect 4663 10013 4672 10047
rect 4620 10004 4672 10013
rect 8024 10004 8076 10056
rect 9772 10047 9824 10056
rect 9772 10013 9781 10047
rect 9781 10013 9815 10047
rect 9815 10013 9824 10047
rect 9772 10004 9824 10013
rect 2136 9936 2188 9988
rect 1400 9868 1452 9920
rect 2596 9868 2648 9920
rect 4528 9936 4580 9988
rect 5080 9936 5132 9988
rect 9220 9936 9272 9988
rect 13544 10004 13596 10056
rect 15292 10004 15344 10056
rect 16212 10004 16264 10056
rect 17960 10004 18012 10056
rect 19064 10047 19116 10056
rect 19064 10013 19073 10047
rect 19073 10013 19107 10047
rect 19107 10013 19116 10047
rect 19064 10004 19116 10013
rect 21180 10004 21232 10056
rect 11980 9936 12032 9988
rect 14004 9936 14056 9988
rect 21640 9936 21692 9988
rect 23664 9936 23716 9988
rect 10968 9868 11020 9920
rect 12164 9868 12216 9920
rect 16580 9868 16632 9920
rect 20444 9911 20496 9920
rect 20444 9877 20453 9911
rect 20453 9877 20487 9911
rect 20487 9877 20496 9911
rect 20444 9868 20496 9877
rect 21364 9868 21416 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 2412 9707 2464 9716
rect 2412 9673 2421 9707
rect 2421 9673 2455 9707
rect 2455 9673 2464 9707
rect 2412 9664 2464 9673
rect 4160 9664 4212 9716
rect 5264 9664 5316 9716
rect 6092 9707 6144 9716
rect 1860 9596 1912 9648
rect 6092 9673 6101 9707
rect 6101 9673 6135 9707
rect 6135 9673 6144 9707
rect 6092 9664 6144 9673
rect 6276 9664 6328 9716
rect 6552 9664 6604 9716
rect 10140 9707 10192 9716
rect 10140 9673 10149 9707
rect 10149 9673 10183 9707
rect 10183 9673 10192 9707
rect 10140 9664 10192 9673
rect 10784 9664 10836 9716
rect 11888 9639 11940 9648
rect 11888 9605 11897 9639
rect 11897 9605 11931 9639
rect 11931 9605 11940 9639
rect 11888 9596 11940 9605
rect 13636 9664 13688 9716
rect 15292 9664 15344 9716
rect 2688 9528 2740 9580
rect 3148 9528 3200 9580
rect 4620 9528 4672 9580
rect 4896 9571 4948 9580
rect 4896 9537 4905 9571
rect 4905 9537 4939 9571
rect 4939 9537 4948 9571
rect 4896 9528 4948 9537
rect 9220 9571 9272 9580
rect 9220 9537 9229 9571
rect 9229 9537 9263 9571
rect 9263 9537 9272 9571
rect 9220 9528 9272 9537
rect 9680 9571 9732 9580
rect 9680 9537 9689 9571
rect 9689 9537 9723 9571
rect 9723 9537 9732 9571
rect 9680 9528 9732 9537
rect 2596 9460 2648 9512
rect 10784 9503 10836 9512
rect 10784 9469 10793 9503
rect 10793 9469 10827 9503
rect 10827 9469 10836 9503
rect 10784 9460 10836 9469
rect 10968 9460 11020 9512
rect 11244 9503 11296 9512
rect 11244 9469 11253 9503
rect 11253 9469 11287 9503
rect 11287 9469 11296 9503
rect 11244 9460 11296 9469
rect 13084 9596 13136 9648
rect 13452 9639 13504 9648
rect 13452 9605 13461 9639
rect 13461 9605 13495 9639
rect 13495 9605 13504 9639
rect 13452 9596 13504 9605
rect 13820 9639 13872 9648
rect 13820 9605 13829 9639
rect 13829 9605 13863 9639
rect 13863 9605 13872 9639
rect 13820 9596 13872 9605
rect 21088 9664 21140 9716
rect 17960 9596 18012 9648
rect 21180 9596 21232 9648
rect 24032 9664 24084 9716
rect 12624 9528 12676 9580
rect 12716 9503 12768 9512
rect 12716 9469 12725 9503
rect 12725 9469 12759 9503
rect 12759 9469 12768 9503
rect 12716 9460 12768 9469
rect 21364 9571 21416 9580
rect 21364 9537 21373 9571
rect 21373 9537 21407 9571
rect 21407 9537 21416 9571
rect 21364 9528 21416 9537
rect 21640 9571 21692 9580
rect 21640 9537 21649 9571
rect 21649 9537 21683 9571
rect 21683 9537 21692 9571
rect 21640 9528 21692 9537
rect 15108 9503 15160 9512
rect 15108 9469 15117 9503
rect 15117 9469 15151 9503
rect 15151 9469 15160 9503
rect 15108 9460 15160 9469
rect 16764 9460 16816 9512
rect 19524 9503 19576 9512
rect 19524 9469 19533 9503
rect 19533 9469 19567 9503
rect 19567 9469 19576 9503
rect 19524 9460 19576 9469
rect 2136 9435 2188 9444
rect 2136 9401 2145 9435
rect 2145 9401 2179 9435
rect 2179 9401 2188 9435
rect 2136 9392 2188 9401
rect 3056 9435 3108 9444
rect 3056 9401 3065 9435
rect 3065 9401 3099 9435
rect 3099 9401 3108 9435
rect 3056 9392 3108 9401
rect 1676 9324 1728 9376
rect 3240 9392 3292 9444
rect 3884 9392 3936 9444
rect 4712 9435 4764 9444
rect 4712 9401 4721 9435
rect 4721 9401 4755 9435
rect 4755 9401 4764 9435
rect 4712 9392 4764 9401
rect 7288 9392 7340 9444
rect 4068 9367 4120 9376
rect 4068 9333 4077 9367
rect 4077 9333 4111 9367
rect 4111 9333 4120 9367
rect 4068 9324 4120 9333
rect 4252 9324 4304 9376
rect 7012 9367 7064 9376
rect 7012 9333 7021 9367
rect 7021 9333 7055 9367
rect 7055 9333 7064 9367
rect 7012 9324 7064 9333
rect 7748 9435 7800 9444
rect 7748 9401 7757 9435
rect 7757 9401 7791 9435
rect 7791 9401 7800 9435
rect 7748 9392 7800 9401
rect 9312 9435 9364 9444
rect 9312 9401 9321 9435
rect 9321 9401 9355 9435
rect 9355 9401 9364 9435
rect 9312 9392 9364 9401
rect 10048 9392 10100 9444
rect 15752 9392 15804 9444
rect 16396 9392 16448 9444
rect 19432 9392 19484 9444
rect 8576 9367 8628 9376
rect 8576 9333 8585 9367
rect 8585 9333 8619 9367
rect 8619 9333 8628 9367
rect 8576 9324 8628 9333
rect 10784 9367 10836 9376
rect 10784 9333 10793 9367
rect 10793 9333 10827 9367
rect 10827 9333 10836 9367
rect 10784 9324 10836 9333
rect 14188 9367 14240 9376
rect 14188 9333 14197 9367
rect 14197 9333 14231 9367
rect 14231 9333 14240 9367
rect 14188 9324 14240 9333
rect 16120 9324 16172 9376
rect 17684 9324 17736 9376
rect 17960 9324 18012 9376
rect 18512 9367 18564 9376
rect 18512 9333 18521 9367
rect 18521 9333 18555 9367
rect 18555 9333 18564 9367
rect 18512 9324 18564 9333
rect 20812 9367 20864 9376
rect 20812 9333 20821 9367
rect 20821 9333 20855 9367
rect 20855 9333 20864 9367
rect 20812 9324 20864 9333
rect 24768 9639 24820 9648
rect 24768 9605 24777 9639
rect 24777 9605 24811 9639
rect 24811 9605 24820 9639
rect 24768 9596 24820 9605
rect 25320 9596 25372 9648
rect 23572 9324 23624 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 1860 9163 1912 9172
rect 1860 9129 1869 9163
rect 1869 9129 1903 9163
rect 1903 9129 1912 9163
rect 1860 9120 1912 9129
rect 3884 9163 3936 9172
rect 3884 9129 3893 9163
rect 3893 9129 3927 9163
rect 3927 9129 3936 9163
rect 3884 9120 3936 9129
rect 7012 9120 7064 9172
rect 7748 9163 7800 9172
rect 7748 9129 7757 9163
rect 7757 9129 7791 9163
rect 7791 9129 7800 9163
rect 7748 9120 7800 9129
rect 8484 9120 8536 9172
rect 9312 9120 9364 9172
rect 11980 9120 12032 9172
rect 12716 9120 12768 9172
rect 16028 9120 16080 9172
rect 17960 9120 18012 9172
rect 19064 9163 19116 9172
rect 19064 9129 19073 9163
rect 19073 9129 19107 9163
rect 19107 9129 19116 9163
rect 19064 9120 19116 9129
rect 20904 9120 20956 9172
rect 2780 9052 2832 9104
rect 3148 9095 3200 9104
rect 3148 9061 3157 9095
rect 3157 9061 3191 9095
rect 3191 9061 3200 9095
rect 3148 9052 3200 9061
rect 5448 9052 5500 9104
rect 7196 9095 7248 9104
rect 7196 9061 7199 9095
rect 7199 9061 7233 9095
rect 7233 9061 7248 9095
rect 7196 9052 7248 9061
rect 10048 9095 10100 9104
rect 10048 9061 10051 9095
rect 10051 9061 10085 9095
rect 10085 9061 10100 9095
rect 10048 9052 10100 9061
rect 15108 9052 15160 9104
rect 15752 9052 15804 9104
rect 17592 9052 17644 9104
rect 19432 9052 19484 9104
rect 20996 9095 21048 9104
rect 20996 9061 21005 9095
rect 21005 9061 21039 9095
rect 21039 9061 21048 9095
rect 20996 9052 21048 9061
rect 21272 9120 21324 9172
rect 22100 9120 22152 9172
rect 22652 9095 22704 9104
rect 22652 9061 22661 9095
rect 22661 9061 22695 9095
rect 22695 9061 22704 9095
rect 22652 9052 22704 9061
rect 2320 8984 2372 9036
rect 4712 8984 4764 9036
rect 8484 8984 8536 9036
rect 2136 8916 2188 8968
rect 2688 8916 2740 8968
rect 4436 8916 4488 8968
rect 5540 8916 5592 8968
rect 7932 8916 7984 8968
rect 10784 8916 10836 8968
rect 12440 8916 12492 8968
rect 13360 8984 13412 9036
rect 14740 8984 14792 9036
rect 14832 8984 14884 9036
rect 16580 8984 16632 9036
rect 19340 9027 19392 9036
rect 19340 8993 19349 9027
rect 19349 8993 19383 9027
rect 19383 8993 19392 9027
rect 19340 8984 19392 8993
rect 19708 9027 19760 9036
rect 19708 8993 19717 9027
rect 19717 8993 19751 9027
rect 19751 8993 19760 9027
rect 19708 8984 19760 8993
rect 25504 8984 25556 9036
rect 12624 8916 12676 8968
rect 13452 8916 13504 8968
rect 17132 8916 17184 8968
rect 21180 8916 21232 8968
rect 22560 8959 22612 8968
rect 22560 8925 22569 8959
rect 22569 8925 22603 8959
rect 22603 8925 22612 8959
rect 22560 8916 22612 8925
rect 11980 8848 12032 8900
rect 19524 8848 19576 8900
rect 21364 8848 21416 8900
rect 2044 8780 2096 8832
rect 2228 8780 2280 8832
rect 3148 8780 3200 8832
rect 8024 8823 8076 8832
rect 8024 8789 8033 8823
rect 8033 8789 8067 8823
rect 8067 8789 8076 8823
rect 8024 8780 8076 8789
rect 9128 8823 9180 8832
rect 9128 8789 9137 8823
rect 9137 8789 9171 8823
rect 9171 8789 9180 8823
rect 9128 8780 9180 8789
rect 9588 8780 9640 8832
rect 11888 8780 11940 8832
rect 13084 8780 13136 8832
rect 14740 8823 14792 8832
rect 14740 8789 14749 8823
rect 14749 8789 14783 8823
rect 14783 8789 14792 8823
rect 14740 8780 14792 8789
rect 24768 8823 24820 8832
rect 24768 8789 24777 8823
rect 24777 8789 24811 8823
rect 24811 8789 24820 8823
rect 24768 8780 24820 8789
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 1584 8619 1636 8628
rect 1584 8585 1593 8619
rect 1593 8585 1627 8619
rect 1627 8585 1636 8619
rect 1584 8576 1636 8585
rect 2228 8576 2280 8628
rect 2780 8576 2832 8628
rect 7288 8576 7340 8628
rect 8484 8576 8536 8628
rect 10048 8576 10100 8628
rect 10784 8576 10836 8628
rect 9956 8508 10008 8560
rect 1308 8440 1360 8492
rect 1584 8440 1636 8492
rect 2780 8483 2832 8492
rect 2780 8449 2789 8483
rect 2789 8449 2823 8483
rect 2823 8449 2832 8483
rect 2780 8440 2832 8449
rect 3148 8440 3200 8492
rect 3884 8440 3936 8492
rect 12072 8576 12124 8628
rect 12624 8576 12676 8628
rect 13360 8576 13412 8628
rect 15752 8576 15804 8628
rect 16580 8619 16632 8628
rect 16580 8585 16589 8619
rect 16589 8585 16623 8619
rect 16623 8585 16632 8619
rect 16580 8576 16632 8585
rect 17592 8619 17644 8628
rect 17592 8585 17601 8619
rect 17601 8585 17635 8619
rect 17635 8585 17644 8619
rect 17592 8576 17644 8585
rect 19340 8576 19392 8628
rect 20628 8576 20680 8628
rect 20996 8619 21048 8628
rect 20996 8585 21005 8619
rect 21005 8585 21039 8619
rect 21039 8585 21048 8619
rect 20996 8576 21048 8585
rect 22100 8619 22152 8628
rect 22100 8585 22109 8619
rect 22109 8585 22143 8619
rect 22143 8585 22152 8619
rect 22100 8576 22152 8585
rect 22652 8576 22704 8628
rect 25504 8619 25556 8628
rect 25504 8585 25513 8619
rect 25513 8585 25547 8619
rect 25547 8585 25556 8619
rect 25504 8576 25556 8585
rect 11796 8508 11848 8560
rect 16212 8551 16264 8560
rect 16212 8517 16221 8551
rect 16221 8517 16255 8551
rect 16255 8517 16264 8551
rect 16212 8508 16264 8517
rect 12440 8483 12492 8492
rect 12440 8449 12449 8483
rect 12449 8449 12483 8483
rect 12483 8449 12492 8483
rect 12440 8440 12492 8449
rect 1952 8372 2004 8424
rect 4988 8372 5040 8424
rect 5540 8372 5592 8424
rect 6828 8415 6880 8424
rect 6828 8381 6837 8415
rect 6837 8381 6871 8415
rect 6871 8381 6880 8415
rect 6828 8372 6880 8381
rect 9128 8372 9180 8424
rect 9588 8372 9640 8424
rect 10140 8372 10192 8424
rect 11336 8372 11388 8424
rect 13084 8415 13136 8424
rect 13084 8381 13093 8415
rect 13093 8381 13127 8415
rect 13127 8381 13136 8415
rect 13084 8372 13136 8381
rect 14648 8440 14700 8492
rect 15292 8440 15344 8492
rect 16396 8440 16448 8492
rect 18236 8415 18288 8424
rect 18236 8381 18245 8415
rect 18245 8381 18279 8415
rect 18279 8381 18288 8415
rect 18236 8372 18288 8381
rect 18696 8372 18748 8424
rect 19708 8508 19760 8560
rect 20536 8551 20588 8560
rect 20536 8517 20545 8551
rect 20545 8517 20579 8551
rect 20579 8517 20588 8551
rect 20536 8508 20588 8517
rect 19524 8440 19576 8492
rect 21364 8440 21416 8492
rect 22560 8440 22612 8492
rect 2228 8279 2280 8288
rect 2228 8245 2237 8279
rect 2237 8245 2271 8279
rect 2271 8245 2280 8279
rect 2228 8236 2280 8245
rect 4068 8304 4120 8356
rect 5448 8304 5500 8356
rect 7196 8347 7248 8356
rect 7196 8313 7199 8347
rect 7199 8313 7233 8347
rect 7233 8313 7248 8347
rect 7196 8304 7248 8313
rect 9220 8304 9272 8356
rect 10048 8304 10100 8356
rect 14740 8304 14792 8356
rect 16120 8304 16172 8356
rect 21180 8347 21232 8356
rect 21180 8313 21189 8347
rect 21189 8313 21223 8347
rect 21223 8313 21232 8347
rect 21180 8304 21232 8313
rect 21272 8347 21324 8356
rect 21272 8313 21281 8347
rect 21281 8313 21315 8347
rect 21315 8313 21324 8347
rect 21272 8304 21324 8313
rect 24768 8304 24820 8356
rect 7932 8236 7984 8288
rect 17132 8279 17184 8288
rect 17132 8245 17141 8279
rect 17141 8245 17175 8279
rect 17175 8245 17184 8279
rect 17132 8236 17184 8245
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 1676 8032 1728 8084
rect 1952 8075 2004 8084
rect 1952 8041 1961 8075
rect 1961 8041 1995 8075
rect 1995 8041 2004 8075
rect 1952 8032 2004 8041
rect 2320 8075 2372 8084
rect 2320 8041 2329 8075
rect 2329 8041 2363 8075
rect 2363 8041 2372 8075
rect 2320 8032 2372 8041
rect 2780 8032 2832 8084
rect 3700 8032 3752 8084
rect 5632 8075 5684 8084
rect 5632 8041 5641 8075
rect 5641 8041 5675 8075
rect 5675 8041 5684 8075
rect 5632 8032 5684 8041
rect 2228 7964 2280 8016
rect 2872 7964 2924 8016
rect 3148 8007 3200 8016
rect 3148 7973 3157 8007
rect 3157 7973 3191 8007
rect 3191 7973 3200 8007
rect 3148 7964 3200 7973
rect 4436 7964 4488 8016
rect 5540 7964 5592 8016
rect 6736 8032 6788 8084
rect 7472 8032 7524 8084
rect 9220 8032 9272 8084
rect 9680 8032 9732 8084
rect 12164 8075 12216 8084
rect 12164 8041 12173 8075
rect 12173 8041 12207 8075
rect 12207 8041 12216 8075
rect 12164 8032 12216 8041
rect 14740 8032 14792 8084
rect 15568 8032 15620 8084
rect 16120 8032 16172 8084
rect 16396 8032 16448 8084
rect 17132 8075 17184 8084
rect 17132 8041 17141 8075
rect 17141 8041 17175 8075
rect 17175 8041 17184 8075
rect 17132 8032 17184 8041
rect 18236 8075 18288 8084
rect 18236 8041 18245 8075
rect 18245 8041 18279 8075
rect 18279 8041 18288 8075
rect 18236 8032 18288 8041
rect 18696 8075 18748 8084
rect 18696 8041 18705 8075
rect 18705 8041 18739 8075
rect 18739 8041 18748 8075
rect 18696 8032 18748 8041
rect 20444 8032 20496 8084
rect 21180 8032 21232 8084
rect 6828 7964 6880 8016
rect 10876 7964 10928 8016
rect 1400 7939 1452 7948
rect 1400 7905 1444 7939
rect 1444 7905 1452 7939
rect 6276 7939 6328 7948
rect 1400 7896 1452 7905
rect 6276 7905 6285 7939
rect 6285 7905 6319 7939
rect 6319 7905 6328 7939
rect 6276 7896 6328 7905
rect 6736 7939 6788 7948
rect 6736 7905 6745 7939
rect 6745 7905 6779 7939
rect 6779 7905 6788 7939
rect 6736 7896 6788 7905
rect 8116 7896 8168 7948
rect 9956 7939 10008 7948
rect 9956 7905 9965 7939
rect 9965 7905 9999 7939
rect 9999 7905 10008 7939
rect 9956 7896 10008 7905
rect 10048 7896 10100 7948
rect 10968 7896 11020 7948
rect 11888 7939 11940 7948
rect 11888 7905 11897 7939
rect 11897 7905 11931 7939
rect 11931 7905 11940 7939
rect 11888 7896 11940 7905
rect 11980 7896 12032 7948
rect 13544 7896 13596 7948
rect 14372 7964 14424 8016
rect 14556 7896 14608 7948
rect 15384 7939 15436 7948
rect 15384 7905 15428 7939
rect 15428 7905 15436 7939
rect 17040 7939 17092 7948
rect 15384 7896 15436 7905
rect 17040 7905 17049 7939
rect 17049 7905 17083 7939
rect 17083 7905 17092 7939
rect 17040 7896 17092 7905
rect 17500 7896 17552 7948
rect 21456 8032 21508 8084
rect 23480 8032 23532 8084
rect 21364 7964 21416 8016
rect 24492 7964 24544 8016
rect 19892 7939 19944 7948
rect 19892 7905 19910 7939
rect 19910 7905 19944 7939
rect 19892 7896 19944 7905
rect 20352 7896 20404 7948
rect 23756 7896 23808 7948
rect 24676 7939 24728 7948
rect 24676 7905 24694 7939
rect 24694 7905 24728 7939
rect 24676 7896 24728 7905
rect 4712 7871 4764 7880
rect 4712 7837 4721 7871
rect 4721 7837 4755 7871
rect 4755 7837 4764 7871
rect 4712 7828 4764 7837
rect 4896 7828 4948 7880
rect 21548 7828 21600 7880
rect 2412 7692 2464 7744
rect 2780 7692 2832 7744
rect 3516 7735 3568 7744
rect 3516 7701 3525 7735
rect 3525 7701 3559 7735
rect 3559 7701 3568 7735
rect 3516 7692 3568 7701
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 1400 7488 1452 7540
rect 2872 7488 2924 7540
rect 4436 7531 4488 7540
rect 4436 7497 4445 7531
rect 4445 7497 4479 7531
rect 4479 7497 4488 7531
rect 4436 7488 4488 7497
rect 4804 7531 4856 7540
rect 4804 7497 4813 7531
rect 4813 7497 4847 7531
rect 4847 7497 4856 7531
rect 4804 7488 4856 7497
rect 6092 7488 6144 7540
rect 1492 7420 1544 7472
rect 2044 7463 2096 7472
rect 2044 7429 2053 7463
rect 2053 7429 2087 7463
rect 2087 7429 2096 7463
rect 2044 7420 2096 7429
rect 6276 7463 6328 7472
rect 6276 7429 6285 7463
rect 6285 7429 6319 7463
rect 6319 7429 6328 7463
rect 6276 7420 6328 7429
rect 3884 7395 3936 7404
rect 3884 7361 3893 7395
rect 3893 7361 3927 7395
rect 3927 7361 3936 7395
rect 3884 7352 3936 7361
rect 4804 7284 4856 7336
rect 8116 7488 8168 7540
rect 8576 7488 8628 7540
rect 9956 7488 10008 7540
rect 10324 7488 10376 7540
rect 11060 7488 11112 7540
rect 11980 7531 12032 7540
rect 11980 7497 11989 7531
rect 11989 7497 12023 7531
rect 12023 7497 12032 7531
rect 11980 7488 12032 7497
rect 12624 7531 12676 7540
rect 12624 7497 12633 7531
rect 12633 7497 12667 7531
rect 12667 7497 12676 7531
rect 12624 7488 12676 7497
rect 13544 7531 13596 7540
rect 13544 7497 13553 7531
rect 13553 7497 13587 7531
rect 13587 7497 13596 7531
rect 13544 7488 13596 7497
rect 14740 7488 14792 7540
rect 17040 7531 17092 7540
rect 17040 7497 17049 7531
rect 17049 7497 17083 7531
rect 17083 7497 17092 7531
rect 17040 7488 17092 7497
rect 17500 7531 17552 7540
rect 17500 7497 17509 7531
rect 17509 7497 17543 7531
rect 17543 7497 17552 7531
rect 17500 7488 17552 7497
rect 19892 7531 19944 7540
rect 19892 7497 19901 7531
rect 19901 7497 19935 7531
rect 19935 7497 19944 7531
rect 19892 7488 19944 7497
rect 21456 7488 21508 7540
rect 23756 7488 23808 7540
rect 24676 7531 24728 7540
rect 24676 7497 24685 7531
rect 24685 7497 24719 7531
rect 24719 7497 24728 7531
rect 24676 7488 24728 7497
rect 6736 7420 6788 7472
rect 10048 7420 10100 7472
rect 7932 7352 7984 7404
rect 2964 7216 3016 7268
rect 3608 7216 3660 7268
rect 8392 7327 8444 7336
rect 8392 7293 8436 7327
rect 8436 7293 8444 7327
rect 8392 7284 8444 7293
rect 9864 7284 9916 7336
rect 12348 7420 12400 7472
rect 14556 7420 14608 7472
rect 24124 7352 24176 7404
rect 24676 7352 24728 7404
rect 12532 7284 12584 7336
rect 13912 7284 13964 7336
rect 15384 7327 15436 7336
rect 15384 7293 15393 7327
rect 15393 7293 15427 7327
rect 15427 7293 15436 7327
rect 15384 7284 15436 7293
rect 6736 7216 6788 7268
rect 4988 7191 5040 7200
rect 4988 7157 4997 7191
rect 4997 7157 5031 7191
rect 5031 7157 5040 7191
rect 4988 7148 5040 7157
rect 21548 7191 21600 7200
rect 21548 7157 21557 7191
rect 21557 7157 21591 7191
rect 21591 7157 21600 7191
rect 21548 7148 21600 7157
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 2964 6987 3016 6996
rect 2964 6953 2973 6987
rect 2973 6953 3007 6987
rect 3007 6953 3016 6987
rect 2964 6944 3016 6953
rect 3516 6944 3568 6996
rect 4712 6944 4764 6996
rect 4804 6944 4856 6996
rect 6736 6944 6788 6996
rect 11888 6987 11940 6996
rect 11888 6953 11897 6987
rect 11897 6953 11931 6987
rect 11931 6953 11940 6987
rect 11888 6944 11940 6953
rect 8116 6876 8168 6928
rect 1584 6808 1636 6860
rect 3608 6808 3660 6860
rect 4160 6851 4212 6860
rect 4160 6817 4178 6851
rect 4178 6817 4212 6851
rect 4160 6808 4212 6817
rect 4528 6808 4580 6860
rect 5080 6851 5132 6860
rect 5080 6817 5124 6851
rect 5124 6817 5132 6851
rect 5080 6808 5132 6817
rect 5264 6808 5316 6860
rect 7380 6851 7432 6860
rect 7380 6817 7398 6851
rect 7398 6817 7432 6851
rect 7380 6808 7432 6817
rect 8300 6851 8352 6860
rect 8300 6817 8344 6851
rect 8344 6817 8352 6851
rect 8300 6808 8352 6817
rect 10324 6851 10376 6860
rect 10324 6817 10342 6851
rect 10342 6817 10376 6851
rect 10324 6808 10376 6817
rect 11336 6851 11388 6860
rect 11336 6817 11380 6851
rect 11380 6817 11388 6851
rect 11336 6808 11388 6817
rect 11520 6808 11572 6860
rect 2872 6672 2924 6724
rect 8024 6672 8076 6724
rect 9588 6672 9640 6724
rect 9772 6672 9824 6724
rect 2412 6647 2464 6656
rect 2412 6613 2421 6647
rect 2421 6613 2455 6647
rect 2455 6613 2464 6647
rect 2412 6604 2464 6613
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 1768 6400 1820 6452
rect 2044 6443 2096 6452
rect 2044 6409 2053 6443
rect 2053 6409 2087 6443
rect 2087 6409 2096 6443
rect 2044 6400 2096 6409
rect 3700 6400 3752 6452
rect 4160 6443 4212 6452
rect 4160 6409 4169 6443
rect 4169 6409 4203 6443
rect 4203 6409 4212 6443
rect 4160 6400 4212 6409
rect 5080 6443 5132 6452
rect 5080 6409 5089 6443
rect 5089 6409 5123 6443
rect 5123 6409 5132 6443
rect 5080 6400 5132 6409
rect 7380 6443 7432 6452
rect 7380 6409 7389 6443
rect 7389 6409 7423 6443
rect 7423 6409 7432 6443
rect 7380 6400 7432 6409
rect 8300 6443 8352 6452
rect 8300 6409 8309 6443
rect 8309 6409 8343 6443
rect 8343 6409 8352 6443
rect 8300 6400 8352 6409
rect 10324 6443 10376 6452
rect 10324 6409 10333 6443
rect 10333 6409 10367 6443
rect 10367 6409 10376 6443
rect 10324 6400 10376 6409
rect 11336 6443 11388 6452
rect 11336 6409 11345 6443
rect 11345 6409 11379 6443
rect 11379 6409 11388 6443
rect 11336 6400 11388 6409
rect 1584 6264 1636 6316
rect 2504 6307 2556 6316
rect 2504 6273 2513 6307
rect 2513 6273 2547 6307
rect 2547 6273 2556 6307
rect 2504 6264 2556 6273
rect 2044 6196 2096 6248
rect 3332 6103 3384 6112
rect 3332 6069 3341 6103
rect 3341 6069 3375 6103
rect 3375 6069 3384 6103
rect 3332 6060 3384 6069
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 1400 5856 1452 5908
rect 2596 5856 2648 5908
rect 1400 5763 1452 5772
rect 1400 5729 1444 5763
rect 1444 5729 1452 5763
rect 1400 5720 1452 5729
rect 2504 5763 2556 5772
rect 2504 5729 2522 5763
rect 2522 5729 2556 5763
rect 2504 5720 2556 5729
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 1400 5312 1452 5364
rect 2504 5312 2556 5364
rect 2412 5244 2464 5296
rect 1492 5151 1544 5160
rect 1492 5117 1510 5151
rect 1510 5117 1544 5151
rect 1492 5108 1544 5117
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 2136 4768 2188 4820
rect 1400 4675 1452 4684
rect 1400 4641 1444 4675
rect 1444 4641 1452 4675
rect 1400 4632 1452 4641
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 1400 4224 1452 4276
rect 10692 4156 10744 4208
rect 10876 4156 10928 4208
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 1860 3136 1912 3188
rect 24676 3136 24728 3188
rect 1492 2975 1544 2984
rect 1492 2941 1510 2975
rect 1510 2941 1544 2975
rect 1492 2932 1544 2941
rect 25136 2839 25188 2848
rect 25136 2805 25145 2839
rect 25145 2805 25179 2839
rect 25179 2805 25188 2839
rect 25136 2796 25188 2805
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 1952 2592 2004 2644
rect 2688 2592 2740 2644
rect 24216 2592 24268 2644
rect 24860 2592 24912 2644
rect 1400 2499 1452 2508
rect 1400 2465 1444 2499
rect 1444 2465 1452 2499
rect 1400 2456 1452 2465
rect 2780 2456 2832 2508
rect 25596 2456 25648 2508
rect 24676 2252 24728 2304
rect 25596 2295 25648 2304
rect 25596 2261 25605 2295
rect 25605 2261 25639 2295
rect 25639 2261 25648 2295
rect 25596 2252 25648 2261
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 7656 552 7708 604
rect 7840 552 7892 604
rect 10784 552 10836 604
rect 10876 552 10928 604
<< metal2 >>
rect 662 27520 718 28000
rect 2042 27520 2098 28000
rect 3422 27520 3478 28000
rect 4802 27520 4858 28000
rect 6182 27520 6238 28000
rect 7654 27520 7710 28000
rect 9034 27520 9090 28000
rect 10414 27520 10470 28000
rect 11794 27520 11850 28000
rect 13174 27520 13230 28000
rect 14646 27520 14702 28000
rect 16026 27520 16082 28000
rect 17406 27520 17462 28000
rect 18786 27520 18842 28000
rect 20166 27520 20222 28000
rect 21638 27520 21694 28000
rect 23018 27520 23074 28000
rect 24398 27520 24454 28000
rect 25778 27520 25834 28000
rect 27158 27520 27214 28000
rect 676 24274 704 27520
rect 1490 26344 1546 26353
rect 1490 26279 1546 26288
rect 1398 25392 1454 25401
rect 1398 25327 1454 25336
rect 664 24268 716 24274
rect 664 24210 716 24216
rect 1412 23662 1440 25327
rect 1400 23656 1452 23662
rect 1400 23598 1452 23604
rect 1504 21486 1532 26279
rect 2056 23497 2084 27520
rect 2502 27432 2558 27441
rect 2502 27367 2558 27376
rect 2228 24268 2280 24274
rect 2228 24210 2280 24216
rect 2240 23866 2268 24210
rect 2228 23860 2280 23866
rect 2228 23802 2280 23808
rect 2042 23488 2098 23497
rect 2042 23423 2098 23432
rect 1492 21480 1544 21486
rect 1492 21422 1544 21428
rect 1768 21344 1820 21350
rect 1768 21286 1820 21292
rect 1398 21176 1454 21185
rect 1398 21111 1454 21120
rect 1412 19310 1440 21111
rect 1780 21049 1808 21286
rect 1766 21040 1822 21049
rect 1766 20975 1822 20984
rect 1400 19304 1452 19310
rect 1400 19246 1452 19252
rect 1768 19168 1820 19174
rect 1768 19110 1820 19116
rect 1780 17921 1808 19110
rect 1766 17912 1822 17921
rect 1766 17847 1822 17856
rect 2136 17740 2188 17746
rect 2136 17682 2188 17688
rect 1400 17604 1452 17610
rect 1400 17546 1452 17552
rect 1412 17134 1440 17546
rect 1400 17128 1452 17134
rect 2148 17105 2176 17682
rect 2412 17536 2464 17542
rect 2412 17478 2464 17484
rect 1400 17070 1452 17076
rect 1582 17096 1638 17105
rect 1582 17031 1638 17040
rect 2134 17096 2190 17105
rect 2134 17031 2190 17040
rect 1492 16992 1544 16998
rect 1492 16934 1544 16940
rect 1400 16788 1452 16794
rect 1400 16730 1452 16736
rect 1412 14929 1440 16730
rect 1398 14920 1454 14929
rect 1398 14855 1454 14864
rect 1400 14000 1452 14006
rect 1504 13977 1532 16934
rect 1596 16250 1624 17031
rect 2148 16998 2176 17031
rect 2136 16992 2188 16998
rect 2136 16934 2188 16940
rect 2044 16652 2096 16658
rect 2044 16594 2096 16600
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 1676 16040 1728 16046
rect 1582 16008 1638 16017
rect 1676 15982 1728 15988
rect 1582 15943 1638 15952
rect 1596 14074 1624 15943
rect 1688 15366 1716 15982
rect 2056 15910 2084 16594
rect 2044 15904 2096 15910
rect 2044 15846 2096 15852
rect 2056 15745 2084 15846
rect 2042 15736 2098 15745
rect 2042 15671 2098 15680
rect 1860 15564 1912 15570
rect 1860 15506 1912 15512
rect 1676 15360 1728 15366
rect 1676 15302 1728 15308
rect 1584 14068 1636 14074
rect 1584 14010 1636 14016
rect 1400 13942 1452 13948
rect 1490 13968 1546 13977
rect 1412 12186 1440 13942
rect 1490 13903 1546 13912
rect 1584 13728 1636 13734
rect 1584 13670 1636 13676
rect 1596 13530 1624 13670
rect 1584 13524 1636 13530
rect 1584 13466 1636 13472
rect 1320 12158 1440 12186
rect 1320 8498 1348 12158
rect 1400 12096 1452 12102
rect 1400 12038 1452 12044
rect 1412 10130 1440 12038
rect 1584 11144 1636 11150
rect 1584 11086 1636 11092
rect 1400 10124 1452 10130
rect 1400 10066 1452 10072
rect 1400 9920 1452 9926
rect 1400 9862 1452 9868
rect 1308 8492 1360 8498
rect 1308 8434 1360 8440
rect 1412 8072 1440 9862
rect 1490 9752 1546 9761
rect 1490 9687 1546 9696
rect 1320 8044 1440 8072
rect 1320 7426 1348 8044
rect 1400 7948 1452 7954
rect 1400 7890 1452 7896
rect 1412 7721 1440 7890
rect 1398 7712 1454 7721
rect 1398 7647 1454 7656
rect 1412 7546 1440 7647
rect 1400 7540 1452 7546
rect 1400 7482 1452 7488
rect 1504 7478 1532 9687
rect 1596 9194 1624 11086
rect 1688 9382 1716 15302
rect 1872 14618 1900 15506
rect 1952 15428 2004 15434
rect 1952 15370 2004 15376
rect 1860 14612 1912 14618
rect 1860 14554 1912 14560
rect 1872 14346 1900 14554
rect 1860 14340 1912 14346
rect 1860 14282 1912 14288
rect 1768 14272 1820 14278
rect 1768 14214 1820 14220
rect 1780 11762 1808 14214
rect 1860 12232 1912 12238
rect 1860 12174 1912 12180
rect 1768 11756 1820 11762
rect 1768 11698 1820 11704
rect 1872 11354 1900 12174
rect 1860 11348 1912 11354
rect 1860 11290 1912 11296
rect 1766 10840 1822 10849
rect 1766 10775 1822 10784
rect 1676 9376 1728 9382
rect 1676 9318 1728 9324
rect 1596 9166 1716 9194
rect 1582 8800 1638 8809
rect 1582 8735 1638 8744
rect 1596 8634 1624 8735
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 1492 7472 1544 7478
rect 1320 7398 1440 7426
rect 1492 7414 1544 7420
rect 1412 5914 1440 7398
rect 1596 6866 1624 8434
rect 1688 8090 1716 9166
rect 1676 8084 1728 8090
rect 1676 8026 1728 8032
rect 1584 6860 1636 6866
rect 1584 6802 1636 6808
rect 1490 6624 1546 6633
rect 1490 6559 1546 6568
rect 1400 5908 1452 5914
rect 1400 5850 1452 5856
rect 1400 5772 1452 5778
rect 1400 5714 1452 5720
rect 1412 5681 1440 5714
rect 1398 5672 1454 5681
rect 1398 5607 1454 5616
rect 1412 5370 1440 5607
rect 1400 5364 1452 5370
rect 1400 5306 1452 5312
rect 1504 5166 1532 6559
rect 1596 6322 1624 6802
rect 1780 6458 1808 10775
rect 1860 9648 1912 9654
rect 1860 9590 1912 9596
rect 1872 9178 1900 9590
rect 1860 9172 1912 9178
rect 1860 9114 1912 9120
rect 1858 9072 1914 9081
rect 1858 9007 1914 9016
rect 1768 6452 1820 6458
rect 1768 6394 1820 6400
rect 1584 6316 1636 6322
rect 1584 6258 1636 6264
rect 1492 5160 1544 5166
rect 1492 5102 1544 5108
rect 1400 4684 1452 4690
rect 1400 4626 1452 4632
rect 1412 4593 1440 4626
rect 1398 4584 1454 4593
rect 1398 4519 1454 4528
rect 1412 4282 1440 4519
rect 1400 4276 1452 4282
rect 1400 4218 1452 4224
rect 1582 3496 1638 3505
rect 1582 3431 1638 3440
rect 1492 2984 1544 2990
rect 1492 2926 1544 2932
rect 1398 2544 1454 2553
rect 1398 2479 1400 2488
rect 1452 2479 1454 2488
rect 1400 2450 1452 2456
rect 1504 1465 1532 2926
rect 1490 1456 1546 1465
rect 1490 1391 1546 1400
rect 1596 1306 1624 3431
rect 1872 3194 1900 9007
rect 1964 8430 1992 15370
rect 2148 14618 2176 16934
rect 2424 16794 2452 17478
rect 2412 16788 2464 16794
rect 2412 16730 2464 16736
rect 2320 16720 2372 16726
rect 2320 16662 2372 16668
rect 2228 15972 2280 15978
rect 2228 15914 2280 15920
rect 2136 14612 2188 14618
rect 2136 14554 2188 14560
rect 2136 14476 2188 14482
rect 2136 14418 2188 14424
rect 2148 14006 2176 14418
rect 2136 14000 2188 14006
rect 2134 13968 2136 13977
rect 2188 13968 2190 13977
rect 2134 13903 2190 13912
rect 2136 13456 2188 13462
rect 2136 13398 2188 13404
rect 2044 13252 2096 13258
rect 2044 13194 2096 13200
rect 2056 12374 2084 13194
rect 2148 12442 2176 13398
rect 2240 12986 2268 15914
rect 2332 15026 2360 16662
rect 2424 16114 2452 16730
rect 2516 16658 2544 27367
rect 3436 24834 3464 27520
rect 4816 24857 4844 27520
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 2976 24806 3464 24834
rect 4802 24848 4858 24857
rect 2688 24064 2740 24070
rect 2688 24006 2740 24012
rect 2700 23769 2728 24006
rect 2686 23760 2742 23769
rect 2686 23695 2742 23704
rect 2686 23624 2742 23633
rect 2686 23559 2688 23568
rect 2740 23559 2742 23568
rect 2688 23530 2740 23536
rect 2596 16992 2648 16998
rect 2596 16934 2648 16940
rect 2872 16992 2924 16998
rect 2872 16934 2924 16940
rect 2504 16652 2556 16658
rect 2504 16594 2556 16600
rect 2516 16250 2544 16594
rect 2504 16244 2556 16250
rect 2504 16186 2556 16192
rect 2412 16108 2464 16114
rect 2412 16050 2464 16056
rect 2504 15632 2556 15638
rect 2424 15580 2504 15586
rect 2424 15574 2556 15580
rect 2424 15558 2544 15574
rect 2320 15020 2372 15026
rect 2320 14962 2372 14968
rect 2332 14618 2360 14962
rect 2424 14793 2452 15558
rect 2504 15496 2556 15502
rect 2504 15438 2556 15444
rect 2516 15162 2544 15438
rect 2504 15156 2556 15162
rect 2504 15098 2556 15104
rect 2410 14784 2466 14793
rect 2410 14719 2466 14728
rect 2320 14612 2372 14618
rect 2320 14554 2372 14560
rect 2320 14476 2372 14482
rect 2320 14418 2372 14424
rect 2228 12980 2280 12986
rect 2228 12922 2280 12928
rect 2332 12730 2360 14418
rect 2424 13462 2452 14719
rect 2608 14414 2636 16934
rect 2780 16652 2832 16658
rect 2780 16594 2832 16600
rect 2792 15978 2820 16594
rect 2780 15972 2832 15978
rect 2780 15914 2832 15920
rect 2884 15502 2912 16934
rect 2872 15496 2924 15502
rect 2872 15438 2924 15444
rect 2688 14884 2740 14890
rect 2688 14826 2740 14832
rect 2700 14657 2728 14826
rect 2686 14648 2742 14657
rect 2686 14583 2742 14592
rect 2700 14550 2728 14583
rect 2688 14544 2740 14550
rect 2688 14486 2740 14492
rect 2596 14408 2648 14414
rect 2596 14350 2648 14356
rect 2872 14408 2924 14414
rect 2872 14350 2924 14356
rect 2608 14074 2636 14350
rect 2596 14068 2648 14074
rect 2596 14010 2648 14016
rect 2884 13938 2912 14350
rect 2872 13932 2924 13938
rect 2872 13874 2924 13880
rect 2884 13818 2912 13874
rect 2700 13790 2912 13818
rect 2412 13456 2464 13462
rect 2412 13398 2464 13404
rect 2700 13258 2728 13790
rect 2688 13252 2740 13258
rect 2688 13194 2740 13200
rect 2700 12918 2728 13194
rect 2688 12912 2740 12918
rect 2688 12854 2740 12860
rect 2412 12844 2464 12850
rect 2412 12786 2464 12792
rect 2240 12702 2360 12730
rect 2136 12436 2188 12442
rect 2136 12378 2188 12384
rect 2044 12368 2096 12374
rect 2044 12310 2096 12316
rect 2044 12164 2096 12170
rect 2044 12106 2096 12112
rect 2056 11558 2084 12106
rect 2044 11552 2096 11558
rect 2044 11494 2096 11500
rect 2056 11286 2084 11494
rect 2044 11280 2096 11286
rect 2044 11222 2096 11228
rect 2056 10742 2084 11222
rect 2044 10736 2096 10742
rect 2042 10704 2044 10713
rect 2096 10704 2098 10713
rect 2042 10639 2098 10648
rect 2136 10532 2188 10538
rect 2136 10474 2188 10480
rect 2044 10056 2096 10062
rect 2044 9998 2096 10004
rect 2056 8922 2084 9998
rect 2148 9994 2176 10474
rect 2136 9988 2188 9994
rect 2136 9930 2188 9936
rect 2148 9625 2176 9930
rect 2134 9616 2190 9625
rect 2134 9551 2190 9560
rect 2136 9444 2188 9450
rect 2136 9386 2188 9392
rect 2148 9081 2176 9386
rect 2134 9072 2190 9081
rect 2134 9007 2190 9016
rect 2136 8968 2188 8974
rect 2056 8916 2136 8922
rect 2056 8910 2188 8916
rect 2056 8894 2176 8910
rect 2044 8832 2096 8838
rect 2044 8774 2096 8780
rect 1952 8424 2004 8430
rect 1952 8366 2004 8372
rect 1964 8090 1992 8366
rect 1952 8084 2004 8090
rect 1952 8026 2004 8032
rect 2056 7478 2084 8774
rect 2044 7472 2096 7478
rect 2044 7414 2096 7420
rect 2042 6896 2098 6905
rect 2042 6831 2098 6840
rect 2056 6458 2084 6831
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 2056 6254 2084 6394
rect 2044 6248 2096 6254
rect 2044 6190 2096 6196
rect 2148 4826 2176 8894
rect 2240 8838 2268 12702
rect 2424 12594 2452 12786
rect 2502 12744 2558 12753
rect 2502 12679 2504 12688
rect 2556 12679 2558 12688
rect 2504 12650 2556 12656
rect 2332 12566 2452 12594
rect 2332 9330 2360 12566
rect 2410 12472 2466 12481
rect 2976 12458 3004 24806
rect 4802 24783 4858 24792
rect 3514 24304 3570 24313
rect 3514 24239 3570 24248
rect 3422 22264 3478 22273
rect 3422 22199 3478 22208
rect 3436 21457 3464 22199
rect 3422 21448 3478 21457
rect 3422 21383 3478 21392
rect 3528 20505 3556 24239
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 5538 23760 5594 23769
rect 5538 23695 5594 23704
rect 4250 23488 4306 23497
rect 4250 23423 4306 23432
rect 3514 20496 3570 20505
rect 3514 20431 3570 20440
rect 4066 17776 4122 17785
rect 4066 17711 4122 17720
rect 4080 17610 4108 17711
rect 4068 17604 4120 17610
rect 4068 17546 4120 17552
rect 4080 17338 4108 17546
rect 4068 17332 4120 17338
rect 4068 17274 4120 17280
rect 4080 17134 4108 17274
rect 4068 17128 4120 17134
rect 4068 17070 4120 17076
rect 4264 16046 4292 23423
rect 5448 18216 5500 18222
rect 5448 18158 5500 18164
rect 5460 17746 5488 18158
rect 5552 17882 5580 23695
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 6196 18426 6224 27520
rect 7668 24834 7696 27520
rect 8206 24848 8262 24857
rect 7668 24806 7972 24834
rect 7378 19544 7434 19553
rect 7378 19479 7434 19488
rect 7288 19168 7340 19174
rect 7288 19110 7340 19116
rect 6368 18828 6420 18834
rect 6368 18770 6420 18776
rect 6380 18578 6408 18770
rect 6458 18592 6514 18601
rect 6380 18550 6458 18578
rect 6184 18420 6236 18426
rect 6184 18362 6236 18368
rect 5540 17876 5592 17882
rect 5540 17818 5592 17824
rect 4620 17740 4672 17746
rect 4620 17682 4672 17688
rect 5448 17740 5500 17746
rect 5448 17682 5500 17688
rect 4632 17338 4660 17682
rect 5080 17536 5132 17542
rect 5080 17478 5132 17484
rect 5264 17536 5316 17542
rect 5264 17478 5316 17484
rect 4620 17332 4672 17338
rect 4620 17274 4672 17280
rect 4528 16652 4580 16658
rect 4528 16594 4580 16600
rect 4540 16250 4568 16594
rect 4528 16244 4580 16250
rect 4528 16186 4580 16192
rect 4252 16040 4304 16046
rect 4252 15982 4304 15988
rect 4988 16040 5040 16046
rect 4988 15982 5040 15988
rect 3240 15972 3292 15978
rect 3240 15914 3292 15920
rect 3252 15638 3280 15914
rect 4896 15904 4948 15910
rect 4896 15846 4948 15852
rect 4436 15700 4488 15706
rect 4436 15642 4488 15648
rect 3240 15632 3292 15638
rect 3240 15574 3292 15580
rect 3252 15026 3280 15574
rect 3240 15020 3292 15026
rect 3240 14962 3292 14968
rect 3884 15020 3936 15026
rect 3884 14962 3936 14968
rect 4160 15020 4212 15026
rect 4160 14962 4212 14968
rect 3240 14816 3292 14822
rect 3238 14784 3240 14793
rect 3292 14784 3294 14793
rect 3238 14719 3294 14728
rect 3054 14648 3110 14657
rect 3896 14618 3924 14962
rect 3976 14884 4028 14890
rect 3976 14826 4028 14832
rect 3988 14618 4016 14826
rect 3054 14583 3110 14592
rect 3884 14612 3936 14618
rect 3068 13530 3096 14583
rect 3884 14554 3936 14560
rect 3976 14612 4028 14618
rect 3976 14554 4028 14560
rect 4172 14346 4200 14962
rect 4448 14482 4476 15642
rect 4804 15564 4856 15570
rect 4804 15506 4856 15512
rect 4816 15094 4844 15506
rect 4908 15473 4936 15846
rect 4894 15464 4950 15473
rect 4894 15399 4950 15408
rect 4804 15088 4856 15094
rect 4804 15030 4856 15036
rect 4528 14952 4580 14958
rect 4528 14894 4580 14900
rect 4436 14476 4488 14482
rect 4436 14418 4488 14424
rect 4160 14340 4212 14346
rect 4160 14282 4212 14288
rect 3516 14000 3568 14006
rect 3516 13942 3568 13948
rect 3528 13818 3556 13942
rect 4172 13870 4200 14282
rect 4344 14272 4396 14278
rect 4344 14214 4396 14220
rect 4356 13870 4384 14214
rect 4448 14074 4476 14418
rect 4436 14068 4488 14074
rect 4436 14010 4488 14016
rect 3344 13802 3556 13818
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 4344 13864 4396 13870
rect 4344 13806 4396 13812
rect 3332 13796 3556 13802
rect 3384 13790 3556 13796
rect 3332 13738 3384 13744
rect 3528 13530 3556 13790
rect 4172 13705 4200 13806
rect 4158 13696 4214 13705
rect 4158 13631 4214 13640
rect 4356 13530 4384 13806
rect 4436 13796 4488 13802
rect 4436 13738 4488 13744
rect 3056 13524 3108 13530
rect 3056 13466 3108 13472
rect 3516 13524 3568 13530
rect 3516 13466 3568 13472
rect 4344 13524 4396 13530
rect 4344 13466 4396 13472
rect 4448 13462 4476 13738
rect 4540 13734 4568 14894
rect 4816 14822 4844 15030
rect 4804 14816 4856 14822
rect 4804 14758 4856 14764
rect 4528 13728 4580 13734
rect 4528 13670 4580 13676
rect 4436 13456 4488 13462
rect 4488 13416 4660 13444
rect 4436 13398 4488 13404
rect 4436 12912 4488 12918
rect 4436 12854 4488 12860
rect 3884 12708 3936 12714
rect 3884 12650 3936 12656
rect 2410 12407 2466 12416
rect 2792 12430 3004 12458
rect 3896 12442 3924 12650
rect 4344 12640 4396 12646
rect 4344 12582 4396 12588
rect 3884 12436 3936 12442
rect 2424 12238 2452 12407
rect 2792 12356 2820 12430
rect 3884 12378 3936 12384
rect 3056 12368 3108 12374
rect 2792 12328 2912 12356
rect 2412 12232 2464 12238
rect 2412 12174 2464 12180
rect 2412 11756 2464 11762
rect 2412 11698 2464 11704
rect 2780 11756 2832 11762
rect 2780 11698 2832 11704
rect 2424 11354 2452 11698
rect 2792 11642 2820 11698
rect 2504 11620 2556 11626
rect 2504 11562 2556 11568
rect 2700 11614 2820 11642
rect 2516 11529 2544 11562
rect 2502 11520 2558 11529
rect 2502 11455 2558 11464
rect 2412 11348 2464 11354
rect 2412 11290 2464 11296
rect 2516 11234 2544 11455
rect 2424 11206 2544 11234
rect 2424 10198 2452 11206
rect 2504 11144 2556 11150
rect 2504 11086 2556 11092
rect 2412 10192 2464 10198
rect 2412 10134 2464 10140
rect 2424 9722 2452 10134
rect 2516 10062 2544 11086
rect 2700 10742 2728 11614
rect 2780 11552 2832 11558
rect 2780 11494 2832 11500
rect 2688 10736 2740 10742
rect 2688 10678 2740 10684
rect 2792 10588 2820 11494
rect 2700 10560 2820 10588
rect 2504 10056 2556 10062
rect 2504 9998 2556 10004
rect 2596 9920 2648 9926
rect 2502 9888 2558 9897
rect 2596 9862 2648 9868
rect 2502 9823 2558 9832
rect 2412 9716 2464 9722
rect 2412 9658 2464 9664
rect 2332 9302 2452 9330
rect 2318 9208 2374 9217
rect 2318 9143 2374 9152
rect 2332 9042 2360 9143
rect 2320 9036 2372 9042
rect 2320 8978 2372 8984
rect 2228 8832 2280 8838
rect 2228 8774 2280 8780
rect 2228 8628 2280 8634
rect 2228 8570 2280 8576
rect 2240 8294 2268 8570
rect 2228 8288 2280 8294
rect 2228 8230 2280 8236
rect 2240 8022 2268 8230
rect 2332 8090 2360 8978
rect 2320 8084 2372 8090
rect 2320 8026 2372 8032
rect 2228 8016 2280 8022
rect 2228 7958 2280 7964
rect 2424 7868 2452 9302
rect 2240 7840 2452 7868
rect 2136 4820 2188 4826
rect 2136 4762 2188 4768
rect 1860 3188 1912 3194
rect 1860 3130 1912 3136
rect 2240 2802 2268 7840
rect 2412 7744 2464 7750
rect 2412 7686 2464 7692
rect 2424 6662 2452 7686
rect 2412 6656 2464 6662
rect 2412 6598 2464 6604
rect 2424 5302 2452 6598
rect 2516 6322 2544 9823
rect 2608 9518 2636 9862
rect 2700 9586 2728 10560
rect 2688 9580 2740 9586
rect 2688 9522 2740 9528
rect 2596 9512 2648 9518
rect 2596 9454 2648 9460
rect 2608 7041 2636 9454
rect 2778 9344 2834 9353
rect 2778 9279 2834 9288
rect 2792 9110 2820 9279
rect 2780 9104 2832 9110
rect 2780 9046 2832 9052
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 2700 7970 2728 8910
rect 2792 8634 2820 9046
rect 2780 8628 2832 8634
rect 2780 8570 2832 8576
rect 2884 8537 2912 12328
rect 3056 12310 3108 12316
rect 4252 12368 4304 12374
rect 4252 12310 4304 12316
rect 2962 11792 3018 11801
rect 3068 11762 3096 12310
rect 4160 12232 4212 12238
rect 4160 12174 4212 12180
rect 2962 11727 3018 11736
rect 3056 11756 3108 11762
rect 2870 8528 2926 8537
rect 2780 8492 2832 8498
rect 2870 8463 2926 8472
rect 2780 8434 2832 8440
rect 2792 8090 2820 8434
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 2872 8016 2924 8022
rect 2700 7942 2820 7970
rect 2872 7958 2924 7964
rect 2792 7750 2820 7942
rect 2780 7744 2832 7750
rect 2780 7686 2832 7692
rect 2884 7546 2912 7958
rect 2872 7540 2924 7546
rect 2872 7482 2924 7488
rect 2976 7426 3004 11727
rect 3056 11698 3108 11704
rect 4172 11354 4200 12174
rect 4264 11830 4292 12310
rect 4252 11824 4304 11830
rect 4252 11766 4304 11772
rect 4356 11354 4384 12582
rect 4448 12238 4476 12854
rect 4528 12436 4580 12442
rect 4528 12378 4580 12384
rect 4436 12232 4488 12238
rect 4436 12174 4488 12180
rect 4160 11348 4212 11354
rect 4160 11290 4212 11296
rect 4344 11348 4396 11354
rect 4344 11290 4396 11296
rect 4172 10674 4200 11290
rect 3792 10668 3844 10674
rect 3792 10610 3844 10616
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 3804 10577 3832 10610
rect 3790 10568 3846 10577
rect 3790 10503 3792 10512
rect 3844 10503 3846 10512
rect 3792 10474 3844 10480
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3436 9897 3464 10406
rect 3804 10266 3832 10474
rect 3792 10260 3844 10266
rect 3792 10202 3844 10208
rect 4252 10192 4304 10198
rect 4252 10134 4304 10140
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 3422 9888 3478 9897
rect 3422 9823 3478 9832
rect 4172 9722 4200 9998
rect 4160 9716 4212 9722
rect 4160 9658 4212 9664
rect 3148 9580 3200 9586
rect 3148 9522 3200 9528
rect 3056 9444 3108 9450
rect 3056 9386 3108 9392
rect 2884 7398 3004 7426
rect 3068 8786 3096 9386
rect 3160 9110 3188 9522
rect 4264 9489 4292 10134
rect 4250 9480 4306 9489
rect 3240 9444 3292 9450
rect 3240 9386 3292 9392
rect 3884 9444 3936 9450
rect 4250 9415 4306 9424
rect 3884 9386 3936 9392
rect 3148 9104 3200 9110
rect 3148 9046 3200 9052
rect 3252 8945 3280 9386
rect 3896 9178 3924 9386
rect 4264 9382 4292 9415
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 4252 9376 4304 9382
rect 4252 9318 4304 9324
rect 3884 9172 3936 9178
rect 3884 9114 3936 9120
rect 3238 8936 3294 8945
rect 3238 8871 3294 8880
rect 3606 8936 3662 8945
rect 3606 8871 3662 8880
rect 3148 8832 3200 8838
rect 3068 8780 3148 8786
rect 3068 8774 3200 8780
rect 3068 8758 3188 8774
rect 2594 7032 2650 7041
rect 2594 6967 2650 6976
rect 2884 6730 2912 7398
rect 2964 7268 3016 7274
rect 2964 7210 3016 7216
rect 2976 7002 3004 7210
rect 2964 6996 3016 7002
rect 2964 6938 3016 6944
rect 2872 6724 2924 6730
rect 2872 6666 2924 6672
rect 3068 6610 3096 8758
rect 3148 8492 3200 8498
rect 3148 8434 3200 8440
rect 3160 8022 3188 8434
rect 3148 8016 3200 8022
rect 3148 7958 3200 7964
rect 3516 7744 3568 7750
rect 3516 7686 3568 7692
rect 3528 7002 3556 7686
rect 3620 7274 3648 8871
rect 3896 8498 3924 9114
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 3700 8084 3752 8090
rect 3700 8026 3752 8032
rect 3608 7268 3660 7274
rect 3608 7210 3660 7216
rect 3516 6996 3568 7002
rect 3516 6938 3568 6944
rect 3620 6866 3648 7210
rect 3608 6860 3660 6866
rect 3608 6802 3660 6808
rect 2792 6582 3096 6610
rect 2504 6316 2556 6322
rect 2504 6258 2556 6264
rect 2594 5944 2650 5953
rect 2594 5879 2596 5888
rect 2648 5879 2650 5888
rect 2596 5850 2648 5856
rect 2502 5808 2558 5817
rect 2502 5743 2504 5752
rect 2556 5743 2558 5752
rect 2504 5714 2556 5720
rect 2516 5370 2544 5714
rect 2504 5364 2556 5370
rect 2504 5306 2556 5312
rect 2412 5296 2464 5302
rect 2412 5238 2464 5244
rect 2792 4026 2820 6582
rect 3712 6458 3740 8026
rect 3896 7410 3924 8434
rect 4080 8362 4108 9318
rect 4448 9217 4476 12174
rect 4540 11762 4568 12378
rect 4632 11898 4660 13416
rect 4620 11892 4672 11898
rect 4620 11834 4672 11840
rect 4528 11756 4580 11762
rect 4528 11698 4580 11704
rect 4632 11626 4660 11834
rect 4620 11620 4672 11626
rect 4620 11562 4672 11568
rect 4632 11286 4660 11562
rect 4620 11280 4672 11286
rect 4620 11222 4672 11228
rect 4632 10810 4660 11222
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 4816 10470 4844 14758
rect 4896 14544 4948 14550
rect 4896 14486 4948 14492
rect 4908 13802 4936 14486
rect 4896 13796 4948 13802
rect 4896 13738 4948 13744
rect 4896 13388 4948 13394
rect 4896 13330 4948 13336
rect 4908 12646 4936 13330
rect 4896 12640 4948 12646
rect 4896 12582 4948 12588
rect 4804 10464 4856 10470
rect 4804 10406 4856 10412
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 4528 9988 4580 9994
rect 4528 9930 4580 9936
rect 4434 9208 4490 9217
rect 4434 9143 4490 9152
rect 4434 9072 4490 9081
rect 4434 9007 4490 9016
rect 4448 8974 4476 9007
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 4436 8016 4488 8022
rect 4436 7958 4488 7964
rect 4448 7546 4476 7958
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 4540 6866 4568 9930
rect 4632 9586 4660 9998
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 4632 7868 4660 9522
rect 4712 9444 4764 9450
rect 4712 9386 4764 9392
rect 4724 9042 4752 9386
rect 4712 9036 4764 9042
rect 4712 8978 4764 8984
rect 4712 7880 4764 7886
rect 4632 7840 4712 7868
rect 4712 7822 4764 7828
rect 4724 7002 4752 7822
rect 4816 7546 4844 10406
rect 5000 9738 5028 15982
rect 5092 14385 5120 17478
rect 5276 17134 5304 17478
rect 5264 17128 5316 17134
rect 5264 17070 5316 17076
rect 5276 16454 5304 17070
rect 5552 16794 5580 17818
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 6276 17060 6328 17066
rect 6276 17002 6328 17008
rect 5540 16788 5592 16794
rect 5540 16730 5592 16736
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 5264 16448 5316 16454
rect 5264 16390 5316 16396
rect 5276 16046 5304 16390
rect 5172 16040 5224 16046
rect 5172 15982 5224 15988
rect 5264 16040 5316 16046
rect 5264 15982 5316 15988
rect 5184 15609 5212 15982
rect 5170 15600 5226 15609
rect 5170 15535 5226 15544
rect 5172 15496 5224 15502
rect 5276 15484 5304 15982
rect 5354 15736 5410 15745
rect 5354 15671 5410 15680
rect 5224 15456 5304 15484
rect 5172 15438 5224 15444
rect 5184 14822 5212 15438
rect 5172 14816 5224 14822
rect 5172 14758 5224 14764
rect 5264 14816 5316 14822
rect 5264 14758 5316 14764
rect 5078 14376 5134 14385
rect 5078 14311 5134 14320
rect 5080 14272 5132 14278
rect 5080 14214 5132 14220
rect 5092 9994 5120 14214
rect 5184 13394 5212 14758
rect 5172 13388 5224 13394
rect 5172 13330 5224 13336
rect 5184 13297 5212 13330
rect 5170 13288 5226 13297
rect 5170 13223 5226 13232
rect 5184 12850 5212 13223
rect 5172 12844 5224 12850
rect 5172 12786 5224 12792
rect 5276 12481 5304 14758
rect 5368 14278 5396 15671
rect 5356 14272 5408 14278
rect 5356 14214 5408 14220
rect 5460 13920 5488 16594
rect 6092 16584 6144 16590
rect 6092 16526 6144 16532
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 6104 15706 6132 16526
rect 6184 16176 6236 16182
rect 6184 16118 6236 16124
rect 6092 15700 6144 15706
rect 6092 15642 6144 15648
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5540 13932 5592 13938
rect 5460 13892 5540 13920
rect 5540 13874 5592 13880
rect 6196 13546 6224 16118
rect 6288 14482 6316 17002
rect 6276 14476 6328 14482
rect 6276 14418 6328 14424
rect 6288 14074 6316 14418
rect 6276 14068 6328 14074
rect 6276 14010 6328 14016
rect 6196 13518 6316 13546
rect 6184 13456 6236 13462
rect 6184 13398 6236 13404
rect 6000 13184 6052 13190
rect 6000 13126 6052 13132
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5540 12912 5592 12918
rect 5538 12880 5540 12889
rect 5592 12880 5594 12889
rect 5538 12815 5594 12824
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 5262 12472 5318 12481
rect 5262 12407 5318 12416
rect 5368 12102 5396 12718
rect 6012 12646 6040 13126
rect 6196 12646 6224 13398
rect 6288 13025 6316 13518
rect 6274 13016 6330 13025
rect 6274 12951 6330 12960
rect 6000 12640 6052 12646
rect 6184 12640 6236 12646
rect 6000 12582 6052 12588
rect 6182 12608 6184 12617
rect 6236 12608 6238 12617
rect 6012 12306 6040 12582
rect 6182 12543 6238 12552
rect 6000 12300 6052 12306
rect 6000 12242 6052 12248
rect 5356 12096 5408 12102
rect 5356 12038 5408 12044
rect 5264 10600 5316 10606
rect 5264 10542 5316 10548
rect 5276 10266 5304 10542
rect 5264 10260 5316 10266
rect 5264 10202 5316 10208
rect 5080 9988 5132 9994
rect 5080 9930 5132 9936
rect 5000 9710 5120 9738
rect 4894 9616 4950 9625
rect 4894 9551 4896 9560
rect 4948 9551 4950 9560
rect 4896 9522 4948 9528
rect 4908 7886 4936 9522
rect 4988 8424 5040 8430
rect 4988 8366 5040 8372
rect 4896 7880 4948 7886
rect 4896 7822 4948 7828
rect 4804 7540 4856 7546
rect 4804 7482 4856 7488
rect 4816 7342 4844 7482
rect 4804 7336 4856 7342
rect 4804 7278 4856 7284
rect 4802 7032 4858 7041
rect 4712 6996 4764 7002
rect 4802 6967 4804 6976
rect 4712 6938 4764 6944
rect 4856 6967 4858 6976
rect 4804 6938 4856 6944
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 4528 6860 4580 6866
rect 4528 6802 4580 6808
rect 4172 6458 4200 6802
rect 3700 6452 3752 6458
rect 3700 6394 3752 6400
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 3332 6112 3384 6118
rect 3332 6054 3384 6060
rect 1964 2774 2268 2802
rect 2700 3998 2820 4026
rect 1964 2650 1992 2774
rect 2700 2650 2728 3998
rect 3344 3641 3372 6054
rect 4908 5817 4936 7822
rect 5000 7206 5028 8366
rect 5092 7313 5120 9710
rect 5264 9716 5316 9722
rect 5264 9658 5316 9664
rect 5078 7304 5134 7313
rect 5078 7239 5134 7248
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 5078 6896 5134 6905
rect 5276 6866 5304 9658
rect 5078 6831 5080 6840
rect 5132 6831 5134 6840
rect 5264 6860 5316 6866
rect 5080 6802 5132 6808
rect 5264 6802 5316 6808
rect 5092 6458 5120 6802
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 5368 5953 5396 12038
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 6012 11558 6040 12242
rect 6000 11552 6052 11558
rect 6000 11494 6052 11500
rect 5540 11008 5592 11014
rect 5540 10950 5592 10956
rect 5552 10674 5580 10950
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 6288 10130 6316 12951
rect 6276 10124 6328 10130
rect 6276 10066 6328 10072
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 6288 9722 6316 10066
rect 6092 9716 6144 9722
rect 6092 9658 6144 9664
rect 6276 9716 6328 9722
rect 6276 9658 6328 9664
rect 5448 9104 5500 9110
rect 5448 9046 5500 9052
rect 5460 8362 5488 9046
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5552 8514 5580 8910
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5552 8486 5672 8514
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5448 8356 5500 8362
rect 5448 8298 5500 8304
rect 5552 8022 5580 8366
rect 5644 8090 5672 8486
rect 5632 8084 5684 8090
rect 5632 8026 5684 8032
rect 5540 8016 5592 8022
rect 5540 7958 5592 7964
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 6104 7546 6132 9658
rect 6276 7948 6328 7954
rect 6276 7890 6328 7896
rect 6092 7540 6144 7546
rect 6092 7482 6144 7488
rect 6288 7478 6316 7890
rect 6276 7472 6328 7478
rect 6276 7414 6328 7420
rect 6380 6905 6408 18550
rect 6458 18527 6514 18536
rect 6472 18426 6500 18527
rect 6460 18420 6512 18426
rect 6460 18362 6512 18368
rect 7300 18290 7328 19110
rect 7288 18284 7340 18290
rect 7288 18226 7340 18232
rect 6828 18148 6880 18154
rect 6828 18090 6880 18096
rect 7012 18148 7064 18154
rect 7012 18090 7064 18096
rect 6644 17060 6696 17066
rect 6644 17002 6696 17008
rect 6552 16992 6604 16998
rect 6552 16934 6604 16940
rect 6564 15570 6592 16934
rect 6656 16726 6684 17002
rect 6644 16720 6696 16726
rect 6644 16662 6696 16668
rect 6656 16250 6684 16662
rect 6644 16244 6696 16250
rect 6644 16186 6696 16192
rect 6552 15564 6604 15570
rect 6552 15506 6604 15512
rect 6564 14822 6592 15506
rect 6552 14816 6604 14822
rect 6552 14758 6604 14764
rect 6564 12782 6592 14758
rect 6656 14550 6684 16186
rect 6736 15972 6788 15978
rect 6736 15914 6788 15920
rect 6644 14544 6696 14550
rect 6644 14486 6696 14492
rect 6656 14074 6684 14486
rect 6748 14113 6776 15914
rect 6840 15722 6868 18090
rect 7024 17814 7052 18090
rect 7194 17912 7250 17921
rect 7194 17847 7250 17856
rect 7208 17814 7236 17847
rect 7012 17808 7064 17814
rect 7012 17750 7064 17756
rect 7196 17808 7248 17814
rect 7196 17750 7248 17756
rect 6920 17536 6972 17542
rect 6920 17478 6972 17484
rect 6932 17134 6960 17478
rect 7024 17338 7052 17750
rect 7012 17332 7064 17338
rect 7012 17274 7064 17280
rect 6920 17128 6972 17134
rect 6920 17070 6972 17076
rect 6932 15910 6960 17070
rect 7024 16794 7052 17274
rect 7208 16794 7236 17750
rect 7012 16788 7064 16794
rect 7012 16730 7064 16736
rect 7196 16788 7248 16794
rect 7196 16730 7248 16736
rect 7288 16448 7340 16454
rect 7288 16390 7340 16396
rect 7300 16046 7328 16390
rect 7288 16040 7340 16046
rect 7288 15982 7340 15988
rect 6920 15904 6972 15910
rect 6920 15846 6972 15852
rect 6840 15706 6960 15722
rect 6840 15700 6972 15706
rect 6840 15694 6920 15700
rect 6920 15642 6972 15648
rect 6932 15026 6960 15642
rect 7300 15570 7328 15982
rect 7288 15564 7340 15570
rect 7288 15506 7340 15512
rect 7102 15464 7158 15473
rect 7102 15399 7158 15408
rect 6920 15020 6972 15026
rect 6920 14962 6972 14968
rect 7012 14884 7064 14890
rect 7012 14826 7064 14832
rect 7024 14793 7052 14826
rect 7010 14784 7066 14793
rect 7010 14719 7066 14728
rect 7024 14618 7052 14719
rect 7012 14612 7064 14618
rect 7012 14554 7064 14560
rect 6734 14104 6790 14113
rect 6644 14068 6696 14074
rect 6734 14039 6790 14048
rect 6644 14010 6696 14016
rect 6736 13932 6788 13938
rect 6736 13874 6788 13880
rect 6748 13530 6776 13874
rect 6736 13524 6788 13530
rect 6736 13466 6788 13472
rect 7116 13326 7144 15399
rect 7196 14816 7248 14822
rect 7194 14784 7196 14793
rect 7248 14784 7250 14793
rect 7194 14719 7250 14728
rect 7196 14272 7248 14278
rect 7196 14214 7248 14220
rect 7208 13462 7236 14214
rect 7196 13456 7248 13462
rect 7196 13398 7248 13404
rect 7104 13320 7156 13326
rect 7104 13262 7156 13268
rect 7116 12986 7144 13262
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 6552 12776 6604 12782
rect 6604 12736 6684 12764
rect 6552 12718 6604 12724
rect 6552 12300 6604 12306
rect 6552 12242 6604 12248
rect 6564 12102 6592 12242
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 6564 11694 6592 12038
rect 6552 11688 6604 11694
rect 6552 11630 6604 11636
rect 6564 11218 6592 11630
rect 6552 11212 6604 11218
rect 6552 11154 6604 11160
rect 6564 10606 6592 11154
rect 6656 10690 6684 12736
rect 7104 12640 7156 12646
rect 7104 12582 7156 12588
rect 6736 11824 6788 11830
rect 6736 11766 6788 11772
rect 6748 11286 6776 11766
rect 6828 11688 6880 11694
rect 6828 11630 6880 11636
rect 6736 11280 6788 11286
rect 6736 11222 6788 11228
rect 6748 10810 6776 11222
rect 6840 11132 6868 11630
rect 6920 11144 6972 11150
rect 6840 11104 6920 11132
rect 6736 10804 6788 10810
rect 6736 10746 6788 10752
rect 6656 10662 6776 10690
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 6564 10130 6592 10542
rect 6552 10124 6604 10130
rect 6552 10066 6604 10072
rect 6564 9722 6592 10066
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 6748 8090 6776 10662
rect 6840 10198 6868 11104
rect 6920 11086 6972 11092
rect 7116 11014 7144 12582
rect 7196 12368 7248 12374
rect 7196 12310 7248 12316
rect 7208 11762 7236 12310
rect 7196 11756 7248 11762
rect 7196 11698 7248 11704
rect 7208 11529 7236 11698
rect 7194 11520 7250 11529
rect 7194 11455 7250 11464
rect 7208 11354 7236 11455
rect 7196 11348 7248 11354
rect 7196 11290 7248 11296
rect 7104 11008 7156 11014
rect 7104 10950 7156 10956
rect 7116 10810 7144 10950
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 6828 10192 6880 10198
rect 6828 10134 6880 10140
rect 7196 10192 7248 10198
rect 7196 10134 7248 10140
rect 7208 9466 7236 10134
rect 7286 9480 7342 9489
rect 7208 9438 7286 9466
rect 7286 9415 7288 9424
rect 7340 9415 7342 9424
rect 7288 9386 7340 9392
rect 7012 9376 7064 9382
rect 7010 9344 7012 9353
rect 7064 9344 7066 9353
rect 7010 9279 7066 9288
rect 7024 9178 7052 9279
rect 7012 9172 7064 9178
rect 7012 9114 7064 9120
rect 7196 9104 7248 9110
rect 7196 9046 7248 9052
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6736 8084 6788 8090
rect 6736 8026 6788 8032
rect 6840 8022 6868 8366
rect 7208 8362 7236 9046
rect 7300 8634 7328 9386
rect 7288 8628 7340 8634
rect 7288 8570 7340 8576
rect 7196 8356 7248 8362
rect 7196 8298 7248 8304
rect 6828 8016 6880 8022
rect 6828 7958 6880 7964
rect 6736 7948 6788 7954
rect 6736 7890 6788 7896
rect 6748 7478 6776 7890
rect 6736 7472 6788 7478
rect 6736 7414 6788 7420
rect 6748 7274 6776 7414
rect 6736 7268 6788 7274
rect 6736 7210 6788 7216
rect 6748 7002 6776 7210
rect 6736 6996 6788 7002
rect 6736 6938 6788 6944
rect 6366 6896 6422 6905
rect 7392 6866 7420 19479
rect 7656 19168 7708 19174
rect 7656 19110 7708 19116
rect 7564 18896 7616 18902
rect 7564 18838 7616 18844
rect 7472 18760 7524 18766
rect 7472 18702 7524 18708
rect 7484 17882 7512 18702
rect 7576 18426 7604 18838
rect 7564 18420 7616 18426
rect 7564 18362 7616 18368
rect 7472 17876 7524 17882
rect 7472 17818 7524 17824
rect 7576 17814 7604 18362
rect 7668 18057 7696 19110
rect 7748 18760 7800 18766
rect 7748 18702 7800 18708
rect 7760 18465 7788 18702
rect 7746 18456 7802 18465
rect 7746 18391 7802 18400
rect 7654 18048 7710 18057
rect 7654 17983 7710 17992
rect 7564 17808 7616 17814
rect 7564 17750 7616 17756
rect 7576 17338 7604 17750
rect 7564 17332 7616 17338
rect 7564 17274 7616 17280
rect 7668 16153 7696 17983
rect 7760 17610 7788 18391
rect 7840 18148 7892 18154
rect 7840 18090 7892 18096
rect 7852 17814 7880 18090
rect 7840 17808 7892 17814
rect 7840 17750 7892 17756
rect 7748 17604 7800 17610
rect 7748 17546 7800 17552
rect 7654 16144 7710 16153
rect 7654 16079 7710 16088
rect 7656 14884 7708 14890
rect 7656 14826 7708 14832
rect 7668 13462 7696 14826
rect 7748 14612 7800 14618
rect 7748 14554 7800 14560
rect 7760 14074 7788 14554
rect 7748 14068 7800 14074
rect 7748 14010 7800 14016
rect 7656 13456 7708 13462
rect 7656 13398 7708 13404
rect 7838 13424 7894 13433
rect 7838 13359 7894 13368
rect 7564 12776 7616 12782
rect 7564 12718 7616 12724
rect 7472 12708 7524 12714
rect 7472 12650 7524 12656
rect 7484 12073 7512 12650
rect 7576 12102 7604 12718
rect 7564 12096 7616 12102
rect 7470 12064 7526 12073
rect 7564 12038 7616 12044
rect 7470 11999 7526 12008
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7472 11008 7524 11014
rect 7472 10950 7524 10956
rect 7484 10538 7512 10950
rect 7576 10713 7604 11494
rect 7562 10704 7618 10713
rect 7562 10639 7618 10648
rect 7576 10538 7604 10639
rect 7472 10532 7524 10538
rect 7472 10474 7524 10480
rect 7564 10532 7616 10538
rect 7564 10474 7616 10480
rect 7484 8090 7512 10474
rect 7576 10266 7604 10474
rect 7564 10260 7616 10266
rect 7564 10202 7616 10208
rect 7748 9444 7800 9450
rect 7748 9386 7800 9392
rect 7760 9178 7788 9386
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 6366 6831 6422 6840
rect 7380 6860 7432 6866
rect 7380 6802 7432 6808
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 7392 6458 7420 6802
rect 7380 6452 7432 6458
rect 7380 6394 7432 6400
rect 5354 5944 5410 5953
rect 5354 5879 5410 5888
rect 4894 5808 4950 5817
rect 4894 5743 4950 5752
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 4526 4040 4582 4049
rect 4526 3975 4582 3984
rect 3330 3632 3386 3641
rect 3330 3567 3386 3576
rect 1952 2644 2004 2650
rect 1952 2586 2004 2592
rect 2688 2644 2740 2650
rect 2688 2586 2740 2592
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 1504 1278 1624 1306
rect 1504 480 1532 1278
rect 2792 513 2820 2450
rect 2778 504 2834 513
rect 1490 0 1546 480
rect 4540 480 4568 3975
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 7852 610 7880 13359
rect 7944 10588 7972 24806
rect 8206 24783 8262 24792
rect 8220 19553 8248 24783
rect 8206 19544 8262 19553
rect 8206 19479 8262 19488
rect 9048 19310 9076 27520
rect 10428 25786 10456 27520
rect 9692 25758 10456 25786
rect 8392 19304 8444 19310
rect 8392 19246 8444 19252
rect 9036 19304 9088 19310
rect 9036 19246 9088 19252
rect 9588 19304 9640 19310
rect 9692 19292 9720 25758
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 11808 24834 11836 27520
rect 13188 24834 13216 27520
rect 11808 24806 12112 24834
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10784 21072 10836 21078
rect 10690 21040 10746 21049
rect 10784 21014 10836 21020
rect 11888 21072 11940 21078
rect 11888 21014 11940 21020
rect 10690 20975 10746 20984
rect 10704 20942 10732 20975
rect 10692 20936 10744 20942
rect 10692 20878 10744 20884
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10704 20058 10732 20878
rect 10796 20466 10824 21014
rect 11900 20602 11928 21014
rect 11888 20596 11940 20602
rect 11888 20538 11940 20544
rect 10784 20460 10836 20466
rect 10784 20402 10836 20408
rect 11900 20398 11928 20538
rect 11888 20392 11940 20398
rect 11888 20334 11940 20340
rect 11900 20058 11928 20334
rect 11980 20324 12032 20330
rect 11980 20266 12032 20272
rect 10692 20052 10744 20058
rect 10692 19994 10744 20000
rect 11888 20052 11940 20058
rect 11888 19994 11940 20000
rect 11992 19990 12020 20266
rect 11980 19984 12032 19990
rect 11980 19926 12032 19932
rect 9864 19916 9916 19922
rect 9864 19858 9916 19864
rect 10968 19916 11020 19922
rect 10968 19858 11020 19864
rect 9876 19553 9904 19858
rect 10048 19712 10100 19718
rect 10048 19654 10100 19660
rect 9862 19544 9918 19553
rect 9862 19479 9864 19488
rect 9916 19479 9918 19488
rect 9864 19450 9916 19456
rect 9640 19264 9720 19292
rect 9588 19246 9640 19252
rect 8208 17060 8260 17066
rect 8208 17002 8260 17008
rect 8220 16726 8248 17002
rect 8208 16720 8260 16726
rect 8208 16662 8260 16668
rect 8220 16114 8248 16662
rect 8300 16652 8352 16658
rect 8300 16594 8352 16600
rect 8312 16250 8340 16594
rect 8300 16244 8352 16250
rect 8300 16186 8352 16192
rect 8208 16108 8260 16114
rect 8208 16050 8260 16056
rect 8116 16040 8168 16046
rect 8116 15982 8168 15988
rect 8128 15570 8156 15982
rect 8312 15706 8340 16186
rect 8300 15700 8352 15706
rect 8300 15642 8352 15648
rect 8024 15564 8076 15570
rect 8024 15506 8076 15512
rect 8116 15564 8168 15570
rect 8116 15506 8168 15512
rect 8036 15094 8064 15506
rect 8024 15088 8076 15094
rect 8024 15030 8076 15036
rect 8300 15088 8352 15094
rect 8300 15030 8352 15036
rect 8206 14512 8262 14521
rect 8206 14447 8208 14456
rect 8260 14447 8262 14456
rect 8208 14418 8260 14424
rect 8220 14074 8248 14418
rect 8312 14249 8340 15030
rect 8298 14240 8354 14249
rect 8298 14175 8354 14184
rect 8208 14068 8260 14074
rect 8208 14010 8260 14016
rect 8024 12640 8076 12646
rect 8024 12582 8076 12588
rect 8036 12374 8064 12582
rect 8024 12368 8076 12374
rect 8024 12310 8076 12316
rect 8036 10742 8064 12310
rect 8208 11212 8260 11218
rect 8208 11154 8260 11160
rect 8220 11098 8248 11154
rect 8220 11070 8340 11098
rect 8312 10810 8340 11070
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 8024 10736 8076 10742
rect 8024 10678 8076 10684
rect 7944 10560 8156 10588
rect 8024 10056 8076 10062
rect 8024 9998 8076 10004
rect 7932 8968 7984 8974
rect 7932 8910 7984 8916
rect 7944 8294 7972 8910
rect 8036 8838 8064 9998
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 7932 8288 7984 8294
rect 7932 8230 7984 8236
rect 7944 7410 7972 8230
rect 7932 7404 7984 7410
rect 7932 7346 7984 7352
rect 8036 6730 8064 8774
rect 8128 7954 8156 10560
rect 8116 7948 8168 7954
rect 8116 7890 8168 7896
rect 8128 7546 8156 7890
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 8128 6934 8156 7482
rect 8404 7342 8432 19246
rect 8944 19168 8996 19174
rect 8944 19110 8996 19116
rect 9128 19168 9180 19174
rect 9128 19110 9180 19116
rect 8956 17649 8984 19110
rect 8942 17640 8998 17649
rect 8942 17575 8998 17584
rect 9036 16992 9088 16998
rect 9036 16934 9088 16940
rect 9048 16697 9076 16934
rect 9034 16688 9090 16697
rect 9034 16623 9090 16632
rect 8668 15904 8720 15910
rect 8668 15846 8720 15852
rect 8944 15904 8996 15910
rect 8944 15846 8996 15852
rect 8680 15201 8708 15846
rect 8666 15192 8722 15201
rect 8666 15127 8722 15136
rect 8484 14476 8536 14482
rect 8484 14418 8536 14424
rect 8668 14476 8720 14482
rect 8668 14418 8720 14424
rect 8496 13870 8524 14418
rect 8680 14113 8708 14418
rect 8760 14408 8812 14414
rect 8760 14350 8812 14356
rect 8666 14104 8722 14113
rect 8666 14039 8668 14048
rect 8720 14039 8722 14048
rect 8668 14010 8720 14016
rect 8772 13938 8800 14350
rect 8956 13977 8984 15846
rect 9140 15706 9168 19110
rect 9402 18184 9458 18193
rect 9402 18119 9458 18128
rect 9416 18086 9444 18119
rect 9404 18080 9456 18086
rect 9404 18022 9456 18028
rect 9404 17808 9456 17814
rect 9404 17750 9456 17756
rect 9416 16794 9444 17750
rect 9496 16992 9548 16998
rect 9496 16934 9548 16940
rect 9404 16788 9456 16794
rect 9404 16730 9456 16736
rect 9508 16017 9536 16934
rect 9494 16008 9550 16017
rect 9494 15943 9550 15952
rect 9128 15700 9180 15706
rect 9128 15642 9180 15648
rect 9036 15496 9088 15502
rect 9036 15438 9088 15444
rect 9048 15162 9076 15438
rect 9036 15156 9088 15162
rect 9036 15098 9088 15104
rect 9140 15026 9168 15642
rect 9692 15042 9720 19264
rect 9864 17808 9916 17814
rect 9864 17750 9916 17756
rect 9876 16998 9904 17750
rect 9956 17128 10008 17134
rect 9956 17070 10008 17076
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9864 16992 9916 16998
rect 9864 16934 9916 16940
rect 9784 16726 9812 16934
rect 9772 16720 9824 16726
rect 9772 16662 9824 16668
rect 9784 15978 9812 16662
rect 9876 16658 9904 16934
rect 9864 16652 9916 16658
rect 9864 16594 9916 16600
rect 9968 16454 9996 17070
rect 9956 16448 10008 16454
rect 9956 16390 10008 16396
rect 9772 15972 9824 15978
rect 9772 15914 9824 15920
rect 9968 15706 9996 16390
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 9770 15600 9826 15609
rect 9770 15535 9772 15544
rect 9824 15535 9826 15544
rect 9772 15506 9824 15512
rect 9784 15162 9812 15506
rect 9772 15156 9824 15162
rect 9772 15098 9824 15104
rect 10060 15065 10088 19654
rect 10980 19174 11008 19858
rect 11888 19848 11940 19854
rect 11888 19790 11940 19796
rect 11336 19780 11388 19786
rect 11336 19722 11388 19728
rect 10140 19168 10192 19174
rect 10140 19110 10192 19116
rect 10968 19168 11020 19174
rect 11020 19128 11192 19156
rect 10968 19110 11020 19116
rect 10152 17241 10180 19110
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10508 18896 10560 18902
rect 10506 18864 10508 18873
rect 10784 18896 10836 18902
rect 10560 18864 10562 18873
rect 10784 18838 10836 18844
rect 10874 18864 10930 18873
rect 10506 18799 10562 18808
rect 10324 18760 10376 18766
rect 10324 18702 10376 18708
rect 10336 18465 10364 18702
rect 10692 18624 10744 18630
rect 10692 18566 10744 18572
rect 10322 18456 10378 18465
rect 10322 18391 10378 18400
rect 10336 18290 10364 18391
rect 10324 18284 10376 18290
rect 10324 18226 10376 18232
rect 10704 18154 10732 18566
rect 10692 18148 10744 18154
rect 10692 18090 10744 18096
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10138 17232 10194 17241
rect 10138 17167 10194 17176
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10140 16652 10192 16658
rect 10140 16594 10192 16600
rect 10152 16182 10180 16594
rect 10704 16250 10732 18090
rect 10796 18086 10824 18838
rect 10874 18799 10930 18808
rect 10784 18080 10836 18086
rect 10784 18022 10836 18028
rect 10796 17338 10824 18022
rect 10888 17882 10916 18799
rect 11060 18284 11112 18290
rect 11060 18226 11112 18232
rect 10968 18216 11020 18222
rect 10968 18158 11020 18164
rect 10876 17876 10928 17882
rect 10876 17818 10928 17824
rect 10980 17814 11008 18158
rect 11072 17882 11100 18226
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 10968 17808 11020 17814
rect 10968 17750 11020 17756
rect 10784 17332 10836 17338
rect 10784 17274 10836 17280
rect 10968 16788 11020 16794
rect 10968 16730 11020 16736
rect 10980 16697 11008 16730
rect 10966 16688 11022 16697
rect 10966 16623 11022 16632
rect 10968 16448 11020 16454
rect 11020 16396 11100 16402
rect 10968 16390 11100 16396
rect 10980 16374 11100 16390
rect 10692 16244 10744 16250
rect 10692 16186 10744 16192
rect 10140 16176 10192 16182
rect 10140 16118 10192 16124
rect 10152 15473 10180 16118
rect 10968 16108 11020 16114
rect 11072 16096 11100 16374
rect 11020 16068 11100 16096
rect 10968 16050 11020 16056
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10874 15736 10930 15745
rect 10874 15671 10930 15680
rect 10138 15464 10194 15473
rect 10138 15399 10194 15408
rect 10046 15056 10102 15065
rect 9128 15020 9180 15026
rect 9692 15014 9996 15042
rect 9128 14962 9180 14968
rect 9128 14884 9180 14890
rect 9048 14844 9128 14872
rect 9048 14657 9076 14844
rect 9128 14826 9180 14832
rect 9772 14816 9824 14822
rect 9772 14758 9824 14764
rect 9034 14648 9090 14657
rect 9034 14583 9036 14592
rect 9088 14583 9090 14592
rect 9036 14554 9088 14560
rect 8942 13968 8998 13977
rect 8760 13932 8812 13938
rect 8942 13903 8998 13912
rect 9312 13932 9364 13938
rect 8760 13874 8812 13880
rect 9312 13874 9364 13880
rect 8484 13864 8536 13870
rect 8484 13806 8536 13812
rect 8574 13832 8630 13841
rect 8496 13297 8524 13806
rect 8574 13767 8630 13776
rect 8588 13394 8616 13767
rect 9324 13530 9352 13874
rect 9312 13524 9364 13530
rect 9312 13466 9364 13472
rect 8576 13388 8628 13394
rect 8576 13330 8628 13336
rect 8482 13288 8538 13297
rect 8482 13223 8538 13232
rect 8588 12986 8616 13330
rect 9784 13326 9812 14758
rect 9864 13728 9916 13734
rect 9864 13670 9916 13676
rect 9876 13462 9904 13670
rect 9864 13456 9916 13462
rect 9864 13398 9916 13404
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 8576 12980 8628 12986
rect 8576 12922 8628 12928
rect 9036 12708 9088 12714
rect 9036 12650 9088 12656
rect 8852 12368 8904 12374
rect 8852 12310 8904 12316
rect 8484 12164 8536 12170
rect 8484 12106 8536 12112
rect 8496 11558 8524 12106
rect 8864 11898 8892 12310
rect 9048 12170 9076 12650
rect 9508 12442 9536 13262
rect 9876 12986 9904 13398
rect 9864 12980 9916 12986
rect 9864 12922 9916 12928
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9496 12436 9548 12442
rect 9496 12378 9548 12384
rect 9036 12164 9088 12170
rect 9036 12106 9088 12112
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 8852 11892 8904 11898
rect 8852 11834 8904 11840
rect 8758 11656 8814 11665
rect 8758 11591 8814 11600
rect 8484 11552 8536 11558
rect 8484 11494 8536 11500
rect 8496 9178 8524 11494
rect 8772 11286 8800 11591
rect 8760 11280 8812 11286
rect 8760 11222 8812 11228
rect 8576 11212 8628 11218
rect 8576 11154 8628 11160
rect 8588 10810 8616 11154
rect 8576 10804 8628 10810
rect 8576 10746 8628 10752
rect 8864 10577 8892 11834
rect 9600 11762 9628 12038
rect 9692 11898 9720 12582
rect 9968 12356 9996 15014
rect 10046 14991 10102 15000
rect 10784 14952 10836 14958
rect 10784 14894 10836 14900
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10048 14544 10100 14550
rect 10796 14521 10824 14894
rect 10048 14486 10100 14492
rect 10782 14512 10838 14521
rect 10060 13870 10088 14486
rect 10782 14447 10838 14456
rect 10048 13864 10100 13870
rect 10048 13806 10100 13812
rect 10692 13728 10744 13734
rect 10046 13696 10102 13705
rect 10692 13670 10744 13676
rect 10046 13631 10102 13640
rect 10060 13326 10088 13631
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10048 13320 10100 13326
rect 10048 13262 10100 13268
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 9876 12328 9996 12356
rect 10140 12368 10192 12374
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9588 11756 9640 11762
rect 9640 11716 9812 11744
rect 9588 11698 9640 11704
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9404 11008 9456 11014
rect 9404 10950 9456 10956
rect 9218 10704 9274 10713
rect 9218 10639 9274 10648
rect 9232 10606 9260 10639
rect 9416 10606 9444 10950
rect 9692 10690 9720 11086
rect 9600 10674 9720 10690
rect 9588 10668 9720 10674
rect 9640 10662 9720 10668
rect 9588 10610 9640 10616
rect 9220 10600 9272 10606
rect 8850 10568 8906 10577
rect 9220 10542 9272 10548
rect 9404 10600 9456 10606
rect 9404 10542 9456 10548
rect 8850 10503 8906 10512
rect 9232 10266 9260 10542
rect 9600 10266 9628 10610
rect 9784 10538 9812 11716
rect 9772 10532 9824 10538
rect 9772 10474 9824 10480
rect 9220 10260 9272 10266
rect 9220 10202 9272 10208
rect 9588 10260 9640 10266
rect 9588 10202 9640 10208
rect 9772 10056 9824 10062
rect 9772 9998 9824 10004
rect 9220 9988 9272 9994
rect 9220 9930 9272 9936
rect 9232 9586 9260 9930
rect 9678 9616 9734 9625
rect 9220 9580 9272 9586
rect 9678 9551 9680 9560
rect 9220 9522 9272 9528
rect 9732 9551 9734 9560
rect 9680 9522 9732 9528
rect 9312 9444 9364 9450
rect 9312 9386 9364 9392
rect 8576 9376 8628 9382
rect 8576 9318 8628 9324
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 8484 9036 8536 9042
rect 8484 8978 8536 8984
rect 8496 8634 8524 8978
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 8496 8537 8524 8570
rect 8482 8528 8538 8537
rect 8482 8463 8538 8472
rect 8588 7546 8616 9318
rect 9324 9178 9352 9386
rect 9312 9172 9364 9178
rect 9312 9114 9364 9120
rect 9128 8832 9180 8838
rect 9128 8774 9180 8780
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9140 8430 9168 8774
rect 9600 8514 9628 8774
rect 9784 8514 9812 9998
rect 9600 8486 9812 8514
rect 9128 8424 9180 8430
rect 9128 8366 9180 8372
rect 9588 8424 9640 8430
rect 9640 8372 9720 8378
rect 9588 8366 9720 8372
rect 9220 8356 9272 8362
rect 9600 8350 9720 8366
rect 9220 8298 9272 8304
rect 9232 8090 9260 8298
rect 9692 8090 9720 8350
rect 9220 8084 9272 8090
rect 9220 8026 9272 8032
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 8392 7336 8444 7342
rect 8392 7278 8444 7284
rect 8116 6928 8168 6934
rect 8116 6870 8168 6876
rect 8300 6860 8352 6866
rect 8300 6802 8352 6808
rect 8024 6724 8076 6730
rect 8024 6666 8076 6672
rect 8312 6458 8340 6802
rect 9586 6760 9642 6769
rect 9784 6730 9812 8486
rect 9876 7342 9904 12328
rect 10140 12310 10192 12316
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 9968 11082 9996 12174
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 10060 11286 10088 11494
rect 10152 11354 10180 12310
rect 10600 12300 10652 12306
rect 10600 12242 10652 12248
rect 10612 12073 10640 12242
rect 10598 12064 10654 12073
rect 10598 11999 10654 12008
rect 10612 11898 10640 11999
rect 10600 11892 10652 11898
rect 10600 11834 10652 11840
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 10048 11280 10100 11286
rect 10048 11222 10100 11228
rect 9956 11076 10008 11082
rect 9956 11018 10008 11024
rect 9968 8566 9996 11018
rect 10060 10470 10088 11222
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 10060 9450 10088 10406
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10140 10192 10192 10198
rect 10140 10134 10192 10140
rect 10152 9722 10180 10134
rect 10704 9761 10732 13670
rect 10796 11393 10824 14447
rect 10782 11384 10838 11393
rect 10782 11319 10838 11328
rect 10796 10606 10824 11319
rect 10888 10713 10916 15671
rect 11072 15094 11100 16068
rect 11060 15088 11112 15094
rect 11060 15030 11112 15036
rect 10966 14512 11022 14521
rect 10966 14447 11022 14456
rect 10980 14249 11008 14447
rect 10966 14240 11022 14249
rect 10966 14175 11022 14184
rect 11164 13530 11192 19128
rect 11244 18420 11296 18426
rect 11244 18362 11296 18368
rect 11152 13524 11204 13530
rect 11152 13466 11204 13472
rect 11152 13388 11204 13394
rect 11152 13330 11204 13336
rect 11058 13288 11114 13297
rect 11058 13223 11114 13232
rect 10874 10704 10930 10713
rect 10874 10639 10930 10648
rect 10784 10600 10836 10606
rect 10784 10542 10836 10548
rect 10690 9752 10746 9761
rect 10140 9716 10192 9722
rect 10796 9722 10824 10542
rect 10888 9761 10916 10639
rect 10968 9920 11020 9926
rect 10968 9862 11020 9868
rect 10874 9752 10930 9761
rect 10690 9687 10746 9696
rect 10784 9716 10836 9722
rect 10140 9658 10192 9664
rect 10874 9687 10930 9696
rect 10784 9658 10836 9664
rect 10048 9444 10100 9450
rect 10048 9386 10100 9392
rect 10060 9110 10088 9386
rect 10048 9104 10100 9110
rect 10048 9046 10100 9052
rect 10060 8634 10088 9046
rect 10152 8945 10180 9658
rect 10690 9616 10746 9625
rect 10690 9551 10746 9560
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10138 8936 10194 8945
rect 10138 8871 10194 8880
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 9956 8560 10008 8566
rect 9956 8502 10008 8508
rect 10060 8362 10088 8570
rect 10152 8430 10180 8871
rect 10140 8424 10192 8430
rect 10140 8366 10192 8372
rect 10048 8356 10100 8362
rect 10048 8298 10100 8304
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10322 7984 10378 7993
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 10048 7948 10100 7954
rect 10322 7919 10378 7928
rect 10048 7890 10100 7896
rect 9968 7546 9996 7890
rect 9956 7540 10008 7546
rect 9956 7482 10008 7488
rect 10060 7478 10088 7890
rect 10336 7546 10364 7919
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 10048 7472 10100 7478
rect 10048 7414 10100 7420
rect 9864 7336 9916 7342
rect 9864 7278 9916 7284
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10322 6896 10378 6905
rect 10322 6831 10324 6840
rect 10376 6831 10378 6840
rect 10324 6802 10376 6808
rect 9586 6695 9588 6704
rect 9640 6695 9642 6704
rect 9772 6724 9824 6730
rect 9588 6666 9640 6672
rect 9772 6666 9824 6672
rect 10336 6458 10364 6802
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10704 4214 10732 9551
rect 10796 9518 10824 9658
rect 10784 9512 10836 9518
rect 10784 9454 10836 9460
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10796 8974 10824 9318
rect 10784 8968 10836 8974
rect 10784 8910 10836 8916
rect 10796 8634 10824 8910
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 10888 8022 10916 9687
rect 10980 9518 11008 9862
rect 10968 9512 11020 9518
rect 10968 9454 11020 9460
rect 10876 8016 10928 8022
rect 10876 7958 10928 7964
rect 10980 7954 11008 9454
rect 10968 7948 11020 7954
rect 10968 7890 11020 7896
rect 11072 7546 11100 13223
rect 11164 11801 11192 13330
rect 11256 13326 11284 18362
rect 11348 15706 11376 19722
rect 11428 19712 11480 19718
rect 11428 19654 11480 19660
rect 11440 19310 11468 19654
rect 11428 19304 11480 19310
rect 11428 19246 11480 19252
rect 11428 19168 11480 19174
rect 11428 19110 11480 19116
rect 11440 15881 11468 19110
rect 11900 18630 11928 19790
rect 11992 19514 12020 19926
rect 11980 19508 12032 19514
rect 11980 19450 12032 19456
rect 11888 18624 11940 18630
rect 11794 18592 11850 18601
rect 11888 18566 11940 18572
rect 11794 18527 11850 18536
rect 11808 18193 11836 18527
rect 11978 18456 12034 18465
rect 11978 18391 12034 18400
rect 11992 18193 12020 18391
rect 11794 18184 11850 18193
rect 11794 18119 11850 18128
rect 11978 18184 12034 18193
rect 11978 18119 12034 18128
rect 11520 18080 11572 18086
rect 11520 18022 11572 18028
rect 11532 17338 11560 18022
rect 11808 17814 11836 18119
rect 11796 17808 11848 17814
rect 11796 17750 11848 17756
rect 11808 17338 11836 17750
rect 11520 17332 11572 17338
rect 11520 17274 11572 17280
rect 11796 17332 11848 17338
rect 11796 17274 11848 17280
rect 11612 16992 11664 16998
rect 11612 16934 11664 16940
rect 11520 16584 11572 16590
rect 11520 16526 11572 16532
rect 11532 16250 11560 16526
rect 11520 16244 11572 16250
rect 11520 16186 11572 16192
rect 11426 15872 11482 15881
rect 11426 15807 11482 15816
rect 11336 15700 11388 15706
rect 11336 15642 11388 15648
rect 11440 15502 11468 15807
rect 11532 15706 11560 16186
rect 11520 15700 11572 15706
rect 11520 15642 11572 15648
rect 11428 15496 11480 15502
rect 11428 15438 11480 15444
rect 11440 14618 11468 15438
rect 11428 14612 11480 14618
rect 11428 14554 11480 14560
rect 11334 13968 11390 13977
rect 11334 13903 11390 13912
rect 11348 13870 11376 13903
rect 11336 13864 11388 13870
rect 11440 13841 11468 14554
rect 11520 14000 11572 14006
rect 11520 13942 11572 13948
rect 11336 13806 11388 13812
rect 11426 13832 11482 13841
rect 11348 13394 11376 13806
rect 11426 13767 11482 13776
rect 11428 13728 11480 13734
rect 11428 13670 11480 13676
rect 11336 13388 11388 13394
rect 11336 13330 11388 13336
rect 11244 13320 11296 13326
rect 11440 13274 11468 13670
rect 11244 13262 11296 13268
rect 11348 13246 11468 13274
rect 11150 11792 11206 11801
rect 11150 11727 11206 11736
rect 11348 11694 11376 13246
rect 11532 13025 11560 13942
rect 11518 13016 11574 13025
rect 11518 12951 11574 12960
rect 11532 12850 11560 12951
rect 11520 12844 11572 12850
rect 11520 12786 11572 12792
rect 11428 12776 11480 12782
rect 11428 12718 11480 12724
rect 11440 12170 11468 12718
rect 11624 12714 11652 16934
rect 11794 16280 11850 16289
rect 11794 16215 11850 16224
rect 11808 15609 11836 16215
rect 11794 15600 11850 15609
rect 11704 15564 11756 15570
rect 11794 15535 11850 15544
rect 11704 15506 11756 15512
rect 11716 15162 11744 15506
rect 11704 15156 11756 15162
rect 11704 15098 11756 15104
rect 11716 14958 11744 15098
rect 11704 14952 11756 14958
rect 11704 14894 11756 14900
rect 11704 14816 11756 14822
rect 11704 14758 11756 14764
rect 11716 13734 11744 14758
rect 11980 14340 12032 14346
rect 11980 14282 12032 14288
rect 11704 13728 11756 13734
rect 11704 13670 11756 13676
rect 11796 13728 11848 13734
rect 11796 13670 11848 13676
rect 11808 13462 11836 13670
rect 11796 13456 11848 13462
rect 11794 13424 11796 13433
rect 11848 13424 11850 13433
rect 11794 13359 11850 13368
rect 11888 13388 11940 13394
rect 11808 13333 11836 13359
rect 11888 13330 11940 13336
rect 11796 13252 11848 13258
rect 11796 13194 11848 13200
rect 11612 12708 11664 12714
rect 11612 12650 11664 12656
rect 11428 12164 11480 12170
rect 11428 12106 11480 12112
rect 11336 11688 11388 11694
rect 11336 11630 11388 11636
rect 11152 11008 11204 11014
rect 11152 10950 11204 10956
rect 11164 10606 11192 10950
rect 11152 10600 11204 10606
rect 11152 10542 11204 10548
rect 11164 8537 11192 10542
rect 11244 9512 11296 9518
rect 11242 9480 11244 9489
rect 11296 9480 11298 9489
rect 11242 9415 11298 9424
rect 11348 9330 11376 11630
rect 11624 11218 11652 12650
rect 11808 12646 11836 13194
rect 11900 12782 11928 13330
rect 11888 12776 11940 12782
rect 11888 12718 11940 12724
rect 11796 12640 11848 12646
rect 11796 12582 11848 12588
rect 11808 12424 11836 12582
rect 11716 12396 11836 12424
rect 11716 11558 11744 12396
rect 11992 11898 12020 14282
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11980 11552 12032 11558
rect 11980 11494 12032 11500
rect 11992 11354 12020 11494
rect 11980 11348 12032 11354
rect 11980 11290 12032 11296
rect 11992 11218 12020 11290
rect 11612 11212 11664 11218
rect 11612 11154 11664 11160
rect 11980 11212 12032 11218
rect 11980 11154 12032 11160
rect 11518 11112 11574 11121
rect 11518 11047 11574 11056
rect 11256 9302 11376 9330
rect 11150 8528 11206 8537
rect 11150 8463 11206 8472
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 10692 4208 10744 4214
rect 10692 4150 10744 4156
rect 10876 4208 10928 4214
rect 10876 4150 10928 4156
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10888 610 10916 4150
rect 11256 4049 11284 9302
rect 11336 8424 11388 8430
rect 11336 8366 11388 8372
rect 11348 6866 11376 8366
rect 11532 6866 11560 11047
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 11900 10266 11928 10950
rect 11992 10742 12020 11154
rect 11980 10736 12032 10742
rect 11980 10678 12032 10684
rect 11992 10470 12020 10678
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 11888 10260 11940 10266
rect 11888 10202 11940 10208
rect 11900 9654 11928 10202
rect 11992 9994 12020 10406
rect 11980 9988 12032 9994
rect 11980 9930 12032 9936
rect 11888 9648 11940 9654
rect 11888 9590 11940 9596
rect 11980 9172 12032 9178
rect 11980 9114 12032 9120
rect 11992 8906 12020 9114
rect 11980 8900 12032 8906
rect 11980 8842 12032 8848
rect 11888 8832 11940 8838
rect 11888 8774 11940 8780
rect 11796 8560 11848 8566
rect 11796 8502 11848 8508
rect 11336 6860 11388 6866
rect 11336 6802 11388 6808
rect 11520 6860 11572 6866
rect 11520 6802 11572 6808
rect 11348 6458 11376 6802
rect 11336 6452 11388 6458
rect 11336 6394 11388 6400
rect 11242 4040 11298 4049
rect 11242 3975 11298 3984
rect 11808 3505 11836 8502
rect 11900 7954 11928 8774
rect 11992 7954 12020 8842
rect 12084 8634 12112 24806
rect 13096 24806 13216 24834
rect 12990 23896 13046 23905
rect 12990 23831 12992 23840
rect 13044 23831 13046 23840
rect 12992 23802 13044 23808
rect 12440 23656 12492 23662
rect 12360 23604 12440 23610
rect 12360 23598 12492 23604
rect 12360 23582 12480 23598
rect 12256 19304 12308 19310
rect 12256 19246 12308 19252
rect 12268 18850 12296 19246
rect 12360 18970 12388 23582
rect 12532 20936 12584 20942
rect 12532 20878 12584 20884
rect 12438 19408 12494 19417
rect 12438 19343 12494 19352
rect 12452 19310 12480 19343
rect 12440 19304 12492 19310
rect 12440 19246 12492 19252
rect 12544 19174 12572 20878
rect 12716 20392 12768 20398
rect 12716 20334 12768 20340
rect 12728 19718 12756 20334
rect 12716 19712 12768 19718
rect 12716 19654 12768 19660
rect 12532 19168 12584 19174
rect 12532 19110 12584 19116
rect 12348 18964 12400 18970
rect 12348 18906 12400 18912
rect 12164 18828 12216 18834
rect 12268 18822 12572 18850
rect 12164 18770 12216 18776
rect 12176 18222 12204 18770
rect 12348 18624 12400 18630
rect 12440 18624 12492 18630
rect 12348 18566 12400 18572
rect 12438 18592 12440 18601
rect 12492 18592 12494 18601
rect 12164 18216 12216 18222
rect 12164 18158 12216 18164
rect 12176 17542 12204 18158
rect 12256 18080 12308 18086
rect 12256 18022 12308 18028
rect 12268 17746 12296 18022
rect 12360 17882 12388 18566
rect 12438 18527 12494 18536
rect 12544 18442 12572 18822
rect 12452 18414 12572 18442
rect 12348 17876 12400 17882
rect 12348 17818 12400 17824
rect 12256 17740 12308 17746
rect 12256 17682 12308 17688
rect 12164 17536 12216 17542
rect 12164 17478 12216 17484
rect 12176 17202 12204 17478
rect 12164 17196 12216 17202
rect 12164 17138 12216 17144
rect 12268 16998 12296 17682
rect 12348 17264 12400 17270
rect 12348 17206 12400 17212
rect 12360 16998 12388 17206
rect 12256 16992 12308 16998
rect 12256 16934 12308 16940
rect 12348 16992 12400 16998
rect 12348 16934 12400 16940
rect 12164 15904 12216 15910
rect 12164 15846 12216 15852
rect 12176 14346 12204 15846
rect 12348 14476 12400 14482
rect 12348 14418 12400 14424
rect 12164 14340 12216 14346
rect 12164 14282 12216 14288
rect 12176 13802 12204 14282
rect 12164 13796 12216 13802
rect 12164 13738 12216 13744
rect 12360 13734 12388 14418
rect 12452 13938 12480 18414
rect 12728 18086 12756 19654
rect 13096 19281 13124 24806
rect 14660 23905 14688 27520
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14646 23896 14702 23905
rect 14956 23888 15252 23908
rect 16040 23866 16068 27520
rect 17420 24449 17448 27520
rect 16394 24440 16450 24449
rect 16394 24375 16396 24384
rect 16448 24375 16450 24384
rect 17406 24440 17462 24449
rect 17406 24375 17462 24384
rect 16396 24346 16448 24352
rect 17406 24304 17462 24313
rect 16120 24268 16172 24274
rect 17406 24239 17408 24248
rect 16120 24210 16172 24216
rect 17460 24239 17462 24248
rect 17408 24210 17460 24216
rect 14646 23831 14702 23840
rect 16028 23860 16080 23866
rect 16028 23802 16080 23808
rect 15292 23656 15344 23662
rect 15292 23598 15344 23604
rect 15304 23322 15332 23598
rect 16132 23526 16160 24210
rect 16488 24064 16540 24070
rect 16488 24006 16540 24012
rect 16500 23633 16528 24006
rect 17420 23866 17448 24210
rect 17500 24064 17552 24070
rect 17500 24006 17552 24012
rect 17408 23860 17460 23866
rect 17408 23802 17460 23808
rect 16486 23624 16542 23633
rect 17130 23624 17186 23633
rect 16486 23559 16488 23568
rect 16540 23559 16542 23568
rect 16948 23588 17000 23594
rect 16488 23530 16540 23536
rect 17130 23559 17132 23568
rect 16948 23530 17000 23536
rect 17184 23559 17186 23568
rect 17132 23530 17184 23536
rect 16120 23520 16172 23526
rect 16120 23462 16172 23468
rect 15292 23316 15344 23322
rect 15292 23258 15344 23264
rect 15476 23180 15528 23186
rect 15476 23122 15528 23128
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 15488 22234 15516 23122
rect 15660 22568 15712 22574
rect 15660 22510 15712 22516
rect 15568 22500 15620 22506
rect 15568 22442 15620 22448
rect 15476 22228 15528 22234
rect 15476 22170 15528 22176
rect 15580 22166 15608 22442
rect 13268 22160 13320 22166
rect 13188 22108 13268 22114
rect 13188 22102 13320 22108
rect 15568 22160 15620 22166
rect 15568 22102 15620 22108
rect 13188 22086 13308 22102
rect 13188 21690 13216 22086
rect 13268 22024 13320 22030
rect 13268 21966 13320 21972
rect 13912 22024 13964 22030
rect 13912 21966 13964 21972
rect 13176 21684 13228 21690
rect 13176 21626 13228 21632
rect 13188 20602 13216 21626
rect 13280 21146 13308 21966
rect 13924 21554 13952 21966
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 13912 21548 13964 21554
rect 13912 21490 13964 21496
rect 15672 21418 15700 22510
rect 15752 22432 15804 22438
rect 15752 22374 15804 22380
rect 15764 22137 15792 22374
rect 16132 22273 16160 23462
rect 16580 23248 16632 23254
rect 16580 23190 16632 23196
rect 16592 22506 16620 23190
rect 16672 23112 16724 23118
rect 16672 23054 16724 23060
rect 16580 22500 16632 22506
rect 16580 22442 16632 22448
rect 16684 22386 16712 23054
rect 16764 22636 16816 22642
rect 16764 22578 16816 22584
rect 16316 22358 16712 22386
rect 16118 22264 16174 22273
rect 16118 22199 16174 22208
rect 15936 22160 15988 22166
rect 15750 22128 15806 22137
rect 15936 22102 15988 22108
rect 15750 22063 15806 22072
rect 13636 21412 13688 21418
rect 13636 21354 13688 21360
rect 13728 21412 13780 21418
rect 13728 21354 13780 21360
rect 15660 21412 15712 21418
rect 15660 21354 15712 21360
rect 13648 21146 13676 21354
rect 13268 21140 13320 21146
rect 13268 21082 13320 21088
rect 13636 21140 13688 21146
rect 13636 21082 13688 21088
rect 13740 20754 13768 21354
rect 14832 20800 14884 20806
rect 13740 20726 13860 20754
rect 14832 20742 14884 20748
rect 13176 20596 13228 20602
rect 13176 20538 13228 20544
rect 13188 20058 13216 20538
rect 13452 20256 13504 20262
rect 13452 20198 13504 20204
rect 13176 20052 13228 20058
rect 13176 19994 13228 20000
rect 13082 19272 13138 19281
rect 13082 19207 13138 19216
rect 12900 18624 12952 18630
rect 12900 18566 12952 18572
rect 12912 18222 12940 18566
rect 12900 18216 12952 18222
rect 12900 18158 12952 18164
rect 12716 18080 12768 18086
rect 12716 18022 12768 18028
rect 12912 17746 12940 18158
rect 12900 17740 12952 17746
rect 12900 17682 12952 17688
rect 12530 17232 12586 17241
rect 12530 17167 12586 17176
rect 12544 17066 12572 17167
rect 12532 17060 12584 17066
rect 12532 17002 12584 17008
rect 12624 17060 12676 17066
rect 12624 17002 12676 17008
rect 12544 16726 12572 17002
rect 12636 16794 12664 17002
rect 12624 16788 12676 16794
rect 12624 16730 12676 16736
rect 12532 16720 12584 16726
rect 12532 16662 12584 16668
rect 12912 16658 12940 17682
rect 12900 16652 12952 16658
rect 12900 16594 12952 16600
rect 12530 15192 12586 15201
rect 12530 15127 12586 15136
rect 12544 14618 12572 15127
rect 12808 15020 12860 15026
rect 12808 14962 12860 14968
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 12820 14550 12848 14962
rect 12808 14544 12860 14550
rect 12808 14486 12860 14492
rect 12440 13932 12492 13938
rect 12440 13874 12492 13880
rect 12820 13870 12848 14486
rect 12808 13864 12860 13870
rect 12808 13806 12860 13812
rect 12348 13728 12400 13734
rect 12348 13670 12400 13676
rect 12624 13184 12676 13190
rect 12624 13126 12676 13132
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 12176 11830 12204 12242
rect 12256 12232 12308 12238
rect 12254 12200 12256 12209
rect 12308 12200 12310 12209
rect 12254 12135 12310 12144
rect 12256 12096 12308 12102
rect 12256 12038 12308 12044
rect 12164 11824 12216 11830
rect 12164 11766 12216 11772
rect 12268 11626 12296 12038
rect 12256 11620 12308 11626
rect 12176 11580 12256 11608
rect 12176 11286 12204 11580
rect 12256 11562 12308 11568
rect 12348 11552 12400 11558
rect 12348 11494 12400 11500
rect 12164 11280 12216 11286
rect 12164 11222 12216 11228
rect 12256 11280 12308 11286
rect 12256 11222 12308 11228
rect 12176 10538 12204 11222
rect 12268 11150 12296 11222
rect 12256 11144 12308 11150
rect 12256 11086 12308 11092
rect 12164 10532 12216 10538
rect 12164 10474 12216 10480
rect 12176 9926 12204 10474
rect 12164 9920 12216 9926
rect 12164 9862 12216 9868
rect 12072 8628 12124 8634
rect 12072 8570 12124 8576
rect 12176 8090 12204 9862
rect 12164 8084 12216 8090
rect 12164 8026 12216 8032
rect 11888 7948 11940 7954
rect 11888 7890 11940 7896
rect 11980 7948 12032 7954
rect 11980 7890 12032 7896
rect 11900 7002 11928 7890
rect 11992 7546 12020 7890
rect 11980 7540 12032 7546
rect 11980 7482 12032 7488
rect 12360 7478 12388 11494
rect 12532 11144 12584 11150
rect 12532 11086 12584 11092
rect 12440 10124 12492 10130
rect 12440 10066 12492 10072
rect 12452 8974 12480 10066
rect 12440 8968 12492 8974
rect 12440 8910 12492 8916
rect 12452 8498 12480 8910
rect 12440 8492 12492 8498
rect 12440 8434 12492 8440
rect 12348 7472 12400 7478
rect 12348 7414 12400 7420
rect 12544 7342 12572 11086
rect 12636 9586 12664 13126
rect 12912 12918 12940 16594
rect 13096 14362 13124 19207
rect 13464 19174 13492 20198
rect 13832 20058 13860 20726
rect 14844 20398 14872 20742
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 15764 20602 15792 22063
rect 15948 21690 15976 22102
rect 15936 21684 15988 21690
rect 15936 21626 15988 21632
rect 15752 20596 15804 20602
rect 15752 20538 15804 20544
rect 14832 20392 14884 20398
rect 14832 20334 14884 20340
rect 13820 20052 13872 20058
rect 13820 19994 13872 20000
rect 14740 19712 14792 19718
rect 14740 19654 14792 19660
rect 14752 19310 14780 19654
rect 14844 19446 14872 20334
rect 15568 20324 15620 20330
rect 15568 20266 15620 20272
rect 15580 19990 15608 20266
rect 15568 19984 15620 19990
rect 15568 19926 15620 19932
rect 15476 19848 15528 19854
rect 15476 19790 15528 19796
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 14832 19440 14884 19446
rect 14832 19382 14884 19388
rect 14188 19304 14240 19310
rect 14188 19246 14240 19252
rect 14740 19304 14792 19310
rect 14740 19246 14792 19252
rect 13636 19236 13688 19242
rect 13636 19178 13688 19184
rect 13912 19236 13964 19242
rect 13912 19178 13964 19184
rect 13452 19168 13504 19174
rect 13452 19110 13504 19116
rect 13544 18828 13596 18834
rect 13544 18770 13596 18776
rect 13176 18284 13228 18290
rect 13176 18226 13228 18232
rect 13188 16658 13216 18226
rect 13556 18086 13584 18770
rect 13544 18080 13596 18086
rect 13544 18022 13596 18028
rect 13544 17740 13596 17746
rect 13544 17682 13596 17688
rect 13556 16998 13584 17682
rect 13268 16992 13320 16998
rect 13268 16934 13320 16940
rect 13544 16992 13596 16998
rect 13544 16934 13596 16940
rect 13176 16652 13228 16658
rect 13176 16594 13228 16600
rect 13188 15366 13216 16594
rect 13280 15570 13308 16934
rect 13360 15972 13412 15978
rect 13360 15914 13412 15920
rect 13372 15570 13400 15914
rect 13268 15564 13320 15570
rect 13268 15506 13320 15512
rect 13360 15564 13412 15570
rect 13360 15506 13412 15512
rect 13544 15564 13596 15570
rect 13544 15506 13596 15512
rect 13176 15360 13228 15366
rect 13176 15302 13228 15308
rect 13188 15026 13216 15302
rect 13280 15094 13308 15506
rect 13268 15088 13320 15094
rect 13268 15030 13320 15036
rect 13176 15020 13228 15026
rect 13176 14962 13228 14968
rect 13280 14482 13308 15030
rect 13372 14618 13400 15506
rect 13556 14822 13584 15506
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 13360 14612 13412 14618
rect 13360 14554 13412 14560
rect 13268 14476 13320 14482
rect 13268 14418 13320 14424
rect 13096 14334 13308 14362
rect 13280 13410 13308 14334
rect 13372 14006 13400 14554
rect 13360 14000 13412 14006
rect 13360 13942 13412 13948
rect 13372 13530 13400 13942
rect 13360 13524 13412 13530
rect 13360 13466 13412 13472
rect 13176 13388 13228 13394
rect 13280 13382 13400 13410
rect 13176 13330 13228 13336
rect 12900 12912 12952 12918
rect 12900 12854 12952 12860
rect 12808 12776 12860 12782
rect 12728 12724 12808 12730
rect 12728 12718 12860 12724
rect 12728 12714 12848 12718
rect 12716 12708 12848 12714
rect 12768 12702 12848 12708
rect 12716 12650 12768 12656
rect 12808 12640 12860 12646
rect 12808 12582 12860 12588
rect 12820 12170 12848 12582
rect 12808 12164 12860 12170
rect 12808 12106 12860 12112
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 12728 11354 12756 11834
rect 12820 11762 12848 12106
rect 12808 11756 12860 11762
rect 12808 11698 12860 11704
rect 12716 11348 12768 11354
rect 12716 11290 12768 11296
rect 12820 11014 12848 11698
rect 12912 11150 12940 12854
rect 13188 12102 13216 13330
rect 13268 13252 13320 13258
rect 13268 13194 13320 13200
rect 13280 12714 13308 13194
rect 13268 12708 13320 12714
rect 13268 12650 13320 12656
rect 13372 12594 13400 13382
rect 13452 13388 13504 13394
rect 13452 13330 13504 13336
rect 13464 12646 13492 13330
rect 13280 12566 13400 12594
rect 13452 12640 13504 12646
rect 13452 12582 13504 12588
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 12900 11144 12952 11150
rect 12900 11086 12952 11092
rect 12808 11008 12860 11014
rect 12808 10950 12860 10956
rect 12820 10674 12848 10950
rect 12912 10810 12940 11086
rect 12900 10804 12952 10810
rect 12900 10746 12952 10752
rect 12808 10668 12860 10674
rect 12808 10610 12860 10616
rect 12912 10266 12940 10746
rect 12900 10260 12952 10266
rect 12900 10202 12952 10208
rect 13084 9648 13136 9654
rect 13084 9590 13136 9596
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 12728 9178 12756 9454
rect 12716 9172 12768 9178
rect 12716 9114 12768 9120
rect 12624 8968 12676 8974
rect 12624 8910 12676 8916
rect 12636 8634 12664 8910
rect 13096 8838 13124 9590
rect 13084 8832 13136 8838
rect 13084 8774 13136 8780
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12622 8528 12678 8537
rect 12622 8463 12678 8472
rect 12636 7546 12664 8463
rect 13096 8430 13124 8774
rect 13084 8424 13136 8430
rect 13084 8366 13136 8372
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 12532 7336 12584 7342
rect 12532 7278 12584 7284
rect 11888 6996 11940 7002
rect 11888 6938 11940 6944
rect 13096 3505 13124 8366
rect 13280 6905 13308 12566
rect 13358 12200 13414 12209
rect 13358 12135 13414 12144
rect 13372 9042 13400 12135
rect 13544 12096 13596 12102
rect 13544 12038 13596 12044
rect 13556 11218 13584 12038
rect 13648 11642 13676 19178
rect 13924 18834 13952 19178
rect 14200 19174 14228 19246
rect 14188 19168 14240 19174
rect 14188 19110 14240 19116
rect 13912 18828 13964 18834
rect 13912 18770 13964 18776
rect 13820 18760 13872 18766
rect 13820 18702 13872 18708
rect 13832 17746 13860 18702
rect 13924 18426 13952 18770
rect 13912 18420 13964 18426
rect 13912 18362 13964 18368
rect 13924 18154 13952 18362
rect 14200 18222 14228 19110
rect 14752 18834 14780 19246
rect 14740 18828 14792 18834
rect 14740 18770 14792 18776
rect 15488 18630 15516 19790
rect 15580 19514 15608 19926
rect 15568 19508 15620 19514
rect 15568 19450 15620 19456
rect 16028 19508 16080 19514
rect 16028 19450 16080 19456
rect 15752 19304 15804 19310
rect 15752 19246 15804 19252
rect 14740 18624 14792 18630
rect 14740 18566 14792 18572
rect 15476 18624 15528 18630
rect 15476 18566 15528 18572
rect 14752 18222 14780 18566
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 15488 18358 15516 18566
rect 15476 18352 15528 18358
rect 15476 18294 15528 18300
rect 14188 18216 14240 18222
rect 14188 18158 14240 18164
rect 14740 18216 14792 18222
rect 14740 18158 14792 18164
rect 15568 18216 15620 18222
rect 15568 18158 15620 18164
rect 13912 18148 13964 18154
rect 13912 18090 13964 18096
rect 13924 17882 13952 18090
rect 13912 17876 13964 17882
rect 13912 17818 13964 17824
rect 13820 17740 13872 17746
rect 13820 17682 13872 17688
rect 13924 17338 13952 17818
rect 13912 17332 13964 17338
rect 13912 17274 13964 17280
rect 13820 17060 13872 17066
rect 13820 17002 13872 17008
rect 13832 16658 13860 17002
rect 14200 16946 14228 18158
rect 14464 18080 14516 18086
rect 14464 18022 14516 18028
rect 14280 17536 14332 17542
rect 14280 17478 14332 17484
rect 14292 17066 14320 17478
rect 14476 17134 14504 18022
rect 15580 17542 15608 18158
rect 15660 17672 15712 17678
rect 15660 17614 15712 17620
rect 15568 17536 15620 17542
rect 15568 17478 15620 17484
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 14464 17128 14516 17134
rect 15200 17128 15252 17134
rect 14464 17070 14516 17076
rect 14844 17076 15200 17082
rect 14844 17070 15252 17076
rect 14280 17060 14332 17066
rect 14280 17002 14332 17008
rect 14370 16960 14426 16969
rect 14200 16918 14320 16946
rect 13820 16652 13872 16658
rect 13820 16594 13872 16600
rect 13728 16516 13780 16522
rect 13728 16458 13780 16464
rect 13740 16046 13768 16458
rect 13728 16040 13780 16046
rect 14188 16040 14240 16046
rect 13728 15982 13780 15988
rect 13818 16008 13874 16017
rect 14188 15982 14240 15988
rect 13818 15943 13874 15952
rect 13832 15502 13860 15943
rect 14096 15904 14148 15910
rect 14200 15881 14228 15982
rect 14096 15846 14148 15852
rect 14186 15872 14242 15881
rect 13820 15496 13872 15502
rect 13820 15438 13872 15444
rect 13912 14816 13964 14822
rect 13912 14758 13964 14764
rect 13924 14482 13952 14758
rect 13912 14476 13964 14482
rect 13912 14418 13964 14424
rect 13924 13870 13952 14418
rect 14004 14340 14056 14346
rect 14004 14282 14056 14288
rect 14016 14074 14044 14282
rect 14004 14068 14056 14074
rect 14004 14010 14056 14016
rect 13912 13864 13964 13870
rect 13912 13806 13964 13812
rect 14016 13530 14044 14010
rect 14004 13524 14056 13530
rect 14004 13466 14056 13472
rect 14004 13320 14056 13326
rect 14004 13262 14056 13268
rect 13910 12336 13966 12345
rect 13910 12271 13912 12280
rect 13964 12271 13966 12280
rect 13912 12242 13964 12248
rect 13648 11614 13768 11642
rect 13636 11552 13688 11558
rect 13636 11494 13688 11500
rect 13544 11212 13596 11218
rect 13544 11154 13596 11160
rect 13556 10713 13584 11154
rect 13542 10704 13598 10713
rect 13542 10639 13598 10648
rect 13452 10124 13504 10130
rect 13452 10066 13504 10072
rect 13464 9654 13492 10066
rect 13556 10062 13584 10639
rect 13648 10470 13676 11494
rect 13740 10577 13768 11614
rect 13924 11393 13952 12242
rect 13910 11384 13966 11393
rect 13910 11319 13912 11328
rect 13964 11319 13966 11328
rect 13912 11290 13964 11296
rect 13820 11280 13872 11286
rect 13924 11259 13952 11290
rect 13820 11222 13872 11228
rect 13832 10810 13860 11222
rect 13912 11144 13964 11150
rect 13912 11086 13964 11092
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 13820 10600 13872 10606
rect 13726 10568 13782 10577
rect 13820 10542 13872 10548
rect 13726 10503 13782 10512
rect 13636 10464 13688 10470
rect 13636 10406 13688 10412
rect 13726 10432 13782 10441
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13452 9648 13504 9654
rect 13452 9590 13504 9596
rect 13360 9036 13412 9042
rect 13360 8978 13412 8984
rect 13372 8634 13400 8978
rect 13464 8974 13492 9590
rect 13452 8968 13504 8974
rect 13452 8910 13504 8916
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 13556 7954 13584 9998
rect 13648 9722 13676 10406
rect 13726 10367 13782 10376
rect 13740 10266 13768 10367
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 13636 9716 13688 9722
rect 13636 9658 13688 9664
rect 13648 9625 13676 9658
rect 13832 9654 13860 10542
rect 13820 9648 13872 9654
rect 13634 9616 13690 9625
rect 13820 9590 13872 9596
rect 13634 9551 13690 9560
rect 13544 7948 13596 7954
rect 13544 7890 13596 7896
rect 13556 7546 13584 7890
rect 13544 7540 13596 7546
rect 13544 7482 13596 7488
rect 13924 7342 13952 11086
rect 14016 10130 14044 13262
rect 14108 10266 14136 15846
rect 14186 15807 14242 15816
rect 14200 15706 14228 15807
rect 14188 15700 14240 15706
rect 14188 15642 14240 15648
rect 14292 14396 14320 16918
rect 14370 16895 14426 16904
rect 14384 16726 14412 16895
rect 14476 16810 14504 17070
rect 14844 17054 15240 17070
rect 14476 16782 14596 16810
rect 14372 16720 14424 16726
rect 14372 16662 14424 16668
rect 14464 16652 14516 16658
rect 14464 16594 14516 16600
rect 14370 16008 14426 16017
rect 14370 15943 14426 15952
rect 14384 14550 14412 15943
rect 14476 15162 14504 16594
rect 14464 15156 14516 15162
rect 14464 15098 14516 15104
rect 14476 14618 14504 15098
rect 14464 14612 14516 14618
rect 14464 14554 14516 14560
rect 14372 14544 14424 14550
rect 14372 14486 14424 14492
rect 14292 14368 14412 14396
rect 14280 13184 14332 13190
rect 14280 13126 14332 13132
rect 14292 12850 14320 13126
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 14292 10606 14320 12786
rect 14384 12617 14412 14368
rect 14476 13870 14504 14554
rect 14464 13864 14516 13870
rect 14464 13806 14516 13812
rect 14370 12608 14426 12617
rect 14370 12543 14426 12552
rect 14568 11665 14596 16782
rect 14844 16114 14872 17054
rect 15672 16998 15700 17614
rect 15764 17338 15792 19246
rect 16040 19242 16068 19450
rect 16028 19236 16080 19242
rect 16028 19178 16080 19184
rect 16040 18902 16068 19178
rect 16028 18896 16080 18902
rect 16028 18838 16080 18844
rect 16040 18426 16068 18838
rect 16028 18420 16080 18426
rect 16028 18362 16080 18368
rect 16040 17814 16068 18362
rect 16028 17808 16080 17814
rect 16132 17785 16160 22199
rect 16316 22030 16344 22358
rect 16488 22160 16540 22166
rect 16488 22102 16540 22108
rect 16500 22030 16528 22102
rect 16304 22024 16356 22030
rect 16302 21992 16304 22001
rect 16488 22024 16540 22030
rect 16356 21992 16358 22001
rect 16212 21956 16264 21962
rect 16488 21966 16540 21972
rect 16302 21927 16358 21936
rect 16212 21898 16264 21904
rect 16224 21554 16252 21898
rect 16212 21548 16264 21554
rect 16212 21490 16264 21496
rect 16212 21412 16264 21418
rect 16212 21354 16264 21360
rect 16224 20058 16252 21354
rect 16316 20874 16344 21927
rect 16396 21616 16448 21622
rect 16394 21584 16396 21593
rect 16448 21584 16450 21593
rect 16500 21554 16528 21966
rect 16776 21962 16804 22578
rect 16764 21956 16816 21962
rect 16764 21898 16816 21904
rect 16394 21519 16450 21528
rect 16488 21548 16540 21554
rect 16488 21490 16540 21496
rect 16396 21344 16448 21350
rect 16396 21286 16448 21292
rect 16408 21078 16436 21286
rect 16396 21072 16448 21078
rect 16396 21014 16448 21020
rect 16304 20868 16356 20874
rect 16304 20810 16356 20816
rect 16408 20602 16436 21014
rect 16580 20936 16632 20942
rect 16580 20878 16632 20884
rect 16592 20602 16620 20878
rect 16776 20874 16804 21898
rect 16764 20868 16816 20874
rect 16764 20810 16816 20816
rect 16396 20596 16448 20602
rect 16396 20538 16448 20544
rect 16580 20596 16632 20602
rect 16580 20538 16632 20544
rect 16672 20392 16724 20398
rect 16672 20334 16724 20340
rect 16684 20233 16712 20334
rect 16670 20224 16726 20233
rect 16670 20159 16726 20168
rect 16212 20052 16264 20058
rect 16212 19994 16264 20000
rect 16672 19712 16724 19718
rect 16672 19654 16724 19660
rect 16684 19378 16712 19654
rect 16672 19372 16724 19378
rect 16672 19314 16724 19320
rect 16488 18760 16540 18766
rect 16488 18702 16540 18708
rect 16500 18426 16528 18702
rect 16488 18420 16540 18426
rect 16488 18362 16540 18368
rect 16580 18216 16632 18222
rect 16580 18158 16632 18164
rect 16028 17750 16080 17756
rect 16118 17776 16174 17785
rect 15844 17536 15896 17542
rect 15844 17478 15896 17484
rect 15752 17332 15804 17338
rect 15752 17274 15804 17280
rect 15856 17134 15884 17478
rect 16040 17338 16068 17750
rect 16118 17711 16174 17720
rect 16028 17332 16080 17338
rect 16028 17274 16080 17280
rect 15844 17128 15896 17134
rect 15844 17070 15896 17076
rect 16040 17048 16068 17274
rect 16120 17060 16172 17066
rect 16040 17020 16120 17048
rect 15660 16992 15712 16998
rect 15660 16934 15712 16940
rect 15384 16788 15436 16794
rect 15384 16730 15436 16736
rect 15290 16688 15346 16697
rect 15290 16623 15292 16632
rect 15344 16623 15346 16632
rect 15292 16594 15344 16600
rect 15292 16516 15344 16522
rect 15292 16458 15344 16464
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15304 16250 15332 16458
rect 15292 16244 15344 16250
rect 15292 16186 15344 16192
rect 15396 16182 15424 16730
rect 15476 16448 15528 16454
rect 15476 16390 15528 16396
rect 15384 16176 15436 16182
rect 15384 16118 15436 16124
rect 14832 16108 14884 16114
rect 14832 16050 14884 16056
rect 15488 15745 15516 16390
rect 15672 15910 15700 16934
rect 15750 16824 15806 16833
rect 16040 16794 16068 17020
rect 16120 17002 16172 17008
rect 16592 16833 16620 18158
rect 16856 18080 16908 18086
rect 16856 18022 16908 18028
rect 16578 16824 16634 16833
rect 15750 16759 15806 16768
rect 16028 16788 16080 16794
rect 15764 16046 15792 16759
rect 16578 16759 16634 16768
rect 16028 16730 16080 16736
rect 16396 16652 16448 16658
rect 16396 16594 16448 16600
rect 16408 16266 16436 16594
rect 16408 16250 16620 16266
rect 16408 16244 16632 16250
rect 16408 16238 16580 16244
rect 16580 16186 16632 16192
rect 15752 16040 15804 16046
rect 15752 15982 15804 15988
rect 16396 16040 16448 16046
rect 16396 15982 16448 15988
rect 15660 15904 15712 15910
rect 15660 15846 15712 15852
rect 15474 15736 15530 15745
rect 15764 15706 15792 15982
rect 15474 15671 15530 15680
rect 15752 15700 15804 15706
rect 15752 15642 15804 15648
rect 14738 15464 14794 15473
rect 14738 15399 14794 15408
rect 14648 15088 14700 15094
rect 14648 15030 14700 15036
rect 14660 14550 14688 15030
rect 14648 14544 14700 14550
rect 14648 14486 14700 14492
rect 14660 13802 14688 14486
rect 14752 13938 14780 15399
rect 15292 15360 15344 15366
rect 15292 15302 15344 15308
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15304 14074 15332 15302
rect 15764 15162 15792 15642
rect 16408 15570 16436 15982
rect 16592 15570 16620 16186
rect 16028 15564 16080 15570
rect 16028 15506 16080 15512
rect 16120 15564 16172 15570
rect 16120 15506 16172 15512
rect 16396 15564 16448 15570
rect 16396 15506 16448 15512
rect 16580 15564 16632 15570
rect 16580 15506 16632 15512
rect 15752 15156 15804 15162
rect 15752 15098 15804 15104
rect 16040 14958 16068 15506
rect 16028 14952 16080 14958
rect 16028 14894 16080 14900
rect 15936 14544 15988 14550
rect 16040 14532 16068 14894
rect 15988 14504 16068 14532
rect 15936 14486 15988 14492
rect 15844 14476 15896 14482
rect 15844 14418 15896 14424
rect 15292 14068 15344 14074
rect 15292 14010 15344 14016
rect 14740 13932 14792 13938
rect 14740 13874 14792 13880
rect 14648 13796 14700 13802
rect 14648 13738 14700 13744
rect 14660 13530 14688 13738
rect 15856 13530 15884 14418
rect 16040 14006 16068 14504
rect 16132 14074 16160 15506
rect 16488 15496 16540 15502
rect 16486 15464 16488 15473
rect 16540 15464 16542 15473
rect 16486 15399 16542 15408
rect 16488 14476 16540 14482
rect 16592 14464 16620 15506
rect 16672 14952 16724 14958
rect 16672 14894 16724 14900
rect 16540 14436 16620 14464
rect 16488 14418 16540 14424
rect 16684 14414 16712 14894
rect 16868 14521 16896 18022
rect 16960 17882 16988 23530
rect 17316 23044 17368 23050
rect 17316 22986 17368 22992
rect 17328 22234 17356 22986
rect 17512 22778 17540 24006
rect 18800 23866 18828 27520
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 18788 23860 18840 23866
rect 18788 23802 18840 23808
rect 18696 23520 18748 23526
rect 18696 23462 18748 23468
rect 18708 23225 18736 23462
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 18694 23216 18750 23225
rect 18604 23180 18656 23186
rect 18694 23151 18750 23160
rect 18604 23122 18656 23128
rect 18616 22817 18644 23122
rect 18602 22808 18658 22817
rect 17500 22772 17552 22778
rect 18602 22743 18604 22752
rect 17500 22714 17552 22720
rect 18656 22743 18658 22752
rect 18604 22714 18656 22720
rect 17868 22432 17920 22438
rect 17868 22374 17920 22380
rect 17316 22228 17368 22234
rect 17316 22170 17368 22176
rect 17880 22030 17908 22374
rect 17960 22160 18012 22166
rect 17960 22102 18012 22108
rect 18050 22128 18106 22137
rect 17868 22024 17920 22030
rect 17868 21966 17920 21972
rect 17880 21690 17908 21966
rect 17868 21684 17920 21690
rect 17868 21626 17920 21632
rect 17972 21350 18000 22102
rect 18050 22063 18106 22072
rect 18064 21486 18092 22063
rect 18144 22024 18196 22030
rect 18142 21992 18144 22001
rect 18196 21992 18198 22001
rect 18142 21927 18198 21936
rect 18052 21480 18104 21486
rect 18052 21422 18104 21428
rect 17960 21344 18012 21350
rect 17960 21286 18012 21292
rect 17776 21004 17828 21010
rect 17776 20946 17828 20952
rect 17788 20058 17816 20946
rect 17960 20800 18012 20806
rect 17960 20742 18012 20748
rect 17972 20602 18000 20742
rect 17960 20596 18012 20602
rect 17960 20538 18012 20544
rect 17972 20262 18000 20538
rect 18604 20460 18656 20466
rect 18604 20402 18656 20408
rect 17960 20256 18012 20262
rect 17960 20198 18012 20204
rect 17776 20052 17828 20058
rect 17776 19994 17828 20000
rect 17788 19514 17816 19994
rect 18616 19990 18644 20402
rect 18604 19984 18656 19990
rect 18604 19926 18656 19932
rect 18420 19848 18472 19854
rect 18420 19790 18472 19796
rect 17776 19508 17828 19514
rect 17776 19450 17828 19456
rect 17590 19408 17646 19417
rect 18432 19378 18460 19790
rect 17590 19343 17646 19352
rect 18420 19372 18472 19378
rect 17500 18964 17552 18970
rect 17500 18906 17552 18912
rect 17512 17882 17540 18906
rect 17604 18902 17632 19343
rect 18420 19314 18472 19320
rect 18144 19236 18196 19242
rect 18144 19178 18196 19184
rect 18328 19236 18380 19242
rect 18328 19178 18380 19184
rect 18156 18970 18184 19178
rect 18144 18964 18196 18970
rect 18144 18906 18196 18912
rect 17592 18896 17644 18902
rect 17592 18838 17644 18844
rect 18052 18896 18104 18902
rect 18340 18850 18368 19178
rect 18432 18902 18460 19314
rect 18104 18844 18368 18850
rect 18052 18838 18368 18844
rect 18420 18896 18472 18902
rect 18420 18838 18472 18844
rect 18064 18822 18368 18838
rect 18420 18216 18472 18222
rect 18420 18158 18472 18164
rect 18052 18080 18104 18086
rect 18052 18022 18104 18028
rect 16948 17876 17000 17882
rect 16948 17818 17000 17824
rect 17500 17876 17552 17882
rect 17500 17818 17552 17824
rect 17776 17740 17828 17746
rect 17776 17682 17828 17688
rect 17222 17232 17278 17241
rect 17222 17167 17278 17176
rect 16948 16992 17000 16998
rect 16948 16934 17000 16940
rect 16960 16726 16988 16934
rect 16948 16720 17000 16726
rect 16948 16662 17000 16668
rect 16960 15706 16988 16662
rect 17236 16590 17264 17167
rect 17788 16998 17816 17682
rect 17960 17536 18012 17542
rect 17960 17478 18012 17484
rect 17972 17066 18000 17478
rect 17960 17060 18012 17066
rect 17960 17002 18012 17008
rect 17776 16992 17828 16998
rect 17774 16960 17776 16969
rect 17828 16960 17830 16969
rect 17774 16895 17830 16904
rect 17224 16584 17276 16590
rect 17130 16552 17186 16561
rect 17224 16526 17276 16532
rect 17130 16487 17132 16496
rect 17184 16487 17186 16496
rect 17132 16458 17184 16464
rect 17236 16250 17264 16526
rect 17224 16244 17276 16250
rect 17224 16186 17276 16192
rect 18064 15978 18092 18022
rect 18432 17542 18460 18158
rect 18420 17536 18472 17542
rect 18420 17478 18472 17484
rect 18328 17060 18380 17066
rect 18328 17002 18380 17008
rect 18236 16992 18288 16998
rect 18236 16934 18288 16940
rect 17500 15972 17552 15978
rect 17500 15914 17552 15920
rect 18052 15972 18104 15978
rect 18052 15914 18104 15920
rect 17512 15706 17540 15914
rect 16948 15700 17000 15706
rect 16948 15642 17000 15648
rect 17500 15700 17552 15706
rect 17500 15642 17552 15648
rect 17512 15162 17540 15642
rect 17868 15564 17920 15570
rect 17868 15506 17920 15512
rect 17880 15178 17908 15506
rect 17880 15162 18000 15178
rect 17500 15156 17552 15162
rect 17880 15156 18012 15162
rect 17880 15150 17960 15156
rect 17500 15098 17552 15104
rect 17960 15098 18012 15104
rect 17130 14920 17186 14929
rect 17130 14855 17132 14864
rect 17184 14855 17186 14864
rect 17132 14826 17184 14832
rect 16854 14512 16910 14521
rect 17408 14476 17460 14482
rect 16910 14456 16988 14464
rect 16854 14447 16988 14456
rect 16868 14436 16988 14447
rect 16672 14408 16724 14414
rect 16868 14387 16896 14436
rect 16672 14350 16724 14356
rect 16762 14376 16818 14385
rect 16762 14311 16764 14320
rect 16816 14311 16818 14320
rect 16764 14282 16816 14288
rect 16120 14068 16172 14074
rect 16120 14010 16172 14016
rect 16028 14000 16080 14006
rect 16028 13942 16080 13948
rect 16776 13938 16804 14282
rect 16764 13932 16816 13938
rect 16764 13874 16816 13880
rect 16580 13796 16632 13802
rect 16580 13738 16632 13744
rect 14648 13524 14700 13530
rect 14648 13466 14700 13472
rect 15844 13524 15896 13530
rect 15844 13466 15896 13472
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 14740 13184 14792 13190
rect 14740 13126 14792 13132
rect 14752 12782 14780 13126
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15304 12986 15332 13330
rect 16592 13190 16620 13738
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 16580 13184 16632 13190
rect 16580 13126 16632 13132
rect 16592 13025 16620 13126
rect 16578 13016 16634 13025
rect 15292 12980 15344 12986
rect 16578 12951 16580 12960
rect 15292 12922 15344 12928
rect 16632 12951 16634 12960
rect 16580 12922 16632 12928
rect 14740 12776 14792 12782
rect 14740 12718 14792 12724
rect 14752 12306 14780 12718
rect 14740 12300 14792 12306
rect 14740 12242 14792 12248
rect 14752 12084 14780 12242
rect 14832 12096 14884 12102
rect 14752 12056 14832 12084
rect 14832 12038 14884 12044
rect 14648 11688 14700 11694
rect 14554 11656 14610 11665
rect 14844 11676 14872 12038
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 14924 11688 14976 11694
rect 14844 11656 14924 11676
rect 14976 11656 14978 11665
rect 14844 11648 14922 11656
rect 14648 11630 14700 11636
rect 14554 11591 14610 11600
rect 14370 11248 14426 11257
rect 14370 11183 14426 11192
rect 14280 10600 14332 10606
rect 14280 10542 14332 10548
rect 14096 10260 14148 10266
rect 14096 10202 14148 10208
rect 14292 10130 14320 10542
rect 14004 10124 14056 10130
rect 14004 10066 14056 10072
rect 14280 10124 14332 10130
rect 14280 10066 14332 10072
rect 14004 9988 14056 9994
rect 14004 9930 14056 9936
rect 13912 7336 13964 7342
rect 13912 7278 13964 7284
rect 13266 6896 13322 6905
rect 13266 6831 13322 6840
rect 11794 3496 11850 3505
rect 11794 3431 11850 3440
rect 13082 3496 13138 3505
rect 13082 3431 13138 3440
rect 14016 626 14044 9930
rect 14186 9480 14242 9489
rect 14186 9415 14242 9424
rect 14200 9382 14228 9415
rect 14188 9376 14240 9382
rect 14188 9318 14240 9324
rect 14384 8022 14412 11183
rect 14372 8016 14424 8022
rect 14372 7958 14424 7964
rect 14568 7954 14596 11591
rect 14660 11354 14688 11630
rect 14922 11591 14978 11600
rect 14648 11348 14700 11354
rect 14648 11290 14700 11296
rect 14660 9761 14688 11290
rect 15304 11257 15332 12922
rect 15752 12912 15804 12918
rect 15752 12854 15804 12860
rect 15764 12714 15792 12854
rect 15752 12708 15804 12714
rect 15752 12650 15804 12656
rect 15764 12374 15792 12650
rect 15752 12368 15804 12374
rect 15752 12310 15804 12316
rect 15764 11626 15792 12310
rect 16776 12102 16804 13262
rect 16764 12096 16816 12102
rect 16764 12038 16816 12044
rect 15936 11688 15988 11694
rect 15936 11630 15988 11636
rect 15752 11620 15804 11626
rect 15752 11562 15804 11568
rect 15948 11354 15976 11630
rect 15936 11348 15988 11354
rect 15936 11290 15988 11296
rect 16028 11280 16080 11286
rect 15290 11248 15346 11257
rect 16028 11222 16080 11228
rect 15290 11183 15346 11192
rect 15842 11112 15898 11121
rect 15842 11047 15898 11056
rect 15856 11014 15884 11047
rect 15292 11008 15344 11014
rect 15292 10950 15344 10956
rect 15844 11008 15896 11014
rect 15844 10950 15896 10956
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 14832 10532 14884 10538
rect 14832 10474 14884 10480
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14646 9752 14702 9761
rect 14646 9687 14702 9696
rect 14660 8498 14688 9687
rect 14752 9042 14780 10406
rect 14844 9042 14872 10474
rect 15304 10470 15332 10950
rect 15658 10840 15714 10849
rect 15658 10775 15660 10784
rect 15712 10775 15714 10784
rect 15660 10746 15712 10752
rect 15856 10674 15884 10950
rect 15844 10668 15896 10674
rect 15844 10610 15896 10616
rect 16040 10577 16068 11222
rect 16212 11144 16264 11150
rect 16212 11086 16264 11092
rect 16224 10674 16252 11086
rect 16396 11076 16448 11082
rect 16396 11018 16448 11024
rect 16212 10668 16264 10674
rect 16212 10610 16264 10616
rect 16026 10568 16082 10577
rect 16026 10503 16082 10512
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 15752 10192 15804 10198
rect 15566 10160 15622 10169
rect 15752 10134 15804 10140
rect 15566 10095 15622 10104
rect 15292 10056 15344 10062
rect 15292 9998 15344 10004
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15304 9722 15332 9998
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 15108 9512 15160 9518
rect 15108 9454 15160 9460
rect 15120 9110 15148 9454
rect 15108 9104 15160 9110
rect 15108 9046 15160 9052
rect 14740 9036 14792 9042
rect 14740 8978 14792 8984
rect 14832 9036 14884 9042
rect 14832 8978 14884 8984
rect 14752 8838 14780 8978
rect 14740 8832 14792 8838
rect 14740 8774 14792 8780
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14752 8362 14780 8774
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15304 8498 15332 9658
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 14740 8356 14792 8362
rect 14740 8298 14792 8304
rect 14752 8265 14780 8298
rect 14738 8256 14794 8265
rect 14738 8191 14794 8200
rect 14752 8090 14780 8191
rect 15580 8090 15608 10095
rect 15764 9450 15792 10134
rect 15752 9444 15804 9450
rect 15752 9386 15804 9392
rect 15764 9110 15792 9386
rect 16040 9178 16068 10503
rect 16224 10062 16252 10610
rect 16304 10532 16356 10538
rect 16304 10474 16356 10480
rect 16316 10266 16344 10474
rect 16304 10260 16356 10266
rect 16304 10202 16356 10208
rect 16212 10056 16264 10062
rect 16212 9998 16264 10004
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 16028 9172 16080 9178
rect 16028 9114 16080 9120
rect 15752 9104 15804 9110
rect 15752 9046 15804 9052
rect 15764 8634 15792 9046
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 16132 8362 16160 9318
rect 16224 8566 16252 9998
rect 16316 9761 16344 10202
rect 16408 9874 16436 11018
rect 16776 10826 16804 12038
rect 16856 11212 16908 11218
rect 16856 11154 16908 11160
rect 16684 10798 16804 10826
rect 16580 9920 16632 9926
rect 16408 9868 16580 9874
rect 16408 9862 16632 9868
rect 16408 9846 16620 9862
rect 16302 9752 16358 9761
rect 16302 9687 16358 9696
rect 16396 9444 16448 9450
rect 16396 9386 16448 9392
rect 16212 8560 16264 8566
rect 16212 8502 16264 8508
rect 16408 8498 16436 9386
rect 16396 8492 16448 8498
rect 16396 8434 16448 8440
rect 16120 8356 16172 8362
rect 16120 8298 16172 8304
rect 16132 8090 16160 8298
rect 16408 8090 16436 8434
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 15568 8084 15620 8090
rect 15568 8026 15620 8032
rect 16120 8084 16172 8090
rect 16120 8026 16172 8032
rect 16396 8084 16448 8090
rect 16396 8026 16448 8032
rect 14556 7948 14608 7954
rect 14556 7890 14608 7896
rect 14568 7478 14596 7890
rect 14752 7546 14780 8026
rect 16132 7993 16160 8026
rect 16118 7984 16174 7993
rect 15384 7948 15436 7954
rect 16118 7919 16174 7928
rect 15384 7890 15436 7896
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14740 7540 14792 7546
rect 14740 7482 14792 7488
rect 14556 7472 14608 7478
rect 14556 7414 14608 7420
rect 15396 7342 15424 7890
rect 15384 7336 15436 7342
rect 15382 7304 15384 7313
rect 15436 7304 15438 7313
rect 15382 7239 15438 7248
rect 16500 6769 16528 9846
rect 16580 9036 16632 9042
rect 16580 8978 16632 8984
rect 16592 8634 16620 8978
rect 16580 8628 16632 8634
rect 16580 8570 16632 8576
rect 16684 8129 16712 10798
rect 16868 10470 16896 11154
rect 16960 10810 16988 14436
rect 17408 14418 17460 14424
rect 17592 14476 17644 14482
rect 17592 14418 17644 14424
rect 17316 13796 17368 13802
rect 17316 13738 17368 13744
rect 17328 13462 17356 13738
rect 17420 13734 17448 14418
rect 17604 14006 17632 14418
rect 17776 14408 17828 14414
rect 17774 14376 17776 14385
rect 17828 14376 17830 14385
rect 17774 14311 17830 14320
rect 17592 14000 17644 14006
rect 17592 13942 17644 13948
rect 17408 13728 17460 13734
rect 17408 13670 17460 13676
rect 17592 13728 17644 13734
rect 17592 13670 17644 13676
rect 17132 13456 17184 13462
rect 17132 13398 17184 13404
rect 17316 13456 17368 13462
rect 17316 13398 17368 13404
rect 17144 12986 17172 13398
rect 17604 13258 17632 13670
rect 18052 13456 18104 13462
rect 18052 13398 18104 13404
rect 17592 13252 17644 13258
rect 17592 13194 17644 13200
rect 17132 12980 17184 12986
rect 17132 12922 17184 12928
rect 17316 12980 17368 12986
rect 17316 12922 17368 12928
rect 17038 12336 17094 12345
rect 17038 12271 17094 12280
rect 16948 10804 17000 10810
rect 16948 10746 17000 10752
rect 16856 10464 16908 10470
rect 16854 10432 16856 10441
rect 16948 10464 17000 10470
rect 16908 10432 16910 10441
rect 16948 10406 17000 10412
rect 16854 10367 16910 10376
rect 16764 9512 16816 9518
rect 16764 9454 16816 9460
rect 16776 8401 16804 9454
rect 16762 8392 16818 8401
rect 16762 8327 16818 8336
rect 16670 8120 16726 8129
rect 16670 8055 16726 8064
rect 16486 6760 16542 6769
rect 16486 6695 16542 6704
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 7656 604 7708 610
rect 7656 546 7708 552
rect 7840 604 7892 610
rect 7840 546 7892 552
rect 10784 604 10836 610
rect 10784 546 10836 552
rect 10876 604 10928 610
rect 10876 546 10928 552
rect 13924 598 14044 626
rect 7668 480 7696 546
rect 10796 480 10824 546
rect 13924 480 13952 598
rect 16960 480 16988 10406
rect 17052 7954 17080 12271
rect 17328 12073 17356 12922
rect 17498 12608 17554 12617
rect 17498 12543 17554 12552
rect 17408 12368 17460 12374
rect 17408 12310 17460 12316
rect 17314 12064 17370 12073
rect 17314 11999 17370 12008
rect 17328 11898 17356 11999
rect 17316 11892 17368 11898
rect 17316 11834 17368 11840
rect 17420 11830 17448 12310
rect 17408 11824 17460 11830
rect 17406 11792 17408 11801
rect 17460 11792 17462 11801
rect 17406 11727 17462 11736
rect 17420 11626 17448 11727
rect 17408 11620 17460 11626
rect 17408 11562 17460 11568
rect 17512 11354 17540 12543
rect 17500 11348 17552 11354
rect 17500 11290 17552 11296
rect 17604 11218 17632 13194
rect 17960 13184 18012 13190
rect 17960 13126 18012 13132
rect 17408 11212 17460 11218
rect 17408 11154 17460 11160
rect 17592 11212 17644 11218
rect 17592 11154 17644 11160
rect 17420 10470 17448 11154
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 17684 10192 17736 10198
rect 17972 10169 18000 13126
rect 18064 12646 18092 13398
rect 18052 12640 18104 12646
rect 18052 12582 18104 12588
rect 18064 12306 18092 12582
rect 18248 12345 18276 16934
rect 18340 16454 18368 17002
rect 18328 16448 18380 16454
rect 18328 16390 18380 16396
rect 18340 16046 18368 16390
rect 18328 16040 18380 16046
rect 18328 15982 18380 15988
rect 18328 13864 18380 13870
rect 18328 13806 18380 13812
rect 18234 12336 18290 12345
rect 18052 12300 18104 12306
rect 18234 12271 18290 12280
rect 18052 12242 18104 12248
rect 18064 12209 18092 12242
rect 18050 12200 18106 12209
rect 18050 12135 18106 12144
rect 18144 11688 18196 11694
rect 18144 11630 18196 11636
rect 18156 11354 18184 11630
rect 18340 11558 18368 13806
rect 18432 12442 18460 17478
rect 18708 15609 18736 23151
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19432 22092 19484 22098
rect 19432 22034 19484 22040
rect 19444 21690 19472 22034
rect 20180 21962 20208 27520
rect 21546 23624 21602 23633
rect 21546 23559 21602 23568
rect 20904 23180 20956 23186
rect 20904 23122 20956 23128
rect 20916 22545 20944 23122
rect 20902 22536 20958 22545
rect 20902 22471 20904 22480
rect 20956 22471 20958 22480
rect 20904 22442 20956 22448
rect 20168 21956 20220 21962
rect 20168 21898 20220 21904
rect 19432 21684 19484 21690
rect 19432 21626 19484 21632
rect 19444 21146 19472 21626
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19432 21140 19484 21146
rect 19432 21082 19484 21088
rect 19340 21004 19392 21010
rect 19340 20946 19392 20952
rect 18788 20800 18840 20806
rect 18788 20742 18840 20748
rect 18800 20641 18828 20742
rect 18786 20632 18842 20641
rect 18786 20567 18842 20576
rect 18800 20534 18828 20567
rect 18788 20528 18840 20534
rect 18788 20470 18840 20476
rect 19352 20466 19380 20946
rect 20810 20632 20866 20641
rect 20810 20567 20866 20576
rect 19798 20496 19854 20505
rect 19340 20460 19392 20466
rect 20824 20466 20852 20567
rect 19798 20431 19854 20440
rect 20812 20460 20864 20466
rect 19340 20402 19392 20408
rect 19812 20398 19840 20431
rect 20812 20402 20864 20408
rect 19800 20392 19852 20398
rect 19800 20334 19852 20340
rect 20260 20392 20312 20398
rect 20260 20334 20312 20340
rect 19432 20256 19484 20262
rect 19432 20198 19484 20204
rect 19340 19712 19392 19718
rect 19340 19654 19392 19660
rect 19352 19417 19380 19654
rect 19338 19408 19394 19417
rect 19338 19343 19394 19352
rect 19444 19258 19472 20198
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19522 19952 19578 19961
rect 19522 19887 19524 19896
rect 19576 19887 19578 19896
rect 19524 19858 19576 19864
rect 19260 19230 19472 19258
rect 19260 18970 19288 19230
rect 19536 19174 19564 19858
rect 19524 19168 19576 19174
rect 19524 19110 19576 19116
rect 19248 18964 19300 18970
rect 19536 18952 19564 19110
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19248 18906 19300 18912
rect 19444 18924 19564 18952
rect 18880 18828 18932 18834
rect 18880 18770 18932 18776
rect 18892 17882 18920 18770
rect 19340 18760 19392 18766
rect 19340 18702 19392 18708
rect 19064 18216 19116 18222
rect 19064 18158 19116 18164
rect 19248 18216 19300 18222
rect 19248 18158 19300 18164
rect 18972 18080 19024 18086
rect 18972 18022 19024 18028
rect 18880 17876 18932 17882
rect 18880 17818 18932 17824
rect 18694 15600 18750 15609
rect 18694 15535 18750 15544
rect 18696 15360 18748 15366
rect 18696 15302 18748 15308
rect 18602 15056 18658 15065
rect 18602 14991 18604 15000
rect 18656 14991 18658 15000
rect 18604 14962 18656 14968
rect 18616 14618 18644 14962
rect 18708 14890 18736 15302
rect 18696 14884 18748 14890
rect 18696 14826 18748 14832
rect 18604 14612 18656 14618
rect 18604 14554 18656 14560
rect 18892 14113 18920 17818
rect 18984 17814 19012 18022
rect 18972 17808 19024 17814
rect 18972 17750 19024 17756
rect 18984 17338 19012 17750
rect 19076 17678 19104 18158
rect 19064 17672 19116 17678
rect 19062 17640 19064 17649
rect 19116 17640 19118 17649
rect 19062 17575 19118 17584
rect 18972 17332 19024 17338
rect 18972 17274 19024 17280
rect 18984 17202 19012 17274
rect 18972 17196 19024 17202
rect 18972 17138 19024 17144
rect 18984 16726 19012 17138
rect 18972 16720 19024 16726
rect 18972 16662 19024 16668
rect 18972 16584 19024 16590
rect 18972 16526 19024 16532
rect 18984 15638 19012 16526
rect 19260 16114 19288 18158
rect 19248 16108 19300 16114
rect 19248 16050 19300 16056
rect 18972 15632 19024 15638
rect 19352 15586 19380 18702
rect 19444 17785 19472 18924
rect 19524 18828 19576 18834
rect 19524 18770 19576 18776
rect 19536 18426 19564 18770
rect 20076 18624 20128 18630
rect 20076 18566 20128 18572
rect 19524 18420 19576 18426
rect 19524 18362 19576 18368
rect 19430 17776 19486 17785
rect 19430 17711 19486 17720
rect 19432 16720 19484 16726
rect 19536 16697 19564 18362
rect 20088 18222 20116 18566
rect 20076 18216 20128 18222
rect 20076 18158 20128 18164
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 20166 17504 20222 17513
rect 20166 17439 20222 17448
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 20180 16726 20208 17439
rect 20168 16720 20220 16726
rect 19432 16662 19484 16668
rect 19522 16688 19578 16697
rect 19444 16250 19472 16662
rect 20168 16662 20220 16668
rect 19522 16623 19578 16632
rect 19892 16652 19944 16658
rect 19892 16594 19944 16600
rect 19432 16244 19484 16250
rect 19484 16204 19564 16232
rect 19432 16186 19484 16192
rect 19432 16108 19484 16114
rect 19432 16050 19484 16056
rect 18972 15574 19024 15580
rect 19260 15570 19380 15586
rect 19248 15564 19380 15570
rect 19300 15558 19380 15564
rect 19248 15506 19300 15512
rect 18972 15156 19024 15162
rect 18972 15098 19024 15104
rect 18984 14550 19012 15098
rect 19352 14618 19380 15558
rect 19444 15502 19472 16050
rect 19536 15638 19564 16204
rect 19904 15978 19932 16594
rect 19892 15972 19944 15978
rect 19892 15914 19944 15920
rect 19984 15972 20036 15978
rect 19984 15914 20036 15920
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19524 15632 19576 15638
rect 19524 15574 19576 15580
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 19444 15094 19472 15438
rect 19536 15162 19564 15574
rect 19996 15450 20024 15914
rect 20272 15609 20300 20334
rect 20720 18828 20772 18834
rect 20720 18770 20772 18776
rect 20732 18329 20760 18770
rect 20812 18624 20864 18630
rect 20812 18566 20864 18572
rect 20718 18320 20774 18329
rect 20718 18255 20720 18264
rect 20772 18255 20774 18264
rect 20720 18226 20772 18232
rect 20548 18154 20760 18170
rect 20548 18148 20772 18154
rect 20548 18142 20720 18148
rect 20548 17882 20576 18142
rect 20720 18090 20772 18096
rect 20628 18080 20680 18086
rect 20628 18022 20680 18028
rect 20536 17876 20588 17882
rect 20536 17818 20588 17824
rect 20640 17796 20668 18022
rect 20720 17808 20772 17814
rect 20640 17768 20720 17796
rect 20720 17750 20772 17756
rect 20824 17678 20852 18566
rect 20812 17672 20864 17678
rect 20718 17640 20774 17649
rect 20812 17614 20864 17620
rect 20718 17575 20774 17584
rect 20732 17338 20760 17575
rect 20720 17332 20772 17338
rect 20720 17274 20772 17280
rect 20824 17202 20852 17614
rect 20812 17196 20864 17202
rect 20812 17138 20864 17144
rect 20628 16992 20680 16998
rect 20812 16992 20864 16998
rect 20680 16952 20760 16980
rect 20628 16934 20680 16940
rect 20732 15978 20760 16952
rect 20812 16934 20864 16940
rect 20824 16794 20852 16934
rect 20812 16788 20864 16794
rect 20812 16730 20864 16736
rect 20720 15972 20772 15978
rect 20720 15914 20772 15920
rect 20258 15600 20314 15609
rect 20314 15558 20392 15586
rect 20258 15535 20314 15544
rect 19904 15422 20024 15450
rect 20074 15464 20130 15473
rect 19904 15178 19932 15422
rect 20074 15399 20130 15408
rect 19984 15360 20036 15366
rect 19982 15328 19984 15337
rect 20036 15328 20038 15337
rect 19982 15263 20038 15272
rect 19524 15156 19576 15162
rect 19904 15150 20024 15178
rect 19524 15098 19576 15104
rect 19432 15088 19484 15094
rect 19432 15030 19484 15036
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19340 14612 19392 14618
rect 19340 14554 19392 14560
rect 18972 14544 19024 14550
rect 19996 14498 20024 15150
rect 20088 15026 20116 15399
rect 20076 15020 20128 15026
rect 20076 14962 20128 14968
rect 20088 14618 20116 14962
rect 20076 14612 20128 14618
rect 20076 14554 20128 14560
rect 18972 14486 19024 14492
rect 18878 14104 18934 14113
rect 18984 14074 19012 14486
rect 19904 14470 20024 14498
rect 20168 14476 20220 14482
rect 19524 14272 19576 14278
rect 19524 14214 19576 14220
rect 19536 14074 19564 14214
rect 18878 14039 18934 14048
rect 18972 14068 19024 14074
rect 18892 14006 18920 14039
rect 18972 14010 19024 14016
rect 19524 14068 19576 14074
rect 19524 14010 19576 14016
rect 18880 14000 18932 14006
rect 18880 13942 18932 13948
rect 18512 13728 18564 13734
rect 18512 13670 18564 13676
rect 18524 12918 18552 13670
rect 18604 13524 18656 13530
rect 18604 13466 18656 13472
rect 18512 12912 18564 12918
rect 18512 12854 18564 12860
rect 18420 12436 18472 12442
rect 18420 12378 18472 12384
rect 18524 12374 18552 12854
rect 18616 12850 18644 13466
rect 18604 12844 18656 12850
rect 18604 12786 18656 12792
rect 18616 12374 18644 12786
rect 18788 12640 18840 12646
rect 18788 12582 18840 12588
rect 18800 12442 18828 12582
rect 18788 12436 18840 12442
rect 18788 12378 18840 12384
rect 18512 12368 18564 12374
rect 18512 12310 18564 12316
rect 18604 12368 18656 12374
rect 18604 12310 18656 12316
rect 18420 12232 18472 12238
rect 18420 12174 18472 12180
rect 18328 11552 18380 11558
rect 18328 11494 18380 11500
rect 18432 11354 18460 12174
rect 18892 11762 18920 13942
rect 18984 13734 19012 14010
rect 19904 14006 19932 14470
rect 20168 14418 20220 14424
rect 20180 14006 20208 14418
rect 19892 14000 19944 14006
rect 19890 13968 19892 13977
rect 20168 14000 20220 14006
rect 19944 13968 19946 13977
rect 20168 13942 20220 13948
rect 19890 13903 19946 13912
rect 18972 13728 19024 13734
rect 18972 13670 19024 13676
rect 18984 13530 19012 13670
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 18972 13524 19024 13530
rect 18972 13466 19024 13472
rect 19800 13388 19852 13394
rect 19800 13330 19852 13336
rect 19812 12986 19840 13330
rect 19800 12980 19852 12986
rect 19800 12922 19852 12928
rect 19340 12776 19392 12782
rect 19340 12718 19392 12724
rect 19248 12708 19300 12714
rect 19248 12650 19300 12656
rect 19260 12345 19288 12650
rect 19352 12617 19380 12718
rect 20260 12640 20312 12646
rect 19338 12608 19394 12617
rect 20260 12582 20312 12588
rect 19338 12543 19394 12552
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 20272 12442 20300 12582
rect 20260 12436 20312 12442
rect 20180 12396 20260 12424
rect 19246 12336 19302 12345
rect 19246 12271 19302 12280
rect 19892 12300 19944 12306
rect 19892 12242 19944 12248
rect 19904 11898 19932 12242
rect 19892 11892 19944 11898
rect 19892 11834 19944 11840
rect 19432 11824 19484 11830
rect 19432 11766 19484 11772
rect 18880 11756 18932 11762
rect 18880 11698 18932 11704
rect 19062 11656 19118 11665
rect 19062 11591 19118 11600
rect 18144 11348 18196 11354
rect 18144 11290 18196 11296
rect 18420 11348 18472 11354
rect 18420 11290 18472 11296
rect 19076 11218 19104 11591
rect 19340 11552 19392 11558
rect 19340 11494 19392 11500
rect 19352 11286 19380 11494
rect 19340 11280 19392 11286
rect 19246 11248 19302 11257
rect 19064 11212 19116 11218
rect 19340 11222 19392 11228
rect 19246 11183 19302 11192
rect 19064 11154 19116 11160
rect 19076 10606 19104 11154
rect 19260 10674 19288 11183
rect 19340 11144 19392 11150
rect 19340 11086 19392 11092
rect 19352 10810 19380 11086
rect 19444 11014 19472 11766
rect 20076 11620 20128 11626
rect 20076 11562 20128 11568
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 20088 11014 20116 11562
rect 19432 11008 19484 11014
rect 19432 10950 19484 10956
rect 20076 11008 20128 11014
rect 20076 10950 20128 10956
rect 19340 10804 19392 10810
rect 19340 10746 19392 10752
rect 19248 10668 19300 10674
rect 19248 10610 19300 10616
rect 18236 10600 18288 10606
rect 18236 10542 18288 10548
rect 19064 10600 19116 10606
rect 19064 10542 19116 10548
rect 17684 10134 17736 10140
rect 17958 10160 18014 10169
rect 17696 9382 17724 10134
rect 17958 10095 18014 10104
rect 17960 10056 18012 10062
rect 17960 9998 18012 10004
rect 17972 9654 18000 9998
rect 17960 9648 18012 9654
rect 17960 9590 18012 9596
rect 17684 9376 17736 9382
rect 17684 9318 17736 9324
rect 17960 9376 18012 9382
rect 17960 9318 18012 9324
rect 17972 9178 18000 9318
rect 17960 9172 18012 9178
rect 17960 9114 18012 9120
rect 17592 9104 17644 9110
rect 17592 9046 17644 9052
rect 17132 8968 17184 8974
rect 17132 8910 17184 8916
rect 17144 8294 17172 8910
rect 17604 8634 17632 9046
rect 17592 8628 17644 8634
rect 17592 8570 17644 8576
rect 18248 8430 18276 10542
rect 18604 10464 18656 10470
rect 18604 10406 18656 10412
rect 18616 10266 18644 10406
rect 18604 10260 18656 10266
rect 18604 10202 18656 10208
rect 19064 10056 19116 10062
rect 19064 9998 19116 10004
rect 18512 9376 18564 9382
rect 18512 9318 18564 9324
rect 18524 9081 18552 9318
rect 19076 9178 19104 9998
rect 19064 9172 19116 9178
rect 19064 9114 19116 9120
rect 18510 9072 18566 9081
rect 19352 9042 19380 10746
rect 19444 10198 19472 10950
rect 20180 10849 20208 12396
rect 20260 12378 20312 12384
rect 20166 10840 20222 10849
rect 20166 10775 20222 10784
rect 20258 10568 20314 10577
rect 20258 10503 20260 10512
rect 20312 10503 20314 10512
rect 20260 10474 20312 10480
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19432 10192 19484 10198
rect 19432 10134 19484 10140
rect 19444 9450 19472 10134
rect 20074 9616 20130 9625
rect 20074 9551 20130 9560
rect 19524 9512 19576 9518
rect 19524 9454 19576 9460
rect 19432 9444 19484 9450
rect 19432 9386 19484 9392
rect 19444 9110 19472 9386
rect 19432 9104 19484 9110
rect 19432 9046 19484 9052
rect 18510 9007 18566 9016
rect 19340 9036 19392 9042
rect 19340 8978 19392 8984
rect 19352 8634 19380 8978
rect 19536 8906 19564 9454
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19708 9036 19760 9042
rect 19708 8978 19760 8984
rect 19524 8900 19576 8906
rect 19524 8842 19576 8848
rect 19340 8628 19392 8634
rect 19340 8570 19392 8576
rect 19536 8498 19564 8842
rect 19720 8566 19748 8978
rect 19708 8560 19760 8566
rect 19708 8502 19760 8508
rect 19524 8492 19576 8498
rect 19524 8434 19576 8440
rect 18236 8424 18288 8430
rect 18236 8366 18288 8372
rect 18696 8424 18748 8430
rect 18696 8366 18748 8372
rect 17132 8288 17184 8294
rect 17132 8230 17184 8236
rect 17498 8256 17554 8265
rect 17144 8090 17172 8230
rect 17498 8191 17554 8200
rect 17132 8084 17184 8090
rect 17132 8026 17184 8032
rect 17512 7954 17540 8191
rect 18248 8090 18276 8366
rect 18708 8090 18736 8366
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 18236 8084 18288 8090
rect 18236 8026 18288 8032
rect 18696 8084 18748 8090
rect 18696 8026 18748 8032
rect 17040 7948 17092 7954
rect 17040 7890 17092 7896
rect 17500 7948 17552 7954
rect 17500 7890 17552 7896
rect 19892 7948 19944 7954
rect 19892 7890 19944 7896
rect 17052 7546 17080 7890
rect 17512 7546 17540 7890
rect 19904 7546 19932 7890
rect 17040 7540 17092 7546
rect 17040 7482 17092 7488
rect 17500 7540 17552 7546
rect 17500 7482 17552 7488
rect 19892 7540 19944 7546
rect 19892 7482 19944 7488
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 20088 480 20116 9551
rect 20364 7954 20392 15558
rect 20916 14226 20944 22442
rect 21180 19304 21232 19310
rect 21178 19272 21180 19281
rect 21232 19272 21234 19281
rect 21178 19207 21234 19216
rect 20996 19168 21048 19174
rect 20996 19110 21048 19116
rect 20824 14198 20944 14226
rect 20626 13832 20682 13841
rect 20626 13767 20682 13776
rect 20640 12850 20668 13767
rect 20824 13394 20852 14198
rect 20904 14068 20956 14074
rect 20904 14010 20956 14016
rect 20916 13802 20944 14010
rect 21008 13938 21036 19110
rect 21456 18624 21508 18630
rect 21456 18566 21508 18572
rect 21272 18284 21324 18290
rect 21272 18226 21324 18232
rect 21178 17368 21234 17377
rect 21178 17303 21234 17312
rect 21088 17264 21140 17270
rect 21088 17206 21140 17212
rect 21100 16726 21128 17206
rect 21088 16720 21140 16726
rect 21192 16697 21220 17303
rect 21088 16662 21140 16668
rect 21178 16688 21234 16697
rect 21100 15706 21128 16662
rect 21178 16623 21234 16632
rect 21192 16250 21220 16623
rect 21180 16244 21232 16250
rect 21180 16186 21232 16192
rect 21192 16046 21220 16186
rect 21180 16040 21232 16046
rect 21180 15982 21232 15988
rect 21284 15722 21312 18226
rect 21468 18154 21496 18566
rect 21456 18148 21508 18154
rect 21456 18090 21508 18096
rect 21560 17610 21588 23559
rect 21652 23322 21680 27520
rect 22468 23656 22520 23662
rect 22466 23624 22468 23633
rect 22520 23624 22522 23633
rect 22466 23559 22522 23568
rect 23032 23497 23060 27520
rect 24412 27418 24440 27520
rect 24320 27390 24440 27418
rect 25318 27432 25374 27441
rect 23478 26344 23534 26353
rect 23478 26279 23534 26288
rect 22006 23488 22062 23497
rect 22006 23423 22062 23432
rect 23018 23488 23074 23497
rect 23018 23423 23074 23432
rect 21640 23316 21692 23322
rect 21640 23258 21692 23264
rect 21824 22092 21876 22098
rect 21824 22034 21876 22040
rect 21836 21486 21864 22034
rect 22020 21962 22048 23423
rect 22650 23352 22706 23361
rect 22650 23287 22652 23296
rect 22704 23287 22706 23296
rect 22652 23258 22704 23264
rect 22468 23180 22520 23186
rect 22468 23122 22520 23128
rect 22480 22438 22508 23122
rect 23492 22817 23520 26279
rect 24320 25242 24348 27390
rect 25318 27367 25374 27376
rect 24674 25392 24730 25401
rect 24674 25327 24730 25336
rect 24228 25214 24348 25242
rect 23570 24440 23626 24449
rect 23570 24375 23626 24384
rect 23478 22808 23534 22817
rect 23478 22743 23534 22752
rect 22468 22432 22520 22438
rect 22468 22374 22520 22380
rect 22008 21956 22060 21962
rect 22008 21898 22060 21904
rect 22480 21593 22508 22374
rect 22466 21584 22522 21593
rect 22466 21519 22522 21528
rect 21824 21480 21876 21486
rect 21822 21448 21824 21457
rect 21876 21448 21878 21457
rect 21822 21383 21878 21392
rect 23584 19961 23612 24375
rect 23846 24168 23902 24177
rect 23846 24103 23902 24112
rect 23860 23866 23888 24103
rect 23848 23860 23900 23866
rect 23848 23802 23900 23808
rect 24228 23361 24256 25214
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24214 23352 24270 23361
rect 24214 23287 24270 23296
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 23662 21448 23718 21457
rect 23662 21383 23718 21392
rect 23570 19952 23626 19961
rect 23570 19887 23626 19896
rect 23480 19168 23532 19174
rect 23480 19110 23532 19116
rect 23492 19009 23520 19110
rect 21822 19000 21878 19009
rect 21822 18935 21824 18944
rect 21876 18935 21878 18944
rect 23478 19000 23534 19009
rect 23478 18935 23534 18944
rect 21824 18906 21876 18912
rect 21836 18358 21864 18906
rect 23480 18896 23532 18902
rect 23478 18864 23480 18873
rect 23532 18864 23534 18873
rect 23478 18799 23534 18808
rect 21824 18352 21876 18358
rect 21824 18294 21876 18300
rect 21640 18284 21692 18290
rect 21640 18226 21692 18232
rect 21652 17678 21680 18226
rect 23478 18048 23534 18057
rect 23478 17983 23534 17992
rect 22284 17808 22336 17814
rect 22284 17750 22336 17756
rect 21640 17672 21692 17678
rect 21640 17614 21692 17620
rect 21548 17604 21600 17610
rect 21548 17546 21600 17552
rect 21560 16561 21588 17546
rect 21652 17202 21680 17614
rect 22296 17338 22324 17750
rect 22468 17672 22520 17678
rect 22468 17614 22520 17620
rect 22284 17332 22336 17338
rect 22284 17274 22336 17280
rect 22480 17241 22508 17614
rect 22650 17368 22706 17377
rect 23492 17354 23520 17983
rect 23400 17338 23520 17354
rect 22650 17303 22706 17312
rect 23388 17332 23520 17338
rect 22466 17232 22522 17241
rect 21640 17196 21692 17202
rect 22466 17167 22522 17176
rect 21640 17138 21692 17144
rect 21652 16726 21680 17138
rect 22560 17128 22612 17134
rect 22558 17096 22560 17105
rect 22612 17096 22614 17105
rect 22558 17031 22614 17040
rect 22376 16992 22428 16998
rect 22376 16934 22428 16940
rect 22388 16794 22416 16934
rect 22664 16794 22692 17303
rect 23440 17326 23520 17332
rect 23388 17274 23440 17280
rect 23676 17134 23704 21383
rect 24122 20904 24178 20913
rect 24122 20839 24178 20848
rect 23664 17128 23716 17134
rect 23664 17070 23716 17076
rect 23940 17128 23992 17134
rect 23940 17070 23992 17076
rect 24030 17096 24086 17105
rect 23848 16992 23900 16998
rect 23848 16934 23900 16940
rect 22376 16788 22428 16794
rect 22376 16730 22428 16736
rect 22652 16788 22704 16794
rect 22652 16730 22704 16736
rect 23756 16788 23808 16794
rect 23756 16730 23808 16736
rect 21640 16720 21692 16726
rect 21640 16662 21692 16668
rect 22468 16652 22520 16658
rect 22468 16594 22520 16600
rect 21546 16552 21602 16561
rect 21546 16487 21602 16496
rect 22480 16046 22508 16594
rect 23112 16584 23164 16590
rect 23112 16526 23164 16532
rect 22468 16040 22520 16046
rect 22466 16008 22468 16017
rect 22520 16008 22522 16017
rect 22466 15943 22522 15952
rect 21088 15700 21140 15706
rect 21088 15642 21140 15648
rect 21192 15694 21312 15722
rect 21192 15586 21220 15694
rect 23124 15638 23152 16526
rect 23480 15904 23532 15910
rect 23480 15846 23532 15852
rect 21100 15558 21220 15586
rect 21272 15632 21324 15638
rect 21272 15574 21324 15580
rect 23112 15632 23164 15638
rect 23112 15574 23164 15580
rect 23204 15632 23256 15638
rect 23204 15574 23256 15580
rect 20996 13932 21048 13938
rect 20996 13874 21048 13880
rect 20904 13796 20956 13802
rect 20904 13738 20956 13744
rect 21008 13530 21036 13874
rect 20996 13524 21048 13530
rect 20996 13466 21048 13472
rect 20812 13388 20864 13394
rect 20812 13330 20864 13336
rect 20720 13320 20772 13326
rect 20720 13262 20772 13268
rect 20628 12844 20680 12850
rect 20628 12786 20680 12792
rect 20732 12442 20760 13262
rect 20824 12889 20852 13330
rect 20810 12880 20866 12889
rect 20810 12815 20866 12824
rect 20720 12436 20772 12442
rect 20720 12378 20772 12384
rect 20812 12368 20864 12374
rect 20812 12310 20864 12316
rect 20720 12232 20772 12238
rect 20720 12174 20772 12180
rect 20732 11354 20760 12174
rect 20824 11558 20852 12310
rect 21100 11898 21128 15558
rect 21180 15496 21232 15502
rect 21180 15438 21232 15444
rect 21192 14618 21220 15438
rect 21284 15162 21312 15574
rect 21824 15496 21876 15502
rect 21824 15438 21876 15444
rect 21836 15201 21864 15438
rect 21916 15360 21968 15366
rect 21916 15302 21968 15308
rect 21822 15192 21878 15201
rect 21272 15156 21324 15162
rect 21822 15127 21878 15136
rect 21272 15098 21324 15104
rect 21824 14952 21876 14958
rect 21822 14920 21824 14929
rect 21928 14940 21956 15302
rect 23124 15162 23152 15574
rect 23112 15156 23164 15162
rect 23112 15098 23164 15104
rect 21876 14920 21956 14940
rect 21878 14912 21956 14920
rect 21822 14855 21878 14864
rect 21732 14816 21784 14822
rect 21732 14758 21784 14764
rect 22744 14816 22796 14822
rect 23216 14770 23244 15574
rect 23492 15337 23520 15846
rect 23572 15632 23624 15638
rect 23572 15574 23624 15580
rect 23478 15328 23534 15337
rect 23478 15263 23534 15272
rect 23492 15162 23520 15263
rect 23480 15156 23532 15162
rect 23480 15098 23532 15104
rect 23492 14890 23520 15098
rect 23480 14884 23532 14890
rect 23480 14826 23532 14832
rect 22744 14758 22796 14764
rect 21180 14612 21232 14618
rect 21180 14554 21232 14560
rect 21192 13938 21220 14554
rect 21744 14550 21772 14758
rect 22756 14657 22784 14758
rect 23124 14742 23244 14770
rect 22742 14648 22798 14657
rect 22742 14583 22798 14592
rect 21732 14544 21784 14550
rect 21732 14486 21784 14492
rect 21456 14408 21508 14414
rect 21454 14376 21456 14385
rect 21508 14376 21510 14385
rect 21454 14311 21510 14320
rect 21468 14074 21496 14311
rect 21456 14068 21508 14074
rect 21456 14010 21508 14016
rect 21180 13932 21232 13938
rect 21180 13874 21232 13880
rect 21744 13734 21772 14486
rect 23124 14278 23152 14742
rect 23584 14634 23612 15574
rect 23662 15192 23718 15201
rect 23662 15127 23718 15136
rect 23204 14612 23256 14618
rect 23204 14554 23256 14560
rect 23492 14606 23612 14634
rect 23112 14272 23164 14278
rect 23112 14214 23164 14220
rect 22466 14104 22522 14113
rect 22466 14039 22468 14048
rect 22520 14039 22522 14048
rect 22468 14010 22520 14016
rect 23124 14006 23152 14214
rect 23216 14074 23244 14554
rect 23492 14498 23520 14606
rect 23400 14470 23520 14498
rect 23400 14414 23428 14470
rect 23676 14414 23704 15127
rect 23388 14408 23440 14414
rect 23388 14350 23440 14356
rect 23664 14408 23716 14414
rect 23664 14350 23716 14356
rect 23204 14068 23256 14074
rect 23204 14010 23256 14016
rect 23112 14000 23164 14006
rect 23112 13942 23164 13948
rect 23294 13968 23350 13977
rect 22284 13864 22336 13870
rect 22282 13832 22284 13841
rect 23124 13841 23152 13942
rect 23294 13903 23350 13912
rect 22336 13832 22338 13841
rect 22282 13767 22338 13776
rect 23110 13832 23166 13841
rect 23308 13802 23336 13903
rect 23110 13767 23166 13776
rect 23296 13796 23348 13802
rect 23296 13738 23348 13744
rect 21732 13728 21784 13734
rect 21732 13670 21784 13676
rect 21640 13456 21692 13462
rect 21640 13398 21692 13404
rect 21652 13025 21680 13398
rect 21638 13016 21694 13025
rect 21638 12951 21640 12960
rect 21692 12951 21694 12960
rect 21640 12922 21692 12928
rect 21652 12891 21680 12922
rect 21272 12436 21324 12442
rect 21272 12378 21324 12384
rect 21284 12238 21312 12378
rect 21546 12336 21602 12345
rect 21546 12271 21602 12280
rect 21560 12238 21588 12271
rect 21272 12232 21324 12238
rect 21272 12174 21324 12180
rect 21548 12232 21600 12238
rect 21548 12174 21600 12180
rect 21088 11892 21140 11898
rect 21088 11834 21140 11840
rect 21100 11665 21128 11834
rect 21086 11656 21142 11665
rect 21086 11591 21142 11600
rect 20812 11552 20864 11558
rect 20812 11494 20864 11500
rect 21272 11552 21324 11558
rect 21272 11494 21324 11500
rect 20824 11354 20852 11494
rect 20720 11348 20772 11354
rect 20720 11290 20772 11296
rect 20812 11348 20864 11354
rect 20812 11290 20864 11296
rect 21284 11257 21312 11494
rect 21456 11280 21508 11286
rect 21270 11248 21326 11257
rect 21456 11222 21508 11228
rect 21270 11183 21326 11192
rect 20720 11144 20772 11150
rect 20720 11086 20772 11092
rect 21180 11144 21232 11150
rect 21180 11086 21232 11092
rect 20732 10962 20760 11086
rect 20640 10934 20760 10962
rect 20534 10840 20590 10849
rect 20534 10775 20590 10784
rect 20444 10736 20496 10742
rect 20444 10678 20496 10684
rect 20456 9926 20484 10678
rect 20444 9920 20496 9926
rect 20444 9862 20496 9868
rect 20456 8090 20484 9862
rect 20548 8566 20576 10775
rect 20640 8634 20668 10934
rect 20732 10810 20760 10934
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 21192 10674 21220 11086
rect 21468 10742 21496 11222
rect 21560 11200 21588 12174
rect 21744 11762 21772 13670
rect 23308 13462 23336 13738
rect 23400 13462 23428 14350
rect 23296 13456 23348 13462
rect 23296 13398 23348 13404
rect 23388 13456 23440 13462
rect 23388 13398 23440 13404
rect 22192 13320 22244 13326
rect 22192 13262 22244 13268
rect 22204 12850 22232 13262
rect 23308 12986 23336 13398
rect 23296 12980 23348 12986
rect 23296 12922 23348 12928
rect 22008 12844 22060 12850
rect 22008 12786 22060 12792
rect 22192 12844 22244 12850
rect 22192 12786 22244 12792
rect 21916 12708 21968 12714
rect 21916 12650 21968 12656
rect 21928 12102 21956 12650
rect 21916 12096 21968 12102
rect 21914 12064 21916 12073
rect 21968 12064 21970 12073
rect 21914 11999 21970 12008
rect 21928 11973 21956 11999
rect 21732 11756 21784 11762
rect 21732 11698 21784 11704
rect 21640 11212 21692 11218
rect 21560 11172 21640 11200
rect 21640 11154 21692 11160
rect 21456 10736 21508 10742
rect 21456 10678 21508 10684
rect 21180 10668 21232 10674
rect 21180 10610 21232 10616
rect 21088 10192 21140 10198
rect 21088 10134 21140 10140
rect 20902 9752 20958 9761
rect 21100 9722 21128 10134
rect 21192 10062 21220 10610
rect 21180 10056 21232 10062
rect 21180 9998 21232 10004
rect 20902 9687 20958 9696
rect 21088 9716 21140 9722
rect 20812 9376 20864 9382
rect 20810 9344 20812 9353
rect 20864 9344 20866 9353
rect 20810 9279 20866 9288
rect 20916 9178 20944 9687
rect 21088 9658 21140 9664
rect 21192 9654 21220 9998
rect 21364 9920 21416 9926
rect 21364 9862 21416 9868
rect 21180 9648 21232 9654
rect 21180 9590 21232 9596
rect 20904 9172 20956 9178
rect 20904 9114 20956 9120
rect 20996 9104 21048 9110
rect 20994 9072 20996 9081
rect 21048 9072 21050 9081
rect 20994 9007 21050 9016
rect 21008 8634 21036 9007
rect 21192 8974 21220 9590
rect 21376 9586 21404 9862
rect 21364 9580 21416 9586
rect 21364 9522 21416 9528
rect 21272 9172 21324 9178
rect 21272 9114 21324 9120
rect 21180 8968 21232 8974
rect 21180 8910 21232 8916
rect 20628 8628 20680 8634
rect 20628 8570 20680 8576
rect 20996 8628 21048 8634
rect 20996 8570 21048 8576
rect 20536 8560 20588 8566
rect 20536 8502 20588 8508
rect 21284 8362 21312 9114
rect 21376 8906 21404 9522
rect 21364 8900 21416 8906
rect 21364 8842 21416 8848
rect 21376 8498 21404 8842
rect 21364 8492 21416 8498
rect 21364 8434 21416 8440
rect 21180 8356 21232 8362
rect 21180 8298 21232 8304
rect 21272 8356 21324 8362
rect 21272 8298 21324 8304
rect 21192 8265 21220 8298
rect 21178 8256 21234 8265
rect 21178 8191 21234 8200
rect 21192 8090 21220 8191
rect 20444 8084 20496 8090
rect 20444 8026 20496 8032
rect 21180 8084 21232 8090
rect 21180 8026 21232 8032
rect 21376 8022 21404 8434
rect 21468 8090 21496 10678
rect 22020 10266 22048 12786
rect 22204 12442 22232 12786
rect 23388 12708 23440 12714
rect 23440 12668 23520 12696
rect 23388 12650 23440 12656
rect 23492 12594 23520 12668
rect 23492 12566 23612 12594
rect 22192 12436 22244 12442
rect 22192 12378 22244 12384
rect 23584 12374 23612 12566
rect 22836 12368 22888 12374
rect 22836 12310 22888 12316
rect 23572 12368 23624 12374
rect 23572 12310 23624 12316
rect 23768 12322 23796 16730
rect 23860 13326 23888 16934
rect 23848 13320 23900 13326
rect 23848 13262 23900 13268
rect 23860 12986 23888 13262
rect 23848 12980 23900 12986
rect 23848 12922 23900 12928
rect 22848 12209 22876 12310
rect 23768 12294 23888 12322
rect 22928 12232 22980 12238
rect 22834 12200 22890 12209
rect 22928 12174 22980 12180
rect 22834 12135 22890 12144
rect 22848 11898 22876 12135
rect 22836 11892 22888 11898
rect 22836 11834 22888 11840
rect 22940 11286 22968 12174
rect 23756 12164 23808 12170
rect 23756 12106 23808 12112
rect 23664 12096 23716 12102
rect 23664 12038 23716 12044
rect 23572 11892 23624 11898
rect 23572 11834 23624 11840
rect 23480 11824 23532 11830
rect 23400 11772 23480 11778
rect 23400 11766 23532 11772
rect 23400 11750 23520 11766
rect 22928 11280 22980 11286
rect 22928 11222 22980 11228
rect 22376 11212 22428 11218
rect 22376 11154 22428 11160
rect 22388 10810 22416 11154
rect 23400 10810 23428 11750
rect 23584 11642 23612 11834
rect 23492 11614 23612 11642
rect 23492 10810 23520 11614
rect 23676 11286 23704 12038
rect 23768 11762 23796 12106
rect 23860 11937 23888 12294
rect 23846 11928 23902 11937
rect 23846 11863 23902 11872
rect 23756 11756 23808 11762
rect 23756 11698 23808 11704
rect 23664 11280 23716 11286
rect 23664 11222 23716 11228
rect 23572 11144 23624 11150
rect 23572 11086 23624 11092
rect 22376 10804 22428 10810
rect 22376 10746 22428 10752
rect 23388 10804 23440 10810
rect 23388 10746 23440 10752
rect 23480 10804 23532 10810
rect 23480 10746 23532 10752
rect 22650 10568 22706 10577
rect 22650 10503 22706 10512
rect 22008 10260 22060 10266
rect 22008 10202 22060 10208
rect 21640 9988 21692 9994
rect 21640 9930 21692 9936
rect 21652 9761 21680 9930
rect 21638 9752 21694 9761
rect 21638 9687 21694 9696
rect 21652 9586 21680 9687
rect 21640 9580 21692 9586
rect 21640 9522 21692 9528
rect 22100 9172 22152 9178
rect 22100 9114 22152 9120
rect 22112 8634 22140 9114
rect 22664 9110 22692 10503
rect 23020 10464 23072 10470
rect 23020 10406 23072 10412
rect 22652 9104 22704 9110
rect 22652 9046 22704 9052
rect 22560 8968 22612 8974
rect 22560 8910 22612 8916
rect 22100 8628 22152 8634
rect 22100 8570 22152 8576
rect 22572 8498 22600 8910
rect 22664 8634 22692 9046
rect 22652 8628 22704 8634
rect 22652 8570 22704 8576
rect 22560 8492 22612 8498
rect 22560 8434 22612 8440
rect 21456 8084 21508 8090
rect 21456 8026 21508 8032
rect 21364 8016 21416 8022
rect 21468 7993 21496 8026
rect 21364 7958 21416 7964
rect 21454 7984 21510 7993
rect 20352 7948 20404 7954
rect 21454 7919 21510 7928
rect 20352 7890 20404 7896
rect 21468 7546 21496 7919
rect 21548 7880 21600 7886
rect 21548 7822 21600 7828
rect 21456 7540 21508 7546
rect 21456 7482 21508 7488
rect 21560 7206 21588 7822
rect 21548 7200 21600 7206
rect 21546 7168 21548 7177
rect 21600 7168 21602 7177
rect 21546 7103 21602 7112
rect 23032 5250 23060 10406
rect 23584 10266 23612 11086
rect 23572 10260 23624 10266
rect 23572 10202 23624 10208
rect 23572 10124 23624 10130
rect 23572 10066 23624 10072
rect 23584 9382 23612 10066
rect 23676 9994 23704 11222
rect 23768 11150 23796 11698
rect 23756 11144 23808 11150
rect 23756 11086 23808 11092
rect 23768 10674 23796 11086
rect 23848 10804 23900 10810
rect 23848 10746 23900 10752
rect 23756 10668 23808 10674
rect 23756 10610 23808 10616
rect 23860 10538 23888 10746
rect 23848 10532 23900 10538
rect 23848 10474 23900 10480
rect 23664 9988 23716 9994
rect 23664 9930 23716 9936
rect 23754 9752 23810 9761
rect 23754 9687 23810 9696
rect 23572 9376 23624 9382
rect 23572 9318 23624 9324
rect 23478 8256 23534 8265
rect 23478 8191 23534 8200
rect 23492 8090 23520 8191
rect 23480 8084 23532 8090
rect 23480 8026 23532 8032
rect 23584 6905 23612 9318
rect 23768 7954 23796 9687
rect 23756 7948 23808 7954
rect 23756 7890 23808 7896
rect 23768 7546 23796 7890
rect 23756 7540 23808 7546
rect 23756 7482 23808 7488
rect 23570 6896 23626 6905
rect 23570 6831 23626 6840
rect 23952 5681 23980 17070
rect 24030 17031 24086 17040
rect 24044 12209 24072 17031
rect 24136 15706 24164 20839
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24688 18850 24716 25327
rect 25332 23866 25360 27367
rect 25792 24177 25820 27520
rect 27172 24857 27200 27520
rect 26698 24848 26754 24857
rect 26698 24783 26754 24792
rect 27158 24848 27214 24857
rect 27158 24783 27214 24792
rect 26712 24313 26740 24783
rect 26698 24304 26754 24313
rect 26698 24239 26754 24248
rect 25778 24168 25834 24177
rect 25778 24103 25834 24112
rect 25320 23860 25372 23866
rect 25320 23802 25372 23808
rect 25332 23662 25360 23802
rect 25320 23656 25372 23662
rect 25320 23598 25372 23604
rect 24860 23520 24912 23526
rect 24860 23462 24912 23468
rect 24766 21176 24822 21185
rect 24766 21111 24822 21120
rect 24780 19310 24808 21111
rect 24872 20913 24900 23462
rect 24858 20904 24914 20913
rect 24858 20839 24914 20848
rect 24768 19304 24820 19310
rect 24768 19246 24820 19252
rect 24596 18834 24716 18850
rect 24584 18828 24716 18834
rect 24636 18822 24716 18828
rect 24584 18770 24636 18776
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24688 18426 24716 18822
rect 24676 18420 24728 18426
rect 24676 18362 24728 18368
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24952 17060 25004 17066
rect 24952 17002 25004 17008
rect 24676 16992 24728 16998
rect 24676 16934 24728 16940
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24400 15972 24452 15978
rect 24400 15914 24452 15920
rect 24124 15700 24176 15706
rect 24124 15642 24176 15648
rect 24136 15026 24164 15642
rect 24412 15638 24440 15914
rect 24400 15632 24452 15638
rect 24400 15574 24452 15580
rect 24582 15600 24638 15609
rect 24582 15535 24584 15544
rect 24636 15535 24638 15544
rect 24584 15506 24636 15512
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24688 15042 24716 16934
rect 24768 16652 24820 16658
rect 24768 16594 24820 16600
rect 24780 16250 24808 16594
rect 24768 16244 24820 16250
rect 24768 16186 24820 16192
rect 24766 16008 24822 16017
rect 24766 15943 24822 15952
rect 24780 15706 24808 15943
rect 24768 15700 24820 15706
rect 24768 15642 24820 15648
rect 24860 15564 24912 15570
rect 24860 15506 24912 15512
rect 24872 15162 24900 15506
rect 24860 15156 24912 15162
rect 24860 15098 24912 15104
rect 24124 15020 24176 15026
rect 24688 15014 24808 15042
rect 24124 14962 24176 14968
rect 24214 14920 24270 14929
rect 24214 14855 24270 14864
rect 24676 14884 24728 14890
rect 24124 13796 24176 13802
rect 24124 13738 24176 13744
rect 24136 13190 24164 13738
rect 24124 13184 24176 13190
rect 24124 13126 24176 13132
rect 24030 12200 24086 12209
rect 24030 12135 24086 12144
rect 24032 11756 24084 11762
rect 24032 11698 24084 11704
rect 24044 11082 24072 11698
rect 24032 11076 24084 11082
rect 24032 11018 24084 11024
rect 24032 10124 24084 10130
rect 24032 10066 24084 10072
rect 24044 9722 24072 10066
rect 24032 9716 24084 9722
rect 24032 9658 24084 9664
rect 24136 7410 24164 13126
rect 24228 12646 24256 14855
rect 24676 14826 24728 14832
rect 24688 14550 24716 14826
rect 24676 14544 24728 14550
rect 24676 14486 24728 14492
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24688 14006 24716 14486
rect 24676 14000 24728 14006
rect 24676 13942 24728 13948
rect 24780 13462 24808 15014
rect 24964 14958 24992 17002
rect 25226 16144 25282 16153
rect 25226 16079 25282 16088
rect 25240 16046 25268 16079
rect 25228 16040 25280 16046
rect 25228 15982 25280 15988
rect 25240 15178 25268 15982
rect 25240 15150 25360 15178
rect 24952 14952 25004 14958
rect 24952 14894 25004 14900
rect 24950 14648 25006 14657
rect 24950 14583 25006 14592
rect 24964 14550 24992 14583
rect 24952 14544 25004 14550
rect 24952 14486 25004 14492
rect 24964 14074 24992 14486
rect 24952 14068 25004 14074
rect 24952 14010 25004 14016
rect 24858 13832 24914 13841
rect 24858 13767 24914 13776
rect 24872 13462 24900 13767
rect 24768 13456 24820 13462
rect 24768 13398 24820 13404
rect 24860 13456 24912 13462
rect 24860 13398 24912 13404
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24780 12986 24808 13398
rect 24872 12986 24900 13398
rect 24768 12980 24820 12986
rect 24768 12922 24820 12928
rect 24860 12980 24912 12986
rect 24860 12922 24912 12928
rect 24582 12880 24638 12889
rect 24582 12815 24638 12824
rect 25226 12880 25282 12889
rect 25226 12815 25282 12824
rect 24596 12782 24624 12815
rect 24584 12776 24636 12782
rect 24584 12718 24636 12724
rect 24216 12640 24268 12646
rect 24216 12582 24268 12588
rect 24676 12368 24728 12374
rect 24676 12310 24728 12316
rect 24216 12232 24268 12238
rect 24216 12174 24268 12180
rect 24228 11830 24256 12174
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24688 11898 24716 12310
rect 24676 11892 24728 11898
rect 24676 11834 24728 11840
rect 24216 11824 24268 11830
rect 24216 11766 24268 11772
rect 24860 11688 24912 11694
rect 24214 11656 24270 11665
rect 24214 11591 24270 11600
rect 24688 11636 24860 11642
rect 24688 11630 24912 11636
rect 24688 11614 24900 11630
rect 24228 10554 24256 11591
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24228 10526 24348 10554
rect 24216 10464 24268 10470
rect 24216 10406 24268 10412
rect 24124 7404 24176 7410
rect 24124 7346 24176 7352
rect 23938 5672 23994 5681
rect 23938 5607 23994 5616
rect 23032 5222 23520 5250
rect 23492 3505 23520 5222
rect 23202 3496 23258 3505
rect 23202 3431 23258 3440
rect 23478 3496 23534 3505
rect 23478 3431 23534 3440
rect 23216 480 23244 3431
rect 24228 2650 24256 10406
rect 24320 10130 24348 10526
rect 24308 10124 24360 10130
rect 24308 10066 24360 10072
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24688 8548 24716 11614
rect 25240 11354 25268 12815
rect 25228 11348 25280 11354
rect 25228 11290 25280 11296
rect 25136 11212 25188 11218
rect 25136 11154 25188 11160
rect 24766 10840 24822 10849
rect 24766 10775 24822 10784
rect 24780 10266 24808 10775
rect 25044 10464 25096 10470
rect 25044 10406 25096 10412
rect 24768 10260 24820 10266
rect 24768 10202 24820 10208
rect 25056 10198 25084 10406
rect 25148 10266 25176 11154
rect 25226 10704 25282 10713
rect 25226 10639 25282 10648
rect 25240 10606 25268 10639
rect 25228 10600 25280 10606
rect 25228 10542 25280 10548
rect 25136 10260 25188 10266
rect 25136 10202 25188 10208
rect 25044 10192 25096 10198
rect 25044 10134 25096 10140
rect 24766 9752 24822 9761
rect 24766 9687 24822 9696
rect 24780 9654 24808 9687
rect 25332 9654 25360 15150
rect 25688 14816 25740 14822
rect 25688 14758 25740 14764
rect 25596 14408 25648 14414
rect 25596 14350 25648 14356
rect 25412 14000 25464 14006
rect 25412 13942 25464 13948
rect 25424 13462 25452 13942
rect 25504 13932 25556 13938
rect 25504 13874 25556 13880
rect 25412 13456 25464 13462
rect 25412 13398 25464 13404
rect 25410 12200 25466 12209
rect 25410 12135 25466 12144
rect 25424 11898 25452 12135
rect 25412 11892 25464 11898
rect 25412 11834 25464 11840
rect 25410 11792 25466 11801
rect 25410 11727 25466 11736
rect 25424 10810 25452 11727
rect 25412 10804 25464 10810
rect 25412 10746 25464 10752
rect 24768 9648 24820 9654
rect 24768 9590 24820 9596
rect 25320 9648 25372 9654
rect 25320 9590 25372 9596
rect 25516 9042 25544 13874
rect 25608 13870 25636 14350
rect 25700 13977 25728 14758
rect 25686 13968 25742 13977
rect 25686 13903 25742 13912
rect 25596 13864 25648 13870
rect 25596 13806 25648 13812
rect 26330 9344 26386 9353
rect 26330 9279 26386 9288
rect 25504 9036 25556 9042
rect 25504 8978 25556 8984
rect 24768 8832 24820 8838
rect 24766 8800 24768 8809
rect 24820 8800 24822 8809
rect 24766 8735 24822 8744
rect 25516 8634 25544 8978
rect 25504 8628 25556 8634
rect 25504 8570 25556 8576
rect 24504 8520 24716 8548
rect 24504 8022 24532 8520
rect 24768 8356 24820 8362
rect 24768 8298 24820 8304
rect 24492 8016 24544 8022
rect 24492 7958 24544 7964
rect 24676 7948 24728 7954
rect 24676 7890 24728 7896
rect 24688 7721 24716 7890
rect 24674 7712 24730 7721
rect 24289 7644 24585 7664
rect 24674 7647 24730 7656
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24688 7546 24716 7647
rect 24676 7540 24728 7546
rect 24676 7482 24728 7488
rect 24676 7404 24728 7410
rect 24676 7346 24728 7352
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24688 3194 24716 7346
rect 24780 4593 24808 8298
rect 24858 7168 24914 7177
rect 24858 7103 24914 7112
rect 24766 4584 24822 4593
rect 24766 4519 24822 4528
rect 24676 3188 24728 3194
rect 24676 3130 24728 3136
rect 24872 2650 24900 7103
rect 25136 2848 25188 2854
rect 25134 2816 25136 2825
rect 25188 2816 25190 2825
rect 25134 2751 25190 2760
rect 24216 2644 24268 2650
rect 24216 2586 24268 2592
rect 24860 2644 24912 2650
rect 24860 2586 24912 2592
rect 25596 2508 25648 2514
rect 25596 2450 25648 2456
rect 25608 2310 25636 2450
rect 24676 2304 24728 2310
rect 24676 2246 24728 2252
rect 25596 2304 25648 2310
rect 25596 2246 25648 2252
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24688 513 24716 2246
rect 25608 1465 25636 2246
rect 25594 1456 25650 1465
rect 25594 1391 25650 1400
rect 24674 504 24730 513
rect 2778 439 2834 448
rect 4526 0 4582 480
rect 7654 0 7710 480
rect 10782 0 10838 480
rect 13910 0 13966 480
rect 16946 0 17002 480
rect 20074 0 20130 480
rect 23202 0 23258 480
rect 26344 480 26372 9279
rect 24674 439 24730 448
rect 26330 0 26386 480
<< via2 >>
rect 1490 26288 1546 26344
rect 1398 25336 1454 25392
rect 2502 27376 2558 27432
rect 2042 23432 2098 23488
rect 1398 21120 1454 21176
rect 1766 20984 1822 21040
rect 1766 17856 1822 17912
rect 1582 17040 1638 17096
rect 2134 17040 2190 17096
rect 1398 14864 1454 14920
rect 1582 15952 1638 16008
rect 2042 15680 2098 15736
rect 1490 13912 1546 13968
rect 1490 9696 1546 9752
rect 1398 7656 1454 7712
rect 1766 10784 1822 10840
rect 1582 8744 1638 8800
rect 1490 6568 1546 6624
rect 1398 5616 1454 5672
rect 1858 9016 1914 9072
rect 1398 4528 1454 4584
rect 1582 3440 1638 3496
rect 1398 2508 1454 2544
rect 1398 2488 1400 2508
rect 1400 2488 1452 2508
rect 1452 2488 1454 2508
rect 1490 1400 1546 1456
rect 2134 13948 2136 13968
rect 2136 13948 2188 13968
rect 2188 13948 2190 13968
rect 2134 13912 2190 13948
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 2686 23704 2742 23760
rect 2686 23588 2742 23624
rect 2686 23568 2688 23588
rect 2688 23568 2740 23588
rect 2740 23568 2742 23588
rect 2410 14728 2466 14784
rect 2686 14592 2742 14648
rect 2042 10684 2044 10704
rect 2044 10684 2096 10704
rect 2096 10684 2098 10704
rect 2042 10648 2098 10684
rect 2134 9560 2190 9616
rect 2134 9016 2190 9072
rect 2042 6840 2098 6896
rect 2502 12708 2558 12744
rect 2502 12688 2504 12708
rect 2504 12688 2556 12708
rect 2556 12688 2558 12708
rect 2410 12416 2466 12472
rect 4802 24792 4858 24848
rect 3514 24248 3570 24304
rect 3422 22208 3478 22264
rect 3422 21392 3478 21448
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5538 23704 5594 23760
rect 4250 23432 4306 23488
rect 3514 20440 3570 20496
rect 4066 17720 4122 17776
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 7378 19488 7434 19544
rect 3238 14764 3240 14784
rect 3240 14764 3292 14784
rect 3292 14764 3294 14784
rect 3238 14728 3294 14764
rect 3054 14592 3110 14648
rect 4894 15408 4950 15464
rect 4158 13640 4214 13696
rect 2502 11464 2558 11520
rect 2502 9832 2558 9888
rect 2318 9152 2374 9208
rect 2778 9288 2834 9344
rect 2962 11736 3018 11792
rect 2870 8472 2926 8528
rect 3790 10532 3846 10568
rect 3790 10512 3792 10532
rect 3792 10512 3844 10532
rect 3844 10512 3846 10532
rect 3422 9832 3478 9888
rect 4250 9424 4306 9480
rect 3238 8880 3294 8936
rect 3606 8880 3662 8936
rect 2594 6976 2650 7032
rect 2594 5908 2650 5944
rect 2594 5888 2596 5908
rect 2596 5888 2648 5908
rect 2648 5888 2650 5908
rect 2502 5772 2558 5808
rect 2502 5752 2504 5772
rect 2504 5752 2556 5772
rect 2556 5752 2558 5772
rect 4434 9152 4490 9208
rect 4434 9016 4490 9072
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5170 15544 5226 15600
rect 5354 15680 5410 15736
rect 5078 14320 5134 14376
rect 5170 13232 5226 13288
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5538 12860 5540 12880
rect 5540 12860 5592 12880
rect 5592 12860 5594 12880
rect 5538 12824 5594 12860
rect 5262 12416 5318 12472
rect 6274 12960 6330 13016
rect 6182 12588 6184 12608
rect 6184 12588 6236 12608
rect 6236 12588 6238 12608
rect 6182 12552 6238 12588
rect 4894 9580 4950 9616
rect 4894 9560 4896 9580
rect 4896 9560 4948 9580
rect 4948 9560 4950 9580
rect 4802 6996 4858 7032
rect 4802 6976 4804 6996
rect 4804 6976 4856 6996
rect 4856 6976 4858 6996
rect 5078 7248 5134 7304
rect 5078 6860 5134 6896
rect 5078 6840 5080 6860
rect 5080 6840 5132 6860
rect 5132 6840 5134 6860
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 6458 18536 6514 18592
rect 7194 17856 7250 17912
rect 7102 15408 7158 15464
rect 7010 14728 7066 14784
rect 6734 14048 6790 14104
rect 7194 14764 7196 14784
rect 7196 14764 7248 14784
rect 7248 14764 7250 14784
rect 7194 14728 7250 14764
rect 7194 11464 7250 11520
rect 7286 9444 7342 9480
rect 7286 9424 7288 9444
rect 7288 9424 7340 9444
rect 7340 9424 7342 9444
rect 7010 9324 7012 9344
rect 7012 9324 7064 9344
rect 7064 9324 7066 9344
rect 7010 9288 7066 9324
rect 6366 6840 6422 6896
rect 7746 18400 7802 18456
rect 7654 17992 7710 18048
rect 7654 16088 7710 16144
rect 7838 13368 7894 13424
rect 7470 12008 7526 12064
rect 7562 10648 7618 10704
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5354 5888 5410 5944
rect 4894 5752 4950 5808
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 4526 3984 4582 4040
rect 3330 3576 3386 3632
rect 2778 448 2834 504
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 8206 24792 8262 24848
rect 8206 19488 8262 19544
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10690 20984 10746 21040
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 9862 19508 9918 19544
rect 9862 19488 9864 19508
rect 9864 19488 9916 19508
rect 9916 19488 9918 19508
rect 8206 14476 8262 14512
rect 8206 14456 8208 14476
rect 8208 14456 8260 14476
rect 8260 14456 8262 14476
rect 8298 14184 8354 14240
rect 8942 17584 8998 17640
rect 9034 16632 9090 16688
rect 8666 15136 8722 15192
rect 8666 14068 8722 14104
rect 8666 14048 8668 14068
rect 8668 14048 8720 14068
rect 8720 14048 8722 14068
rect 9402 18128 9458 18184
rect 9494 15952 9550 16008
rect 9770 15564 9826 15600
rect 9770 15544 9772 15564
rect 9772 15544 9824 15564
rect 9824 15544 9826 15564
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10506 18844 10508 18864
rect 10508 18844 10560 18864
rect 10560 18844 10562 18864
rect 10506 18808 10562 18844
rect 10322 18400 10378 18456
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10138 17176 10194 17232
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10874 18808 10930 18864
rect 10966 16632 11022 16688
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10874 15680 10930 15736
rect 10138 15408 10194 15464
rect 9034 14612 9090 14648
rect 9034 14592 9036 14612
rect 9036 14592 9088 14612
rect 9088 14592 9090 14612
rect 8942 13912 8998 13968
rect 8574 13776 8630 13832
rect 8482 13232 8538 13288
rect 8758 11600 8814 11656
rect 10046 15000 10102 15056
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10782 14456 10838 14512
rect 10046 13640 10102 13696
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 9218 10648 9274 10704
rect 8850 10512 8906 10568
rect 9678 9580 9734 9616
rect 9678 9560 9680 9580
rect 9680 9560 9732 9580
rect 9732 9560 9734 9580
rect 8482 8472 8538 8528
rect 9586 6724 9642 6760
rect 10598 12008 10654 12064
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10782 11328 10838 11384
rect 10966 14456 11022 14512
rect 10966 14184 11022 14240
rect 11058 13232 11114 13288
rect 10874 10648 10930 10704
rect 10690 9696 10746 9752
rect 10874 9696 10930 9752
rect 10690 9560 10746 9616
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10138 8880 10194 8936
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10322 7928 10378 7984
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10322 6860 10378 6896
rect 10322 6840 10324 6860
rect 10324 6840 10376 6860
rect 10376 6840 10378 6860
rect 9586 6704 9588 6724
rect 9588 6704 9640 6724
rect 9640 6704 9642 6724
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 11794 18536 11850 18592
rect 11978 18400 12034 18456
rect 11794 18128 11850 18184
rect 11978 18128 12034 18184
rect 11426 15816 11482 15872
rect 11334 13912 11390 13968
rect 11426 13776 11482 13832
rect 11150 11736 11206 11792
rect 11518 12960 11574 13016
rect 11794 16224 11850 16280
rect 11794 15544 11850 15600
rect 11794 13404 11796 13424
rect 11796 13404 11848 13424
rect 11848 13404 11850 13424
rect 11794 13368 11850 13404
rect 11242 9460 11244 9480
rect 11244 9460 11296 9480
rect 11296 9460 11298 9480
rect 11242 9424 11298 9460
rect 11518 11056 11574 11112
rect 11150 8472 11206 8528
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 11242 3984 11298 4040
rect 12990 23860 13046 23896
rect 12990 23840 12992 23860
rect 12992 23840 13044 23860
rect 13044 23840 13046 23860
rect 12438 19352 12494 19408
rect 12438 18572 12440 18592
rect 12440 18572 12492 18592
rect 12492 18572 12494 18592
rect 12438 18536 12494 18572
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 14646 23840 14702 23896
rect 16394 24404 16450 24440
rect 16394 24384 16396 24404
rect 16396 24384 16448 24404
rect 16448 24384 16450 24404
rect 17406 24384 17462 24440
rect 17406 24268 17462 24304
rect 17406 24248 17408 24268
rect 17408 24248 17460 24268
rect 17460 24248 17462 24268
rect 16486 23588 16542 23624
rect 16486 23568 16488 23588
rect 16488 23568 16540 23588
rect 16540 23568 16542 23588
rect 17130 23588 17186 23624
rect 17130 23568 17132 23588
rect 17132 23568 17184 23588
rect 17184 23568 17186 23588
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 16118 22208 16174 22264
rect 15750 22072 15806 22128
rect 13082 19216 13138 19272
rect 12530 17176 12586 17232
rect 12530 15136 12586 15192
rect 12254 12180 12256 12200
rect 12256 12180 12308 12200
rect 12308 12180 12310 12200
rect 12254 12144 12310 12180
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 12622 8472 12678 8528
rect 13358 12144 13414 12200
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 13818 15952 13874 16008
rect 13910 12300 13966 12336
rect 13910 12280 13912 12300
rect 13912 12280 13964 12300
rect 13964 12280 13966 12300
rect 13542 10648 13598 10704
rect 13910 11348 13966 11384
rect 13910 11328 13912 11348
rect 13912 11328 13964 11348
rect 13964 11328 13966 11348
rect 13726 10512 13782 10568
rect 13726 10376 13782 10432
rect 13634 9560 13690 9616
rect 14186 15816 14242 15872
rect 14370 16904 14426 16960
rect 14370 15952 14426 16008
rect 14370 12552 14426 12608
rect 16302 21972 16304 21992
rect 16304 21972 16356 21992
rect 16356 21972 16358 21992
rect 16302 21936 16358 21972
rect 16394 21564 16396 21584
rect 16396 21564 16448 21584
rect 16448 21564 16450 21584
rect 16394 21528 16450 21564
rect 16670 20168 16726 20224
rect 16118 17720 16174 17776
rect 15290 16652 15346 16688
rect 15290 16632 15292 16652
rect 15292 16632 15344 16652
rect 15344 16632 15346 16652
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 15750 16768 15806 16824
rect 16578 16768 16634 16824
rect 15474 15680 15530 15736
rect 14738 15408 14794 15464
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 16486 15444 16488 15464
rect 16488 15444 16540 15464
rect 16540 15444 16542 15464
rect 16486 15408 16542 15444
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 18694 23160 18750 23216
rect 18602 22772 18658 22808
rect 18602 22752 18604 22772
rect 18604 22752 18656 22772
rect 18656 22752 18658 22772
rect 18050 22072 18106 22128
rect 18142 21972 18144 21992
rect 18144 21972 18196 21992
rect 18196 21972 18198 21992
rect 18142 21936 18198 21972
rect 17590 19352 17646 19408
rect 17222 17176 17278 17232
rect 17774 16940 17776 16960
rect 17776 16940 17828 16960
rect 17828 16940 17830 16960
rect 17774 16904 17830 16940
rect 17130 16516 17186 16552
rect 17130 16496 17132 16516
rect 17132 16496 17184 16516
rect 17184 16496 17186 16516
rect 17130 14884 17186 14920
rect 17130 14864 17132 14884
rect 17132 14864 17184 14884
rect 17184 14864 17186 14884
rect 16854 14456 16910 14512
rect 16762 14340 16818 14376
rect 16762 14320 16764 14340
rect 16764 14320 16816 14340
rect 16816 14320 16818 14340
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 16578 12980 16634 13016
rect 16578 12960 16580 12980
rect 16580 12960 16632 12980
rect 16632 12960 16634 12980
rect 14554 11600 14610 11656
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14922 11636 14924 11656
rect 14924 11636 14976 11656
rect 14976 11636 14978 11656
rect 14370 11192 14426 11248
rect 13266 6840 13322 6896
rect 11794 3440 11850 3496
rect 13082 3440 13138 3496
rect 14186 9424 14242 9480
rect 14922 11600 14978 11636
rect 15290 11192 15346 11248
rect 15842 11056 15898 11112
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14646 9696 14702 9752
rect 15658 10804 15714 10840
rect 15658 10784 15660 10804
rect 15660 10784 15712 10804
rect 15712 10784 15714 10804
rect 16026 10512 16082 10568
rect 15566 10104 15622 10160
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14738 8200 14794 8256
rect 16302 9696 16358 9752
rect 16118 7928 16174 7984
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 15382 7284 15384 7304
rect 15384 7284 15436 7304
rect 15436 7284 15438 7304
rect 15382 7248 15438 7284
rect 17774 14356 17776 14376
rect 17776 14356 17828 14376
rect 17828 14356 17830 14376
rect 17774 14320 17830 14356
rect 17038 12280 17094 12336
rect 16854 10412 16856 10432
rect 16856 10412 16908 10432
rect 16908 10412 16910 10432
rect 16854 10376 16910 10412
rect 16762 8336 16818 8392
rect 16670 8064 16726 8120
rect 16486 6704 16542 6760
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 17498 12552 17554 12608
rect 17314 12008 17370 12064
rect 17406 11772 17408 11792
rect 17408 11772 17460 11792
rect 17460 11772 17462 11792
rect 17406 11736 17462 11772
rect 18234 12280 18290 12336
rect 18050 12144 18106 12200
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 21546 23568 21602 23624
rect 20902 22500 20958 22536
rect 20902 22480 20904 22500
rect 20904 22480 20956 22500
rect 20956 22480 20958 22500
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 18786 20576 18842 20632
rect 20810 20576 20866 20632
rect 19798 20440 19854 20496
rect 19338 19352 19394 19408
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19522 19916 19578 19952
rect 19522 19896 19524 19916
rect 19524 19896 19576 19916
rect 19576 19896 19578 19916
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 18694 15544 18750 15600
rect 18602 15020 18658 15056
rect 18602 15000 18604 15020
rect 18604 15000 18656 15020
rect 18656 15000 18658 15020
rect 19062 17620 19064 17640
rect 19064 17620 19116 17640
rect 19116 17620 19118 17640
rect 19062 17584 19118 17620
rect 19430 17720 19486 17776
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 20166 17448 20222 17504
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19522 16632 19578 16688
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 20718 18284 20774 18320
rect 20718 18264 20720 18284
rect 20720 18264 20772 18284
rect 20772 18264 20774 18284
rect 20718 17584 20774 17640
rect 20258 15544 20314 15600
rect 20074 15408 20130 15464
rect 19982 15308 19984 15328
rect 19984 15308 20036 15328
rect 20036 15308 20038 15328
rect 19982 15272 20038 15308
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 18878 14048 18934 14104
rect 19890 13948 19892 13968
rect 19892 13948 19944 13968
rect 19944 13948 19946 13968
rect 19890 13912 19946 13948
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19338 12552 19394 12608
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19246 12280 19302 12336
rect 19062 11600 19118 11656
rect 19246 11192 19302 11248
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 17958 10104 18014 10160
rect 18510 9016 18566 9072
rect 20166 10784 20222 10840
rect 20258 10532 20314 10568
rect 20258 10512 20260 10532
rect 20260 10512 20312 10532
rect 20312 10512 20314 10532
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 20074 9560 20130 9616
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 17498 8200 17554 8256
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 21178 19252 21180 19272
rect 21180 19252 21232 19272
rect 21232 19252 21234 19272
rect 21178 19216 21234 19252
rect 20626 13776 20682 13832
rect 21178 17312 21234 17368
rect 21178 16632 21234 16688
rect 22466 23604 22468 23624
rect 22468 23604 22520 23624
rect 22520 23604 22522 23624
rect 22466 23568 22522 23604
rect 23478 26288 23534 26344
rect 22006 23432 22062 23488
rect 23018 23432 23074 23488
rect 22650 23316 22706 23352
rect 22650 23296 22652 23316
rect 22652 23296 22704 23316
rect 22704 23296 22706 23316
rect 25318 27376 25374 27432
rect 24674 25336 24730 25392
rect 23570 24384 23626 24440
rect 23478 22752 23534 22808
rect 22466 21528 22522 21584
rect 21822 21428 21824 21448
rect 21824 21428 21876 21448
rect 21876 21428 21878 21448
rect 21822 21392 21878 21428
rect 23846 24112 23902 24168
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24214 23296 24270 23352
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 23662 21392 23718 21448
rect 23570 19896 23626 19952
rect 21822 18964 21878 19000
rect 21822 18944 21824 18964
rect 21824 18944 21876 18964
rect 21876 18944 21878 18964
rect 23478 18944 23534 19000
rect 23478 18844 23480 18864
rect 23480 18844 23532 18864
rect 23532 18844 23534 18864
rect 23478 18808 23534 18844
rect 23478 17992 23534 18048
rect 22650 17312 22706 17368
rect 22466 17176 22522 17232
rect 22558 17076 22560 17096
rect 22560 17076 22612 17096
rect 22612 17076 22614 17096
rect 22558 17040 22614 17076
rect 24122 20848 24178 20904
rect 21546 16496 21602 16552
rect 22466 15988 22468 16008
rect 22468 15988 22520 16008
rect 22520 15988 22522 16008
rect 22466 15952 22522 15988
rect 20810 12824 20866 12880
rect 21822 15136 21878 15192
rect 21822 14900 21824 14920
rect 21824 14900 21876 14920
rect 21876 14900 21878 14920
rect 21822 14864 21878 14900
rect 23478 15272 23534 15328
rect 22742 14592 22798 14648
rect 21454 14356 21456 14376
rect 21456 14356 21508 14376
rect 21508 14356 21510 14376
rect 21454 14320 21510 14356
rect 23662 15136 23718 15192
rect 22466 14068 22522 14104
rect 22466 14048 22468 14068
rect 22468 14048 22520 14068
rect 22520 14048 22522 14068
rect 23294 13912 23350 13968
rect 22282 13812 22284 13832
rect 22284 13812 22336 13832
rect 22336 13812 22338 13832
rect 22282 13776 22338 13812
rect 23110 13776 23166 13832
rect 21638 12980 21694 13016
rect 21638 12960 21640 12980
rect 21640 12960 21692 12980
rect 21692 12960 21694 12980
rect 21546 12280 21602 12336
rect 21086 11600 21142 11656
rect 21270 11192 21326 11248
rect 20534 10784 20590 10840
rect 21914 12044 21916 12064
rect 21916 12044 21968 12064
rect 21968 12044 21970 12064
rect 21914 12008 21970 12044
rect 20902 9696 20958 9752
rect 20810 9324 20812 9344
rect 20812 9324 20864 9344
rect 20864 9324 20866 9344
rect 20810 9288 20866 9324
rect 20994 9052 20996 9072
rect 20996 9052 21048 9072
rect 21048 9052 21050 9072
rect 20994 9016 21050 9052
rect 21178 8200 21234 8256
rect 22834 12144 22890 12200
rect 23846 11872 23902 11928
rect 22650 10512 22706 10568
rect 21638 9696 21694 9752
rect 21454 7928 21510 7984
rect 21546 7148 21548 7168
rect 21548 7148 21600 7168
rect 21600 7148 21602 7168
rect 21546 7112 21602 7148
rect 23754 9696 23810 9752
rect 23478 8200 23534 8256
rect 23570 6840 23626 6896
rect 24030 17040 24086 17096
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 26698 24792 26754 24848
rect 27158 24792 27214 24848
rect 26698 24248 26754 24304
rect 25778 24112 25834 24168
rect 24766 21120 24822 21176
rect 24858 20848 24914 20904
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24582 15564 24638 15600
rect 24582 15544 24584 15564
rect 24584 15544 24636 15564
rect 24636 15544 24638 15564
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24766 15952 24822 16008
rect 24214 14864 24270 14920
rect 24030 12144 24086 12200
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 25226 16088 25282 16144
rect 24950 14592 25006 14648
rect 24858 13776 24914 13832
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24582 12824 24638 12880
rect 25226 12824 25282 12880
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24214 11600 24270 11656
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 23938 5616 23994 5672
rect 23202 3440 23258 3496
rect 23478 3440 23534 3496
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24766 10784 24822 10840
rect 25226 10648 25282 10704
rect 24766 9696 24822 9752
rect 25410 12144 25466 12200
rect 25410 11736 25466 11792
rect 25686 13912 25742 13968
rect 26330 9288 26386 9344
rect 24766 8780 24768 8800
rect 24768 8780 24820 8800
rect 24820 8780 24822 8800
rect 24766 8744 24822 8780
rect 24674 7656 24730 7712
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24858 7112 24914 7168
rect 24766 4528 24822 4584
rect 25134 2796 25136 2816
rect 25136 2796 25188 2816
rect 25188 2796 25190 2816
rect 25134 2760 25190 2796
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 25594 1400 25650 1456
rect 24674 448 24730 504
<< metal3 >>
rect 0 27434 480 27464
rect 2497 27434 2563 27437
rect 0 27432 2563 27434
rect 0 27376 2502 27432
rect 2558 27376 2563 27432
rect 0 27374 2563 27376
rect 0 27344 480 27374
rect 2497 27371 2563 27374
rect 25313 27434 25379 27437
rect 27520 27434 28000 27464
rect 25313 27432 28000 27434
rect 25313 27376 25318 27432
rect 25374 27376 28000 27432
rect 25313 27374 28000 27376
rect 25313 27371 25379 27374
rect 27520 27344 28000 27374
rect 0 26346 480 26376
rect 1485 26346 1551 26349
rect 0 26344 1551 26346
rect 0 26288 1490 26344
rect 1546 26288 1551 26344
rect 0 26286 1551 26288
rect 0 26256 480 26286
rect 1485 26283 1551 26286
rect 23473 26346 23539 26349
rect 27520 26346 28000 26376
rect 23473 26344 28000 26346
rect 23473 26288 23478 26344
rect 23534 26288 28000 26344
rect 23473 26286 28000 26288
rect 23473 26283 23539 26286
rect 27520 26256 28000 26286
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 0 25394 480 25424
rect 1393 25394 1459 25397
rect 0 25392 1459 25394
rect 0 25336 1398 25392
rect 1454 25336 1459 25392
rect 0 25334 1459 25336
rect 0 25304 480 25334
rect 1393 25331 1459 25334
rect 24669 25394 24735 25397
rect 27520 25394 28000 25424
rect 24669 25392 28000 25394
rect 24669 25336 24674 25392
rect 24730 25336 28000 25392
rect 24669 25334 28000 25336
rect 24669 25331 24735 25334
rect 27520 25304 28000 25334
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 4797 24850 4863 24853
rect 8201 24850 8267 24853
rect 4797 24848 8267 24850
rect 4797 24792 4802 24848
rect 4858 24792 8206 24848
rect 8262 24792 8267 24848
rect 4797 24790 8267 24792
rect 4797 24787 4863 24790
rect 8201 24787 8267 24790
rect 26693 24850 26759 24853
rect 27153 24850 27219 24853
rect 26693 24848 27219 24850
rect 26693 24792 26698 24848
rect 26754 24792 27158 24848
rect 27214 24792 27219 24848
rect 26693 24790 27219 24792
rect 26693 24787 26759 24790
rect 27153 24787 27219 24790
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 16389 24442 16455 24445
rect 17401 24442 17467 24445
rect 16389 24440 17467 24442
rect 16389 24384 16394 24440
rect 16450 24384 17406 24440
rect 17462 24384 17467 24440
rect 16389 24382 17467 24384
rect 16389 24379 16455 24382
rect 17401 24379 17467 24382
rect 23565 24442 23631 24445
rect 23565 24440 26986 24442
rect 23565 24384 23570 24440
rect 23626 24384 26986 24440
rect 23565 24382 26986 24384
rect 23565 24379 23631 24382
rect 0 24306 480 24336
rect 3509 24306 3575 24309
rect 0 24304 3575 24306
rect 0 24248 3514 24304
rect 3570 24248 3575 24304
rect 0 24246 3575 24248
rect 0 24216 480 24246
rect 3509 24243 3575 24246
rect 17401 24306 17467 24309
rect 26693 24306 26759 24309
rect 17401 24304 26759 24306
rect 17401 24248 17406 24304
rect 17462 24248 26698 24304
rect 26754 24248 26759 24304
rect 17401 24246 26759 24248
rect 26926 24306 26986 24382
rect 27520 24306 28000 24336
rect 26926 24246 28000 24306
rect 17401 24243 17467 24246
rect 26693 24243 26759 24246
rect 27520 24216 28000 24246
rect 23841 24170 23907 24173
rect 25773 24170 25839 24173
rect 23841 24168 25839 24170
rect 23841 24112 23846 24168
rect 23902 24112 25778 24168
rect 25834 24112 25839 24168
rect 23841 24110 25839 24112
rect 23841 24107 23907 24110
rect 25773 24107 25839 24110
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 12985 23898 13051 23901
rect 14641 23898 14707 23901
rect 12985 23896 14707 23898
rect 12985 23840 12990 23896
rect 13046 23840 14646 23896
rect 14702 23840 14707 23896
rect 12985 23838 14707 23840
rect 12985 23835 13051 23838
rect 14641 23835 14707 23838
rect 2681 23762 2747 23765
rect 5533 23762 5599 23765
rect 2681 23760 5599 23762
rect 2681 23704 2686 23760
rect 2742 23704 5538 23760
rect 5594 23704 5599 23760
rect 2681 23702 5599 23704
rect 2681 23699 2747 23702
rect 5533 23699 5599 23702
rect 2681 23626 2747 23629
rect 16481 23626 16547 23629
rect 2681 23624 16547 23626
rect 2681 23568 2686 23624
rect 2742 23568 16486 23624
rect 16542 23568 16547 23624
rect 2681 23566 16547 23568
rect 2681 23563 2747 23566
rect 16481 23563 16547 23566
rect 17125 23626 17191 23629
rect 21541 23626 21607 23629
rect 22461 23626 22527 23629
rect 17125 23624 22527 23626
rect 17125 23568 17130 23624
rect 17186 23568 21546 23624
rect 21602 23568 22466 23624
rect 22522 23568 22527 23624
rect 17125 23566 22527 23568
rect 17125 23563 17191 23566
rect 21541 23563 21607 23566
rect 22461 23563 22527 23566
rect 2037 23490 2103 23493
rect 4245 23490 4311 23493
rect 2037 23488 4311 23490
rect 2037 23432 2042 23488
rect 2098 23432 4250 23488
rect 4306 23432 4311 23488
rect 2037 23430 4311 23432
rect 2037 23427 2103 23430
rect 4245 23427 4311 23430
rect 22001 23490 22067 23493
rect 23013 23490 23079 23493
rect 22001 23488 23079 23490
rect 22001 23432 22006 23488
rect 22062 23432 23018 23488
rect 23074 23432 23079 23488
rect 22001 23430 23079 23432
rect 22001 23427 22067 23430
rect 23013 23427 23079 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 22645 23354 22711 23357
rect 24209 23354 24275 23357
rect 22645 23352 24275 23354
rect 22645 23296 22650 23352
rect 22706 23296 24214 23352
rect 24270 23296 24275 23352
rect 22645 23294 24275 23296
rect 22645 23291 22711 23294
rect 24209 23291 24275 23294
rect 0 23218 480 23248
rect 18689 23218 18755 23221
rect 27520 23218 28000 23248
rect 0 23158 674 23218
rect 0 23128 480 23158
rect 614 22538 674 23158
rect 18689 23216 28000 23218
rect 18689 23160 18694 23216
rect 18750 23160 28000 23216
rect 18689 23158 28000 23160
rect 18689 23155 18755 23158
rect 27520 23128 28000 23158
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 18597 22810 18663 22813
rect 23473 22810 23539 22813
rect 18597 22808 23539 22810
rect 18597 22752 18602 22808
rect 18658 22752 23478 22808
rect 23534 22752 23539 22808
rect 18597 22750 23539 22752
rect 18597 22747 18663 22750
rect 23473 22747 23539 22750
rect 20897 22538 20963 22541
rect 614 22536 20963 22538
rect 614 22480 20902 22536
rect 20958 22480 20963 22536
rect 614 22478 20963 22480
rect 20897 22475 20963 22478
rect 10277 22336 10597 22337
rect 0 22266 480 22296
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 3417 22266 3483 22269
rect 0 22264 3483 22266
rect 0 22208 3422 22264
rect 3478 22208 3483 22264
rect 0 22206 3483 22208
rect 0 22176 480 22206
rect 3417 22203 3483 22206
rect 16113 22266 16179 22269
rect 27520 22266 28000 22296
rect 16113 22264 18338 22266
rect 16113 22208 16118 22264
rect 16174 22208 18338 22264
rect 16113 22206 18338 22208
rect 16113 22203 16179 22206
rect 15745 22130 15811 22133
rect 18045 22130 18111 22133
rect 15745 22128 18111 22130
rect 15745 22072 15750 22128
rect 15806 22072 18050 22128
rect 18106 22072 18111 22128
rect 15745 22070 18111 22072
rect 18278 22130 18338 22206
rect 27478 22176 28000 22266
rect 27478 22130 27538 22176
rect 18278 22070 27538 22130
rect 15745 22067 15811 22070
rect 18045 22067 18111 22070
rect 16297 21994 16363 21997
rect 18137 21994 18203 21997
rect 16297 21992 18203 21994
rect 16297 21936 16302 21992
rect 16358 21936 18142 21992
rect 18198 21936 18203 21992
rect 16297 21934 18203 21936
rect 16297 21931 16363 21934
rect 18137 21931 18203 21934
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 16389 21586 16455 21589
rect 22461 21586 22527 21589
rect 16389 21584 22527 21586
rect 16389 21528 16394 21584
rect 16450 21528 22466 21584
rect 22522 21528 22527 21584
rect 16389 21526 22527 21528
rect 16389 21523 16455 21526
rect 22461 21523 22527 21526
rect 3417 21450 3483 21453
rect 21817 21450 21883 21453
rect 23657 21450 23723 21453
rect 3417 21448 23723 21450
rect 3417 21392 3422 21448
rect 3478 21392 21822 21448
rect 21878 21392 23662 21448
rect 23718 21392 23723 21448
rect 3417 21390 23723 21392
rect 3417 21387 3483 21390
rect 21817 21387 21883 21390
rect 23657 21387 23723 21390
rect 10277 21248 10597 21249
rect 0 21178 480 21208
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 1393 21178 1459 21181
rect 0 21176 1459 21178
rect 0 21120 1398 21176
rect 1454 21120 1459 21176
rect 0 21118 1459 21120
rect 0 21088 480 21118
rect 1393 21115 1459 21118
rect 24761 21178 24827 21181
rect 27520 21178 28000 21208
rect 24761 21176 28000 21178
rect 24761 21120 24766 21176
rect 24822 21120 28000 21176
rect 24761 21118 28000 21120
rect 24761 21115 24827 21118
rect 27520 21088 28000 21118
rect 1761 21042 1827 21045
rect 10685 21042 10751 21045
rect 1761 21040 10751 21042
rect 1761 20984 1766 21040
rect 1822 20984 10690 21040
rect 10746 20984 10751 21040
rect 1761 20982 10751 20984
rect 1761 20979 1827 20982
rect 10685 20979 10751 20982
rect 24117 20906 24183 20909
rect 24853 20906 24919 20909
rect 24117 20904 24919 20906
rect 24117 20848 24122 20904
rect 24178 20848 24858 20904
rect 24914 20848 24919 20904
rect 24117 20846 24919 20848
rect 24117 20843 24183 20846
rect 24853 20843 24919 20846
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 18781 20634 18847 20637
rect 20805 20634 20871 20637
rect 18781 20632 20871 20634
rect 18781 20576 18786 20632
rect 18842 20576 20810 20632
rect 20866 20576 20871 20632
rect 18781 20574 20871 20576
rect 18781 20571 18847 20574
rect 20805 20571 20871 20574
rect 3509 20498 3575 20501
rect 19793 20498 19859 20501
rect 3509 20496 19859 20498
rect 3509 20440 3514 20496
rect 3570 20440 19798 20496
rect 19854 20440 19859 20496
rect 3509 20438 19859 20440
rect 3509 20435 3575 20438
rect 19793 20435 19859 20438
rect 19382 20302 27538 20362
rect 16665 20228 16731 20229
rect 16614 20164 16620 20228
rect 16684 20226 16731 20228
rect 19382 20226 19442 20302
rect 16684 20224 19442 20226
rect 16726 20168 19442 20224
rect 16684 20166 19442 20168
rect 16684 20164 16731 20166
rect 16665 20163 16731 20164
rect 10277 20160 10597 20161
rect 0 20090 480 20120
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 27478 20120 27538 20302
rect 0 20030 674 20090
rect 27478 20030 28000 20120
rect 0 20000 480 20030
rect 614 19410 674 20030
rect 27520 20000 28000 20030
rect 19517 19954 19583 19957
rect 23565 19954 23631 19957
rect 19517 19952 23631 19954
rect 19517 19896 19522 19952
rect 19578 19896 23570 19952
rect 23626 19896 23631 19952
rect 19517 19894 23631 19896
rect 19517 19891 19583 19894
rect 23565 19891 23631 19894
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 7373 19546 7439 19549
rect 8201 19546 8267 19549
rect 9857 19546 9923 19549
rect 7373 19544 9923 19546
rect 7373 19488 7378 19544
rect 7434 19488 8206 19544
rect 8262 19488 9862 19544
rect 9918 19488 9923 19544
rect 7373 19486 9923 19488
rect 7373 19483 7439 19486
rect 8201 19483 8267 19486
rect 9857 19483 9923 19486
rect 12433 19410 12499 19413
rect 614 19408 12499 19410
rect 614 19352 12438 19408
rect 12494 19352 12499 19408
rect 614 19350 12499 19352
rect 12433 19347 12499 19350
rect 17585 19410 17651 19413
rect 19333 19410 19399 19413
rect 17585 19408 19399 19410
rect 17585 19352 17590 19408
rect 17646 19352 19338 19408
rect 19394 19352 19399 19408
rect 17585 19350 19399 19352
rect 17585 19347 17651 19350
rect 19333 19347 19399 19350
rect 13077 19274 13143 19277
rect 21173 19274 21239 19277
rect 13077 19272 21239 19274
rect 13077 19216 13082 19272
rect 13138 19216 21178 19272
rect 21234 19216 21239 19272
rect 13077 19214 21239 19216
rect 13077 19211 13143 19214
rect 21173 19211 21239 19214
rect 0 19138 480 19168
rect 27520 19138 28000 19168
rect 0 19078 674 19138
rect 0 19048 480 19078
rect 614 18322 674 19078
rect 24902 19078 28000 19138
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 21817 19002 21883 19005
rect 23473 19002 23539 19005
rect 21817 19000 23539 19002
rect 21817 18944 21822 19000
rect 21878 18944 23478 19000
rect 23534 18944 23539 19000
rect 21817 18942 23539 18944
rect 21817 18939 21883 18942
rect 23473 18939 23539 18942
rect 10501 18866 10567 18869
rect 10869 18866 10935 18869
rect 23473 18866 23539 18869
rect 10501 18864 23539 18866
rect 10501 18808 10506 18864
rect 10562 18808 10874 18864
rect 10930 18808 23478 18864
rect 23534 18808 23539 18864
rect 10501 18806 23539 18808
rect 10501 18803 10567 18806
rect 10869 18803 10935 18806
rect 23473 18803 23539 18806
rect 6453 18594 6519 18597
rect 11789 18594 11855 18597
rect 12433 18594 12499 18597
rect 6453 18592 10610 18594
rect 6453 18536 6458 18592
rect 6514 18536 10610 18592
rect 6453 18534 10610 18536
rect 6453 18531 6519 18534
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 7741 18458 7807 18461
rect 10317 18458 10383 18461
rect 7741 18456 10383 18458
rect 7741 18400 7746 18456
rect 7802 18400 10322 18456
rect 10378 18400 10383 18456
rect 7741 18398 10383 18400
rect 10550 18458 10610 18534
rect 11789 18592 12499 18594
rect 11789 18536 11794 18592
rect 11850 18536 12438 18592
rect 12494 18536 12499 18592
rect 11789 18534 12499 18536
rect 11789 18531 11855 18534
rect 12433 18531 12499 18534
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 11973 18458 12039 18461
rect 10550 18456 12039 18458
rect 10550 18400 11978 18456
rect 12034 18400 12039 18456
rect 10550 18398 12039 18400
rect 7741 18395 7807 18398
rect 10317 18395 10383 18398
rect 11973 18395 12039 18398
rect 20713 18322 20779 18325
rect 614 18320 20779 18322
rect 614 18264 20718 18320
rect 20774 18264 20779 18320
rect 614 18262 20779 18264
rect 20713 18259 20779 18262
rect 9397 18186 9463 18189
rect 11789 18186 11855 18189
rect 9397 18184 11855 18186
rect 9397 18128 9402 18184
rect 9458 18128 11794 18184
rect 11850 18128 11855 18184
rect 9397 18126 11855 18128
rect 9397 18123 9463 18126
rect 11789 18123 11855 18126
rect 11973 18186 12039 18189
rect 24902 18186 24962 19078
rect 27520 19048 28000 19078
rect 11973 18184 24962 18186
rect 11973 18128 11978 18184
rect 12034 18128 24962 18184
rect 11973 18126 24962 18128
rect 11973 18123 12039 18126
rect 0 18050 480 18080
rect 7649 18050 7715 18053
rect 0 18048 7715 18050
rect 0 17992 7654 18048
rect 7710 17992 7715 18048
rect 0 17990 7715 17992
rect 0 17960 480 17990
rect 7649 17987 7715 17990
rect 23473 18050 23539 18053
rect 27520 18050 28000 18080
rect 23473 18048 28000 18050
rect 23473 17992 23478 18048
rect 23534 17992 28000 18048
rect 23473 17990 28000 17992
rect 23473 17987 23539 17990
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 27520 17960 28000 17990
rect 19610 17919 19930 17920
rect 1761 17914 1827 17917
rect 7189 17914 7255 17917
rect 1761 17912 7255 17914
rect 1761 17856 1766 17912
rect 1822 17856 7194 17912
rect 7250 17856 7255 17912
rect 1761 17854 7255 17856
rect 1761 17851 1827 17854
rect 7189 17851 7255 17854
rect 4061 17778 4127 17781
rect 16113 17778 16179 17781
rect 19425 17780 19491 17781
rect 4061 17776 16179 17778
rect 4061 17720 4066 17776
rect 4122 17720 16118 17776
rect 16174 17720 16179 17776
rect 4061 17718 16179 17720
rect 4061 17715 4127 17718
rect 16113 17715 16179 17718
rect 19374 17716 19380 17780
rect 19444 17778 19491 17780
rect 19444 17776 19536 17778
rect 19486 17720 19536 17776
rect 19444 17718 19536 17720
rect 19444 17716 19491 17718
rect 19425 17715 19491 17716
rect 8937 17642 9003 17645
rect 19057 17642 19123 17645
rect 20713 17642 20779 17645
rect 8937 17640 18890 17642
rect 8937 17584 8942 17640
rect 8998 17584 18890 17640
rect 8937 17582 18890 17584
rect 8937 17579 9003 17582
rect 18830 17506 18890 17582
rect 19057 17640 20779 17642
rect 19057 17584 19062 17640
rect 19118 17584 20718 17640
rect 20774 17584 20779 17640
rect 19057 17582 20779 17584
rect 19057 17579 19123 17582
rect 20713 17579 20779 17582
rect 20161 17506 20227 17509
rect 18830 17504 20227 17506
rect 18830 17448 20166 17504
rect 20222 17448 20227 17504
rect 18830 17446 20227 17448
rect 20161 17443 20227 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 21173 17370 21239 17373
rect 22645 17370 22711 17373
rect 21173 17368 22711 17370
rect 21173 17312 21178 17368
rect 21234 17312 22650 17368
rect 22706 17312 22711 17368
rect 21173 17310 22711 17312
rect 21173 17307 21239 17310
rect 22645 17307 22711 17310
rect 10133 17234 10199 17237
rect 12525 17234 12591 17237
rect 10133 17232 12591 17234
rect 10133 17176 10138 17232
rect 10194 17176 12530 17232
rect 12586 17176 12591 17232
rect 10133 17174 12591 17176
rect 10133 17171 10199 17174
rect 12525 17171 12591 17174
rect 17217 17234 17283 17237
rect 22461 17234 22527 17237
rect 17217 17232 22527 17234
rect 17217 17176 17222 17232
rect 17278 17176 22466 17232
rect 22522 17176 22527 17232
rect 17217 17174 22527 17176
rect 17217 17171 17283 17174
rect 22461 17171 22527 17174
rect 0 17098 480 17128
rect 1577 17098 1643 17101
rect 0 17096 1643 17098
rect 0 17040 1582 17096
rect 1638 17040 1643 17096
rect 0 17038 1643 17040
rect 0 17008 480 17038
rect 1577 17035 1643 17038
rect 2129 17098 2195 17101
rect 22553 17098 22619 17101
rect 2129 17096 22619 17098
rect 2129 17040 2134 17096
rect 2190 17040 22558 17096
rect 22614 17040 22619 17096
rect 2129 17038 22619 17040
rect 2129 17035 2195 17038
rect 22553 17035 22619 17038
rect 24025 17098 24091 17101
rect 27520 17098 28000 17128
rect 24025 17096 28000 17098
rect 24025 17040 24030 17096
rect 24086 17040 28000 17096
rect 24025 17038 28000 17040
rect 24025 17035 24091 17038
rect 27520 17008 28000 17038
rect 14365 16962 14431 16965
rect 17769 16962 17835 16965
rect 14365 16960 17835 16962
rect 14365 16904 14370 16960
rect 14426 16904 17774 16960
rect 17830 16904 17835 16960
rect 14365 16902 17835 16904
rect 14365 16899 14431 16902
rect 17769 16899 17835 16902
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 15745 16826 15811 16829
rect 16573 16826 16639 16829
rect 10734 16824 16639 16826
rect 10734 16768 15750 16824
rect 15806 16768 16578 16824
rect 16634 16768 16639 16824
rect 10734 16766 16639 16768
rect 9029 16690 9095 16693
rect 10734 16690 10794 16766
rect 15745 16763 15811 16766
rect 16573 16763 16639 16766
rect 9029 16688 10794 16690
rect 9029 16632 9034 16688
rect 9090 16632 10794 16688
rect 9029 16630 10794 16632
rect 10961 16690 11027 16693
rect 15285 16690 15351 16693
rect 10961 16688 15351 16690
rect 10961 16632 10966 16688
rect 11022 16632 15290 16688
rect 15346 16632 15351 16688
rect 10961 16630 15351 16632
rect 9029 16627 9095 16630
rect 10961 16627 11027 16630
rect 15285 16627 15351 16630
rect 19517 16690 19583 16693
rect 21173 16690 21239 16693
rect 19517 16688 21239 16690
rect 19517 16632 19522 16688
rect 19578 16632 21178 16688
rect 21234 16632 21239 16688
rect 19517 16630 21239 16632
rect 19517 16627 19583 16630
rect 21173 16627 21239 16630
rect 17125 16554 17191 16557
rect 21541 16554 21607 16557
rect 17125 16552 21607 16554
rect 17125 16496 17130 16552
rect 17186 16496 21546 16552
rect 21602 16496 21607 16552
rect 17125 16494 21607 16496
rect 17125 16491 17191 16494
rect 21541 16491 21607 16494
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 11789 16282 11855 16285
rect 6686 16280 11855 16282
rect 6686 16224 11794 16280
rect 11850 16224 11855 16280
rect 6686 16222 11855 16224
rect 0 16010 480 16040
rect 1577 16010 1643 16013
rect 0 16008 1643 16010
rect 0 15952 1582 16008
rect 1638 15952 1643 16008
rect 0 15950 1643 15952
rect 0 15920 480 15950
rect 1577 15947 1643 15950
rect 2037 15738 2103 15741
rect 5349 15738 5415 15741
rect 6686 15738 6746 16222
rect 11789 16219 11855 16222
rect 7649 16146 7715 16149
rect 25221 16146 25287 16149
rect 7649 16144 25287 16146
rect 7649 16088 7654 16144
rect 7710 16088 25226 16144
rect 25282 16088 25287 16144
rect 7649 16086 25287 16088
rect 7649 16083 7715 16086
rect 25221 16083 25287 16086
rect 9489 16010 9555 16013
rect 13813 16010 13879 16013
rect 9489 16008 13879 16010
rect 9489 15952 9494 16008
rect 9550 15952 13818 16008
rect 13874 15952 13879 16008
rect 9489 15950 13879 15952
rect 9489 15947 9555 15950
rect 13813 15947 13879 15950
rect 14365 16010 14431 16013
rect 22461 16010 22527 16013
rect 14365 16008 22527 16010
rect 14365 15952 14370 16008
rect 14426 15952 22466 16008
rect 22522 15952 22527 16008
rect 14365 15950 22527 15952
rect 14365 15947 14431 15950
rect 22461 15947 22527 15950
rect 24761 16010 24827 16013
rect 27520 16010 28000 16040
rect 24761 16008 28000 16010
rect 24761 15952 24766 16008
rect 24822 15952 28000 16008
rect 24761 15950 28000 15952
rect 24761 15947 24827 15950
rect 27520 15920 28000 15950
rect 11421 15874 11487 15877
rect 14181 15874 14247 15877
rect 11421 15872 14247 15874
rect 11421 15816 11426 15872
rect 11482 15816 14186 15872
rect 14242 15816 14247 15872
rect 11421 15814 14247 15816
rect 11421 15811 11487 15814
rect 14181 15811 14247 15814
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 10869 15738 10935 15741
rect 15469 15738 15535 15741
rect 2037 15736 6746 15738
rect 2037 15680 2042 15736
rect 2098 15680 5354 15736
rect 5410 15680 6746 15736
rect 2037 15678 6746 15680
rect 10734 15736 15535 15738
rect 10734 15680 10874 15736
rect 10930 15680 15474 15736
rect 15530 15680 15535 15736
rect 10734 15678 15535 15680
rect 2037 15675 2103 15678
rect 5349 15675 5415 15678
rect 5165 15602 5231 15605
rect 9765 15602 9831 15605
rect 10734 15602 10794 15678
rect 10869 15675 10935 15678
rect 15469 15675 15535 15678
rect 5165 15600 10794 15602
rect 5165 15544 5170 15600
rect 5226 15544 9770 15600
rect 9826 15544 10794 15600
rect 5165 15542 10794 15544
rect 11789 15602 11855 15605
rect 18689 15602 18755 15605
rect 11789 15600 18755 15602
rect 11789 15544 11794 15600
rect 11850 15544 18694 15600
rect 18750 15544 18755 15600
rect 11789 15542 18755 15544
rect 5165 15539 5231 15542
rect 9765 15539 9831 15542
rect 11789 15539 11855 15542
rect 18689 15539 18755 15542
rect 20253 15602 20319 15605
rect 24577 15602 24643 15605
rect 20253 15600 24643 15602
rect 20253 15544 20258 15600
rect 20314 15544 24582 15600
rect 24638 15544 24643 15600
rect 20253 15542 24643 15544
rect 20253 15539 20319 15542
rect 24577 15539 24643 15542
rect 4889 15466 4955 15469
rect 7097 15466 7163 15469
rect 4889 15464 7163 15466
rect 4889 15408 4894 15464
rect 4950 15408 7102 15464
rect 7158 15408 7163 15464
rect 4889 15406 7163 15408
rect 4889 15403 4955 15406
rect 7097 15403 7163 15406
rect 10133 15466 10199 15469
rect 14733 15466 14799 15469
rect 10133 15464 14799 15466
rect 10133 15408 10138 15464
rect 10194 15408 14738 15464
rect 14794 15408 14799 15464
rect 10133 15406 14799 15408
rect 10133 15403 10199 15406
rect 14733 15403 14799 15406
rect 16481 15466 16547 15469
rect 20069 15466 20135 15469
rect 16481 15464 20135 15466
rect 16481 15408 16486 15464
rect 16542 15408 20074 15464
rect 20130 15408 20135 15464
rect 16481 15406 20135 15408
rect 16481 15403 16547 15406
rect 20069 15403 20135 15406
rect 19977 15330 20043 15333
rect 23473 15330 23539 15333
rect 19977 15328 23539 15330
rect 19977 15272 19982 15328
rect 20038 15272 23478 15328
rect 23534 15272 23539 15328
rect 19977 15270 23539 15272
rect 19977 15267 20043 15270
rect 23473 15267 23539 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 8661 15194 8727 15197
rect 12525 15194 12591 15197
rect 8661 15192 12591 15194
rect 8661 15136 8666 15192
rect 8722 15136 12530 15192
rect 12586 15136 12591 15192
rect 8661 15134 12591 15136
rect 8661 15131 8727 15134
rect 12525 15131 12591 15134
rect 21817 15194 21883 15197
rect 23657 15194 23723 15197
rect 21817 15192 23723 15194
rect 21817 15136 21822 15192
rect 21878 15136 23662 15192
rect 23718 15136 23723 15192
rect 21817 15134 23723 15136
rect 21817 15131 21883 15134
rect 23657 15131 23723 15134
rect 10041 15058 10107 15061
rect 18597 15058 18663 15061
rect 10041 15056 18663 15058
rect 10041 15000 10046 15056
rect 10102 15000 18602 15056
rect 18658 15000 18663 15056
rect 10041 14998 18663 15000
rect 10041 14995 10107 14998
rect 18597 14995 18663 14998
rect 0 14922 480 14952
rect 1393 14922 1459 14925
rect 17125 14922 17191 14925
rect 21817 14922 21883 14925
rect 0 14920 1459 14922
rect 0 14864 1398 14920
rect 1454 14864 1459 14920
rect 9768 14888 10794 14922
rect 0 14862 1459 14864
rect 0 14832 480 14862
rect 1393 14859 1459 14862
rect 9492 14862 10794 14888
rect 9492 14828 9828 14862
rect 2405 14786 2471 14789
rect 3233 14786 3299 14789
rect 7005 14786 7071 14789
rect 2405 14784 7071 14786
rect 2405 14728 2410 14784
rect 2466 14728 3238 14784
rect 3294 14728 7010 14784
rect 7066 14728 7071 14784
rect 2405 14726 7071 14728
rect 2405 14723 2471 14726
rect 3233 14723 3299 14726
rect 7005 14723 7071 14726
rect 7189 14786 7255 14789
rect 9492 14786 9552 14828
rect 7189 14784 9552 14786
rect 7189 14728 7194 14784
rect 7250 14728 9552 14784
rect 7189 14726 9552 14728
rect 10734 14786 10794 14862
rect 17125 14920 21883 14922
rect 17125 14864 17130 14920
rect 17186 14864 21822 14920
rect 21878 14864 21883 14920
rect 17125 14862 21883 14864
rect 17125 14859 17191 14862
rect 21817 14859 21883 14862
rect 24209 14922 24275 14925
rect 27520 14922 28000 14952
rect 24209 14920 28000 14922
rect 24209 14864 24214 14920
rect 24270 14864 28000 14920
rect 24209 14862 28000 14864
rect 24209 14859 24275 14862
rect 27520 14832 28000 14862
rect 19328 14786 19334 14788
rect 10734 14726 19334 14786
rect 7189 14723 7255 14726
rect 19328 14724 19334 14726
rect 19398 14724 19404 14788
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 2681 14650 2747 14653
rect 3049 14650 3115 14653
rect 9029 14650 9095 14653
rect 2681 14648 9095 14650
rect 2681 14592 2686 14648
rect 2742 14592 3054 14648
rect 3110 14592 9034 14648
rect 9090 14592 9095 14648
rect 2681 14590 9095 14592
rect 2681 14587 2747 14590
rect 3049 14587 3115 14590
rect 9029 14587 9095 14590
rect 22737 14650 22803 14653
rect 24945 14650 25011 14653
rect 22737 14648 25011 14650
rect 22737 14592 22742 14648
rect 22798 14592 24950 14648
rect 25006 14592 25011 14648
rect 22737 14590 25011 14592
rect 22737 14587 22803 14590
rect 24945 14587 25011 14590
rect 8201 14514 8267 14517
rect 10777 14514 10843 14517
rect 8201 14512 10843 14514
rect 8201 14456 8206 14512
rect 8262 14456 10782 14512
rect 10838 14456 10843 14512
rect 8201 14454 10843 14456
rect 8201 14451 8267 14454
rect 10777 14451 10843 14454
rect 10961 14514 11027 14517
rect 16849 14514 16915 14517
rect 10961 14512 16915 14514
rect 10961 14456 10966 14512
rect 11022 14456 16854 14512
rect 16910 14456 16915 14512
rect 10961 14454 16915 14456
rect 10961 14451 11027 14454
rect 16849 14451 16915 14454
rect 5073 14378 5139 14381
rect 16757 14378 16823 14381
rect 5073 14376 16823 14378
rect 5073 14320 5078 14376
rect 5134 14320 16762 14376
rect 16818 14320 16823 14376
rect 5073 14318 16823 14320
rect 5073 14315 5139 14318
rect 16757 14315 16823 14318
rect 17769 14378 17835 14381
rect 21449 14378 21515 14381
rect 17769 14376 21515 14378
rect 17769 14320 17774 14376
rect 17830 14320 21454 14376
rect 21510 14320 21515 14376
rect 17769 14318 21515 14320
rect 17769 14315 17835 14318
rect 21449 14315 21515 14318
rect 8293 14242 8359 14245
rect 10961 14242 11027 14245
rect 8293 14240 11027 14242
rect 8293 14184 8298 14240
rect 8354 14184 10966 14240
rect 11022 14184 11027 14240
rect 8293 14182 11027 14184
rect 8293 14179 8359 14182
rect 10961 14179 11027 14182
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 6729 14106 6795 14109
rect 8661 14106 8727 14109
rect 6729 14104 8727 14106
rect 6729 14048 6734 14104
rect 6790 14048 8666 14104
rect 8722 14048 8727 14104
rect 6729 14046 8727 14048
rect 6729 14043 6795 14046
rect 8661 14043 8727 14046
rect 18873 14106 18939 14109
rect 22461 14106 22527 14109
rect 18873 14104 22527 14106
rect 18873 14048 18878 14104
rect 18934 14048 22466 14104
rect 22522 14048 22527 14104
rect 18873 14046 22527 14048
rect 18873 14043 18939 14046
rect 22461 14043 22527 14046
rect 0 13970 480 14000
rect 1485 13970 1551 13973
rect 0 13968 1551 13970
rect 0 13912 1490 13968
rect 1546 13912 1551 13968
rect 0 13910 1551 13912
rect 0 13880 480 13910
rect 1485 13907 1551 13910
rect 2129 13970 2195 13973
rect 2262 13970 2268 13972
rect 2129 13968 2268 13970
rect 2129 13912 2134 13968
rect 2190 13912 2268 13968
rect 2129 13910 2268 13912
rect 2129 13907 2195 13910
rect 2262 13908 2268 13910
rect 2332 13908 2338 13972
rect 8937 13970 9003 13973
rect 11329 13970 11395 13973
rect 8937 13968 11395 13970
rect 8937 13912 8942 13968
rect 8998 13912 11334 13968
rect 11390 13912 11395 13968
rect 8937 13910 11395 13912
rect 8937 13907 9003 13910
rect 11329 13907 11395 13910
rect 19885 13970 19951 13973
rect 23289 13970 23355 13973
rect 19885 13968 23355 13970
rect 19885 13912 19890 13968
rect 19946 13912 23294 13968
rect 23350 13912 23355 13968
rect 19885 13910 23355 13912
rect 19885 13907 19951 13910
rect 23289 13907 23355 13910
rect 25681 13970 25747 13973
rect 27520 13970 28000 14000
rect 25681 13968 28000 13970
rect 25681 13912 25686 13968
rect 25742 13912 28000 13968
rect 25681 13910 28000 13912
rect 25681 13907 25747 13910
rect 27520 13880 28000 13910
rect 8569 13834 8635 13837
rect 11421 13834 11487 13837
rect 8569 13832 11487 13834
rect 8569 13776 8574 13832
rect 8630 13776 11426 13832
rect 11482 13776 11487 13832
rect 8569 13774 11487 13776
rect 8569 13771 8635 13774
rect 11421 13771 11487 13774
rect 20621 13834 20687 13837
rect 22277 13834 22343 13837
rect 20621 13832 22343 13834
rect 20621 13776 20626 13832
rect 20682 13776 22282 13832
rect 22338 13776 22343 13832
rect 20621 13774 22343 13776
rect 20621 13771 20687 13774
rect 22277 13771 22343 13774
rect 23105 13834 23171 13837
rect 24853 13834 24919 13837
rect 23105 13832 24919 13834
rect 23105 13776 23110 13832
rect 23166 13776 24858 13832
rect 24914 13776 24919 13832
rect 23105 13774 24919 13776
rect 23105 13771 23171 13774
rect 24853 13771 24919 13774
rect 4153 13698 4219 13701
rect 10041 13698 10107 13701
rect 4153 13696 10107 13698
rect 4153 13640 4158 13696
rect 4214 13640 10046 13696
rect 10102 13640 10107 13696
rect 4153 13638 10107 13640
rect 4153 13635 4219 13638
rect 10041 13635 10107 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 7833 13426 7899 13429
rect 11789 13426 11855 13429
rect 7833 13424 11855 13426
rect 7833 13368 7838 13424
rect 7894 13368 11794 13424
rect 11850 13368 11855 13424
rect 7833 13366 11855 13368
rect 7833 13363 7899 13366
rect 11789 13363 11855 13366
rect 5165 13290 5231 13293
rect 8477 13290 8543 13293
rect 11053 13290 11119 13293
rect 5165 13288 11119 13290
rect 5165 13232 5170 13288
rect 5226 13232 8482 13288
rect 8538 13232 11058 13288
rect 11114 13232 11119 13288
rect 5165 13230 11119 13232
rect 5165 13227 5231 13230
rect 8477 13227 8543 13230
rect 11053 13227 11119 13230
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 6269 13018 6335 13021
rect 11513 13018 11579 13021
rect 6269 13016 9690 13018
rect 6269 12960 6274 13016
rect 6330 12984 9690 13016
rect 9768 13016 11579 13018
rect 9768 12984 11518 13016
rect 6330 12960 11518 12984
rect 11574 12960 11579 13016
rect 6269 12958 11579 12960
rect 6269 12955 6335 12958
rect 9630 12924 9828 12958
rect 11513 12955 11579 12958
rect 16573 13018 16639 13021
rect 21633 13018 21699 13021
rect 16573 13016 21699 13018
rect 16573 12960 16578 13016
rect 16634 12960 21638 13016
rect 21694 12960 21699 13016
rect 16573 12958 21699 12960
rect 16573 12955 16639 12958
rect 21633 12955 21699 12958
rect 0 12882 480 12912
rect 5533 12882 5599 12885
rect 0 12880 5599 12882
rect 0 12824 5538 12880
rect 5594 12824 5599 12880
rect 0 12822 5599 12824
rect 0 12792 480 12822
rect 5533 12819 5599 12822
rect 20805 12882 20871 12885
rect 24577 12882 24643 12885
rect 20805 12880 24643 12882
rect 20805 12824 20810 12880
rect 20866 12824 24582 12880
rect 24638 12824 24643 12880
rect 20805 12822 24643 12824
rect 20805 12819 20871 12822
rect 24577 12819 24643 12822
rect 25221 12882 25287 12885
rect 27520 12882 28000 12912
rect 25221 12880 28000 12882
rect 25221 12824 25226 12880
rect 25282 12824 28000 12880
rect 25221 12822 28000 12824
rect 25221 12819 25287 12822
rect 27520 12792 28000 12822
rect 2497 12746 2563 12749
rect 2497 12744 4354 12746
rect 2497 12688 2502 12744
rect 2558 12688 4354 12744
rect 2497 12686 4354 12688
rect 2497 12683 2563 12686
rect 4294 12610 4354 12686
rect 6177 12610 6243 12613
rect 4294 12608 6243 12610
rect 4294 12552 6182 12608
rect 6238 12552 6243 12608
rect 4294 12550 6243 12552
rect 6177 12547 6243 12550
rect 14365 12610 14431 12613
rect 17493 12610 17559 12613
rect 19333 12610 19399 12613
rect 14365 12608 19399 12610
rect 14365 12552 14370 12608
rect 14426 12552 17498 12608
rect 17554 12552 19338 12608
rect 19394 12552 19399 12608
rect 14365 12550 19399 12552
rect 14365 12547 14431 12550
rect 17493 12547 17559 12550
rect 19333 12547 19399 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 2405 12474 2471 12477
rect 5257 12474 5323 12477
rect 2405 12472 5323 12474
rect 2405 12416 2410 12472
rect 2466 12416 5262 12472
rect 5318 12416 5323 12472
rect 2405 12414 5323 12416
rect 2405 12411 2471 12414
rect 5257 12411 5323 12414
rect 13905 12338 13971 12341
rect 17033 12338 17099 12341
rect 18229 12338 18295 12341
rect 13905 12336 18295 12338
rect 13905 12280 13910 12336
rect 13966 12280 17038 12336
rect 17094 12280 18234 12336
rect 18290 12280 18295 12336
rect 13905 12278 18295 12280
rect 13905 12275 13971 12278
rect 17033 12275 17099 12278
rect 18229 12275 18295 12278
rect 19241 12338 19307 12341
rect 21541 12338 21607 12341
rect 19241 12336 21607 12338
rect 19241 12280 19246 12336
rect 19302 12280 21546 12336
rect 21602 12280 21607 12336
rect 19241 12278 21607 12280
rect 19241 12275 19307 12278
rect 21541 12275 21607 12278
rect 12249 12202 12315 12205
rect 13353 12202 13419 12205
rect 18045 12202 18111 12205
rect 22829 12202 22895 12205
rect 12249 12200 15394 12202
rect 12249 12144 12254 12200
rect 12310 12144 13358 12200
rect 13414 12144 15394 12200
rect 12249 12142 15394 12144
rect 12249 12139 12315 12142
rect 13353 12139 13419 12142
rect 7465 12066 7531 12069
rect 10593 12066 10659 12069
rect 7465 12064 10659 12066
rect 7465 12008 7470 12064
rect 7526 12008 10598 12064
rect 10654 12008 10659 12064
rect 7465 12006 10659 12008
rect 7465 12003 7531 12006
rect 10593 12003 10659 12006
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 15334 11930 15394 12142
rect 18045 12200 22895 12202
rect 18045 12144 18050 12200
rect 18106 12144 22834 12200
rect 22890 12144 22895 12200
rect 18045 12142 22895 12144
rect 18045 12139 18111 12142
rect 22829 12139 22895 12142
rect 24025 12202 24091 12205
rect 25405 12202 25471 12205
rect 24025 12200 25471 12202
rect 24025 12144 24030 12200
rect 24086 12144 25410 12200
rect 25466 12144 25471 12200
rect 24025 12142 25471 12144
rect 24025 12139 24091 12142
rect 25405 12139 25471 12142
rect 17309 12066 17375 12069
rect 21909 12066 21975 12069
rect 17309 12064 21975 12066
rect 17309 12008 17314 12064
rect 17370 12008 21914 12064
rect 21970 12008 21975 12064
rect 17309 12006 21975 12008
rect 17309 12003 17375 12006
rect 21909 12003 21975 12006
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 23841 11930 23907 11933
rect 15334 11928 23907 11930
rect 15334 11872 23846 11928
rect 23902 11872 23907 11928
rect 15334 11870 23907 11872
rect 23841 11867 23907 11870
rect 0 11794 480 11824
rect 2957 11794 3023 11797
rect 0 11792 3023 11794
rect 0 11736 2962 11792
rect 3018 11736 3023 11792
rect 0 11734 3023 11736
rect 0 11704 480 11734
rect 2957 11731 3023 11734
rect 11145 11794 11211 11797
rect 17401 11794 17467 11797
rect 11145 11792 17467 11794
rect 11145 11736 11150 11792
rect 11206 11736 17406 11792
rect 17462 11736 17467 11792
rect 11145 11734 17467 11736
rect 11145 11731 11211 11734
rect 17401 11731 17467 11734
rect 25405 11794 25471 11797
rect 27520 11794 28000 11824
rect 25405 11792 28000 11794
rect 25405 11736 25410 11792
rect 25466 11736 28000 11792
rect 25405 11734 28000 11736
rect 25405 11731 25471 11734
rect 27520 11704 28000 11734
rect 8753 11658 8819 11661
rect 14549 11658 14615 11661
rect 8753 11656 14615 11658
rect 8753 11600 8758 11656
rect 8814 11600 14554 11656
rect 14610 11600 14615 11656
rect 8753 11598 14615 11600
rect 8753 11595 8819 11598
rect 14549 11595 14615 11598
rect 14917 11658 14983 11661
rect 19057 11658 19123 11661
rect 14917 11656 19123 11658
rect 14917 11600 14922 11656
rect 14978 11600 19062 11656
rect 19118 11600 19123 11656
rect 14917 11598 19123 11600
rect 14917 11595 14983 11598
rect 19057 11595 19123 11598
rect 21081 11658 21147 11661
rect 24209 11658 24275 11661
rect 21081 11656 24275 11658
rect 21081 11600 21086 11656
rect 21142 11600 24214 11656
rect 24270 11600 24275 11656
rect 21081 11598 24275 11600
rect 21081 11595 21147 11598
rect 24209 11595 24275 11598
rect 2497 11522 2563 11525
rect 7189 11522 7255 11525
rect 2497 11520 7255 11522
rect 2497 11464 2502 11520
rect 2558 11464 7194 11520
rect 7250 11464 7255 11520
rect 2497 11462 7255 11464
rect 2497 11459 2563 11462
rect 7189 11459 7255 11462
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 10777 11386 10843 11389
rect 13905 11386 13971 11389
rect 10777 11384 13971 11386
rect 10777 11328 10782 11384
rect 10838 11328 13910 11384
rect 13966 11328 13971 11384
rect 10777 11326 13971 11328
rect 10777 11323 10843 11326
rect 13905 11323 13971 11326
rect 14365 11250 14431 11253
rect 15285 11250 15351 11253
rect 14365 11248 15351 11250
rect 14365 11192 14370 11248
rect 14426 11192 15290 11248
rect 15346 11192 15351 11248
rect 14365 11190 15351 11192
rect 14365 11187 14431 11190
rect 15285 11187 15351 11190
rect 19241 11250 19307 11253
rect 21265 11250 21331 11253
rect 19241 11248 21331 11250
rect 19241 11192 19246 11248
rect 19302 11192 21270 11248
rect 21326 11192 21331 11248
rect 19241 11190 21331 11192
rect 19241 11187 19307 11190
rect 21265 11187 21331 11190
rect 11513 11114 11579 11117
rect 15837 11114 15903 11117
rect 11513 11112 15903 11114
rect 11513 11056 11518 11112
rect 11574 11056 15842 11112
rect 15898 11056 15903 11112
rect 11513 11054 15903 11056
rect 11513 11051 11579 11054
rect 15837 11051 15903 11054
rect 5610 10912 5930 10913
rect 0 10842 480 10872
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 1761 10842 1827 10845
rect 15653 10842 15719 10845
rect 20161 10842 20227 10845
rect 20529 10842 20595 10845
rect 24761 10842 24827 10845
rect 27520 10842 28000 10872
rect 0 10840 1827 10842
rect 0 10784 1766 10840
rect 1822 10784 1827 10840
rect 0 10782 1827 10784
rect 0 10752 480 10782
rect 1761 10779 1827 10782
rect 15334 10840 20227 10842
rect 15334 10784 15658 10840
rect 15714 10784 20166 10840
rect 20222 10784 20227 10840
rect 15334 10782 20227 10784
rect 2037 10706 2103 10709
rect 7557 10706 7623 10709
rect 2037 10704 7623 10706
rect 2037 10648 2042 10704
rect 2098 10648 7562 10704
rect 7618 10648 7623 10704
rect 2037 10646 7623 10648
rect 2037 10643 2103 10646
rect 7557 10643 7623 10646
rect 9213 10706 9279 10709
rect 10869 10706 10935 10709
rect 9213 10704 10935 10706
rect 9213 10648 9218 10704
rect 9274 10648 10874 10704
rect 10930 10648 10935 10704
rect 9213 10646 10935 10648
rect 9213 10643 9279 10646
rect 10869 10643 10935 10646
rect 13537 10706 13603 10709
rect 15334 10706 15394 10782
rect 15653 10779 15719 10782
rect 20161 10779 20227 10782
rect 20302 10840 24042 10842
rect 20302 10784 20534 10840
rect 20590 10784 24042 10840
rect 20302 10782 24042 10784
rect 20302 10706 20362 10782
rect 20529 10779 20595 10782
rect 13537 10704 15394 10706
rect 13537 10648 13542 10704
rect 13598 10648 15394 10704
rect 13537 10646 15394 10648
rect 15886 10646 20362 10706
rect 23982 10706 24042 10782
rect 24761 10840 28000 10842
rect 24761 10784 24766 10840
rect 24822 10784 28000 10840
rect 24761 10782 28000 10784
rect 24761 10779 24827 10782
rect 27520 10752 28000 10782
rect 25221 10706 25287 10709
rect 23982 10704 25287 10706
rect 23982 10648 25226 10704
rect 25282 10648 25287 10704
rect 23982 10646 25287 10648
rect 13537 10643 13603 10646
rect 3785 10570 3851 10573
rect 8845 10570 8911 10573
rect 3785 10568 8911 10570
rect 3785 10512 3790 10568
rect 3846 10512 8850 10568
rect 8906 10512 8911 10568
rect 3785 10510 8911 10512
rect 3785 10507 3851 10510
rect 8845 10507 8911 10510
rect 13721 10570 13787 10573
rect 15886 10570 15946 10646
rect 25221 10643 25287 10646
rect 13721 10568 15946 10570
rect 13721 10512 13726 10568
rect 13782 10512 15946 10568
rect 13721 10510 15946 10512
rect 16021 10570 16087 10573
rect 20253 10570 20319 10573
rect 22645 10570 22711 10573
rect 16021 10568 22711 10570
rect 16021 10512 16026 10568
rect 16082 10512 20258 10568
rect 20314 10512 22650 10568
rect 22706 10512 22711 10568
rect 16021 10510 22711 10512
rect 13721 10507 13787 10510
rect 16021 10507 16087 10510
rect 20253 10507 20319 10510
rect 22645 10507 22711 10510
rect 13721 10434 13787 10437
rect 16849 10434 16915 10437
rect 13721 10432 16915 10434
rect 13721 10376 13726 10432
rect 13782 10376 16854 10432
rect 16910 10376 16915 10432
rect 13721 10374 16915 10376
rect 13721 10371 13787 10374
rect 16849 10371 16915 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 15561 10162 15627 10165
rect 17953 10162 18019 10165
rect 15561 10160 18019 10162
rect 15561 10104 15566 10160
rect 15622 10104 17958 10160
rect 18014 10104 18019 10160
rect 15561 10102 18019 10104
rect 15561 10099 15627 10102
rect 17953 10099 18019 10102
rect 2497 9890 2563 9893
rect 3417 9890 3483 9893
rect 2497 9888 3483 9890
rect 2497 9832 2502 9888
rect 2558 9832 3422 9888
rect 3478 9832 3483 9888
rect 2497 9830 3483 9832
rect 2497 9827 2563 9830
rect 3417 9827 3483 9830
rect 5610 9824 5930 9825
rect 0 9754 480 9784
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 1485 9754 1551 9757
rect 0 9752 1551 9754
rect 0 9696 1490 9752
rect 1546 9696 1551 9752
rect 0 9694 1551 9696
rect 0 9664 480 9694
rect 1485 9691 1551 9694
rect 10685 9754 10751 9757
rect 10869 9754 10935 9757
rect 14641 9754 14707 9757
rect 10685 9752 10794 9754
rect 10685 9696 10690 9752
rect 10746 9696 10794 9752
rect 10685 9691 10794 9696
rect 10869 9752 14707 9754
rect 10869 9696 10874 9752
rect 10930 9696 14646 9752
rect 14702 9696 14707 9752
rect 10869 9694 14707 9696
rect 10869 9691 10935 9694
rect 14641 9691 14707 9694
rect 16297 9754 16363 9757
rect 20897 9754 20963 9757
rect 16297 9752 20963 9754
rect 16297 9696 16302 9752
rect 16358 9696 20902 9752
rect 20958 9696 20963 9752
rect 16297 9694 20963 9696
rect 16297 9691 16363 9694
rect 20897 9691 20963 9694
rect 21633 9754 21699 9757
rect 23749 9754 23815 9757
rect 21633 9752 23815 9754
rect 21633 9696 21638 9752
rect 21694 9696 23754 9752
rect 23810 9696 23815 9752
rect 21633 9694 23815 9696
rect 21633 9691 21699 9694
rect 23749 9691 23815 9694
rect 24761 9754 24827 9757
rect 27520 9754 28000 9784
rect 24761 9752 28000 9754
rect 24761 9696 24766 9752
rect 24822 9696 28000 9752
rect 24761 9694 28000 9696
rect 24761 9691 24827 9694
rect 10734 9621 10794 9691
rect 27520 9664 28000 9694
rect 2129 9618 2195 9621
rect 1902 9616 2195 9618
rect 1902 9560 2134 9616
rect 2190 9560 2195 9616
rect 1902 9558 2195 9560
rect 1902 9077 1962 9558
rect 2129 9555 2195 9558
rect 4889 9618 4955 9621
rect 9673 9618 9739 9621
rect 4889 9616 9739 9618
rect 4889 9560 4894 9616
rect 4950 9560 9678 9616
rect 9734 9560 9739 9616
rect 4889 9558 9739 9560
rect 4889 9555 4955 9558
rect 9673 9555 9739 9558
rect 10685 9616 10794 9621
rect 10685 9560 10690 9616
rect 10746 9560 10794 9616
rect 10685 9558 10794 9560
rect 13629 9618 13695 9621
rect 20069 9618 20135 9621
rect 13629 9616 20135 9618
rect 13629 9560 13634 9616
rect 13690 9560 20074 9616
rect 20130 9560 20135 9616
rect 13629 9558 20135 9560
rect 10685 9555 10751 9558
rect 13629 9555 13695 9558
rect 20069 9555 20135 9558
rect 4245 9482 4311 9485
rect 7281 9482 7347 9485
rect 4245 9480 7347 9482
rect 4245 9424 4250 9480
rect 4306 9424 7286 9480
rect 7342 9424 7347 9480
rect 4245 9422 7347 9424
rect 4245 9419 4311 9422
rect 7281 9419 7347 9422
rect 11237 9482 11303 9485
rect 14181 9482 14247 9485
rect 11237 9480 14247 9482
rect 11237 9424 11242 9480
rect 11298 9424 14186 9480
rect 14242 9424 14247 9480
rect 11237 9422 14247 9424
rect 11237 9419 11303 9422
rect 14181 9419 14247 9422
rect 2773 9346 2839 9349
rect 7005 9346 7071 9349
rect 2773 9344 7071 9346
rect 2773 9288 2778 9344
rect 2834 9288 7010 9344
rect 7066 9288 7071 9344
rect 2773 9286 7071 9288
rect 2773 9283 2839 9286
rect 7005 9283 7071 9286
rect 20805 9346 20871 9349
rect 26325 9346 26391 9349
rect 20805 9344 26391 9346
rect 20805 9288 20810 9344
rect 20866 9288 26330 9344
rect 26386 9288 26391 9344
rect 20805 9286 26391 9288
rect 20805 9283 20871 9286
rect 26325 9283 26391 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 2313 9210 2379 9213
rect 4429 9210 4495 9213
rect 2313 9208 4495 9210
rect 2313 9152 2318 9208
rect 2374 9152 4434 9208
rect 4490 9152 4495 9208
rect 2313 9150 4495 9152
rect 2313 9147 2379 9150
rect 4429 9147 4495 9150
rect 1853 9072 1962 9077
rect 1853 9016 1858 9072
rect 1914 9016 1962 9072
rect 1853 9014 1962 9016
rect 2129 9074 2195 9077
rect 4429 9074 4495 9077
rect 2129 9072 4495 9074
rect 2129 9016 2134 9072
rect 2190 9016 4434 9072
rect 4490 9016 4495 9072
rect 2129 9014 4495 9016
rect 1853 9011 1919 9014
rect 2129 9011 2195 9014
rect 4429 9011 4495 9014
rect 18505 9074 18571 9077
rect 20989 9074 21055 9077
rect 18505 9072 21055 9074
rect 18505 9016 18510 9072
rect 18566 9016 20994 9072
rect 21050 9016 21055 9072
rect 18505 9014 21055 9016
rect 18505 9011 18571 9014
rect 20989 9011 21055 9014
rect 3233 8938 3299 8941
rect 3601 8938 3667 8941
rect 10133 8938 10199 8941
rect 3233 8936 10199 8938
rect 3233 8880 3238 8936
rect 3294 8880 3606 8936
rect 3662 8880 10138 8936
rect 10194 8880 10199 8936
rect 3233 8878 10199 8880
rect 3233 8875 3299 8878
rect 3601 8875 3667 8878
rect 10133 8875 10199 8878
rect 0 8802 480 8832
rect 1577 8802 1643 8805
rect 0 8800 1643 8802
rect 0 8744 1582 8800
rect 1638 8744 1643 8800
rect 0 8742 1643 8744
rect 0 8712 480 8742
rect 1577 8739 1643 8742
rect 24761 8802 24827 8805
rect 27520 8802 28000 8832
rect 24761 8800 28000 8802
rect 24761 8744 24766 8800
rect 24822 8744 28000 8800
rect 24761 8742 28000 8744
rect 24761 8739 24827 8742
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 27520 8712 28000 8742
rect 24277 8671 24597 8672
rect 2865 8530 2931 8533
rect 8477 8530 8543 8533
rect 11145 8530 11211 8533
rect 12617 8530 12683 8533
rect 2865 8528 8586 8530
rect 2865 8472 2870 8528
rect 2926 8472 8482 8528
rect 8538 8472 8586 8528
rect 2865 8470 8586 8472
rect 2865 8467 2931 8470
rect 8477 8467 8586 8470
rect 11145 8528 12683 8530
rect 11145 8472 11150 8528
rect 11206 8472 12622 8528
rect 12678 8472 12683 8528
rect 11145 8470 12683 8472
rect 11145 8467 11211 8470
rect 12617 8467 12683 8470
rect 8526 8394 8586 8467
rect 16757 8394 16823 8397
rect 8526 8392 16823 8394
rect 8526 8336 16762 8392
rect 16818 8336 16823 8392
rect 8526 8334 16823 8336
rect 16757 8331 16823 8334
rect 14733 8258 14799 8261
rect 17493 8258 17559 8261
rect 14733 8256 17559 8258
rect 14733 8200 14738 8256
rect 14794 8200 17498 8256
rect 17554 8200 17559 8256
rect 14733 8198 17559 8200
rect 14733 8195 14799 8198
rect 17493 8195 17559 8198
rect 21173 8258 21239 8261
rect 23473 8258 23539 8261
rect 21173 8256 23539 8258
rect 21173 8200 21178 8256
rect 21234 8200 23478 8256
rect 23534 8200 23539 8256
rect 21173 8198 23539 8200
rect 21173 8195 21239 8198
rect 23473 8195 23539 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 16665 8122 16731 8125
rect 15886 8120 16731 8122
rect 15886 8064 16670 8120
rect 16726 8064 16731 8120
rect 15886 8062 16731 8064
rect 10317 7986 10383 7989
rect 15886 7986 15946 8062
rect 16665 8059 16731 8062
rect 10317 7984 15946 7986
rect 10317 7928 10322 7984
rect 10378 7928 15946 7984
rect 10317 7926 15946 7928
rect 16113 7986 16179 7989
rect 21449 7986 21515 7989
rect 16113 7984 21515 7986
rect 16113 7928 16118 7984
rect 16174 7928 21454 7984
rect 21510 7928 21515 7984
rect 16113 7926 21515 7928
rect 10317 7923 10383 7926
rect 16113 7923 16179 7926
rect 21449 7923 21515 7926
rect 0 7714 480 7744
rect 1393 7714 1459 7717
rect 0 7712 1459 7714
rect 0 7656 1398 7712
rect 1454 7656 1459 7712
rect 0 7654 1459 7656
rect 0 7624 480 7654
rect 1393 7651 1459 7654
rect 24669 7714 24735 7717
rect 27520 7714 28000 7744
rect 24669 7712 28000 7714
rect 24669 7656 24674 7712
rect 24730 7656 28000 7712
rect 24669 7654 28000 7656
rect 24669 7651 24735 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 27520 7624 28000 7654
rect 24277 7583 24597 7584
rect 5073 7306 5139 7309
rect 15377 7306 15443 7309
rect 5073 7304 15443 7306
rect 5073 7248 5078 7304
rect 5134 7248 15382 7304
rect 15438 7248 15443 7304
rect 5073 7246 15443 7248
rect 5073 7243 5139 7246
rect 15377 7243 15443 7246
rect 21541 7170 21607 7173
rect 24853 7170 24919 7173
rect 21541 7168 24919 7170
rect 21541 7112 21546 7168
rect 21602 7112 24858 7168
rect 24914 7112 24919 7168
rect 21541 7110 24919 7112
rect 21541 7107 21607 7110
rect 24853 7107 24919 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 2589 7034 2655 7037
rect 4797 7034 4863 7037
rect 2589 7032 4863 7034
rect 2589 6976 2594 7032
rect 2650 6976 4802 7032
rect 4858 6976 4863 7032
rect 2589 6974 4863 6976
rect 2589 6971 2655 6974
rect 4797 6971 4863 6974
rect 2037 6898 2103 6901
rect 5073 6898 5139 6901
rect 6361 6898 6427 6901
rect 2037 6896 6427 6898
rect 2037 6840 2042 6896
rect 2098 6840 5078 6896
rect 5134 6840 6366 6896
rect 6422 6840 6427 6896
rect 2037 6838 6427 6840
rect 2037 6835 2103 6838
rect 5073 6835 5139 6838
rect 6361 6835 6427 6838
rect 10317 6898 10383 6901
rect 13261 6898 13327 6901
rect 10317 6896 13327 6898
rect 10317 6840 10322 6896
rect 10378 6840 13266 6896
rect 13322 6840 13327 6896
rect 10317 6838 13327 6840
rect 10317 6835 10383 6838
rect 13261 6835 13327 6838
rect 23565 6898 23631 6901
rect 23565 6896 24778 6898
rect 23565 6840 23570 6896
rect 23626 6840 24778 6896
rect 23565 6838 24778 6840
rect 23565 6835 23631 6838
rect 9581 6762 9647 6765
rect 16481 6762 16547 6765
rect 9581 6760 16547 6762
rect 9581 6704 9586 6760
rect 9642 6704 16486 6760
rect 16542 6704 16547 6760
rect 9581 6702 16547 6704
rect 9581 6699 9647 6702
rect 16481 6699 16547 6702
rect 0 6626 480 6656
rect 1485 6626 1551 6629
rect 0 6624 1551 6626
rect 0 6568 1490 6624
rect 1546 6568 1551 6624
rect 0 6566 1551 6568
rect 24718 6626 24778 6838
rect 27520 6626 28000 6656
rect 24718 6566 28000 6626
rect 0 6536 480 6566
rect 1485 6563 1551 6566
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 27520 6536 28000 6566
rect 24277 6495 24597 6496
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 2589 5946 2655 5949
rect 5349 5946 5415 5949
rect 2589 5944 5415 5946
rect 2589 5888 2594 5944
rect 2650 5888 5354 5944
rect 5410 5888 5415 5944
rect 2589 5886 5415 5888
rect 2589 5883 2655 5886
rect 5349 5883 5415 5886
rect 2497 5810 2563 5813
rect 4889 5810 4955 5813
rect 2497 5808 4955 5810
rect 2497 5752 2502 5808
rect 2558 5752 4894 5808
rect 4950 5752 4955 5808
rect 2497 5750 4955 5752
rect 2497 5747 2563 5750
rect 4889 5747 4955 5750
rect 0 5674 480 5704
rect 1393 5674 1459 5677
rect 0 5672 1459 5674
rect 0 5616 1398 5672
rect 1454 5616 1459 5672
rect 0 5614 1459 5616
rect 0 5584 480 5614
rect 1393 5611 1459 5614
rect 23933 5674 23999 5677
rect 27520 5674 28000 5704
rect 23933 5672 28000 5674
rect 23933 5616 23938 5672
rect 23994 5616 28000 5672
rect 23933 5614 28000 5616
rect 23933 5611 23999 5614
rect 27520 5584 28000 5614
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 0 4586 480 4616
rect 1393 4586 1459 4589
rect 0 4584 1459 4586
rect 0 4528 1398 4584
rect 1454 4528 1459 4584
rect 0 4526 1459 4528
rect 0 4496 480 4526
rect 1393 4523 1459 4526
rect 24761 4586 24827 4589
rect 27520 4586 28000 4616
rect 24761 4584 28000 4586
rect 24761 4528 24766 4584
rect 24822 4528 28000 4584
rect 24761 4526 28000 4528
rect 24761 4523 24827 4526
rect 27520 4496 28000 4526
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 4521 4042 4587 4045
rect 11237 4042 11303 4045
rect 4521 4040 11303 4042
rect 4521 3984 4526 4040
rect 4582 3984 11242 4040
rect 11298 3984 11303 4040
rect 4521 3982 11303 3984
rect 4521 3979 4587 3982
rect 11237 3979 11303 3982
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 3325 3634 3391 3637
rect 1396 3632 3391 3634
rect 1396 3576 3330 3632
rect 3386 3576 3391 3632
rect 1396 3574 3391 3576
rect 0 3498 480 3528
rect 1396 3498 1456 3574
rect 3325 3571 3391 3574
rect 0 3438 1456 3498
rect 1577 3498 1643 3501
rect 11789 3498 11855 3501
rect 1577 3496 11855 3498
rect 1577 3440 1582 3496
rect 1638 3440 11794 3496
rect 11850 3440 11855 3496
rect 1577 3438 11855 3440
rect 0 3408 480 3438
rect 1577 3435 1643 3438
rect 11789 3435 11855 3438
rect 13077 3498 13143 3501
rect 23197 3498 23263 3501
rect 13077 3496 23263 3498
rect 13077 3440 13082 3496
rect 13138 3440 23202 3496
rect 23258 3440 23263 3496
rect 13077 3438 23263 3440
rect 13077 3435 13143 3438
rect 23197 3435 23263 3438
rect 23473 3498 23539 3501
rect 27520 3498 28000 3528
rect 23473 3496 28000 3498
rect 23473 3440 23478 3496
rect 23534 3440 28000 3496
rect 23473 3438 28000 3440
rect 23473 3435 23539 3438
rect 27520 3408 28000 3438
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 25129 2818 25195 2821
rect 25086 2816 25195 2818
rect 25086 2760 25134 2816
rect 25190 2760 25195 2816
rect 25086 2755 25195 2760
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 0 2546 480 2576
rect 1393 2546 1459 2549
rect 0 2544 1459 2546
rect 0 2488 1398 2544
rect 1454 2488 1459 2544
rect 0 2486 1459 2488
rect 25086 2546 25146 2755
rect 27520 2546 28000 2576
rect 25086 2486 28000 2546
rect 0 2456 480 2486
rect 1393 2483 1459 2486
rect 27520 2456 28000 2486
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 0 1458 480 1488
rect 1485 1458 1551 1461
rect 0 1456 1551 1458
rect 0 1400 1490 1456
rect 1546 1400 1551 1456
rect 0 1398 1551 1400
rect 0 1368 480 1398
rect 1485 1395 1551 1398
rect 25589 1458 25655 1461
rect 27520 1458 28000 1488
rect 25589 1456 28000 1458
rect 25589 1400 25594 1456
rect 25650 1400 28000 1456
rect 25589 1398 28000 1400
rect 25589 1395 25655 1398
rect 27520 1368 28000 1398
rect 0 506 480 536
rect 2773 506 2839 509
rect 0 504 2839 506
rect 0 448 2778 504
rect 2834 448 2839 504
rect 0 446 2839 448
rect 0 416 480 446
rect 2773 443 2839 446
rect 24669 506 24735 509
rect 27520 506 28000 536
rect 24669 504 28000 506
rect 24669 448 24674 504
rect 24730 448 28000 504
rect 24669 446 28000 448
rect 24669 443 24735 446
rect 27520 416 28000 446
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 16620 20224 16684 20228
rect 16620 20168 16670 20224
rect 16670 20168 16684 20224
rect 16620 20164 16684 20168
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 19380 17776 19444 17780
rect 19380 17720 19430 17776
rect 19430 17720 19444 17776
rect 19380 17716 19444 17720
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 19334 14724 19398 14788
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 2268 13908 2332 13972
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 16619 20228 16685 20229
rect 16619 20164 16620 20228
rect 16684 20164 16685 20228
rect 16619 20163 16685 20164
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 16622 14058 16682 20163
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19379 17780 19445 17781
rect 19379 17716 19380 17780
rect 19444 17716 19445 17780
rect 19379 17715 19445 17716
rect 19382 15330 19442 17715
rect 19336 15270 19442 15330
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19336 14789 19396 15270
rect 19333 14788 19399 14789
rect 19333 14724 19334 14788
rect 19398 14724 19399 14788
rect 19333 14723 19399 14724
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
<< via4 >>
rect 2182 13972 2418 14058
rect 2182 13908 2268 13972
rect 2268 13908 2332 13972
rect 2332 13908 2418 13972
rect 2182 13822 2418 13908
rect 16534 13822 16770 14058
<< metal5 >>
rect 2140 14058 16812 14100
rect 2140 13822 2182 14058
rect 2418 13822 16534 14058
rect 16770 13822 16812 14058
rect 2140 13780 16812 13822
use scs8hd_fill_2  FILLER_1_6 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1656 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_6
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_6_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_5_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_17
timestamp 1586364061
transform 1 0 2668 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_10 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_10 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2024 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2852 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_21 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3036 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_29
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_22
timestamp 1586364061
transform 1 0 3128 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_34
timestamp 1586364061
transform 1 0 4232 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_46
timestamp 1586364061
transform 1 0 5336 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_1_58
timestamp 1586364061
transform 1 0 6440 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_87
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_118
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_110
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_211
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_242
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_258
timestamp 1586364061
transform 1 0 24840 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_253
timestamp 1586364061
transform 1 0 24380 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_256
timestamp 1586364061
transform 1 0 24656 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_252
timestamp 1586364061
transform 1 0 24288 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24472 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_0_267
timestamp 1586364061
transform 1 0 25668 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_263
timestamp 1586364061
transform 1 0 25300 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25484 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25024 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_262
timestamp 1586364061
transform 1 0 25208 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_275
timestamp 1586364061
transform 1 0 26404 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_274
timestamp 1586364061
transform 1 0 26312 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_141
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_276 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_7
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_19
timestamp 1586364061
transform 1 0 2852 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_31
timestamp 1586364061
transform 1 0 3956 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_43
timestamp 1586364061
transform 1 0 5060 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_3_55
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 590 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_110
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_171
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_220
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_232
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_6
timestamp 1586364061
transform 1 0 1656 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_18
timestamp 1586364061
transform 1 0 2760 0 -1 4896
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_4_30
timestamp 1586364061
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_141
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_166
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_178
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_190
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_239
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_263
timestamp 1586364061
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2576 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_6
timestamp 1586364061
transform 1 0 1656 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_10
timestamp 1586364061
transform 1 0 2024 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_14
timestamp 1586364061
transform 1 0 2392 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_18
timestamp 1586364061
transform 1 0 2760 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_30
timestamp 1586364061
transform 1 0 3864 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_42
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_decap_6  FILLER_5_54
timestamp 1586364061
transform 1 0 6072 0 1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_5_60
timestamp 1586364061
transform 1 0 6624 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_147
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_159
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_171
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_196
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_220
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_232
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_7
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_6
timestamp 1586364061
transform 1 0 1656 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use scs8hd_buf_2  _190_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_11
timestamp 1586364061
transform 1 0 2116 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 2300 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 -1 5984
box -38 -48 314 592
use scs8hd_conb_1  _174_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_17
timestamp 1586364061
transform 1 0 2668 0 -1 5984
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3496 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3312 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_29
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_7_18
timestamp 1586364061
transform 1 0 2760 0 1 5984
box -38 -48 590 592
use scs8hd_decap_3  FILLER_7_29
timestamp 1586364061
transform 1 0 3772 0 1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_7_34
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5060 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_7_42
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_45
timestamp 1586364061
transform 1 0 5244 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_66
timestamp 1586364061
transform 1 0 7176 0 1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_69
timestamp 1586364061
transform 1 0 7452 0 1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8280 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_7_77
timestamp 1586364061
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_80
timestamp 1586364061
transform 1 0 8464 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_105
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_7_92
timestamp 1586364061
transform 1 0 9568 0 1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_7_98
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_101
timestamp 1586364061
transform 1 0 10396 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11316 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_109
timestamp 1586364061
transform 1 0 11132 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_7_113
timestamp 1586364061
transform 1 0 11500 0 1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_7_121
timestamp 1586364061
transform 1 0 12236 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_147
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_159
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_166
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_178
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_171
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_196
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_220
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_232
timestamp 1586364061
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_263
timestamp 1586364061
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_257
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use scs8hd_buf_2  _189_
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_7
timestamp 1586364061
transform 1 0 1748 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_13
timestamp 1586364061
transform 1 0 2300 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_16
timestamp 1586364061
transform 1 0 2576 0 -1 7072
box -38 -48 406 592
use scs8hd_conb_1  _175_
timestamp 1586364061
transform 1 0 2944 0 -1 7072
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_35
timestamp 1586364061
transform 1 0 4324 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5060 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4508 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_39
timestamp 1586364061
transform 1 0 4692 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_46
timestamp 1586364061
transform 1 0 5336 0 -1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7268 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_54
timestamp 1586364061
transform 1 0 6072 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_58
timestamp 1586364061
transform 1 0 6440 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_3  FILLER_8_64
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_70
timestamp 1586364061
transform 1 0 7544 0 -1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8280 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_81
timestamp 1586364061
transform 1 0 8556 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_8_89
timestamp 1586364061
transform 1 0 9292 0 -1 7072
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10212 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 590 592
use scs8hd_decap_8  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_110
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_114
timestamp 1586364061
transform 1 0 11592 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_119
timestamp 1586364061
transform 1 0 12052 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_131
timestamp 1586364061
transform 1 0 13156 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_143
timestamp 1586364061
transform 1 0 14260 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_151
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_166
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_190
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_202
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_251
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_263
timestamp 1586364061
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_buf_2  _191_
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 1932 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2300 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2668 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_7
timestamp 1586364061
transform 1 0 1748 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_11
timestamp 1586364061
transform 1 0 2116 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3312 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3128 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_19
timestamp 1586364061
transform 1 0 2852 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_33
timestamp 1586364061
transform 1 0 4140 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _130_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4876 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_37
timestamp 1586364061
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_50
timestamp 1586364061
transform 1 0 5704 0 1 7072
box -38 -48 406 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_54
timestamp 1586364061
transform 1 0 6072 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_71
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8832 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 9292 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_75
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_82
timestamp 1586364061
transform 1 0 8648 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_86
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10028 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10488 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_91
timestamp 1586364061
transform 1 0 9476 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_95
timestamp 1586364061
transform 1 0 9844 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_100
timestamp 1586364061
transform 1 0 10304 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_104
timestamp 1586364061
transform 1 0 10672 0 1 7072
box -38 -48 406 592
use scs8hd_buf_1  _120_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11040 0 1 7072
box -38 -48 314 592
use scs8hd_buf_1  _136_
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 11868 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 11500 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_111
timestamp 1586364061
transform 1 0 11316 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_115
timestamp 1586364061
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_119
timestamp 1586364061
transform 1 0 12052 0 1 7072
box -38 -48 314 592
use scs8hd_buf_1  _110_
timestamp 1586364061
transform 1 0 13708 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__096__B
timestamp 1586364061
transform 1 0 14168 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 12880 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_126
timestamp 1586364061
transform 1 0 12696 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_130
timestamp 1586364061
transform 1 0 13064 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_134
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_140
timestamp 1586364061
transform 1 0 13984 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15364 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 14536 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_144
timestamp 1586364061
transform 1 0 14352 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_148
timestamp 1586364061
transform 1 0 14720 0 1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_9_154
timestamp 1586364061
transform 1 0 15272 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_157
timestamp 1586364061
transform 1 0 15548 0 1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 17020 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__B
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_169
timestamp 1586364061
transform 1 0 16652 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_196
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19780 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_202
timestamp 1586364061
transform 1 0 19688 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_205
timestamp 1586364061
transform 1 0 19964 0 1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21068 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21436 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_219
timestamp 1586364061
transform 1 0 21252 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_223
timestamp 1586364061
transform 1 0 21620 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_235
timestamp 1586364061
transform 1 0 22724 0 1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_9_243
timestamp 1586364061
transform 1 0 23460 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_249
timestamp 1586364061
transform 1 0 24012 0 1 7072
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 1840 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_6
timestamp 1586364061
transform 1 0 1656 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_10
timestamp 1586364061
transform 1 0 2024 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_23
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4600 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5612 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_47
timestamp 1586364061
transform 1 0 5428 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_51
timestamp 1586364061
transform 1 0 5796 0 -1 8160
box -38 -48 406 592
use scs8hd_nor2_4  _134_
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7268 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_55
timestamp 1586364061
transform 1 0 6164 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_65
timestamp 1586364061
transform 1 0 7084 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_69
timestamp 1586364061
transform 1 0 7452 0 -1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7820 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_76
timestamp 1586364061
transform 1 0 8096 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_88
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 406 592
use scs8hd_nor2_4  _132_
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_102
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 1142 592
use scs8hd_or2_4  _118_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 682 592
use scs8hd_decap_3  FILLER_10_114
timestamp 1586364061
transform 1 0 11592 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_124
timestamp 1586364061
transform 1 0 12512 0 -1 8160
box -38 -48 1142 592
use scs8hd_or2_4  _096_
timestamp 1586364061
transform 1 0 13616 0 -1 8160
box -38 -48 682 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15364 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_143
timestamp 1586364061
transform 1 0 14260 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_147
timestamp 1586364061
transform 1 0 14628 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_158
timestamp 1586364061
transform 1 0 15640 0 -1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _113_
timestamp 1586364061
transform 1 0 17020 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16192 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_162
timestamp 1586364061
transform 1 0 16008 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_166
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_172
timestamp 1586364061
transform 1 0 16928 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 18216 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 18584 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_182
timestamp 1586364061
transform 1 0 17848 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_188
timestamp 1586364061
transform 1 0 18400 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_192
timestamp 1586364061
transform 1 0 18768 0 -1 8160
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_200
timestamp 1586364061
transform 1 0 19504 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_6  FILLER_10_206
timestamp 1586364061
transform 1 0 20056 0 -1 8160
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21068 0 -1 8160
box -38 -48 866 592
use scs8hd_fill_2  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_226
timestamp 1586364061
transform 1 0 21896 0 -1 8160
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23460 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_10_238
timestamp 1586364061
transform 1 0 23000 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_242
timestamp 1586364061
transform 1 0 23368 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_246
timestamp 1586364061
transform 1 0 23736 0 -1 8160
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_254
timestamp 1586364061
transform 1 0 24472 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_258
timestamp 1586364061
transform 1 0 24840 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_270
timestamp 1586364061
transform 1 0 25944 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_274
timestamp 1586364061
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_buf_2  _192_
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2668 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2116 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_13
timestamp 1586364061
transform 1 0 2300 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 4232 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_26
timestamp 1586364061
transform 1 0 3496 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_32
timestamp 1586364061
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_4_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4784 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 4600 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_36
timestamp 1586364061
transform 1 0 4416 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_51
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_73
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_77
timestamp 1586364061
transform 1 0 8188 0 1 8160
box -38 -48 406 592
use scs8hd_decap_3  FILLER_11_83
timestamp 1586364061
transform 1 0 8740 0 1 8160
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10764 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 10212 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_97
timestamp 1586364061
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_101
timestamp 1586364061
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use scs8hd_inv_8  _072_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_108
timestamp 1586364061
transform 1 0 11040 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_112
timestamp 1586364061
transform 1 0 11408 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _114_
timestamp 1586364061
transform 1 0 13984 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_132
timestamp 1586364061
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_136
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15548 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15272 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_149
timestamp 1586364061
transform 1 0 14812 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_153
timestamp 1586364061
transform 1 0 15180 0 1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_11_156
timestamp 1586364061
transform 1 0 15456 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 17480 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16560 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17112 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_166
timestamp 1586364061
transform 1 0 16376 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_170
timestamp 1586364061
transform 1 0 16744 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_176
timestamp 1586364061
transform 1 0 17296 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 18216 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_11_180
timestamp 1586364061
transform 1 0 17664 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_195
timestamp 1586364061
transform 1 0 19044 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20056 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20516 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 19228 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 19596 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_199
timestamp 1586364061
transform 1 0 19412 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_203
timestamp 1586364061
transform 1 0 19780 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_209
timestamp 1586364061
transform 1 0 20332 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_213
timestamp 1586364061
transform 1 0 20700 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21068 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20884 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22080 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_226
timestamp 1586364061
transform 1 0 21896 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_230
timestamp 1586364061
transform 1 0 22264 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_234
timestamp 1586364061
transform 1 0 22632 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_238
timestamp 1586364061
transform 1 0 23000 0 1 8160
box -38 -48 590 592
use scs8hd_decap_8  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 25392 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_253
timestamp 1586364061
transform 1 0 24380 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_258
timestamp 1586364061
transform 1 0 24840 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_262
timestamp 1586364061
transform 1 0 25208 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_266
timestamp 1586364061
transform 1 0 25576 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_11_274
timestamp 1586364061
transform 1 0 26312 0 1 8160
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 1840 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_6
timestamp 1586364061
transform 1 0 1656 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_10
timestamp 1586364061
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_5_.latch
timestamp 1586364061
transform 1 0 4784 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4508 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_36
timestamp 1586364061
transform 1 0 4416 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_39
timestamp 1586364061
transform 1 0 4692 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_51
timestamp 1586364061
transform 1 0 5796 0 -1 9248
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 -1 9248
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_12_59
timestamp 1586364061
transform 1 0 6532 0 -1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_73
timestamp 1586364061
transform 1 0 7820 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_77
timestamp 1586364061
transform 1 0 8188 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_88
timestamp 1586364061
transform 1 0 9200 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_104
timestamp 1586364061
transform 1 0 10672 0 -1 9248
box -38 -48 774 592
use scs8hd_inv_8  _117_
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__073__B
timestamp 1586364061
transform 1 0 11684 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_112
timestamp 1586364061
transform 1 0 11408 0 -1 9248
box -38 -48 314 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 13616 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 12880 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 13248 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_126
timestamp 1586364061
transform 1 0 12696 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_130
timestamp 1586364061
transform 1 0 13064 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_134
timestamp 1586364061
transform 1 0 13432 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 14628 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_149
timestamp 1586364061
transform 1 0 14812 0 -1 9248
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 1050 592
use scs8hd_decap_12  FILLER_12_165
timestamp 1586364061
transform 1 0 16284 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_12_177
timestamp 1586364061
transform 1 0 17388 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19044 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_189
timestamp 1586364061
transform 1 0 18492 0 -1 9248
box -38 -48 590 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 19228 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20240 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_206
timestamp 1586364061
transform 1 0 20056 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_210
timestamp 1586364061
transform 1 0 20424 0 -1 9248
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21896 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_224
timestamp 1586364061
transform 1 0 21712 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_228
timestamp 1586364061
transform 1 0 22080 0 -1 9248
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22448 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_12  FILLER_12_241
timestamp 1586364061
transform 1 0 23276 0 -1 9248
box -38 -48 1142 592
use scs8hd_buf_2  _201_
timestamp 1586364061
transform 1 0 24564 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_253
timestamp 1586364061
transform 1 0 24380 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_259
timestamp 1586364061
transform 1 0 24932 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_271
timestamp 1586364061
transform 1 0 26036 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_7
timestamp 1586364061
transform 1 0 1748 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 1564 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_16
timestamp 1586364061
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_12
timestamp 1586364061
transform 1 0 2208 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1932 0 -1 10336
box -38 -48 866 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 866 592
use scs8hd_fill_1  FILLER_14_26
timestamp 1586364061
transform 1 0 3496 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_22
timestamp 1586364061
transform 1 0 3128 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_18
timestamp 1586364061
transform 1 0 2760 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2944 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2760 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_29
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_34
timestamp 1586364061
transform 1 0 4232 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_29
timestamp 1586364061
transform 1 0 3772 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4048 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2944 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_3  FILLER_14_41
timestamp 1586364061
transform 1 0 4876 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_52
timestamp 1586364061
transform 1 0 5888 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_14_46
timestamp 1586364061
transform 1 0 5336 0 -1 10336
box -38 -48 590 592
use scs8hd_decap_3  FILLER_13_50
timestamp 1586364061
transform 1 0 5704 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_46
timestamp 1586364061
transform 1 0 5336 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5520 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4508 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 5980 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_6  FILLER_14_62
timestamp 1586364061
transform 1 0 6808 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_59
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_55
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_66
timestamp 1586364061
transform 1 0 7176 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6992 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7360 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7544 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7544 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_79
timestamp 1586364061
transform 1 0 8372 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_79
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_87
timestamp 1586364061
transform 1 0 9108 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_83
timestamp 1586364061
transform 1 0 8740 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_83
timestamp 1586364061
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8556 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 8924 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9108 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_13_96
timestamp 1586364061
transform 1 0 9936 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_14_106
timestamp 1586364061
transform 1 0 10856 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_14_102
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_100
timestamp 1586364061
transform 1 0 10304 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 10488 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 10672 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_114
timestamp 1586364061
transform 1 0 11592 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_113
timestamp 1586364061
transform 1 0 11500 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__135__D
timestamp 1586364061
transform 1 0 11408 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_118
timestamp 1586364061
transform 1 0 11960 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__C
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__C
timestamp 1586364061
transform 1 0 11776 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__C
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_or3_4  _149_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use scs8hd_nand3_4  _073_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12052 0 -1 10336
box -38 -48 1326 592
use scs8hd_fill_2  FILLER_13_132
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_133
timestamp 1586364061
transform 1 0 13340 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_136
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 13524 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_137
timestamp 1586364061
transform 1 0 13708 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 13892 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use scs8hd_buf_1  _128_
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 314 592
use scs8hd_buf_1  _166_
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_148
timestamp 1586364061
transform 1 0 14720 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_144
timestamp 1586364061
transform 1 0 14352 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_148
timestamp 1586364061
transform 1 0 14720 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_143
timestamp 1586364061
transform 1 0 14260 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 14904 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 14536 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 14536 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 14904 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_152
timestamp 1586364061
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_2_.latch
timestamp 1586364061
transform 1 0 15364 0 -1 10336
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15088 0 1 9248
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_14_166
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_167
timestamp 1586364061
transform 1 0 16468 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_163
timestamp 1586364061
transform 1 0 16100 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16652 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16560 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16284 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_174
timestamp 1586364061
transform 1 0 17112 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_170
timestamp 1586364061
transform 1 0 16744 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_178
timestamp 1586364061
transform 1 0 17480 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_174
timestamp 1586364061
transform 1 0 17112 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16928 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17296 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17480 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_3  FILLER_14_187
timestamp 1586364061
transform 1 0 18308 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_182
timestamp 1586364061
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18216 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17664 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_14_192
timestamp 1586364061
transform 1 0 18768 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_192
timestamp 1586364061
transform 1 0 18768 0 1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_13_188
timestamp 1586364061
transform 1 0 18400 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use scs8hd_conb_1  _177_
timestamp 1586364061
transform 1 0 18492 0 1 9248
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 19044 0 -1 10336
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 19504 0 1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 20700 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20424 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_197
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_211
timestamp 1586364061
transform 1 0 20516 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_206
timestamp 1586364061
transform 1 0 20056 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_212
timestamp 1586364061
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21252 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21068 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22264 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_215
timestamp 1586364061
transform 1 0 20884 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_228
timestamp 1586364061
transform 1 0 22080 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_224
timestamp 1586364061
transform 1 0 21712 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_228
timestamp 1586364061
transform 1 0 22080 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_235
timestamp 1586364061
transform 1 0 22724 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_8  FILLER_13_236
timestamp 1586364061
transform 1 0 22816 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_232
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22632 0 1 9248
box -38 -48 222 592
use scs8hd_conb_1  _178_
timestamp 1586364061
transform 1 0 22448 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_247
timestamp 1586364061
transform 1 0 23828 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_243
timestamp 1586364061
transform 1 0 23460 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_249
timestamp 1586364061
transform 1 0 24012 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24012 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23552 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_251
timestamp 1586364061
transform 1 0 24196 0 -1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 24380 0 1 9248
box -38 -48 222 592
use scs8hd_buf_2  _200_
timestamp 1586364061
transform 1 0 24564 0 1 9248
box -38 -48 406 592
use scs8hd_buf_2  _199_
timestamp 1586364061
transform 1 0 24564 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_259
timestamp 1586364061
transform 1 0 24932 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_259
timestamp 1586364061
transform 1 0 24932 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 25116 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 25116 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_263
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_263
timestamp 1586364061
transform 1 0 25300 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_275
timestamp 1586364061
transform 1 0 26404 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2024 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1840 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3036 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_19
timestamp 1586364061
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_23
timestamp 1586364061
transform 1 0 3220 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _138_
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_36
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_40
timestamp 1586364061
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7360 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6440 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6992 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_15_60
timestamp 1586364061
transform 1 0 6624 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_66
timestamp 1586364061
transform 1 0 7176 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _140_
timestamp 1586364061
transform 1 0 8924 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 8372 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 8740 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_77
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_81
timestamp 1586364061
transform 1 0 8556 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _139_
timestamp 1586364061
transform 1 0 10488 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 10304 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_94
timestamp 1586364061
transform 1 0 9752 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_98
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use scs8hd_or4_4  _127_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_111
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_115
timestamp 1586364061
transform 1 0 11684 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _115_
timestamp 1586364061
transform 1 0 14168 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__127__C
timestamp 1586364061
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 13800 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_132
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_136
timestamp 1586364061
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_140
timestamp 1586364061
transform 1 0 13984 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 15180 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__C
timestamp 1586364061
transform 1 0 15548 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_151
timestamp 1586364061
transform 1 0 14996 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_155
timestamp 1586364061
transform 1 0 15364 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__B
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_168
timestamp 1586364061
transform 1 0 16560 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_173
timestamp 1586364061
transform 1 0 17020 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_177
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 406 592
use scs8hd_nor2_4  _100_
timestamp 1586364061
transform 1 0 18492 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__100__B
timestamp 1586364061
transform 1 0 18308 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20424 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 19504 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_198
timestamp 1586364061
transform 1 0 19320 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_202
timestamp 1586364061
transform 1 0 19688 0 1 10336
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21436 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21804 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22356 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_219
timestamp 1586364061
transform 1 0 21252 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_223
timestamp 1586364061
transform 1 0 21620 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_227
timestamp 1586364061
transform 1 0 21988 0 1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_236
timestamp 1586364061
transform 1 0 22816 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_240
timestamp 1586364061
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use scs8hd_buf_2  _198_
timestamp 1586364061
transform 1 0 25208 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24656 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25024 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_254
timestamp 1586364061
transform 1 0 24472 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_258
timestamp 1586364061
transform 1 0 24840 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_266
timestamp 1586364061
transform 1 0 25576 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 25760 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_270
timestamp 1586364061
transform 1 0 25944 0 1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_15_276
timestamp 1586364061
transform 1 0 26496 0 1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1932 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1748 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4324 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2944 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_18
timestamp 1586364061
transform 1 0 2760 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_22
timestamp 1586364061
transform 1 0 3128 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_26
timestamp 1586364061
transform 1 0 3496 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_4_.latch
timestamp 1586364061
transform 1 0 4508 0 -1 11424
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_16_48
timestamp 1586364061
transform 1 0 5520 0 -1 11424
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6440 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7636 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_69
timestamp 1586364061
transform 1 0 7452 0 -1 11424
box -38 -48 222 592
use scs8hd_or2_4  _095_
timestamp 1586364061
transform 1 0 8188 0 -1 11424
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_73
timestamp 1586364061
transform 1 0 7820 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_84
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_88
timestamp 1586364061
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 10856 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_104
timestamp 1586364061
transform 1 0 10672 0 -1 11424
box -38 -48 222 592
use scs8hd_or4_4  _135_
timestamp 1586364061
transform 1 0 11776 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 11592 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_108
timestamp 1586364061
transform 1 0 11040 0 -1 11424
box -38 -48 590 592
use scs8hd_or3_4  _109_
timestamp 1586364061
transform 1 0 13340 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 12788 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__D
timestamp 1586364061
transform 1 0 13156 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_125
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_129
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_142
timestamp 1586364061
transform 1 0 14168 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15640 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 14352 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 14720 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15456 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_146
timestamp 1586364061
transform 1 0 14536 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_150
timestamp 1586364061
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use scs8hd_or2_4  _071_
timestamp 1586364061
transform 1 0 17204 0 -1 11424
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16652 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17020 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_167
timestamp 1586364061
transform 1 0 16468 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_171
timestamp 1586364061
transform 1 0 16836 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _098_
timestamp 1586364061
transform 1 0 18584 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 18032 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18400 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_182
timestamp 1586364061
transform 1 0 17848 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_186
timestamp 1586364061
transform 1 0 18216 0 -1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 19872 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_199
timestamp 1586364061
transform 1 0 19412 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_203
timestamp 1586364061
transform 1 0 19780 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_206
timestamp 1586364061
transform 1 0 20056 0 -1 11424
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21896 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_224
timestamp 1586364061
transform 1 0 21712 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_228
timestamp 1586364061
transform 1 0 22080 0 -1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23460 0 -1 11424
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22908 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_235
timestamp 1586364061
transform 1 0 22724 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 406 592
use scs8hd_buf_2  _197_
timestamp 1586364061
transform 1 0 25024 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_8  FILLER_16_252
timestamp 1586364061
transform 1 0 24288 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_8  FILLER_16_264
timestamp 1586364061
transform 1 0 25392 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_16_272
timestamp 1586364061
transform 1 0 26128 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2300 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2116 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_9
timestamp 1586364061
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 4324 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3956 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_22
timestamp 1586364061
transform 1 0 3128 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_26
timestamp 1586364061
transform 1 0 3496 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_29
timestamp 1586364061
transform 1 0 3772 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_33
timestamp 1586364061
transform 1 0 4140 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_5_.latch
timestamp 1586364061
transform 1 0 4508 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 5704 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_48
timestamp 1586364061
transform 1 0 5520 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_52
timestamp 1586364061
transform 1 0 5888 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 6072 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_56
timestamp 1586364061
transform 1 0 6256 0 1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9292 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8740 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_73
timestamp 1586364061
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_77
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_81
timestamp 1586364061
transform 1 0 8556 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_85
timestamp 1586364061
transform 1 0 8924 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 10764 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_100
timestamp 1586364061
transform 1 0 10304 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_104
timestamp 1586364061
transform 1 0 10672 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_107
timestamp 1586364061
transform 1 0 10948 0 1 11424
box -38 -48 222 592
use scs8hd_buf_1  _077_
timestamp 1586364061
transform 1 0 11316 0 1 11424
box -38 -48 314 592
use scs8hd_or4_4  _119_
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 11132 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__C
timestamp 1586364061
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 14168 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 13800 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_132
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_136
timestamp 1586364061
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_140
timestamp 1586364061
transform 1 0 13984 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _104_
timestamp 1586364061
transform 1 0 14352 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15364 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_153
timestamp 1586364061
transform 1 0 15180 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_157
timestamp 1586364061
transform 1 0 15548 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_2_.latch
timestamp 1586364061
transform 1 0 15916 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__090__B
timestamp 1586364061
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_172
timestamp 1586364061
transform 1 0 16928 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_176
timestamp 1586364061
transform 1 0 17296 0 1 11424
box -38 -48 130 592
use scs8hd_nor2_4  _090_
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_179
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_193
timestamp 1586364061
transform 1 0 18860 0 1 11424
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_5_.latch
timestamp 1586364061
transform 1 0 19872 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19688 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19320 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_197
timestamp 1586364061
transform 1 0 19228 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_200
timestamp 1586364061
transform 1 0 19504 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_4_.latch
timestamp 1586364061
transform 1 0 21804 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 21620 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21252 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_215
timestamp 1586364061
transform 1 0 20884 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_221
timestamp 1586364061
transform 1 0 21436 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_236
timestamp 1586364061
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_240
timestamp 1586364061
transform 1 0 23184 0 1 11424
box -38 -48 222 592
use scs8hd_buf_2  _193_
timestamp 1586364061
transform 1 0 25208 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24656 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25024 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_254
timestamp 1586364061
transform 1 0 24472 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_258
timestamp 1586364061
transform 1 0 24840 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_266
timestamp 1586364061
transform 1 0 25576 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 25760 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_270
timestamp 1586364061
transform 1 0 25944 0 1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_17_276
timestamp 1586364061
transform 1 0 26496 0 1 11424
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2300 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2024 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1656 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_8
timestamp 1586364061
transform 1 0 1840 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_12
timestamp 1586364061
transform 1 0 2208 0 -1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_22
timestamp 1586364061
transform 1 0 3128 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_28
timestamp 1586364061
transform 1 0 3680 0 -1 12512
box -38 -48 130 592
use scs8hd_nor2_4  _137_
timestamp 1586364061
transform 1 0 5612 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 5336 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_41
timestamp 1586364061
transform 1 0 4876 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_45
timestamp 1586364061
transform 1 0 5244 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_48
timestamp 1586364061
transform 1 0 5520 0 -1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_58
timestamp 1586364061
transform 1 0 6440 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_3  FILLER_18_64
timestamp 1586364061
transform 1 0 6992 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9292 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_76
timestamp 1586364061
transform 1 0 8096 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_87
timestamp 1586364061
transform 1 0 9108 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_91
timestamp 1586364061
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 1142 592
use scs8hd_nor2_4  _108_
timestamp 1586364061
transform 1 0 12052 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 11592 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_116
timestamp 1586364061
transform 1 0 11776 0 -1 12512
box -38 -48 314 592
use scs8hd_nor2_4  _102_
timestamp 1586364061
transform 1 0 13616 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__119__D
timestamp 1586364061
transform 1 0 13064 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__C
timestamp 1586364061
transform 1 0 13432 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_128
timestamp 1586364061
transform 1 0 12880 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_132
timestamp 1586364061
transform 1 0 13248 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15640 0 -1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__106__B
timestamp 1586364061
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15456 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_149
timestamp 1586364061
transform 1 0 14812 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_169
timestamp 1586364061
transform 1 0 16652 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_173
timestamp 1586364061
transform 1 0 17020 0 -1 12512
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_3_.latch
timestamp 1586364061
transform 1 0 17848 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_181
timestamp 1586364061
transform 1 0 17756 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_193
timestamp 1586364061
transform 1 0 18860 0 -1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__074__B
timestamp 1586364061
transform 1 0 20240 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_197
timestamp 1586364061
transform 1 0 19228 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_18_206
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_210
timestamp 1586364061
transform 1 0 20424 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21160 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22172 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_231
timestamp 1586364061
transform 1 0 22356 0 -1 12512
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22724 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23736 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_244
timestamp 1586364061
transform 1 0 23552 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_248
timestamp 1586364061
transform 1 0 23920 0 -1 12512
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24288 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_12  FILLER_18_261
timestamp 1586364061
transform 1 0 25116 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_273
timestamp 1586364061
transform 1 0 26220 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_20_7
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1840 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 1564 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2024 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2024 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_19
timestamp 1586364061
transform 1 0 2852 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_23
timestamp 1586364061
transform 1 0 3220 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_19
timestamp 1586364061
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3036 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3772 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _121_
timestamp 1586364061
transform 1 0 4600 0 -1 13600
box -38 -48 866 592
use scs8hd_buf_2  _188_
timestamp 1586364061
transform 1 0 5336 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 4416 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_38
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_42
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_50
timestamp 1586364061
transform 1 0 5704 0 1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_47
timestamp 1586364061
transform 1 0 5428 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_20_59
timestamp 1586364061
transform 1 0 6532 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_54
timestamp 1586364061
transform 1 0 6072 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6716 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_71
timestamp 1586364061
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 866 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use scs8hd_fill_1  FILLER_20_80
timestamp 1586364061
transform 1 0 8464 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_20_72
timestamp 1586364061
transform 1 0 7728 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_79
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_75
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_88
timestamp 1586364061
transform 1 0 9200 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_3  FILLER_19_83
timestamp 1586364061
transform 1 0 8740 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9292 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  _069_
timestamp 1586364061
transform 1 0 8556 0 -1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9200 0 1 12512
box -38 -48 866 592
use scs8hd_inv_8  _094_
timestamp 1586364061
transform 1 0 10764 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_97
timestamp 1586364061
transform 1 0 10028 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_101
timestamp 1586364061
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_91
timestamp 1586364061
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_20_102
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_20_110
timestamp 1586364061
transform 1 0 11224 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 11040 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__C
timestamp 1586364061
transform 1 0 11408 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_123
timestamp 1586364061
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_or3_4  _150_
timestamp 1586364061
transform 1 0 11592 0 -1 13600
box -38 -48 866 592
use scs8hd_inv_8  _070_
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_127
timestamp 1586364061
transform 1 0 12788 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_132
timestamp 1586364061
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__B
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_140
timestamp 1586364061
transform 1 0 13984 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_19_140
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_136
timestamp 1586364061
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__B
timestamp 1586364061
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use scs8hd_or3_4  _165_
timestamp 1586364061
transform 1 0 13156 0 -1 13600
box -38 -48 866 592
use scs8hd_nor2_4  _106_
timestamp 1586364061
transform 1 0 14076 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_149
timestamp 1586364061
transform 1 0 14812 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_150
timestamp 1586364061
transform 1 0 14904 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__C
timestamp 1586364061
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 14628 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 14260 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_157
timestamp 1586364061
transform 1 0 15548 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_154
timestamp 1586364061
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__B
timestamp 1586364061
transform 1 0 15732 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 15088 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15456 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_buf_1  _097_
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15640 0 1 12512
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_20_165
timestamp 1586364061
transform 1 0 16284 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_161
timestamp 1586364061
transform 1 0 15916 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_169
timestamp 1586364061
transform 1 0 16652 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16376 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_177
timestamp 1586364061
transform 1 0 17388 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_4  FILLER_19_177
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_173
timestamp 1586364061
transform 1 0 17020 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16560 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17940 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18216 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_194
timestamp 1586364061
transform 1 0 18952 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_188
timestamp 1586364061
transform 1 0 18400 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 19136 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18492 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18124 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_1  FILLER_20_202
timestamp 1586364061
transform 1 0 19688 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_198
timestamp 1586364061
transform 1 0 19320 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_205
timestamp 1586364061
transform 1 0 19964 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_202
timestamp 1586364061
transform 1 0 19688 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_198
timestamp 1586364061
transform 1 0 19320 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19780 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_206
timestamp 1586364061
transform 1 0 20056 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_213
timestamp 1586364061
transform 1 0 20700 0 1 12512
box -38 -48 222 592
use scs8hd_or2_4  _074_
timestamp 1586364061
transform 1 0 20056 0 1 12512
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_219
timestamp 1586364061
transform 1 0 21252 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_217
timestamp 1586364061
transform 1 0 21068 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21068 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21252 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 20884 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_230
timestamp 1586364061
transform 1 0 22264 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_230
timestamp 1586364061
transform 1 0 22264 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21436 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21436 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_1  FILLER_20_236
timestamp 1586364061
transform 1 0 22816 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_238
timestamp 1586364061
transform 1 0 23000 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_234
timestamp 1586364061
transform 1 0 22632 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22908 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23092 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_248
timestamp 1586364061
transform 1 0 23920 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_249
timestamp 1586364061
transform 1 0 24012 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_241
timestamp 1586364061
transform 1 0 23276 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23828 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23092 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_4  FILLER_20_252
timestamp 1586364061
transform 1 0 24288 0 -1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24380 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24104 0 -1 13600
box -38 -48 222 592
use scs8hd_buf_2  _195_
timestamp 1586364061
transform 1 0 24564 0 1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_20_265
timestamp 1586364061
transform 1 0 25484 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_8  FILLER_19_267
timestamp 1586364061
transform 1 0 25668 0 1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_263
timestamp 1586364061
transform 1 0 25300 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_259
timestamp 1586364061
transform 1 0 24932 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25484 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 25116 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24656 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_275
timestamp 1586364061
transform 1 0 26404 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_273
timestamp 1586364061
transform 1 0 26220 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_buf_2  _185_
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1932 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2392 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_7
timestamp 1586364061
transform 1 0 1748 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_11
timestamp 1586364061
transform 1 0 2116 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_16
timestamp 1586364061
transform 1 0 2576 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 4324 0 1 13600
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2760 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 4140 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_27
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_31
timestamp 1586364061
transform 1 0 3956 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_46
timestamp 1586364061
transform 1 0 5336 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_50
timestamp 1586364061
transform 1 0 5704 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9292 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 9108 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 8372 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8740 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_73
timestamp 1586364061
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_77
timestamp 1586364061
transform 1 0 8188 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_81
timestamp 1586364061
transform 1 0 8556 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_85
timestamp 1586364061
transform 1 0 8924 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 10488 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_100
timestamp 1586364061
transform 1 0 10304 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_104
timestamp 1586364061
transform 1 0 10672 0 1 13600
box -38 -48 406 592
use scs8hd_buf_1  _105_
timestamp 1586364061
transform 1 0 11316 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 12052 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 11132 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_108
timestamp 1586364061
transform 1 0 11040 0 1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_21_121
timestamp 1586364061
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use scs8hd_or3_4  _067_
timestamp 1586364061
transform 1 0 12604 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__B
timestamp 1586364061
transform 1 0 13984 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_134
timestamp 1586364061
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_138
timestamp 1586364061
transform 1 0 13800 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_142
timestamp 1586364061
transform 1 0 14168 0 1 13600
box -38 -48 130 592
use scs8hd_or3_4  _085_
timestamp 1586364061
transform 1 0 14260 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__067__C
timestamp 1586364061
transform 1 0 15272 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 15640 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_152
timestamp 1586364061
transform 1 0 15088 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_156
timestamp 1586364061
transform 1 0 15456 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_160
timestamp 1586364061
transform 1 0 15824 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__B
timestamp 1586364061
transform 1 0 16008 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_164
timestamp 1586364061
transform 1 0 16192 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_175
timestamp 1586364061
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18952 0 1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 18584 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__B
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18216 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_179
timestamp 1586364061
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_188
timestamp 1586364061
transform 1 0 18400 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_192
timestamp 1586364061
transform 1 0 18768 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20700 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20516 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20148 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_205
timestamp 1586364061
transform 1 0 19964 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_209
timestamp 1586364061
transform 1 0 20332 0 1 13600
box -38 -48 222 592
use scs8hd_buf_1  _075_
timestamp 1586364061
transform 1 0 22264 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 21712 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22080 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_222
timestamp 1586364061
transform 1 0 21528 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_226
timestamp 1586364061
transform 1 0 21896 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24012 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 22724 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23828 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_233
timestamp 1586364061
transform 1 0 22540 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_237
timestamp 1586364061
transform 1 0 22908 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_242
timestamp 1586364061
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25576 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25024 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25392 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_258
timestamp 1586364061
transform 1 0 24840 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_262
timestamp 1586364061
transform 1 0 25208 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26036 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_269
timestamp 1586364061
transform 1 0 25852 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_273
timestamp 1586364061
transform 1 0 26220 0 1 13600
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_6
timestamp 1586364061
transform 1 0 1656 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_10
timestamp 1586364061
transform 1 0 2024 0 -1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4232 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_23
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 4416 0 -1 14688
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_22_47
timestamp 1586364061
transform 1 0 5428 0 -1 14688
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7452 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_55
timestamp 1586364061
transform 1 0 6164 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_67
timestamp 1586364061
transform 1 0 7268 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_71
timestamp 1586364061
transform 1 0 7636 0 -1 14688
box -38 -48 406 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 8004 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_84
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_88
timestamp 1586364061
transform 1 0 9200 0 -1 14688
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_6  FILLER_22_104
timestamp 1586364061
transform 1 0 10672 0 -1 14688
box -38 -48 590 592
use scs8hd_or3_4  _088_
timestamp 1586364061
transform 1 0 12052 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__088__C
timestamp 1586364061
transform 1 0 11868 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 11224 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_112
timestamp 1586364061
transform 1 0 11408 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_116
timestamp 1586364061
transform 1 0 11776 0 -1 14688
box -38 -48 130 592
use scs8hd_or3_4  _091_
timestamp 1586364061
transform 1 0 13616 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__078__B
timestamp 1586364061
transform 1 0 13248 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_128
timestamp 1586364061
transform 1 0 12880 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_134
timestamp 1586364061
transform 1 0 13432 0 -1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _087_
timestamp 1586364061
transform 1 0 15456 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__091__C
timestamp 1586364061
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_145
timestamp 1586364061
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_149
timestamp 1586364061
transform 1 0 14812 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _076_
timestamp 1586364061
transform 1 0 17020 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 16468 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_165
timestamp 1586364061
transform 1 0 16284 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_169
timestamp 1586364061
transform 1 0 16652 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 18584 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18400 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_182
timestamp 1586364061
transform 1 0 17848 0 -1 14688
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19780 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20148 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_201
timestamp 1586364061
transform 1 0 19596 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_205
timestamp 1586364061
transform 1 0 19964 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_209
timestamp 1586364061
transform 1 0 20332 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_213
timestamp 1586364061
transform 1 0 20700 0 -1 14688
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 21436 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21068 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_219
timestamp 1586364061
transform 1 0 21252 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23184 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_232
timestamp 1586364061
transform 1 0 22448 0 -1 14688
box -38 -48 590 592
use scs8hd_decap_8  FILLER_22_249
timestamp 1586364061
transform 1 0 24012 0 -1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24748 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_266
timestamp 1586364061
transform 1 0 25576 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_274
timestamp 1586364061
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2208 0 1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2024 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1656 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_8
timestamp 1586364061
transform 1 0 1840 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3772 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3220 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_21
timestamp 1586364061
transform 1 0 3036 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_25
timestamp 1586364061
transform 1 0 3404 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5336 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 5152 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_38
timestamp 1586364061
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_42
timestamp 1586364061
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_49
timestamp 1586364061
transform 1 0 5612 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 6440 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_23_60
timestamp 1586364061
transform 1 0 6624 0 1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_23_71
timestamp 1586364061
transform 1 0 7636 0 1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9016 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__B
timestamp 1586364061
transform 1 0 8832 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 8372 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_77
timestamp 1586364061
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_81
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 314 592
use scs8hd_nor2_4  _154_
timestamp 1586364061
transform 1 0 10580 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_95
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_99
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use scs8hd_inv_8  _066_
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_112
timestamp 1586364061
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_116
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 406 592
use scs8hd_inv_8  _081_
timestamp 1586364061
transform 1 0 13984 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 13800 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 13432 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_132
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_136
timestamp 1586364061
transform 1 0 13616 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__C
timestamp 1586364061
transform 1 0 14996 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__B
timestamp 1586364061
transform 1 0 15548 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_149
timestamp 1586364061
transform 1 0 14812 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_153
timestamp 1586364061
transform 1 0 15180 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_159
timestamp 1586364061
transform 1 0 15732 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _080_
timestamp 1586364061
transform 1 0 16376 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 17480 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 15916 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_163
timestamp 1586364061
transform 1 0 16100 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_175
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18492 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 18216 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_180
timestamp 1586364061
transform 1 0 17664 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_188
timestamp 1586364061
transform 1 0 18400 0 1 14688
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 20056 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 19872 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19504 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_198
timestamp 1586364061
transform 1 0 19320 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_202
timestamp 1586364061
transform 1 0 19688 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 21804 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 21620 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21252 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_217
timestamp 1586364061
transform 1 0 21068 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_221
timestamp 1586364061
transform 1 0 21436 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23920 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_236
timestamp 1586364061
transform 1 0 22816 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_240
timestamp 1586364061
transform 1 0 23184 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 314 592
use scs8hd_buf_2  _196_
timestamp 1586364061
transform 1 0 25484 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 24932 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_257
timestamp 1586364061
transform 1 0 24748 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_261
timestamp 1586364061
transform 1 0 25116 0 1 14688
box -38 -48 406 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 26036 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_269
timestamp 1586364061
transform 1 0 25852 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_273
timestamp 1586364061
transform 1 0 26220 0 1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 15776
box -38 -48 866 592
use scs8hd_inv_1  mux_left_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 1840 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_6
timestamp 1586364061
transform 1 0 1656 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_10
timestamp 1586364061
transform 1 0 2024 0 -1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_6  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 590 592
use scs8hd_nor2_4  _122_
timestamp 1586364061
transform 1 0 4600 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5888 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_47
timestamp 1586364061
transform 1 0 5428 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_51
timestamp 1586364061
transform 1 0 5796 0 -1 15776
box -38 -48 130 592
use scs8hd_nor2_4  _157_
timestamp 1586364061
transform 1 0 6440 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_54
timestamp 1586364061
transform 1 0 6072 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_67
timestamp 1586364061
transform 1 0 7268 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_71
timestamp 1586364061
transform 1 0 7636 0 -1 15776
box -38 -48 406 592
use scs8hd_nor2_4  _153_
timestamp 1586364061
transform 1 0 8004 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_88
timestamp 1586364061
transform 1 0 9200 0 -1 15776
box -38 -48 406 592
use scs8hd_nor2_4  _155_
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_102
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_106
timestamp 1586364061
transform 1 0 10856 0 -1 15776
box -38 -48 406 592
use scs8hd_nor2_4  _152_
timestamp 1586364061
transform 1 0 11224 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_12  FILLER_24_119
timestamp 1586364061
transform 1 0 12052 0 -1 15776
box -38 -48 1142 592
use scs8hd_or3_4  _078_
timestamp 1586364061
transform 1 0 13248 0 -1 15776
box -38 -48 866 592
use scs8hd_fill_1  FILLER_24_131
timestamp 1586364061
transform 1 0 13156 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_141
timestamp 1586364061
transform 1 0 14076 0 -1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__082__C
timestamp 1586364061
transform 1 0 14260 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 14628 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 15732 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_145
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_149
timestamp 1586364061
transform 1 0 14812 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_4  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_158
timestamp 1586364061
transform 1 0 15640 0 -1 15776
box -38 -48 130 592
use scs8hd_nor2_4  _084_
timestamp 1586364061
transform 1 0 15916 0 -1 15776
box -38 -48 866 592
use scs8hd_nor2_4  _170_
timestamp 1586364061
transform 1 0 17480 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16928 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_170
timestamp 1586364061
transform 1 0 16744 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_174
timestamp 1586364061
transform 1 0 17112 0 -1 15776
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 19044 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18492 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18860 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_187
timestamp 1586364061
transform 1 0 18308 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_191
timestamp 1586364061
transform 1 0 18676 0 -1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_206
timestamp 1586364061
transform 1 0 20056 0 -1 15776
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21068 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22080 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_226
timestamp 1586364061
transform 1 0 21896 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_230
timestamp 1586364061
transform 1 0 22264 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23000 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24012 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_247
timestamp 1586364061
transform 1 0 23828 0 -1 15776
box -38 -48 222 592
use scs8hd_buf_2  _194_
timestamp 1586364061
transform 1 0 24564 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_4  FILLER_24_251
timestamp 1586364061
transform 1 0 24196 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_259
timestamp 1586364061
transform 1 0 24932 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_271
timestamp 1586364061
transform 1 0 26036 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_buf_2  _184_
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2300 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_7
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_11
timestamp 1586364061
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 3956 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_24
timestamp 1586364061
transform 1 0 3312 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_29
timestamp 1586364061
transform 1 0 3772 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 5152 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 4968 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_36
timestamp 1586364061
transform 1 0 4416 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_40
timestamp 1586364061
transform 1 0 4784 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _156_
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_71
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use scs8hd_buf_1  _089_
timestamp 1586364061
transform 1 0 8740 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 9200 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 8556 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8188 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_75
timestamp 1586364061
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_79
timestamp 1586364061
transform 1 0 8372 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_86
timestamp 1586364061
transform 1 0 9016 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9752 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 9568 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_90
timestamp 1586364061
transform 1 0 9384 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_105
timestamp 1586364061
transform 1 0 10764 0 1 15776
box -38 -48 406 592
use scs8hd_inv_8  _065_
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 11132 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11500 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_111
timestamp 1586364061
transform 1 0 11316 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_115
timestamp 1586364061
transform 1 0 11684 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_119
timestamp 1586364061
transform 1 0 12052 0 1 15776
box -38 -48 130 592
use scs8hd_nor2_4  _167_
timestamp 1586364061
transform 1 0 14168 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__082__B
timestamp 1586364061
transform 1 0 13616 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__B
timestamp 1586364061
transform 1 0 13984 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_132
timestamp 1586364061
transform 1 0 13248 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_138
timestamp 1586364061
transform 1 0 13800 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _168_
timestamp 1586364061
transform 1 0 15732 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 15548 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 15180 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_151
timestamp 1586364061
transform 1 0 14996 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_155
timestamp 1586364061
transform 1 0 15364 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 16744 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17112 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_168
timestamp 1586364061
transform 1 0 16560 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_172
timestamp 1586364061
transform 1 0 16928 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_176
timestamp 1586364061
transform 1 0 17296 0 1 15776
box -38 -48 406 592
use scs8hd_nor2_4  _169_
timestamp 1586364061
transform 1 0 18216 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_180
timestamp 1586364061
transform 1 0 17664 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_195
timestamp 1586364061
transform 1 0 19044 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19780 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 19228 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__B
timestamp 1586364061
transform 1 0 20792 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19596 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_199
timestamp 1586364061
transform 1 0 19412 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_212
timestamp 1586364061
transform 1 0 20608 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _172_
timestamp 1586364061
transform 1 0 21344 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 21160 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_216
timestamp 1586364061
transform 1 0 20976 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_229
timestamp 1586364061
transform 1 0 22172 0 1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 22448 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_234
timestamp 1586364061
transform 1 0 22632 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_240
timestamp 1586364061
transform 1 0 23184 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 24656 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_254
timestamp 1586364061
transform 1 0 24472 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_258
timestamp 1586364061
transform 1 0 24840 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_265
timestamp 1586364061
transform 1 0 25484 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_25_269
timestamp 1586364061
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  FILLER_27_7
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 314 592
use scs8hd_decap_8  FILLER_26_7
timestamp 1586364061
transform 1 0 1748 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_buf_2  _187_
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use scs8hd_buf_2  _186_
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_3  FILLER_27_12
timestamp 1586364061
transform 1 0 2208 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2024 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 314 592
use scs8hd_conb_1  _173_
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 314 592
use scs8hd_decap_8  FILLER_27_18
timestamp 1586364061
transform 1 0 2760 0 1 16864
box -38 -48 774 592
use scs8hd_decap_4  FILLER_26_26
timestamp 1586364061
transform 1 0 3496 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_22
timestamp 1586364061
transform 1 0 3128 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_18
timestamp 1586364061
transform 1 0 2760 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2944 0 -1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3496 0 1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_27_33
timestamp 1586364061
transform 1 0 4140 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_29
timestamp 1586364061
transform 1 0 3772 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_30
timestamp 1586364061
transform 1 0 3864 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3956 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_26_36
timestamp 1586364061
transform 1 0 4416 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 4968 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4508 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_53
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_50
timestamp 1586364061
transform 1 0 5704 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_46
timestamp 1586364061
transform 1 0 5336 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5888 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 5520 0 -1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _126_
timestamp 1586364061
transform 1 0 5152 0 1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 4508 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_69
timestamp 1586364061
transform 1 0 7452 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_65
timestamp 1586364061
transform 1 0 7084 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7636 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 7268 0 -1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6072 0 -1 16864
box -38 -48 1050 592
use scs8hd_buf_1  _079_
timestamp 1586364061
transform 1 0 8832 0 1 16864
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 9292 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_73
timestamp 1586364061
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_77
timestamp 1586364061
transform 1 0 8188 0 1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_27_83
timestamp 1586364061
transform 1 0 8740 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_87
timestamp 1586364061
transform 1 0 9108 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_91
timestamp 1586364061
transform 1 0 9476 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_97
timestamp 1586364061
transform 1 0 10028 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9844 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_buf_1  _086_
timestamp 1586364061
transform 1 0 10120 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_106
timestamp 1586364061
transform 1 0 10856 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_105
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_101
timestamp 1586364061
transform 1 0 10396 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10580 0 -1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9844 0 1 16864
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_110
timestamp 1586364061
transform 1 0 11224 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11040 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__D
timestamp 1586364061
transform 1 0 11408 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_124
timestamp 1586364061
transform 1 0 12512 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_120
timestamp 1586364061
transform 1 0 12144 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__B
timestamp 1586364061
transform 1 0 12328 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__C
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 11132 0 -1 16864
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_27_132
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_26_132
timestamp 1586364061
transform 1 0 13248 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_128
timestamp 1586364061
transform 1 0 12880 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13064 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12696 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_137
timestamp 1586364061
transform 1 0 13708 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 13892 0 1 16864
box -38 -48 222 592
use scs8hd_nor3_4  _161_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 14076 0 1 16864
box -38 -48 1234 592
use scs8hd_or3_4  _082_
timestamp 1586364061
transform 1 0 13616 0 -1 16864
box -38 -48 866 592
use scs8hd_buf_1  _103_
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 15824 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15456 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_145
timestamp 1586364061
transform 1 0 14444 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_4  FILLER_26_157
timestamp 1586364061
transform 1 0 15548 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_154
timestamp 1586364061
transform 1 0 15272 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_158
timestamp 1586364061
transform 1 0 15640 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 16008 0 1 16864
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16468 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 16008 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_161
timestamp 1586364061
transform 1 0 15916 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_26_164
timestamp 1586364061
transform 1 0 16192 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_8  FILLER_26_176
timestamp 1586364061
transform 1 0 17296 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_4  FILLER_27_173
timestamp 1586364061
transform 1 0 17020 0 1 16864
box -38 -48 406 592
use scs8hd_decap_3  FILLER_27_187
timestamp 1586364061
transform 1 0 18308 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_179
timestamp 1586364061
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_184
timestamp 1586364061
transform 1 0 18032 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 18216 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_buf_1  _101_
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_192
timestamp 1586364061
transform 1 0 18768 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_188
timestamp 1586364061
transform 1 0 18400 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 18584 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 18952 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_2_.latch
timestamp 1586364061
transform 1 0 18952 0 -1 16864
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20332 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20700 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20148 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_205
timestamp 1586364061
transform 1 0 19964 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_209
timestamp 1586364061
transform 1 0 20332 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_207
timestamp 1586364061
transform 1 0 20148 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_211
timestamp 1586364061
transform 1 0 20516 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21896 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22264 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_224
timestamp 1586364061
transform 1 0 21712 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_224
timestamp 1586364061
transform 1 0 21712 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_228
timestamp 1586364061
transform 1 0 22080 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_239
timestamp 1586364061
transform 1 0 23092 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_235
timestamp 1586364061
transform 1 0 22724 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_235
timestamp 1586364061
transform 1 0 22724 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22908 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 1 16864
box -38 -48 314 592
use scs8hd_buf_1  _092_
timestamp 1586364061
transform 1 0 22448 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_248
timestamp 1586364061
transform 1 0 23920 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_243
timestamp 1586364061
transform 1 0 23460 0 1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_246
timestamp 1586364061
transform 1 0 23736 0 -1 16864
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 314 592
use scs8hd_conb_1  _176_
timestamp 1586364061
transform 1 0 23460 0 -1 16864
box -38 -48 314 592
use scs8hd_buf_1  _107_
timestamp 1586364061
transform 1 0 24472 0 -1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24656 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25116 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_257
timestamp 1586364061
transform 1 0 24748 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_27_252
timestamp 1586364061
transform 1 0 24288 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_259
timestamp 1586364061
transform 1 0 24932 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_263
timestamp 1586364061
transform 1 0 25300 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_26_269
timestamp 1586364061
transform 1 0 25852 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_275
timestamp 1586364061
transform 1 0 26404 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2024 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 1564 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_7
timestamp 1586364061
transform 1 0 1748 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_13
timestamp 1586364061
transform 1 0 2300 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_6  FILLER_28_25
timestamp 1586364061
transform 1 0 3404 0 -1 17952
box -38 -48 590 592
use scs8hd_decap_4  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4508 0 -1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5520 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_36
timestamp 1586364061
transform 1 0 4416 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_40
timestamp 1586364061
transform 1 0 4784 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_46
timestamp 1586364061
transform 1 0 5336 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7084 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_57
timestamp 1586364061
transform 1 0 6348 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_61
timestamp 1586364061
transform 1 0 6716 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_64
timestamp 1586364061
transform 1 0 6992 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8096 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_74
timestamp 1586364061
transform 1 0 7912 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_78
timestamp 1586364061
transform 1 0 8280 0 -1 17952
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_90
timestamp 1586364061
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_102
timestamp 1586364061
transform 1 0 10488 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_106
timestamp 1586364061
transform 1 0 10856 0 -1 17952
box -38 -48 222 592
use scs8hd_nor4_4  _164_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12144 0 -1 17952
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11960 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_110
timestamp 1586364061
transform 1 0 11224 0 -1 17952
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 13892 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_137
timestamp 1586364061
transform 1 0 13708 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_141
timestamp 1586364061
transform 1 0 14076 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__161__C
timestamp 1586364061
transform 1 0 14260 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__C
timestamp 1586364061
transform 1 0 14720 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15824 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_145
timestamp 1586364061
transform 1 0 14444 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_150
timestamp 1586364061
transform 1 0 14904 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_6  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 16008 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17480 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_173
timestamp 1586364061
transform 1 0 17020 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_177
timestamp 1586364061
transform 1 0 17388 0 -1 17952
box -38 -48 130 592
use scs8hd_buf_1  _083_
timestamp 1586364061
transform 1 0 17756 0 -1 17952
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 19044 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 18860 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 18216 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_180
timestamp 1586364061
transform 1 0 17664 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_184
timestamp 1586364061
transform 1 0 18032 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_188
timestamp 1586364061
transform 1 0 18400 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_192
timestamp 1586364061
transform 1 0 18768 0 -1 17952
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_206
timestamp 1586364061
transform 1 0 20056 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_210
timestamp 1586364061
transform 1 0 20424 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_8  FILLER_28_224
timestamp 1586364061
transform 1 0 21712 0 -1 17952
box -38 -48 774 592
use scs8hd_conb_1  _181_
timestamp 1586364061
transform 1 0 22448 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_235
timestamp 1586364061
transform 1 0 22724 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_247
timestamp 1586364061
transform 1 0 23828 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_259
timestamp 1586364061
transform 1 0 24932 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_271
timestamp 1586364061
transform 1 0 26036 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_27
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5520 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_39
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_29_47
timestamp 1586364061
transform 1 0 5428 0 1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_29_53
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7360 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7176 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 406 592
use scs8hd_buf_1  _158_
timestamp 1586364061
transform 1 0 9200 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_77
timestamp 1586364061
transform 1 0 8188 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_81
timestamp 1586364061
transform 1 0 8556 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_85
timestamp 1586364061
transform 1 0 8924 0 1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 9660 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_91
timestamp 1586364061
transform 1 0 9476 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_95
timestamp 1586364061
transform 1 0 9844 0 1 17952
box -38 -48 222 592
use scs8hd_nor4_4  _163_
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__D
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__C
timestamp 1586364061
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_108
timestamp 1586364061
transform 1 0 11040 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 14168 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_140
timestamp 1586364061
transform 1 0 13984 0 1 17952
box -38 -48 222 592
use scs8hd_nor3_4  _159_
timestamp 1586364061
transform 1 0 14720 0 1 17952
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 14536 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_144
timestamp 1586364061
transform 1 0 14352 0 1 17952
box -38 -48 222 592
use scs8hd_buf_1  _099_
timestamp 1586364061
transform 1 0 16652 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16100 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 17112 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16468 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_161
timestamp 1586364061
transform 1 0 15916 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_165
timestamp 1586364061
transform 1 0 16284 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_172
timestamp 1586364061
transform 1 0 16928 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_176
timestamp 1586364061
transform 1 0 17296 0 1 17952
box -38 -48 406 592
use scs8hd_nor2_4  _171_
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_180
timestamp 1586364061
transform 1 0 17664 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_193
timestamp 1586364061
transform 1 0 18860 0 1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 19596 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 19412 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_197
timestamp 1586364061
transform 1 0 19228 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_212
timestamp 1586364061
transform 1 0 20608 0 1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21344 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_217
timestamp 1586364061
transform 1 0 21068 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_229
timestamp 1586364061
transform 1 0 22172 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_29_241
timestamp 1586364061
transform 1 0 23276 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_253
timestamp 1586364061
transform 1 0 24380 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_269
timestamp 1586364061
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6348 0 -1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 866 592
use scs8hd_fill_1  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_60
timestamp 1586364061
transform 1 0 6624 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_12  FILLER_30_77
timestamp 1586364061
transform 1 0 8188 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_30_89
timestamp 1586364061
transform 1 0 9292 0 -1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 590 592
use scs8hd_inv_1  mux_top_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11960 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 12420 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_110
timestamp 1586364061
transform 1 0 11224 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_2  FILLER_30_121
timestamp 1586364061
transform 1 0 12236 0 -1 19040
box -38 -48 222 592
use scs8hd_nor3_4  _162_
timestamp 1586364061
transform 1 0 13248 0 -1 19040
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 12788 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_125
timestamp 1586364061
transform 1 0 12604 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_129
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15732 0 -1 19040
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 14720 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15456 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_145
timestamp 1586364061
transform 1 0 14444 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_150
timestamp 1586364061
transform 1 0 14904 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_158
timestamp 1586364061
transform 1 0 15640 0 -1 19040
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17480 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17296 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_170
timestamp 1586364061
transform 1 0 16744 0 -1 19040
box -38 -48 590 592
use scs8hd_nor2_4  _093_
timestamp 1586364061
transform 1 0 19044 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18492 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_187
timestamp 1586364061
transform 1 0 18308 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_191
timestamp 1586364061
transform 1 0 18676 0 -1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20056 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_204
timestamp 1586364061
transform 1 0 19872 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_208
timestamp 1586364061
transform 1 0 20240 0 -1 19040
box -38 -48 590 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21344 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21712 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_218
timestamp 1586364061
transform 1 0 21160 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_222
timestamp 1586364061
transform 1 0 21528 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_226
timestamp 1586364061
transform 1 0 21896 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_238
timestamp 1586364061
transform 1 0 23000 0 -1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_30_250
timestamp 1586364061
transform 1 0 24104 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_254
timestamp 1586364061
transform 1 0 24472 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_258
timestamp 1586364061
transform 1 0 24840 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_270
timestamp 1586364061
transform 1 0 25944 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_274
timestamp 1586364061
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_6
timestamp 1586364061
transform 1 0 1656 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_10
timestamp 1586364061
transform 1 0 2024 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_22
timestamp 1586364061
transform 1 0 3128 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_34
timestamp 1586364061
transform 1 0 4232 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_46
timestamp 1586364061
transform 1 0 5336 0 1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6992 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7452 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_58
timestamp 1586364061
transform 1 0 6440 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_67
timestamp 1586364061
transform 1 0 7268 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_71
timestamp 1586364061
transform 1 0 7636 0 1 19040
box -38 -48 590 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9200 0 1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8188 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8648 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_80
timestamp 1586364061
transform 1 0 8464 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_84
timestamp 1586364061
transform 1 0 8832 0 1 19040
box -38 -48 222 592
use scs8hd_conb_1  _179_
timestamp 1586364061
transform 1 0 10304 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9844 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 10856 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_91
timestamp 1586364061
transform 1 0 9476 0 1 19040
box -38 -48 406 592
use scs8hd_decap_3  FILLER_31_97
timestamp 1586364061
transform 1 0 10028 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_31_103
timestamp 1586364061
transform 1 0 10580 0 1 19040
box -38 -48 314 592
use scs8hd_buf_1  _068_
timestamp 1586364061
transform 1 0 11316 0 1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_14.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11868 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_108
timestamp 1586364061
transform 1 0 11040 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_31_114
timestamp 1586364061
transform 1 0 11592 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_31_119
timestamp 1586364061
transform 1 0 12052 0 1 19040
box -38 -48 314 592
use scs8hd_nor3_4  _160_
timestamp 1586364061
transform 1 0 13984 0 1 19040
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 13800 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 13432 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_126
timestamp 1586364061
transform 1 0 12696 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_130
timestamp 1586364061
transform 1 0 13064 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_136
timestamp 1586364061
transform 1 0 13616 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15364 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_153
timestamp 1586364061
transform 1 0 15180 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_157
timestamp 1586364061
transform 1 0 15548 0 1 19040
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16192 0 1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 16008 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_161
timestamp 1586364061
transform 1 0 15916 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_175
timestamp 1586364061
transform 1 0 17204 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 19044 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_179
timestamp 1586364061
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_193
timestamp 1586364061
transform 1 0 18860 0 1 19040
box -38 -48 222 592
use scs8hd_inv_8  _146_
timestamp 1586364061
transform 1 0 19596 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19412 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_197
timestamp 1586364061
transform 1 0 19228 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_210
timestamp 1586364061
transform 1 0 20424 0 1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_221
timestamp 1586364061
transform 1 0 21436 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_225
timestamp 1586364061
transform 1 0 21804 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_31_237
timestamp 1586364061
transform 1 0 22908 0 1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_31_243
timestamp 1586364061
transform 1 0 23460 0 1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_253
timestamp 1586364061
transform 1 0 24380 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_258
timestamp 1586364061
transform 1 0 24840 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_262
timestamp 1586364061
transform 1 0 25208 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_31_274
timestamp 1586364061
transform 1 0 26312 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use scs8hd_buf_1  _151_
timestamp 1586364061
transform 1 0 10856 0 -1 20128
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9844 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10580 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_98
timestamp 1586364061
transform 1 0 10120 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_102
timestamp 1586364061
transform 1 0 10488 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_105
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_14.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 11316 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_109
timestamp 1586364061
transform 1 0 11132 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_113
timestamp 1586364061
transform 1 0 11500 0 -1 20128
box -38 -48 406 592
use scs8hd_inv_8  _147_
timestamp 1586364061
transform 1 0 13616 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 13432 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13064 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_128
timestamp 1586364061
transform 1 0 12880 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_132
timestamp 1586364061
transform 1 0 13248 0 -1 20128
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__160__C
timestamp 1586364061
transform 1 0 14628 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_145
timestamp 1586364061
transform 1 0 14444 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_149
timestamp 1586364061
transform 1 0 14812 0 -1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16468 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17296 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_165
timestamp 1586364061
transform 1 0 16284 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_169
timestamp 1586364061
transform 1 0 16652 0 -1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_32_175
timestamp 1586364061
transform 1 0 17204 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_178
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17848 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 17664 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_191
timestamp 1586364061
transform 1 0 18676 0 -1 20128
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19412 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_202
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_263
timestamp 1586364061
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_39
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_51
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_8  _148_
timestamp 1586364061
transform 1 0 10764 0 1 20128
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 -1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 10212 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_101
timestamp 1586364061
transform 1 0 10396 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_34_101
timestamp 1586364061
transform 1 0 10396 0 -1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12144 0 -1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_114
timestamp 1586364061
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_118
timestamp 1586364061
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_34_112
timestamp 1586364061
transform 1 0 11408 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_34_133
timestamp 1586364061
transform 1 0 13340 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_129
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13156 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_140
timestamp 1586364061
transform 1 0 13984 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_6  FILLER_33_141
timestamp 1586364061
transform 1 0 14076 0 1 20128
box -38 -48 590 592
use scs8hd_fill_2  FILLER_33_137
timestamp 1586364061
transform 1 0 13708 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13892 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13524 0 -1 21216
box -38 -48 222 592
use scs8hd_conb_1  _180_
timestamp 1586364061
transform 1 0 13708 0 -1 21216
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_14.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12696 0 1 20128
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 14904 0 1 20128
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 14720 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14904 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_147
timestamp 1586364061
transform 1 0 14628 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_148
timestamp 1586364061
transform 1 0 14720 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_152
timestamp 1586364061
transform 1 0 15088 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_34_160
timestamp 1586364061
transform 1 0 15824 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_165
timestamp 1586364061
transform 1 0 16284 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_161
timestamp 1586364061
transform 1 0 15916 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15916 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16100 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16652 0 1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_34_172
timestamp 1586364061
transform 1 0 16928 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_4  FILLER_33_176
timestamp 1586364061
transform 1 0 17296 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_172
timestamp 1586364061
transform 1 0 16928 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17112 0 1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 -1 21216
box -38 -48 866 592
use scs8hd_fill_2  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_180
timestamp 1586364061
transform 1 0 17664 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_34_193
timestamp 1586364061
transform 1 0 18860 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_189
timestamp 1586364061
transform 1 0 18492 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_195
timestamp 1586364061
transform 1 0 19044 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18676 0 -1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18216 0 1 20128
box -38 -48 866 592
use scs8hd_inv_8  _145_
timestamp 1586364061
transform 1 0 17664 0 -1 21216
box -38 -48 866 592
use scs8hd_decap_4  FILLER_33_199
timestamp 1586364061
transform 1 0 19412 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19228 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19228 0 -1 21216
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_212
timestamp 1586364061
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_210
timestamp 1586364061
transform 1 0 20424 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_206
timestamp 1586364061
transform 1 0 20056 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_conb_1  _183_
timestamp 1586364061
transform 1 0 20792 0 1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_34_200
timestamp 1586364061
transform 1 0 19504 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_217
timestamp 1586364061
transform 1 0 21068 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_229
timestamp 1586364061
transform 1 0 22172 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_33_241
timestamp 1586364061
transform 1 0 23276 0 1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_263
timestamp 1586364061
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_14.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_6
timestamp 1586364061
transform 1 0 1656 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_10
timestamp 1586364061
transform 1 0 2024 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_22
timestamp 1586364061
transform 1 0 3128 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_34
timestamp 1586364061
transform 1 0 4232 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_46
timestamp 1586364061
transform 1 0 5336 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_decap_3  FILLER_35_58
timestamp 1586364061
transform 1 0 6440 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_86
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_110
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13340 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12972 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_131
timestamp 1586364061
transform 1 0 13156 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_14.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15088 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15548 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14904 0 1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_144
timestamp 1586364061
transform 1 0 14352 0 1 21216
box -38 -48 590 592
use scs8hd_fill_2  FILLER_35_155
timestamp 1586364061
transform 1 0 15364 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_159
timestamp 1586364061
transform 1 0 15732 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15916 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_172
timestamp 1586364061
transform 1 0 16928 0 1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_35_176
timestamp 1586364061
transform 1 0 17296 0 1 21216
box -38 -48 130 592
use scs8hd_inv_8  _144_
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 19044 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_179
timestamp 1586364061
transform 1 0 17572 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_193
timestamp 1586364061
transform 1 0 18860 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 19412 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_197
timestamp 1586364061
transform 1 0 19228 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_201
timestamp 1586364061
transform 1 0 19596 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_213
timestamp 1586364061
transform 1 0 20700 0 1 21216
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 21804 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_227
timestamp 1586364061
transform 1 0 21988 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_35_239
timestamp 1586364061
transform 1 0 23092 0 1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_35_243
timestamp 1586364061
transform 1 0 23460 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_117
timestamp 1586364061
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13156 0 -1 22304
box -38 -48 866 592
use scs8hd_fill_2  FILLER_36_129
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_36_140
timestamp 1586364061
transform 1 0 13984 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15456 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_152
timestamp 1586364061
transform 1 0 15088 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_158
timestamp 1586364061
transform 1 0 15640 0 -1 22304
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16192 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17204 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16008 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_173
timestamp 1586364061
transform 1 0 17020 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_177
timestamp 1586364061
transform 1 0 17388 0 -1 22304
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17756 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_8  FILLER_36_190
timestamp 1586364061
transform 1 0 18584 0 -1 22304
box -38 -48 774 592
use scs8hd_buf_2  _206_
timestamp 1586364061
transform 1 0 19320 0 -1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_202
timestamp 1586364061
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use scs8hd_buf_2  _204_
timestamp 1586364061
transform 1 0 21804 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_8  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_36_223
timestamp 1586364061
transform 1 0 21620 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_36_229
timestamp 1586364061
transform 1 0 22172 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_241
timestamp 1586364061
transform 1 0 23276 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_253
timestamp 1586364061
transform 1 0 24380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_36_265
timestamp 1586364061
transform 1 0 25484 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_273
timestamp 1586364061
transform 1 0 26220 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_27
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_39
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_51
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_86
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_98
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_110
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 1142 592
use scs8hd_inv_8  _143_
timestamp 1586364061
transform 1 0 14812 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 14628 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_158
timestamp 1586364061
transform 1 0 15640 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_162
timestamp 1586364061
transform 1 0 16008 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_175
timestamp 1586364061
transform 1 0 17204 0 1 22304
box -38 -48 222 592
use scs8hd_conb_1  _182_
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_179
timestamp 1586364061
transform 1 0 17572 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_187
timestamp 1586364061
transform 1 0 18308 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_191
timestamp 1586364061
transform 1 0 18676 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_203
timestamp 1586364061
transform 1 0 19780 0 1 22304
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 20884 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_217
timestamp 1586364061
transform 1 0 21068 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_37_229
timestamp 1586364061
transform 1 0 22172 0 1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 22448 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_234
timestamp 1586364061
transform 1 0 22632 0 1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_37_242
timestamp 1586364061
transform 1 0 23368 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_105
timestamp 1586364061
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_117
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_129
timestamp 1586364061
transform 1 0 12972 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_141
timestamp 1586364061
transform 1 0 14076 0 -1 23392
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15456 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_159
timestamp 1586364061
transform 1 0 15732 0 -1 23392
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16468 0 -1 23392
box -38 -48 866 592
use scs8hd_decap_8  FILLER_38_176
timestamp 1586364061
transform 1 0 17296 0 -1 23392
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_187
timestamp 1586364061
transform 1 0 18308 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_199
timestamp 1586364061
transform 1 0 19412 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_38_211
timestamp 1586364061
transform 1 0 20516 0 -1 23392
box -38 -48 314 592
use scs8hd_buf_2  _205_
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_219
timestamp 1586364061
transform 1 0 21252 0 -1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_38_231
timestamp 1586364061
transform 1 0 22356 0 -1 23392
box -38 -48 130 592
use scs8hd_buf_2  _203_
timestamp 1586364061
transform 1 0 22448 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_236
timestamp 1586364061
transform 1 0 22816 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_248
timestamp 1586364061
transform 1 0 23920 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_260
timestamp 1586364061
transform 1 0 25024 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  FILLER_38_272
timestamp 1586364061
transform 1 0 26128 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_6
timestamp 1586364061
transform 1 0 1656 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_10
timestamp 1586364061
transform 1 0 2024 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_6
timestamp 1586364061
transform 1 0 1656 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_14
timestamp 1586364061
transform 1 0 2392 0 1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_26
timestamp 1586364061
transform 1 0 3496 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_18
timestamp 1586364061
transform 1 0 2760 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_30
timestamp 1586364061
transform 1 0 3864 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_38
timestamp 1586364061
transform 1 0 4600 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_50
timestamp 1586364061
transform 1 0 5704 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_decap_3  FILLER_39_58
timestamp 1586364061
transform 1 0 6440 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_98
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_110
timestamp 1586364061
transform 1 0 11224 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _210_
timestamp 1586364061
transform 1 0 12788 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__210__A
timestamp 1586364061
transform 1 0 13340 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_131
timestamp 1586364061
transform 1 0 13156 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_135
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_129
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_141
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _209_
timestamp 1586364061
transform 1 0 15272 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__209__A
timestamp 1586364061
transform 1 0 15088 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_147
timestamp 1586364061
transform 1 0 14628 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_151
timestamp 1586364061
transform 1 0 14996 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_158
timestamp 1586364061
transform 1 0 15640 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_40_168
timestamp 1586364061
transform 1 0 16560 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_162
timestamp 1586364061
transform 1 0 16008 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_162
timestamp 1586364061
transform 1 0 16008 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__208__A
timestamp 1586364061
transform 1 0 16192 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _208_
timestamp 1586364061
transform 1 0 16192 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_4  FILLER_40_172
timestamp 1586364061
transform 1 0 16928 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_175
timestamp 1586364061
transform 1 0 17204 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 23392
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17296 0 -1 24480
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 23392
box -38 -48 866 592
use scs8hd_buf_2  _207_
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 18584 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_179
timestamp 1586364061
transform 1 0 17572 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_188
timestamp 1586364061
transform 1 0 18400 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_192
timestamp 1586364061
transform 1 0 18768 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_179
timestamp 1586364061
transform 1 0 17572 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_191
timestamp 1586364061
transform 1 0 18676 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_204
timestamp 1586364061
transform 1 0 19872 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_40_203
timestamp 1586364061
transform 1 0 19780 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_3  FILLER_40_211
timestamp 1586364061
transform 1 0 20516 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_216
timestamp 1586364061
transform 1 0 20976 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_39_228
timestamp 1586364061
transform 1 0 22080 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _202_
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22908 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_235
timestamp 1586364061
transform 1 0 22724 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_239
timestamp 1586364061
transform 1 0 23092 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_243
timestamp 1586364061
transform 1 0 23460 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_249
timestamp 1586364061
transform 1 0 24012 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24748 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25208 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 24196 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_253
timestamp 1586364061
transform 1 0 24380 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_260
timestamp 1586364061
transform 1 0 25024 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_264
timestamp 1586364061
transform 1 0 25392 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_251
timestamp 1586364061
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_263
timestamp 1586364061
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_39_276
timestamp 1586364061
transform 1 0 26496 0 1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 4526 0 4582 480 6 address[0]
port 0 nsew default input
rlabel metal2 s 7654 0 7710 480 6 address[1]
port 1 nsew default input
rlabel metal2 s 10782 0 10838 480 6 address[2]
port 2 nsew default input
rlabel metal2 s 13910 0 13966 480 6 address[3]
port 3 nsew default input
rlabel metal2 s 16946 0 17002 480 6 address[4]
port 4 nsew default input
rlabel metal2 s 20074 0 20130 480 6 address[5]
port 5 nsew default input
rlabel metal2 s 23202 0 23258 480 6 address[6]
port 6 nsew default input
rlabel metal3 s 0 17960 480 18080 6 chanx_left_in[0]
port 7 nsew default input
rlabel metal3 s 0 19048 480 19168 6 chanx_left_in[1]
port 8 nsew default input
rlabel metal3 s 0 20000 480 20120 6 chanx_left_in[2]
port 9 nsew default input
rlabel metal3 s 0 21088 480 21208 6 chanx_left_in[3]
port 10 nsew default input
rlabel metal3 s 0 22176 480 22296 6 chanx_left_in[4]
port 11 nsew default input
rlabel metal3 s 0 23128 480 23248 6 chanx_left_in[5]
port 12 nsew default input
rlabel metal3 s 0 24216 480 24336 6 chanx_left_in[6]
port 13 nsew default input
rlabel metal3 s 0 25304 480 25424 6 chanx_left_in[7]
port 14 nsew default input
rlabel metal3 s 0 26256 480 26376 6 chanx_left_in[8]
port 15 nsew default input
rlabel metal3 s 0 8712 480 8832 6 chanx_left_out[0]
port 16 nsew default tristate
rlabel metal3 s 0 9664 480 9784 6 chanx_left_out[1]
port 17 nsew default tristate
rlabel metal3 s 0 10752 480 10872 6 chanx_left_out[2]
port 18 nsew default tristate
rlabel metal3 s 0 11704 480 11824 6 chanx_left_out[3]
port 19 nsew default tristate
rlabel metal3 s 0 12792 480 12912 6 chanx_left_out[4]
port 20 nsew default tristate
rlabel metal3 s 0 13880 480 14000 6 chanx_left_out[5]
port 21 nsew default tristate
rlabel metal3 s 0 14832 480 14952 6 chanx_left_out[6]
port 22 nsew default tristate
rlabel metal3 s 0 15920 480 16040 6 chanx_left_out[7]
port 23 nsew default tristate
rlabel metal3 s 0 17008 480 17128 6 chanx_left_out[8]
port 24 nsew default tristate
rlabel metal3 s 27520 17960 28000 18080 6 chanx_right_in[0]
port 25 nsew default input
rlabel metal3 s 27520 19048 28000 19168 6 chanx_right_in[1]
port 26 nsew default input
rlabel metal3 s 27520 20000 28000 20120 6 chanx_right_in[2]
port 27 nsew default input
rlabel metal3 s 27520 21088 28000 21208 6 chanx_right_in[3]
port 28 nsew default input
rlabel metal3 s 27520 22176 28000 22296 6 chanx_right_in[4]
port 29 nsew default input
rlabel metal3 s 27520 23128 28000 23248 6 chanx_right_in[5]
port 30 nsew default input
rlabel metal3 s 27520 24216 28000 24336 6 chanx_right_in[6]
port 31 nsew default input
rlabel metal3 s 27520 25304 28000 25424 6 chanx_right_in[7]
port 32 nsew default input
rlabel metal3 s 27520 26256 28000 26376 6 chanx_right_in[8]
port 33 nsew default input
rlabel metal3 s 27520 8712 28000 8832 6 chanx_right_out[0]
port 34 nsew default tristate
rlabel metal3 s 27520 9664 28000 9784 6 chanx_right_out[1]
port 35 nsew default tristate
rlabel metal3 s 27520 10752 28000 10872 6 chanx_right_out[2]
port 36 nsew default tristate
rlabel metal3 s 27520 11704 28000 11824 6 chanx_right_out[3]
port 37 nsew default tristate
rlabel metal3 s 27520 12792 28000 12912 6 chanx_right_out[4]
port 38 nsew default tristate
rlabel metal3 s 27520 13880 28000 14000 6 chanx_right_out[5]
port 39 nsew default tristate
rlabel metal3 s 27520 14832 28000 14952 6 chanx_right_out[6]
port 40 nsew default tristate
rlabel metal3 s 27520 15920 28000 16040 6 chanx_right_out[7]
port 41 nsew default tristate
rlabel metal3 s 27520 17008 28000 17128 6 chanx_right_out[8]
port 42 nsew default tristate
rlabel metal2 s 2042 27520 2098 28000 6 chany_top_in[0]
port 43 nsew default input
rlabel metal2 s 3422 27520 3478 28000 6 chany_top_in[1]
port 44 nsew default input
rlabel metal2 s 4802 27520 4858 28000 6 chany_top_in[2]
port 45 nsew default input
rlabel metal2 s 6182 27520 6238 28000 6 chany_top_in[3]
port 46 nsew default input
rlabel metal2 s 7654 27520 7710 28000 6 chany_top_in[4]
port 47 nsew default input
rlabel metal2 s 9034 27520 9090 28000 6 chany_top_in[5]
port 48 nsew default input
rlabel metal2 s 10414 27520 10470 28000 6 chany_top_in[6]
port 49 nsew default input
rlabel metal2 s 11794 27520 11850 28000 6 chany_top_in[7]
port 50 nsew default input
rlabel metal2 s 13174 27520 13230 28000 6 chany_top_in[8]
port 51 nsew default input
rlabel metal2 s 14646 27520 14702 28000 6 chany_top_out[0]
port 52 nsew default tristate
rlabel metal2 s 16026 27520 16082 28000 6 chany_top_out[1]
port 53 nsew default tristate
rlabel metal2 s 17406 27520 17462 28000 6 chany_top_out[2]
port 54 nsew default tristate
rlabel metal2 s 18786 27520 18842 28000 6 chany_top_out[3]
port 55 nsew default tristate
rlabel metal2 s 20166 27520 20222 28000 6 chany_top_out[4]
port 56 nsew default tristate
rlabel metal2 s 21638 27520 21694 28000 6 chany_top_out[5]
port 57 nsew default tristate
rlabel metal2 s 23018 27520 23074 28000 6 chany_top_out[6]
port 58 nsew default tristate
rlabel metal2 s 24398 27520 24454 28000 6 chany_top_out[7]
port 59 nsew default tristate
rlabel metal2 s 25778 27520 25834 28000 6 chany_top_out[8]
port 60 nsew default tristate
rlabel metal2 s 26330 0 26386 480 6 data_in
port 61 nsew default input
rlabel metal2 s 1490 0 1546 480 6 enable
port 62 nsew default input
rlabel metal3 s 0 5584 480 5704 6 left_bottom_grid_pin_11_
port 63 nsew default input
rlabel metal3 s 0 6536 480 6656 6 left_bottom_grid_pin_13_
port 64 nsew default input
rlabel metal3 s 0 7624 480 7744 6 left_bottom_grid_pin_15_
port 65 nsew default input
rlabel metal3 s 0 416 480 536 6 left_bottom_grid_pin_1_
port 66 nsew default input
rlabel metal3 s 0 1368 480 1488 6 left_bottom_grid_pin_3_
port 67 nsew default input
rlabel metal3 s 0 2456 480 2576 6 left_bottom_grid_pin_5_
port 68 nsew default input
rlabel metal3 s 0 3408 480 3528 6 left_bottom_grid_pin_7_
port 69 nsew default input
rlabel metal3 s 0 4496 480 4616 6 left_bottom_grid_pin_9_
port 70 nsew default input
rlabel metal3 s 0 27344 480 27464 6 left_top_grid_pin_10_
port 71 nsew default input
rlabel metal3 s 27520 5584 28000 5704 6 right_bottom_grid_pin_11_
port 72 nsew default input
rlabel metal3 s 27520 6536 28000 6656 6 right_bottom_grid_pin_13_
port 73 nsew default input
rlabel metal3 s 27520 7624 28000 7744 6 right_bottom_grid_pin_15_
port 74 nsew default input
rlabel metal3 s 27520 416 28000 536 6 right_bottom_grid_pin_1_
port 75 nsew default input
rlabel metal3 s 27520 1368 28000 1488 6 right_bottom_grid_pin_3_
port 76 nsew default input
rlabel metal3 s 27520 2456 28000 2576 6 right_bottom_grid_pin_5_
port 77 nsew default input
rlabel metal3 s 27520 3408 28000 3528 6 right_bottom_grid_pin_7_
port 78 nsew default input
rlabel metal3 s 27520 4496 28000 4616 6 right_bottom_grid_pin_9_
port 79 nsew default input
rlabel metal3 s 27520 27344 28000 27464 6 right_top_grid_pin_10_
port 80 nsew default input
rlabel metal2 s 662 27520 718 28000 6 top_left_grid_pin_13_
port 81 nsew default input
rlabel metal2 s 27158 27520 27214 28000 6 top_right_grid_pin_11_
port 82 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 83 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 84 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
