* NGSPICE file created from sb_0__1_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor4_4 abstract view
.subckt scs8hd_nor4_4 A B C D Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

.subckt sb_0__1_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] bottom_left_grid_pin_11_ bottom_left_grid_pin_13_ bottom_left_grid_pin_15_
+ bottom_left_grid_pin_1_ bottom_left_grid_pin_3_ bottom_left_grid_pin_5_ bottom_left_grid_pin_7_
+ bottom_left_grid_pin_9_ bottom_right_grid_pin_11_ chanx_right_in[0] chanx_right_in[1]
+ chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6]
+ chanx_right_in[7] chanx_right_in[8] chanx_right_out[0] chanx_right_out[1] chanx_right_out[2]
+ chanx_right_out[3] chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7]
+ chanx_right_out[8] chany_bottom_in[0] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_out[0] chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3]
+ chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7]
+ chany_bottom_out[8] chany_top_in[0] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_out[0] chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4]
+ chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8] data_in enable
+ right_bottom_grid_pin_12_ right_top_grid_pin_10_ top_left_grid_pin_11_ top_left_grid_pin_13_
+ top_left_grid_pin_15_ top_left_grid_pin_1_ top_left_grid_pin_3_ top_left_grid_pin_5_
+ top_left_grid_pin_7_ top_left_grid_pin_9_ top_right_grid_pin_11_ vpwr vgnd
Xmem_right_track_12.LATCH_1_.latch data_in _181_/A _167_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_199 vpwr vgnd scs8hd_fill_2
XFILLER_22_144 vgnd vpwr scs8hd_decap_4
XFILLER_22_100 vgnd vpwr scs8hd_decap_6
Xmux_bottom_track_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[4] mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_74 vgnd vpwr scs8hd_fill_1
XFILLER_13_177 vgnd vpwr scs8hd_decap_4
Xmux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__113__B _110_/B vgnd vpwr scs8hd_diode_2
XFILLER_3_23 vgnd vpwr scs8hd_decap_3
Xmux_top_track_8.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_3_ mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_32 vgnd vpwr scs8hd_decap_12
XFILLER_10_125 vgnd vpwr scs8hd_decap_6
Xmux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _181_/A mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__214__A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_51 vgnd vpwr scs8hd_decap_8
XFILLER_37_62 vgnd vpwr scs8hd_decap_12
XANTENNA__108__B _110_/B vgnd vpwr scs8hd_diode_2
XFILLER_33_206 vgnd vpwr scs8hd_decap_4
XFILLER_33_217 vgnd vpwr scs8hd_decap_12
XFILLER_41_272 vgnd vpwr scs8hd_decap_4
XANTENNA__124__A _113_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _194_/HI _176_/Y mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_184 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _188_/HI mem_bottom_track_17.LATCH_2_.latch/Q
+ mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_24_206 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_200_ _200_/A chanx_right_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_23_261 vgnd vpwr scs8hd_decap_3
XFILLER_15_217 vpwr vgnd scs8hd_fill_2
XANTENNA__209__A _209_/A vgnd vpwr scs8hd_diode_2
X_131_ _110_/A _128_/X _131_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_97 vpwr vgnd scs8hd_fill_2
XFILLER_2_154 vpwr vgnd scs8hd_fill_2
XFILLER_2_132 vpwr vgnd scs8hd_fill_2
XFILLER_0_68 vpwr vgnd scs8hd_fill_2
XANTENNA__119__A _085_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_261 vgnd vpwr scs8hd_decap_12
XFILLER_9_99 vpwr vgnd scs8hd_fill_2
XFILLER_9_88 vgnd vpwr scs8hd_decap_4
Xmem_bottom_track_17.LATCH_2_.latch data_in mem_bottom_track_17.LATCH_2_.latch/Q _151_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _213_/A vgnd vpwr scs8hd_inv_1
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_97 vpwr vgnd scs8hd_fill_2
XFILLER_18_64 vgnd vpwr scs8hd_decap_8
XFILLER_11_231 vpwr vgnd scs8hd_fill_2
X_114_ address[4] _115_/B vgnd vpwr scs8hd_inv_8
XANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB _095_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_6_.scs8hd_inv_1 bottom_left_grid_pin_7_ mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__121__B _119_/B vgnd vpwr scs8hd_diode_2
XFILLER_38_117 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_top_track_0.LATCH_4_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_20_32 vgnd vpwr scs8hd_decap_12
XFILLER_29_74 vgnd vpwr scs8hd_decap_12
XANTENNA__222__A _222_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.INVTX1_7_.scs8hd_inv_1 chany_bottom_in[6] mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_28_150 vgnd vpwr scs8hd_decap_3
XANTENNA__132__A _095_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_67 vpwr vgnd scs8hd_fill_2
XFILLER_6_56 vpwr vgnd scs8hd_fill_2
XFILLER_6_45 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_3 vgnd vpwr scs8hd_decap_12
Xmem_right_track_8.LATCH_1_.latch data_in _183_/A _169_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_208 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_175 vpwr vgnd scs8hd_fill_2
XFILLER_25_131 vpwr vgnd scs8hd_fill_2
XFILLER_40_178 vgnd vpwr scs8hd_decap_8
XANTENNA__217__A _217_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ _178_/A mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_31_86 vgnd vpwr scs8hd_decap_12
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__A _106_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_123 vgnd vpwr scs8hd_decap_12
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _180_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_39_212 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _188_/HI vgnd
+ vpwr scs8hd_diode_2
XFILLER_39_245 vgnd vpwr scs8hd_decap_8
XFILLER_22_123 vgnd vpwr scs8hd_fill_1
Xmux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _191_/HI _182_/Y mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_26_97 vgnd vpwr scs8hd_decap_8
XFILLER_13_167 vpwr vgnd scs8hd_fill_2
XFILLER_13_134 vpwr vgnd scs8hd_fill_2
XFILLER_42_63 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_57 vpwr vgnd scs8hd_fill_2
XFILLER_3_46 vgnd vpwr scs8hd_fill_1
XFILLER_3_35 vpwr vgnd scs8hd_fill_2
XFILLER_36_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_3_.scs8hd_inv_1 chanx_right_in[1] mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _195_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_182 vgnd vpwr scs8hd_decap_8
XFILLER_27_226 vpwr vgnd scs8hd_fill_2
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
XFILLER_12_88 vgnd vpwr scs8hd_decap_4
XFILLER_12_44 vgnd vpwr scs8hd_decap_3
XFILLER_37_74 vgnd vpwr scs8hd_decap_12
XFILLER_18_215 vpwr vgnd scs8hd_fill_2
XFILLER_33_229 vgnd vpwr scs8hd_decap_12
XFILLER_41_251 vgnd vpwr scs8hd_fill_1
XANTENNA__124__B _119_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_163 vgnd vpwr scs8hd_fill_1
XANTENNA__140__A _109_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_1_ vgnd vpwr scs8hd_diode_2
X_130_ _109_/A _128_/X _130_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_240 vpwr vgnd scs8hd_fill_2
XANTENNA__225__A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_23_76 vpwr vgnd scs8hd_fill_2
XANTENNA__119__B _119_/B vgnd vpwr scs8hd_diode_2
XFILLER_0_58 vpwr vgnd scs8hd_fill_2
XFILLER_0_47 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_2_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__135__A _103_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_273 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_2_.scs8hd_inv_1_A top_left_grid_pin_15_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_32 vgnd vpwr scs8hd_decap_12
X_113_ _113_/A _110_/B _113_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_265 vpwr vgnd scs8hd_fill_2
XFILLER_11_254 vpwr vgnd scs8hd_fill_2
XFILLER_11_210 vpwr vgnd scs8hd_fill_2
XFILLER_7_236 vgnd vpwr scs8hd_decap_4
XFILLER_7_269 vgnd vpwr scs8hd_decap_8
XFILLER_7_258 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _182_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_38_129 vgnd vpwr scs8hd_decap_12
Xmux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ _186_/A mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1_A bottom_right_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_37_184 vgnd vpwr scs8hd_decap_12
XFILLER_20_44 vgnd vpwr scs8hd_decap_12
XFILLER_4_206 vgnd vpwr scs8hd_decap_3
XFILLER_29_86 vgnd vpwr scs8hd_decap_12
XFILLER_28_184 vpwr vgnd scs8hd_fill_2
XANTENNA__132__B _128_/X vgnd vpwr scs8hd_diode_2
XFILLER_19_184 vpwr vgnd scs8hd_fill_2
XFILLER_34_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1_A bottom_left_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_165 vpwr vgnd scs8hd_fill_2
XFILLER_25_110 vgnd vpwr scs8hd_fill_1
XFILLER_15_88 vpwr vgnd scs8hd_fill_2
XFILLER_31_98 vgnd vpwr scs8hd_decap_12
XFILLER_0_242 vgnd vpwr scs8hd_decap_4
XFILLER_0_231 vgnd vpwr scs8hd_decap_4
XFILLER_16_132 vpwr vgnd scs8hd_fill_2
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__B _167_/B vgnd vpwr scs8hd_diode_2
XFILLER_31_135 vgnd vpwr scs8hd_decap_12
XFILLER_16_176 vpwr vgnd scs8hd_fill_2
XANTENNA__143__A _098_/B vgnd vpwr scs8hd_diode_2
XFILLER_39_224 vgnd vpwr scs8hd_decap_8
XFILLER_22_157 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _173_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_32 vgnd vpwr scs8hd_decap_12
XFILLER_13_146 vgnd vpwr scs8hd_fill_1
XFILLER_13_113 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _180_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_42_75 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _209_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1_A bottom_left_grid_pin_3_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.INVTX1_2_.scs8hd_inv_1_A right_bottom_grid_pin_12_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA__138__A _137_/X vgnd vpwr scs8hd_diode_2
XFILLER_36_227 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_205 vgnd vpwr scs8hd_decap_4
XFILLER_12_67 vpwr vgnd scs8hd_fill_2
XFILLER_37_86 vgnd vpwr scs8hd_decap_12
XFILLER_5_175 vpwr vgnd scs8hd_fill_2
XFILLER_5_142 vpwr vgnd scs8hd_fill_2
XANTENNA__140__B _138_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_260 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_14.LATCH_1_.latch_SLEEPB _171_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_230 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_145 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_189_ _189_/HI _189_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_right_track_12.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr
+ scs8hd_diode_2
XANTENNA__135__B _115_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_57 vpwr vgnd scs8hd_fill_2
XANTENNA__151__A _095_/B vgnd vpwr scs8hd_diode_2
XFILLER_36_3 vgnd vpwr scs8hd_decap_12
XFILLER_20_266 vgnd vpwr scs8hd_decap_8
XFILLER_20_255 vgnd vpwr scs8hd_decap_8
XFILLER_18_44 vgnd vpwr scs8hd_decap_12
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
XFILLER_18_88 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
X_112_ _098_/B _110_/B _112_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__146__A _160_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _175_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_196 vgnd vpwr scs8hd_decap_12
XFILLER_1_80 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_track_1.LATCH_5_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _173_/A mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_20_56 vgnd vpwr scs8hd_decap_12
XFILLER_4_229 vpwr vgnd scs8hd_fill_2
XFILLER_4_218 vgnd vpwr scs8hd_decap_3
XFILLER_29_98 vgnd vpwr scs8hd_decap_12
XFILLER_28_163 vgnd vpwr scs8hd_decap_3
XFILLER_34_166 vgnd vpwr scs8hd_decap_12
XFILLER_25_100 vgnd vpwr scs8hd_decap_8
XFILLER_15_67 vpwr vgnd scs8hd_fill_2
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__C _169_/C vgnd vpwr scs8hd_diode_2
XFILLER_31_147 vgnd vpwr scs8hd_decap_12
XANTENNA__143__B _138_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_236 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
Xmem_right_track_4.LATCH_1_.latch data_in _175_/A _161_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_2.LATCH_0_.latch_SLEEPB _159_/Y vgnd vpwr scs8hd_diode_2
XFILLER_26_44 vgnd vpwr scs8hd_decap_12
XFILLER_42_87 vgnd vpwr scs8hd_decap_6
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XFILLER_9_118 vpwr vgnd scs8hd_fill_2
Xmux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ _177_/Y mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_3_15 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_17.INVTX1_4_.scs8hd_inv_1 chanx_right_in[8] mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_36_239 vgnd vpwr scs8hd_decap_12
XANTENNA__154__A _106_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_14.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[0] mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_10_106 vgnd vpwr scs8hd_decap_4
XFILLER_5_7 vgnd vpwr scs8hd_decap_12
XFILLER_18_206 vgnd vpwr scs8hd_decap_6
XFILLER_37_98 vgnd vpwr scs8hd_decap_12
XFILLER_41_220 vgnd vpwr scs8hd_decap_12
XFILLER_26_250 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmem_top_track_0.LATCH_0_.latch data_in mem_top_track_0.LATCH_0_.latch/Q _101_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_132 vgnd vpwr scs8hd_decap_4
XANTENNA__149__A _109_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_track_17.LATCH_3_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_113 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.INVTX1_7_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_9_69 vpwr vgnd scs8hd_fill_2
XFILLER_9_47 vgnd vpwr scs8hd_fill_1
X_188_ _188_/HI _188_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__135__C _081_/C vgnd vpwr scs8hd_diode_2
Xmux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _179_/A mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__151__B _149_/B vgnd vpwr scs8hd_diode_2
XFILLER_29_3 vgnd vpwr scs8hd_decap_12
Xmux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _193_/HI _174_/Y mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_56 vgnd vpwr scs8hd_decap_6
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
X_111_ _095_/B _110_/B _111_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA__146__B _125_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__162__A _163_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_14.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_68 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _196_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_197 vpwr vgnd scs8hd_fill_2
XFILLER_3_230 vpwr vgnd scs8hd_fill_2
XANTENNA__157__A _157_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_178 vgnd vpwr scs8hd_decap_12
XFILLER_19_164 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_1.LATCH_2_.latch data_in mem_bottom_track_1.LATCH_2_.latch/Q _132_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _192_/HI _185_/Y mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_3_.latch_SLEEPB _110_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_200 vpwr vgnd scs8hd_fill_2
XFILLER_16_189 vpwr vgnd scs8hd_fill_2
XFILLER_16_167 vgnd vpwr scs8hd_decap_6
XFILLER_16_145 vgnd vpwr scs8hd_decap_6
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_159 vgnd vpwr scs8hd_decap_4
XFILLER_39_259 vpwr vgnd scs8hd_fill_2
XFILLER_11_3 vgnd vpwr scs8hd_decap_12
XFILLER_22_148 vgnd vpwr scs8hd_fill_1
XFILLER_22_126 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_91 vpwr vgnd scs8hd_fill_2
XFILLER_26_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XFILLER_21_192 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_270 vgnd vpwr scs8hd_decap_6
XFILLER_3_49 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ _176_/A mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_8_152 vgnd vpwr scs8hd_fill_1
XANTENNA__170__A _160_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__080__A enable vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_41_232 vgnd vpwr scs8hd_decap_12
XFILLER_26_262 vgnd vpwr scs8hd_decap_12
XFILLER_41_276 vgnd vpwr scs8hd_fill_1
XFILLER_5_155 vpwr vgnd scs8hd_fill_2
Xmux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _190_/HI _180_/Y mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_188 vgnd vpwr scs8hd_fill_1
XANTENNA__149__B _149_/B vgnd vpwr scs8hd_diode_2
XANTENNA__165__A _163_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_243 vgnd vpwr scs8hd_fill_1
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XANTENNA__075__A address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_12.INVTX1_0_.scs8hd_inv_1 chany_top_in[6] mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_169 vgnd vpwr scs8hd_decap_8
XFILLER_2_158 vpwr vgnd scs8hd_fill_2
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
XFILLER_14_232 vgnd vpwr scs8hd_decap_3
XFILLER_9_15 vgnd vpwr scs8hd_decap_12
X_187_ _187_/HI _187_/LO vgnd vpwr scs8hd_conb_1
Xmux_bottom_track_9.INVTX1_3_.scs8hd_inv_1 chanx_right_in[3] mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ _184_/Y mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_110_ _110_/A _110_/B _110_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_34_56 vgnd vpwr scs8hd_decap_12
XFILLER_11_235 vgnd vpwr scs8hd_decap_3
XFILLER_7_217 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _179_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA__146__C _162_/C vgnd vpwr scs8hd_diode_2
XANTENNA__162__B _155_/X vgnd vpwr scs8hd_diode_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XFILLER_6_272 vgnd vpwr scs8hd_decap_3
Xmux_top_track_16.INVTX1_4_.scs8hd_inv_1 chanx_right_in[3] mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_37_110 vgnd vpwr scs8hd_decap_12
XFILLER_1_60 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_154 vgnd vpwr scs8hd_decap_6
XFILLER_10_91 vgnd vpwr scs8hd_fill_1
XANTENNA__157__B _155_/X vgnd vpwr scs8hd_diode_2
XANTENNA__173__A _173_/A vgnd vpwr scs8hd_diode_2
XFILLER_25_135 vpwr vgnd scs8hd_fill_2
Xmux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ _182_/A mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__083__A _106_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_105 vgnd vpwr scs8hd_decap_12
XFILLER_25_179 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_102 vpwr vgnd scs8hd_fill_2
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__168__A _157_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_182 vgnd vpwr scs8hd_decap_4
Xmux_top_track_0.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_1_ mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__078__A _077_/X vgnd vpwr scs8hd_diode_2
XFILLER_38_271 vgnd vpwr scs8hd_decap_4
XFILLER_26_68 vgnd vpwr scs8hd_decap_6
XFILLER_13_138 vpwr vgnd scs8hd_fill_2
XFILLER_42_56 vgnd vpwr scs8hd_decap_6
XANTENNA__170__B _155_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A top_right_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_263 vgnd vpwr scs8hd_decap_12
XFILLER_12_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[4] mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_230 vgnd vpwr scs8hd_decap_6
XFILLER_18_219 vgnd vpwr scs8hd_fill_1
XFILLER_26_274 vgnd vpwr scs8hd_fill_1
Xmem_top_track_8.LATCH_1_.latch data_in mem_top_track_8.LATCH_1_.latch/Q _112_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _181_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_241 vgnd vpwr scs8hd_decap_3
XFILLER_17_230 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__165__B _155_/A vgnd vpwr scs8hd_diode_2
XANTENNA__181__A _181_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_93 vgnd vpwr scs8hd_fill_1
XFILLER_4_71 vpwr vgnd scs8hd_fill_2
XANTENNA__091__A _090_/X vgnd vpwr scs8hd_diode_2
XFILLER_2_104 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_3_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_244 vgnd vpwr scs8hd_decap_8
XFILLER_9_27 vgnd vpwr scs8hd_decap_12
X_186_ _186_/A _186_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _176_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_181 vpwr vgnd scs8hd_fill_2
XANTENNA__176__A _176_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_6_.scs8hd_inv_1 bottom_left_grid_pin_5_ mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__086__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_34_68 vgnd vpwr scs8hd_decap_12
XFILLER_11_269 vgnd vpwr scs8hd_decap_8
XFILLER_11_258 vgnd vpwr scs8hd_decap_4
XFILLER_1_3 vgnd vpwr scs8hd_decap_8
Xmux_top_track_8.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_169_ _160_/A _155_/A _169_/C _163_/D _169_/Y vgnd vpwr scs8hd_nor4_4
Xmux_right_track_10.INVTX1_0_.scs8hd_inv_1 chany_top_in[5] mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__162__C _162_/C vgnd vpwr scs8hd_diode_2
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB _119_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_265 vpwr vgnd scs8hd_fill_2
XFILLER_3_254 vpwr vgnd scs8hd_fill_2
XFILLER_19_90 vpwr vgnd scs8hd_fill_2
XANTENNA__157__C _136_/X vgnd vpwr scs8hd_diode_2
XFILLER_42_180 vgnd vpwr scs8hd_decap_6
Xmem_bottom_track_9.LATCH_3_.latch data_in mem_bottom_track_9.LATCH_3_.latch/Q _141_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_40_117 vgnd vpwr scs8hd_decap_12
XFILLER_25_169 vgnd vpwr scs8hd_decap_4
XFILLER_25_114 vpwr vgnd scs8hd_fill_2
XFILLER_15_15 vgnd vpwr scs8hd_decap_12
XANTENNA__083__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_0_213 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _174_/Y vgnd vpwr
+ scs8hd_diode_2
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA__168__B _167_/B vgnd vpwr scs8hd_diode_2
XANTENNA__184__A _184_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_7_71 vpwr vgnd scs8hd_fill_2
XANTENNA__094__A _093_/X vgnd vpwr scs8hd_diode_2
XFILLER_13_117 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _178_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_194 vpwr vgnd scs8hd_fill_2
XFILLER_12_150 vgnd vpwr scs8hd_fill_1
XANTENNA__170__C _169_/C vgnd vpwr scs8hd_diode_2
XFILLER_8_165 vpwr vgnd scs8hd_fill_2
XANTENNA__179__A _179_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_220 vgnd vpwr scs8hd_decap_12
XFILLER_35_253 vpwr vgnd scs8hd_fill_2
XFILLER_35_275 vpwr vgnd scs8hd_fill_2
XFILLER_12_27 vgnd vpwr scs8hd_decap_4
Xmux_right_track_12.tap_buf4_0_.scs8hd_inv_1 mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ _202_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_track_17.LATCH_4_.latch_SLEEPB _149_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_3_.latch data_in mem_top_track_16.LATCH_3_.latch/Q _121_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__089__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_41_256 vpwr vgnd scs8hd_fill_2
XFILLER_41_245 vgnd vpwr scs8hd_decap_6
XFILLER_5_179 vpwr vgnd scs8hd_fill_2
XANTENNA__165__C _136_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _175_/Y mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_4_50 vgnd vpwr scs8hd_decap_3
XFILLER_23_267 vpwr vgnd scs8hd_fill_2
XFILLER_23_256 vgnd vpwr scs8hd_decap_3
XFILLER_23_234 vgnd vpwr scs8hd_decap_4
XFILLER_23_223 vpwr vgnd scs8hd_fill_2
XFILLER_23_59 vpwr vgnd scs8hd_fill_2
XFILLER_23_15 vgnd vpwr scs8hd_decap_12
XFILLER_2_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_14_201 vpwr vgnd scs8hd_fill_2
X_185_ _185_/A _185_/Y vgnd vpwr scs8hd_inv_8
XFILLER_13_92 vpwr vgnd scs8hd_fill_2
XFILLER_9_39 vgnd vpwr scs8hd_decap_8
Xmux_right_track_6.INVTX1_1_.scs8hd_inv_1 chany_top_in[8] mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_193 vgnd vpwr scs8hd_decap_4
XFILLER_1_171 vgnd vpwr scs8hd_decap_4
XFILLER_20_215 vgnd vpwr scs8hd_decap_4
XFILLER_9_271 vgnd vpwr scs8hd_decap_6
XFILLER_9_260 vpwr vgnd scs8hd_fill_2
XFILLER_18_15 vgnd vpwr scs8hd_decap_12
XANTENNA__086__B _075_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _176_/A vgnd vpwr
+ scs8hd_diode_2
X_168_ _157_/A _167_/B _162_/C _162_/D _168_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__162__D _162_/D vgnd vpwr scs8hd_diode_2
X_099_ address[1] address[2] address[0] _099_/X vgnd vpwr scs8hd_or3_4
XFILLER_27_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_123 vgnd vpwr scs8hd_decap_12
XFILLER_1_95 vpwr vgnd scs8hd_fill_2
XFILLER_1_62 vpwr vgnd scs8hd_fill_2
XFILLER_20_27 vgnd vpwr scs8hd_decap_4
XANTENNA__097__A _096_/X vgnd vpwr scs8hd_diode_2
XFILLER_6_18 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_189 vpwr vgnd scs8hd_fill_2
XFILLER_19_123 vgnd vpwr scs8hd_decap_3
XANTENNA__157__D _163_/D vgnd vpwr scs8hd_diode_2
XFILLER_40_129 vgnd vpwr scs8hd_decap_12
XFILLER_25_148 vpwr vgnd scs8hd_fill_2
XFILLER_25_126 vgnd vpwr scs8hd_decap_3
XFILLER_15_27 vgnd vpwr scs8hd_decap_12
XANTENNA__083__C _162_/C vgnd vpwr scs8hd_diode_2
XFILLER_31_15 vgnd vpwr scs8hd_decap_12
XFILLER_31_59 vpwr vgnd scs8hd_fill_2
XFILLER_0_269 vpwr vgnd scs8hd_fill_2
XFILLER_0_258 vgnd vpwr scs8hd_decap_8
Xmem_bottom_track_17.LATCH_3_.latch data_in mem_bottom_track_17.LATCH_3_.latch/Q _150_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_181 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_70 vpwr vgnd scs8hd_fill_2
XPHY_1 vgnd vpwr scs8hd_decap_3
XANTENNA__168__C _162_/C vgnd vpwr scs8hd_diode_2
XFILLER_7_83 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_17.INVTX1_1_.scs8hd_inv_1 chany_top_in[6] mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_6.tap_buf4_0_.scs8hd_inv_1 mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ _205_/A vgnd vpwr scs8hd_inv_1
XFILLER_38_251 vgnd vpwr scs8hd_decap_4
XFILLER_26_15 vgnd vpwr scs8hd_decap_12
XFILLER_21_162 vpwr vgnd scs8hd_fill_2
Xmux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ _181_/Y mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_21_184 vgnd vpwr scs8hd_fill_1
XFILLER_29_240 vpwr vgnd scs8hd_fill_2
XFILLER_32_80 vgnd vpwr scs8hd_decap_12
XFILLER_12_184 vpwr vgnd scs8hd_fill_2
XFILLER_8_144 vpwr vgnd scs8hd_fill_2
XFILLER_8_111 vgnd vpwr scs8hd_fill_1
XANTENNA__170__D _162_/D vgnd vpwr scs8hd_diode_2
XFILLER_35_232 vgnd vpwr scs8hd_decap_12
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
XFILLER_5_114 vpwr vgnd scs8hd_fill_2
XANTENNA__165__D _163_/D vgnd vpwr scs8hd_diode_2
XFILLER_32_213 vgnd vpwr scs8hd_fill_1
XFILLER_32_224 vgnd vpwr scs8hd_decap_8
XFILLER_32_235 vgnd vpwr scs8hd_decap_8
XFILLER_17_265 vpwr vgnd scs8hd_fill_2
XFILLER_17_254 vgnd vpwr scs8hd_decap_4
XFILLER_4_84 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_2_.latch/Q mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ _174_/A mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_10.LATCH_0_.latch_SLEEPB _166_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_27 vgnd vpwr scs8hd_decap_12
XFILLER_2_128 vpwr vgnd scs8hd_fill_2
XFILLER_14_224 vpwr vgnd scs8hd_fill_2
X_184_ _184_/A _184_/Y vgnd vpwr scs8hd_inv_8
Xmux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_0.LATCH_5_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_20_238 vgnd vpwr scs8hd_decap_8
XFILLER_20_205 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_27 vgnd vpwr scs8hd_decap_4
XANTENNA__086__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_098_ _085_/B _098_/B _098_/Y vgnd vpwr scs8hd_nor2_4
X_167_ _157_/A _167_/B _162_/C _163_/D _167_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_40_91 vgnd vpwr scs8hd_fill_1
XFILLER_6_264 vgnd vpwr scs8hd_decap_8
XFILLER_6_253 vpwr vgnd scs8hd_fill_2
XFILLER_37_135 vgnd vpwr scs8hd_decap_12
Xmux_right_track_4.INVTX1_1_.scs8hd_inv_1 chany_top_in[7] mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_59 vpwr vgnd scs8hd_fill_2
XFILLER_28_168 vgnd vpwr scs8hd_decap_3
Xmux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ _178_/Y mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB _113_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_234 vpwr vgnd scs8hd_fill_2
XFILLER_3_201 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_102 vgnd vpwr scs8hd_fill_1
XFILLER_10_83 vpwr vgnd scs8hd_fill_2
XFILLER_34_105 vgnd vpwr scs8hd_decap_12
XFILLER_19_179 vpwr vgnd scs8hd_fill_2
X_219_ chany_bottom_in[6] chany_top_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_33_171 vgnd vpwr scs8hd_decap_12
XFILLER_15_39 vgnd vpwr scs8hd_decap_12
XFILLER_31_27 vgnd vpwr scs8hd_decap_12
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _198_/HI mem_top_track_16.LATCH_2_.latch/Q
+ mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_208 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XANTENNA__168__D _162_/D vgnd vpwr scs8hd_diode_2
XFILLER_22_119 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_141 vgnd vpwr scs8hd_decap_12
XFILLER_26_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_8.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _182_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XFILLER_21_141 vgnd vpwr scs8hd_fill_1
Xmux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ _180_/A mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A top_left_grid_pin_7_ vgnd vpwr scs8hd_diode_2
XFILLER_37_15 vgnd vpwr scs8hd_decap_12
XFILLER_37_59 vpwr vgnd scs8hd_fill_2
XFILLER_26_211 vgnd vpwr scs8hd_fill_1
XFILLER_5_159 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_247 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_23_39 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_183_ _183_/A _183_/Y vgnd vpwr scs8hd_inv_8
XFILLER_38_80 vgnd vpwr scs8hd_decap_12
Xmux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ _186_/Y mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1_A bottom_left_grid_pin_5_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _180_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
XFILLER_11_206 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.INVTX1_1_.scs8hd_inv_1 top_left_grid_pin_11_ mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_210 vpwr vgnd scs8hd_fill_2
X_097_ _096_/X _098_/B vgnd vpwr scs8hd_buf_1
X_166_ _163_/A _155_/A _136_/X _162_/D _166_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
XFILLER_6_243 vgnd vpwr scs8hd_fill_1
XFILLER_37_147 vgnd vpwr scs8hd_decap_12
XFILLER_1_53 vgnd vpwr scs8hd_decap_4
XFILLER_1_42 vpwr vgnd scs8hd_fill_2
XFILLER_1_31 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.LATCH_4_.latch_SLEEPB _140_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _186_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_29_27 vgnd vpwr scs8hd_decap_12
XFILLER_10_62 vpwr vgnd scs8hd_fill_2
XFILLER_10_51 vgnd vpwr scs8hd_decap_8
XFILLER_3_213 vpwr vgnd scs8hd_fill_2
XFILLER_19_147 vpwr vgnd scs8hd_fill_2
XFILLER_19_114 vpwr vgnd scs8hd_fill_2
XFILLER_19_71 vpwr vgnd scs8hd_fill_2
XFILLER_34_117 vgnd vpwr scs8hd_decap_12
X_149_ _109_/A _149_/B _149_/Y vgnd vpwr scs8hd_nor2_4
X_218_ _218_/A chany_top_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_32_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_39 vgnd vpwr scs8hd_decap_12
XFILLER_0_238 vpwr vgnd scs8hd_fill_2
XFILLER_0_227 vpwr vgnd scs8hd_fill_2
Xmux_right_track_2.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_128 vpwr vgnd scs8hd_fill_2
XFILLER_16_106 vgnd vpwr scs8hd_decap_12
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1_A bottom_left_grid_pin_9_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_83 vpwr vgnd scs8hd_fill_2
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_15_161 vpwr vgnd scs8hd_fill_2
XFILLER_30_186 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _189_/HI mem_bottom_track_9.LATCH_2_.latch/Q
+ mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_13_109 vpwr vgnd scs8hd_fill_2
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XFILLER_21_175 vpwr vgnd scs8hd_fill_2
XFILLER_21_153 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_142 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _175_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_93 vgnd vpwr scs8hd_decap_12
XFILLER_35_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _182_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_37_27 vgnd vpwr scs8hd_decap_12
XFILLER_26_245 vgnd vpwr scs8hd_decap_3
XFILLER_5_138 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_234 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_12.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB _134_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_259 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_108 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_182_ _182_/A _182_/Y vgnd vpwr scs8hd_inv_8
Xmux_bottom_track_1.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_73 vpwr vgnd scs8hd_fill_2
XFILLER_13_62 vpwr vgnd scs8hd_fill_2
XANTENNA__100__A _099_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_2_.scs8hd_inv_1 top_left_grid_pin_15_ mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _173_/Y mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_165_ _163_/A _155_/A _136_/X _163_/D _165_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB _122_/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_72 vgnd vpwr scs8hd_fill_1
XFILLER_10_273 vpwr vgnd scs8hd_fill_2
X_096_ address[1] address[2] _156_/A _096_/X vgnd vpwr scs8hd_or3_4
XFILLER_40_93 vgnd vpwr scs8hd_decap_12
XFILLER_40_71 vgnd vpwr scs8hd_decap_12
XFILLER_37_159 vgnd vpwr scs8hd_decap_12
XFILLER_1_76 vpwr vgnd scs8hd_fill_2
Xmem_top_track_0.LATCH_1_.latch data_in mem_top_track_0.LATCH_1_.latch/Q _098_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_39 vgnd vpwr scs8hd_decap_12
XFILLER_3_269 vgnd vpwr scs8hd_decap_8
XFILLER_3_258 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _177_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_94 vpwr vgnd scs8hd_fill_2
XFILLER_34_129 vgnd vpwr scs8hd_decap_12
X_148_ _085_/A _149_/B _148_/Y vgnd vpwr scs8hd_nor2_4
X_217_ _217_/A chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
X_079_ address[5] _106_/A vgnd vpwr scs8hd_buf_1
XFILLER_25_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.INVTX1_1_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_25_118 vpwr vgnd scs8hd_fill_2
XFILLER_33_184 vgnd vpwr scs8hd_decap_12
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_151 vpwr vgnd scs8hd_fill_2
XFILLER_16_118 vgnd vpwr scs8hd_fill_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_62 vgnd vpwr scs8hd_decap_8
XFILLER_21_51 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB _088_/Y vgnd vpwr scs8hd_diode_2
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_30_154 vgnd vpwr scs8hd_decap_8
XFILLER_30_165 vgnd vpwr scs8hd_decap_8
XFILLER_15_195 vpwr vgnd scs8hd_fill_2
XFILLER_7_75 vpwr vgnd scs8hd_fill_2
XFILLER_7_53 vpwr vgnd scs8hd_fill_2
XFILLER_7_42 vgnd vpwr scs8hd_decap_3
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_21_110 vgnd vpwr scs8hd_fill_1
XFILLER_29_232 vgnd vpwr scs8hd_decap_6
XFILLER_29_254 vpwr vgnd scs8hd_fill_2
XFILLER_29_276 vgnd vpwr scs8hd_fill_1
XFILLER_16_84 vpwr vgnd scs8hd_fill_2
XFILLER_12_165 vpwr vgnd scs8hd_fill_2
XFILLER_8_114 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB _152_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_169 vpwr vgnd scs8hd_fill_2
XANTENNA__103__A address[3] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_track_17.LATCH_4_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_14.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_191 vpwr vgnd scs8hd_fill_2
XFILLER_37_39 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_1.LATCH_3_.latch data_in mem_bottom_track_1.LATCH_3_.latch/Q _131_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
Xmux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ _179_/Y mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_40_271 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_183 vgnd vpwr scs8hd_fill_1
XFILLER_4_32 vgnd vpwr scs8hd_decap_4
XFILLER_14_205 vpwr vgnd scs8hd_fill_2
X_181_ _181_/A _181_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
Xmem_right_track_14.LATCH_0_.latch data_in _186_/A _172_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_96 vpwr vgnd scs8hd_fill_2
XFILLER_1_142 vgnd vpwr scs8hd_fill_1
XFILLER_38_93 vgnd vpwr scs8hd_decap_12
XFILLER_1_197 vgnd vpwr scs8hd_fill_1
XFILLER_9_231 vpwr vgnd scs8hd_fill_2
XFILLER_9_220 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.INVTX1_5_.scs8hd_inv_1 chanx_right_in[7] mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__201__A _201_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_190 vpwr vgnd scs8hd_fill_2
X_095_ _085_/B _095_/B _095_/Y vgnd vpwr scs8hd_nor2_4
X_164_ _163_/A _155_/X _163_/C _162_/D _164_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_24_84 vgnd vpwr scs8hd_decap_8
XFILLER_10_252 vpwr vgnd scs8hd_fill_2
XFILLER_40_83 vgnd vpwr scs8hd_decap_8
XANTENNA__111__A _095_/B vgnd vpwr scs8hd_diode_2
XFILLER_1_99 vgnd vpwr scs8hd_decap_4
XFILLER_1_66 vgnd vpwr scs8hd_fill_1
XFILLER_1_22 vgnd vpwr scs8hd_decap_6
XFILLER_1_11 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_12.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_138 vgnd vpwr scs8hd_decap_12
XFILLER_28_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_51 vgnd vpwr scs8hd_decap_8
X_078_ _077_/X _085_/A vgnd vpwr scs8hd_buf_1
X_147_ _146_/X _149_/B vgnd vpwr scs8hd_buf_1
X_216_ chany_top_in[0] chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA__106__A _106_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_270 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_33_196 vgnd vpwr scs8hd_decap_3
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_185 vpwr vgnd scs8hd_fill_2
XFILLER_24_163 vgnd vpwr scs8hd_decap_3
Xmux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_top_track_16.LATCH_3_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XPHY_5 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_2_.latch/Q mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ _176_/Y mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_15_174 vgnd vpwr scs8hd_decap_3
XFILLER_7_87 vpwr vgnd scs8hd_fill_2
XFILLER_21_133 vpwr vgnd scs8hd_fill_2
XFILLER_21_188 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_266 vpwr vgnd scs8hd_fill_2
XFILLER_12_188 vgnd vpwr scs8hd_decap_4
XFILLER_8_148 vgnd vpwr scs8hd_decap_4
XFILLER_8_137 vgnd vpwr scs8hd_decap_3
XFILLER_26_203 vpwr vgnd scs8hd_fill_2
XFILLER_5_118 vpwr vgnd scs8hd_fill_2
XANTENNA__204__A _204_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_62 vgnd vpwr scs8hd_decap_12
XFILLER_27_51 vgnd vpwr scs8hd_decap_8
XFILLER_17_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_6.LATCH_0_.latch_SLEEPB _164_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__114__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_4_88 vpwr vgnd scs8hd_fill_2
XFILLER_4_55 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_228 vpwr vgnd scs8hd_fill_2
X_180_ _180_/A _180_/Y vgnd vpwr scs8hd_inv_8
XFILLER_13_53 vpwr vgnd scs8hd_fill_2
XFILLER_13_42 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_154 vpwr vgnd scs8hd_fill_2
XFILLER_1_132 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__109__A _109_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_209 vgnd vpwr scs8hd_decap_3
X_094_ _093_/X _095_/B vgnd vpwr scs8hd_buf_1
X_163_ _163_/A _155_/X _163_/C _163_/D _163_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_24_96 vgnd vpwr scs8hd_decap_4
XFILLER_6_257 vgnd vpwr scs8hd_decap_4
XFILLER_6_235 vpwr vgnd scs8hd_fill_2
XFILLER_6_224 vgnd vpwr scs8hd_decap_3
XFILLER_6_202 vpwr vgnd scs8hd_fill_2
XANTENNA__111__B _110_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _199_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.LATCH_2_.latch data_in mem_top_track_8.LATCH_2_.latch/Q _111_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _181_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_28_117 vgnd vpwr scs8hd_decap_12
Xmux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ _182_/Y mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__212__A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_10_87 vgnd vpwr scs8hd_decap_4
XFILLER_10_32 vgnd vpwr scs8hd_decap_12
XFILLER_3_238 vgnd vpwr scs8hd_decap_4
Xmux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_35_51 vgnd vpwr scs8hd_decap_8
XFILLER_19_139 vgnd vpwr scs8hd_decap_8
X_215_ chany_top_in[1] chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_35_62 vgnd vpwr scs8hd_decap_12
X_077_ address[1] _075_/Y _156_/A _077_/X vgnd vpwr scs8hd_or3_4
X_146_ _160_/A _125_/Y _162_/C _146_/X vgnd vpwr scs8hd_or3_4
XANTENNA__122__A _095_/B vgnd vpwr scs8hd_diode_2
XANTENNA__106__B _155_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_4.LATCH_1_.latch_SLEEPB _161_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_208 vgnd vpwr scs8hd_decap_3
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__207__A _207_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_15_142 vgnd vpwr scs8hd_decap_4
XANTENNA__117__A _106_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_189 vgnd vpwr scs8hd_decap_6
X_129_ _085_/A _128_/X _129_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_30_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_track_9.LATCH_3_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_123 vgnd vpwr scs8hd_fill_1
Xmux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_2_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_35_259 vpwr vgnd scs8hd_fill_2
XFILLER_7_182 vgnd vpwr scs8hd_fill_1
XFILLER_26_226 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_9.LATCH_4_.latch data_in mem_bottom_track_9.LATCH_4_.latch/Q _140_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__220__A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _190_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_17_204 vpwr vgnd scs8hd_fill_2
XFILLER_32_207 vgnd vpwr scs8hd_decap_6
XFILLER_27_74 vgnd vpwr scs8hd_decap_12
XANTENNA__130__A _109_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_152 vgnd vpwr scs8hd_fill_1
XFILLER_4_67 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _185_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA__215__A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_8_3 vgnd vpwr scs8hd_decap_12
XFILLER_1_177 vpwr vgnd scs8hd_fill_2
XANTENNA__109__B _110_/B vgnd vpwr scs8hd_diode_2
XFILLER_13_262 vpwr vgnd scs8hd_fill_2
XFILLER_13_240 vpwr vgnd scs8hd_fill_2
XANTENNA__125__A address[6] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_6_.scs8hd_inv_1 bottom_left_grid_pin_9_ mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _178_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB _143_/Y vgnd vpwr scs8hd_diode_2
XFILLER_39_170 vgnd vpwr scs8hd_fill_1
X_162_ _163_/A _155_/X _162_/C _162_/D _162_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_10_210 vpwr vgnd scs8hd_fill_2
X_093_ _090_/A address[2] address[0] _093_/X vgnd vpwr scs8hd_or3_4
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
XFILLER_10_265 vgnd vpwr scs8hd_decap_8
Xmem_top_track_16.LATCH_4_.latch data_in mem_top_track_16.LATCH_4_.latch/Q _120_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_46 vpwr vgnd scs8hd_fill_2
XFILLER_1_35 vpwr vgnd scs8hd_fill_2
Xmem_right_track_10.LATCH_0_.latch data_in _180_/A _166_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_57 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_44 vgnd vpwr scs8hd_decap_4
XFILLER_3_217 vpwr vgnd scs8hd_fill_2
XFILLER_19_118 vpwr vgnd scs8hd_fill_2
XFILLER_10_66 vpwr vgnd scs8hd_fill_2
XFILLER_35_74 vgnd vpwr scs8hd_decap_12
XFILLER_27_184 vpwr vgnd scs8hd_fill_2
XFILLER_27_162 vpwr vgnd scs8hd_fill_2
XFILLER_19_75 vpwr vgnd scs8hd_fill_2
X_145_ address[5] _160_/A vgnd vpwr scs8hd_inv_8
X_214_ chany_top_in[2] chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA__106__C _163_/C vgnd vpwr scs8hd_diode_2
XFILLER_42_187 vgnd vpwr scs8hd_decap_12
X_076_ address[0] _156_/A vgnd vpwr scs8hd_inv_8
XANTENNA__122__B _119_/B vgnd vpwr scs8hd_diode_2
XFILLER_18_140 vgnd vpwr scs8hd_decap_8
XFILLER_33_110 vgnd vpwr scs8hd_decap_12
XFILLER_18_184 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_10.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_132 vpwr vgnd scs8hd_fill_2
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__223__A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_21_87 vpwr vgnd scs8hd_fill_2
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_132 vgnd vpwr scs8hd_decap_4
X_128_ _127_/X _128_/X vgnd vpwr scs8hd_buf_1
XANTENNA__117__B address[6] vgnd vpwr scs8hd_diode_2
XANTENNA__133__A _098_/B vgnd vpwr scs8hd_diode_2
XFILLER_38_202 vgnd vpwr scs8hd_decap_12
XFILLER_23_3 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _176_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_179 vpwr vgnd scs8hd_fill_2
XFILLER_21_157 vgnd vpwr scs8hd_decap_3
XFILLER_21_102 vpwr vgnd scs8hd_fill_2
XFILLER_16_32 vgnd vpwr scs8hd_decap_12
XFILLER_12_102 vpwr vgnd scs8hd_fill_2
XANTENNA__218__A _218_/A vgnd vpwr scs8hd_diode_2
XANTENNA__128__A _127_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _184_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_41_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_8.LATCH_5_.latch_SLEEPB _108_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_7_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_27_86 vgnd vpwr scs8hd_decap_12
XFILLER_17_238 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_17.LATCH_4_.latch data_in mem_bottom_track_17.LATCH_4_.latch/Q _149_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_1.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__130__B _128_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_186 vgnd vpwr scs8hd_decap_3
XFILLER_23_219 vpwr vgnd scs8hd_fill_2
XFILLER_16_260 vgnd vpwr scs8hd_decap_12
XFILLER_31_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_77 vpwr vgnd scs8hd_fill_2
XFILLER_13_66 vpwr vgnd scs8hd_fill_2
Xmem_right_track_6.LATCH_0_.latch data_in _178_/A _164_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_274 vgnd vpwr scs8hd_decap_3
XFILLER_9_267 vpwr vgnd scs8hd_fill_2
XFILLER_9_256 vpwr vgnd scs8hd_fill_2
XFILLER_9_245 vpwr vgnd scs8hd_fill_2
XANTENNA__141__A _110_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_161_ _163_/A _155_/X _162_/C _163_/D _161_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_24_32 vgnd vpwr scs8hd_decap_12
XFILLER_10_233 vgnd vpwr scs8hd_decap_6
XFILLER_10_222 vpwr vgnd scs8hd_fill_2
XANTENNA__226__A _226_/A vgnd vpwr scs8hd_diode_2
X_092_ _085_/B _110_/A _092_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__136__A _135_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _178_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_141 vgnd vpwr scs8hd_decap_12
XFILLER_19_98 vgnd vpwr scs8hd_decap_4
Xmux_right_track_12.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[7] mux_right_track_12.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_86 vgnd vpwr scs8hd_decap_12
XFILLER_27_152 vgnd vpwr scs8hd_fill_1
X_075_ address[2] _075_/Y vgnd vpwr scs8hd_inv_8
X_144_ _113_/A _138_/X _144_/Y vgnd vpwr scs8hd_nor2_4
X_213_ _213_/A chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
Xmux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _199_/HI mem_top_track_8.LATCH_2_.latch/Q
+ mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_42_199 vgnd vpwr scs8hd_decap_12
Xmux_right_track_2.tap_buf4_0_.scs8hd_inv_1 mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ _207_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB _098_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_5_.scs8hd_inv_1 bottom_left_grid_pin_1_ mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_100 vgnd vpwr scs8hd_fill_1
XPHY_8 vgnd vpwr scs8hd_decap_3
XANTENNA__117__C _169_/C vgnd vpwr scs8hd_diode_2
XFILLER_15_199 vpwr vgnd scs8hd_fill_2
X_127_ _106_/A _167_/B _169_/C _127_/X vgnd vpwr scs8hd_or3_4
XANTENNA_mem_bottom_track_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__133__B _128_/X vgnd vpwr scs8hd_diode_2
XFILLER_7_79 vgnd vpwr scs8hd_decap_4
XFILLER_7_57 vpwr vgnd scs8hd_fill_2
XFILLER_7_35 vpwr vgnd scs8hd_fill_2
XFILLER_16_3 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _217_/A vgnd vpwr scs8hd_inv_1
Xmux_top_track_16.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[2] mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_114 vpwr vgnd scs8hd_fill_2
XFILLER_29_203 vgnd vpwr scs8hd_fill_1
XFILLER_29_258 vgnd vpwr scs8hd_decap_4
XFILLER_16_88 vpwr vgnd scs8hd_fill_2
XFILLER_16_44 vgnd vpwr scs8hd_decap_12
XFILLER_12_169 vpwr vgnd scs8hd_fill_2
XFILLER_12_125 vgnd vpwr scs8hd_decap_8
XFILLER_8_107 vgnd vpwr scs8hd_decap_4
XFILLER_32_32 vgnd vpwr scs8hd_decap_12
XFILLER_8_129 vgnd vpwr scs8hd_decap_8
XANTENNA__144__A _113_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_191 vgnd vpwr scs8hd_decap_4
XFILLER_7_195 vgnd vpwr scs8hd_decap_3
Xmux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ _174_/Y mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_27_98 vgnd vpwr scs8hd_decap_12
XFILLER_4_198 vpwr vgnd scs8hd_fill_2
XFILLER_4_165 vpwr vgnd scs8hd_fill_2
XANTENNA__139__A _085_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_231 vpwr vgnd scs8hd_fill_2
XFILLER_16_272 vgnd vpwr scs8hd_decap_3
XFILLER_31_275 vpwr vgnd scs8hd_fill_2
XFILLER_14_209 vgnd vpwr scs8hd_decap_3
Xmux_top_track_0.INVTX1_2_.scs8hd_inv_1 top_left_grid_pin_13_ mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_14.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_9_235 vpwr vgnd scs8hd_fill_2
XFILLER_9_224 vpwr vgnd scs8hd_fill_2
XANTENNA__141__B _138_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_39_194 vpwr vgnd scs8hd_fill_2
X_091_ _090_/X _110_/A vgnd vpwr scs8hd_buf_1
X_160_ _160_/A _163_/A vgnd vpwr scs8hd_buf_1
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
XFILLER_24_44 vgnd vpwr scs8hd_decap_12
XANTENNA__152__A _098_/B vgnd vpwr scs8hd_diode_2
XFILLER_10_79 vpwr vgnd scs8hd_fill_2
XFILLER_27_142 vpwr vgnd scs8hd_fill_2
X_212_ chany_top_in[4] chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_bottom_track_1.LATCH_5_.latch_SLEEPB _129_/Y vgnd vpwr scs8hd_diode_2
XFILLER_35_98 vgnd vpwr scs8hd_decap_12
XFILLER_42_156 vgnd vpwr scs8hd_decap_12
XFILLER_27_197 vpwr vgnd scs8hd_fill_2
XFILLER_27_175 vpwr vgnd scs8hd_fill_2
X_143_ _098_/B _138_/X _143_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_274 vgnd vpwr scs8hd_fill_1
XFILLER_2_241 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_33_123 vgnd vpwr scs8hd_decap_12
XANTENNA__147__A _146_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_145 vgnd vpwr scs8hd_decap_4
XFILLER_24_123 vpwr vgnd scs8hd_fill_2
Xmux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ _180_/Y mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_15_101 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_126_ _125_/Y _167_/B vgnd vpwr scs8hd_buf_1
Xmux_top_track_8.INVTX1_7_.scs8hd_inv_1 chany_bottom_in[5] mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_7_47 vgnd vpwr scs8hd_decap_3
Xmux_right_track_10.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[8] mux_right_track_10.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A top_left_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_38_215 vgnd vpwr scs8hd_decap_12
XFILLER_38_259 vgnd vpwr scs8hd_decap_12
XFILLER_21_137 vgnd vpwr scs8hd_decap_4
XFILLER_29_215 vpwr vgnd scs8hd_fill_2
XFILLER_32_44 vgnd vpwr scs8hd_decap_12
XFILLER_16_67 vgnd vpwr scs8hd_decap_8
XFILLER_16_56 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_170 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _186_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA__144__B _138_/X vgnd vpwr scs8hd_diode_2
XFILLER_11_181 vpwr vgnd scs8hd_fill_2
XFILLER_7_174 vpwr vgnd scs8hd_fill_2
X_109_ _109_/A _110_/B _109_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__160__A _160_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_207 vgnd vpwr scs8hd_decap_4
XFILLER_19_270 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_240 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
XFILLER_40_243 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_177 vgnd vpwr scs8hd_decap_6
XFILLER_4_122 vpwr vgnd scs8hd_fill_2
XFILLER_4_15 vgnd vpwr scs8hd_decap_12
XANTENNA__155__A _155_/A vgnd vpwr scs8hd_diode_2
XANTENNA__139__B _138_/X vgnd vpwr scs8hd_diode_2
XFILLER_31_243 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1_A bottom_left_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_22_243 vpwr vgnd scs8hd_fill_2
XFILLER_13_57 vpwr vgnd scs8hd_fill_2
XFILLER_13_46 vgnd vpwr scs8hd_decap_4
XFILLER_1_158 vpwr vgnd scs8hd_fill_2
XFILLER_1_114 vgnd vpwr scs8hd_decap_3
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XFILLER_13_221 vpwr vgnd scs8hd_fill_2
XFILLER_13_210 vgnd vpwr scs8hd_decap_4
XFILLER_9_203 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_91 vpwr vgnd scs8hd_fill_2
XFILLER_39_184 vpwr vgnd scs8hd_fill_2
XFILLER_24_56 vgnd vpwr scs8hd_decap_12
X_090_ _090_/A address[2] _156_/A _090_/X vgnd vpwr scs8hd_or3_4
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
XFILLER_10_202 vpwr vgnd scs8hd_fill_2
XFILLER_6_239 vpwr vgnd scs8hd_fill_2
XFILLER_6_206 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _182_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_track_14.LATCH_0_.latch_SLEEPB _172_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__152__B _149_/B vgnd vpwr scs8hd_diode_2
Xmem_right_track_2.LATCH_0_.latch data_in _174_/A _159_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_36_154 vgnd vpwr scs8hd_decap_12
XFILLER_27_110 vgnd vpwr scs8hd_decap_8
X_142_ _095_/B _138_/X _142_/Y vgnd vpwr scs8hd_nor2_4
X_211_ chany_top_in[5] chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_42_168 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1_A bottom_left_grid_pin_15_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_2_231 vgnd vpwr scs8hd_fill_1
XFILLER_33_135 vgnd vpwr scs8hd_decap_12
XFILLER_18_165 vgnd vpwr scs8hd_decap_8
XFILLER_18_121 vpwr vgnd scs8hd_fill_2
XANTENNA__163__A _163_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_168 vpwr vgnd scs8hd_fill_2
XFILLER_15_157 vpwr vgnd scs8hd_fill_2
X_125_ address[6] _125_/Y vgnd vpwr scs8hd_inv_8
XFILLER_30_105 vgnd vpwr scs8hd_decap_12
XFILLER_15_179 vpwr vgnd scs8hd_fill_2
XFILLER_7_15 vgnd vpwr scs8hd_decap_12
XFILLER_38_227 vgnd vpwr scs8hd_decap_12
XANTENNA__158__A address[0] vgnd vpwr scs8hd_diode_2
Xmem_top_track_0.LATCH_2_.latch data_in mem_top_track_0.LATCH_2_.latch/Q _095_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_56 vgnd vpwr scs8hd_decap_12
XFILLER_20_182 vgnd vpwr scs8hd_fill_1
XFILLER_35_208 vgnd vpwr scs8hd_decap_12
XFILLER_28_271 vgnd vpwr scs8hd_decap_4
X_108_ _085_/A _110_/B _108_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_160 vpwr vgnd scs8hd_fill_2
XFILLER_7_142 vpwr vgnd scs8hd_fill_2
XFILLER_7_120 vpwr vgnd scs8hd_fill_2
XFILLER_21_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_12.LATCH_1_.latch_SLEEPB _167_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_230 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _177_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_34_274 vgnd vpwr scs8hd_fill_1
Xmux_top_track_8.tap_buf4_0_.scs8hd_inv_1 mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _222_/A vgnd vpwr scs8hd_inv_1
XFILLER_17_208 vgnd vpwr scs8hd_decap_3
XFILLER_25_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _191_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_145 vgnd vpwr scs8hd_fill_1
XFILLER_4_27 vgnd vpwr scs8hd_decap_4
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_200 vgnd vpwr scs8hd_decap_3
XANTENNA__171__A _157_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_3_.scs8hd_inv_1 chanx_right_in[5] mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__081__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_44 vgnd vpwr scs8hd_decap_12
XFILLER_13_266 vgnd vpwr scs8hd_decap_8
XANTENNA__166__A _163_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_130 vgnd vpwr scs8hd_decap_12
XANTENNA__076__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_24_68 vgnd vpwr scs8hd_decap_4
XFILLER_40_56 vgnd vpwr scs8hd_decap_12
XFILLER_6_229 vgnd vpwr scs8hd_decap_3
XFILLER_1_17 vgnd vpwr scs8hd_decap_3
Xmem_bottom_track_1.LATCH_4_.latch data_in mem_bottom_track_1.LATCH_4_.latch/Q _130_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_240 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_4.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_36_166 vgnd vpwr scs8hd_decap_12
XFILLER_10_15 vgnd vpwr scs8hd_decap_12
XFILLER_42_125 vgnd vpwr scs8hd_decap_12
X_141_ _110_/A _138_/X _141_/Y vgnd vpwr scs8hd_nor2_4
X_210_ chany_top_in[6] chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
Xmux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_top_track_8.LATCH_3_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_147 vgnd vpwr scs8hd_decap_12
XANTENNA__163__B _155_/X vgnd vpwr scs8hd_diode_2
Xmem_right_track_14.LATCH_1_.latch data_in _185_/A _171_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _183_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_103 vgnd vpwr scs8hd_decap_3
XFILLER_2_71 vpwr vgnd scs8hd_fill_2
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_117 vgnd vpwr scs8hd_decap_12
XFILLER_15_114 vpwr vgnd scs8hd_fill_2
X_124_ _113_/A _119_/B _124_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_10.INVTX1_0_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_27 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_91 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_track_17.LATCH_5_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_38_239 vgnd vpwr scs8hd_decap_12
XANTENNA__174__A _174_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_106 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_106 vpwr vgnd scs8hd_fill_2
XANTENNA__084__A _084_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_68 vgnd vpwr scs8hd_decap_12
XFILLER_20_194 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_2_.latch_SLEEPB _111_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_150 vgnd vpwr scs8hd_fill_1
X_107_ _106_/X _110_/B vgnd vpwr scs8hd_buf_1
XFILLER_7_187 vpwr vgnd scs8hd_fill_2
XFILLER_7_132 vgnd vpwr scs8hd_decap_4
XFILLER_14_3 vgnd vpwr scs8hd_decap_12
XANTENNA__169__A _160_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_242 vgnd vpwr scs8hd_decap_12
XANTENNA__079__A address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_25_275 vpwr vgnd scs8hd_fill_2
XFILLER_4_39 vgnd vpwr scs8hd_decap_8
XFILLER_16_253 vpwr vgnd scs8hd_fill_2
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_245 vpwr vgnd scs8hd_fill_2
XANTENNA__171__B _167_/B vgnd vpwr scs8hd_diode_2
XFILLER_22_267 vgnd vpwr scs8hd_decap_8
XFILLER_22_256 vgnd vpwr scs8hd_decap_8
XFILLER_22_212 vpwr vgnd scs8hd_fill_2
XFILLER_13_15 vgnd vpwr scs8hd_decap_12
XANTENNA__081__B address[4] vgnd vpwr scs8hd_diode_2
XFILLER_1_138 vgnd vpwr scs8hd_decap_4
XFILLER_38_56 vgnd vpwr scs8hd_decap_12
XFILLER_13_245 vpwr vgnd scs8hd_fill_2
XFILLER_0_182 vpwr vgnd scs8hd_fill_2
XANTENNA__166__B _155_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr
+ scs8hd_diode_2
XANTENNA__182__A _182_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_142 vgnd vpwr scs8hd_decap_12
XFILLER_39_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_248 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA__092__A _085_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_10.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__177__A _177_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_178 vgnd vpwr scs8hd_decap_12
XFILLER_10_27 vgnd vpwr scs8hd_decap_4
XANTENNA__087__A _086_/X vgnd vpwr scs8hd_diode_2
XFILLER_42_137 vgnd vpwr scs8hd_decap_12
XFILLER_27_123 vgnd vpwr scs8hd_decap_4
X_140_ _109_/A _138_/X _140_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_2_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_top_track_16.LATCH_4_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_18_101 vgnd vpwr scs8hd_fill_1
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_159 vgnd vpwr scs8hd_decap_12
XFILLER_18_189 vpwr vgnd scs8hd_fill_2
XANTENNA__163__C _163_/C vgnd vpwr scs8hd_diode_2
XFILLER_2_50 vpwr vgnd scs8hd_fill_2
XFILLER_24_115 vgnd vpwr scs8hd_decap_8
XFILLER_21_15 vgnd vpwr scs8hd_decap_12
XFILLER_21_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.INVTX1_3_.scs8hd_inv_1 chanx_right_in[0] mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_30_129 vgnd vpwr scs8hd_decap_12
X_123_ _098_/B _119_/B _123_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_21_118 vpwr vgnd scs8hd_fill_2
Xmem_top_track_8.LATCH_3_.latch data_in mem_top_track_8.LATCH_3_.latch/Q _110_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_37_262 vpwr vgnd scs8hd_fill_2
XFILLER_16_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_140 vpwr vgnd scs8hd_fill_2
XFILLER_28_251 vgnd vpwr scs8hd_decap_4
XFILLER_11_173 vpwr vgnd scs8hd_fill_2
X_106_ _106_/A _155_/A _163_/C _106_/X vgnd vpwr scs8hd_or3_4
XFILLER_22_80 vgnd vpwr scs8hd_fill_1
XFILLER_7_155 vpwr vgnd scs8hd_fill_2
XANTENNA__169__B _155_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_240 vpwr vgnd scs8hd_fill_2
XANTENNA__185__A _185_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_254 vgnd vpwr scs8hd_decap_12
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XFILLER_8_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__095__A _085_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_169 vpwr vgnd scs8hd_fill_2
XFILLER_4_103 vpwr vgnd scs8hd_fill_2
XFILLER_31_235 vgnd vpwr scs8hd_decap_8
XFILLER_17_91 vpwr vgnd scs8hd_fill_2
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XFILLER_16_232 vpwr vgnd scs8hd_fill_2
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__171__C _163_/C vgnd vpwr scs8hd_diode_2
XFILLER_13_27 vgnd vpwr scs8hd_decap_12
XANTENNA__081__C _081_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_68 vgnd vpwr scs8hd_decap_12
XFILLER_9_239 vgnd vpwr scs8hd_decap_3
XFILLER_0_150 vgnd vpwr scs8hd_decap_3
Xmux_right_track_8.INVTX1_0_.scs8hd_inv_1 chany_top_in[4] mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__166__C _136_/X vgnd vpwr scs8hd_diode_2
XFILLER_39_110 vpwr vgnd scs8hd_fill_2
XFILLER_5_72 vpwr vgnd scs8hd_fill_2
XFILLER_39_154 vgnd vpwr scs8hd_decap_12
XFILLER_39_198 vgnd vpwr scs8hd_decap_4
XFILLER_24_15 vgnd vpwr scs8hd_decap_12
XANTENNA__092__B _110_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_6 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_2_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_17.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_9.LATCH_5_.latch data_in mem_bottom_track_9.LATCH_5_.latch/Q _139_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_30_80 vgnd vpwr scs8hd_decap_12
XFILLER_39_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_2_.latch_SLEEPB _132_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_15 vgnd vpwr scs8hd_decap_12
XFILLER_42_149 vgnd vpwr scs8hd_decap_6
XFILLER_27_179 vpwr vgnd scs8hd_fill_2
XFILLER_27_146 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _185_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_4_3 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.INVTX1_5_.scs8hd_inv_1 bottom_right_grid_pin_11_ mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_track_8.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_113 vgnd vpwr scs8hd_decap_8
XPHY_80 vgnd vpwr scs8hd_decap_3
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_171 vgnd vpwr scs8hd_decap_12
X_199_ _199_/HI _199_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__163__D _163_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _192_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_84 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_track_9.LATCH_4_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_8.INVTX1_4_.scs8hd_inv_1 chanx_right_in[5] mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_32_193 vgnd vpwr scs8hd_fill_1
XFILLER_21_27 vgnd vpwr scs8hd_decap_12
XANTENNA__098__A _085_/B vgnd vpwr scs8hd_diode_2
XFILLER_15_105 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_193 vgnd vpwr scs8hd_decap_3
XFILLER_15_138 vpwr vgnd scs8hd_fill_2
X_122_ _095_/B _119_/B _122_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_60 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB _120_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_5_.latch data_in mem_top_track_16.LATCH_5_.latch/Q _119_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_219 vpwr vgnd scs8hd_fill_2
XFILLER_37_274 vgnd vpwr scs8hd_decap_3
Xmem_right_track_10.LATCH_1_.latch data_in _179_/A _165_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_15 vgnd vpwr scs8hd_decap_12
XFILLER_16_27 vgnd vpwr scs8hd_decap_4
XFILLER_12_119 vgnd vpwr scs8hd_decap_4
XFILLER_20_174 vgnd vpwr scs8hd_decap_8
XFILLER_28_230 vgnd vpwr scs8hd_decap_8
X_105_ _104_/X _163_/C vgnd vpwr scs8hd_buf_1
XFILLER_7_112 vpwr vgnd scs8hd_fill_2
XFILLER_7_178 vpwr vgnd scs8hd_fill_2
XANTENNA__169__C _169_/C vgnd vpwr scs8hd_diode_2
XFILLER_34_266 vgnd vpwr scs8hd_decap_8
XFILLER_8_72 vgnd vpwr scs8hd_fill_1
XFILLER_27_59 vpwr vgnd scs8hd_fill_2
XFILLER_27_15 vgnd vpwr scs8hd_decap_12
XANTENNA__095__B _095_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_148 vgnd vpwr scs8hd_decap_4
XFILLER_4_126 vpwr vgnd scs8hd_fill_2
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_214 vpwr vgnd scs8hd_fill_2
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__171__D _156_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_236 vpwr vgnd scs8hd_fill_2
XFILLER_13_214 vgnd vpwr scs8hd_fill_1
XFILLER_9_207 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_3_.latch_SLEEPB _150_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_80 vgnd vpwr scs8hd_decap_12
XFILLER_0_173 vgnd vpwr scs8hd_fill_1
XANTENNA__166__D _162_/D vgnd vpwr scs8hd_diode_2
XFILLER_8_262 vgnd vpwr scs8hd_decap_12
XFILLER_8_251 vpwr vgnd scs8hd_fill_2
XFILLER_5_62 vgnd vpwr scs8hd_fill_1
XFILLER_39_166 vgnd vpwr scs8hd_decap_4
XFILLER_5_95 vpwr vgnd scs8hd_fill_2
XFILLER_24_27 vgnd vpwr scs8hd_decap_4
XFILLER_40_15 vgnd vpwr scs8hd_decap_12
XFILLER_10_206 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _184_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_93 vpwr vgnd scs8hd_fill_2
XFILLER_5_265 vpwr vgnd scs8hd_fill_2
XFILLER_5_254 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_2_.latch/Q mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_bottom_track_17.LATCH_5_.latch data_in mem_bottom_track_17.LATCH_5_.latch/Q _148_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_6.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
XFILLER_27_158 vpwr vgnd scs8hd_fill_2
XFILLER_19_27 vgnd vpwr scs8hd_decap_12
XFILLER_35_59 vpwr vgnd scs8hd_fill_2
XFILLER_42_106 vgnd vpwr scs8hd_decap_12
XFILLER_2_202 vpwr vgnd scs8hd_fill_2
XFILLER_2_224 vgnd vpwr scs8hd_decap_4
XFILLER_18_125 vgnd vpwr scs8hd_decap_4
XPHY_70 vgnd vpwr scs8hd_decap_3
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _187_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_25_70 vpwr vgnd scs8hd_fill_2
X_198_ _198_/HI _198_/LO vgnd vpwr scs8hd_conb_1
Xmux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_128 vpwr vgnd scs8hd_fill_2
Xmem_right_track_6.LATCH_1_.latch data_in _177_/A _163_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_track_0.INVTX1_7_.scs8hd_inv_1 chany_bottom_in[4] mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_39 vgnd vpwr scs8hd_decap_12
XANTENNA__098__B _098_/B vgnd vpwr scs8hd_diode_2
X_121_ _110_/A _119_/B _121_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_72 vpwr vgnd scs8hd_fill_2
XFILLER_36_80 vgnd vpwr scs8hd_decap_12
XFILLER_14_150 vgnd vpwr scs8hd_decap_3
XFILLER_37_220 vgnd vpwr scs8hd_decap_12
XFILLER_37_253 vpwr vgnd scs8hd_fill_2
XFILLER_32_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _178_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB _169_/Y vgnd vpwr scs8hd_diode_2
X_104_ _103_/Y address[4] _081_/C _104_/X vgnd vpwr scs8hd_or3_4
XFILLER_11_142 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__169__D _163_/D vgnd vpwr scs8hd_diode_2
XFILLER_8_84 vpwr vgnd scs8hd_fill_2
XFILLER_27_27 vgnd vpwr scs8hd_decap_12
XFILLER_40_215 vgnd vpwr scs8hd_decap_12
XFILLER_25_245 vgnd vpwr scs8hd_decap_3
XFILLER_25_223 vpwr vgnd scs8hd_fill_2
XFILLER_40_259 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_259 vpwr vgnd scs8hd_fill_2
XFILLER_12_3 vgnd vpwr scs8hd_decap_12
XFILLER_3_193 vpwr vgnd scs8hd_fill_2
XFILLER_22_215 vpwr vgnd scs8hd_fill_2
XFILLER_22_204 vpwr vgnd scs8hd_fill_2
XFILLER_1_119 vgnd vpwr scs8hd_decap_3
XFILLER_38_15 vgnd vpwr scs8hd_decap_12
XFILLER_0_196 vpwr vgnd scs8hd_fill_2
XFILLER_8_274 vgnd vpwr scs8hd_fill_1
XFILLER_40_27 vgnd vpwr scs8hd_decap_4
XFILLER_10_229 vpwr vgnd scs8hd_fill_2
XFILLER_10_218 vpwr vgnd scs8hd_fill_2
XFILLER_30_93 vgnd vpwr scs8hd_decap_12
XFILLER_5_222 vgnd vpwr scs8hd_decap_3
XFILLER_35_27 vgnd vpwr scs8hd_decap_12
XFILLER_42_118 vgnd vpwr scs8hd_decap_6
XFILLER_19_39 vgnd vpwr scs8hd_decap_12
XFILLER_2_247 vpwr vgnd scs8hd_fill_2
Xmux_right_track_14.tap_buf4_0_.scs8hd_inv_1 mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ _201_/A vgnd vpwr scs8hd_inv_1
XFILLER_2_258 vgnd vpwr scs8hd_decap_12
XPHY_60 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_82 vgnd vpwr scs8hd_decap_3
XFILLER_18_148 vgnd vpwr scs8hd_decap_3
X_197_ _197_/HI _197_/LO vgnd vpwr scs8hd_conb_1
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_184 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.tap_buf4_0_.scs8hd_inv_1 mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _218_/A vgnd vpwr scs8hd_inv_1
XFILLER_17_170 vpwr vgnd scs8hd_fill_2
XFILLER_15_118 vpwr vgnd scs8hd_fill_2
X_120_ _109_/A _119_/B _120_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_162 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_95 vpwr vgnd scs8hd_fill_2
XFILLER_11_62 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_184 vpwr vgnd scs8hd_fill_2
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_37_232 vgnd vpwr scs8hd_decap_12
XFILLER_20_154 vgnd vpwr scs8hd_decap_3
XFILLER_20_132 vpwr vgnd scs8hd_fill_2
XFILLER_20_121 vpwr vgnd scs8hd_fill_2
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
X_103_ address[3] _103_/Y vgnd vpwr scs8hd_inv_8
XFILLER_11_187 vpwr vgnd scs8hd_fill_2
XFILLER_34_202 vgnd vpwr scs8hd_decap_12
XFILLER_19_276 vgnd vpwr scs8hd_fill_1
XFILLER_27_39 vgnd vpwr scs8hd_decap_12
XFILLER_40_227 vgnd vpwr scs8hd_decap_12
XFILLER_4_139 vgnd vpwr scs8hd_decap_6
XFILLER_17_72 vpwr vgnd scs8hd_fill_2
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_249 vgnd vpwr scs8hd_decap_6
XFILLER_3_161 vpwr vgnd scs8hd_fill_2
XFILLER_38_27 vgnd vpwr scs8hd_decap_4
XFILLER_13_249 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_12.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_120 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_93 vgnd vpwr scs8hd_decap_12
XFILLER_5_53 vpwr vgnd scs8hd_fill_2
XFILLER_5_42 vpwr vgnd scs8hd_fill_2
XFILLER_39_179 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_190 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.tap_buf4_0_.scs8hd_inv_1 mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _204_/A vgnd vpwr scs8hd_inv_1
XFILLER_14_84 vgnd vpwr scs8hd_decap_6
XFILLER_5_201 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_2_.latch/Q mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__101__A _085_/B vgnd vpwr scs8hd_diode_2
XFILLER_36_105 vgnd vpwr scs8hd_decap_12
XFILLER_39_70 vpwr vgnd scs8hd_fill_2
XFILLER_39_81 vpwr vgnd scs8hd_fill_2
XFILLER_35_39 vgnd vpwr scs8hd_decap_12
XFILLER_35_171 vgnd vpwr scs8hd_decap_12
XFILLER_27_138 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_25_83 vpwr vgnd scs8hd_fill_2
X_196_ _196_/HI _196_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_41_196 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_5_ mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_32 vgnd vpwr scs8hd_decap_4
XFILLER_17_182 vgnd vpwr scs8hd_fill_1
XFILLER_2_54 vpwr vgnd scs8hd_fill_2
XFILLER_32_141 vgnd vpwr scs8hd_decap_12
XFILLER_17_193 vgnd vpwr scs8hd_decap_4
XFILLER_23_141 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _187_/HI mem_bottom_track_1.LATCH_2_.latch/Q
+ mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_9.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_3_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_93 vgnd vpwr scs8hd_decap_12
XFILLER_14_130 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_179_ _179_/A _179_/Y vgnd vpwr scs8hd_inv_8
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_266 vgnd vpwr scs8hd_decap_8
XFILLER_20_199 vgnd vpwr scs8hd_decap_3
XFILLER_20_166 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_2.LATCH_1_.latch data_in _173_/A _157_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_7_104 vpwr vgnd scs8hd_fill_2
X_102_ address[6] _155_/A vgnd vpwr scs8hd_buf_1
XFILLER_22_84 vgnd vpwr scs8hd_decap_8
XFILLER_22_73 vgnd vpwr scs8hd_fill_1
XFILLER_11_177 vpwr vgnd scs8hd_fill_2
XFILLER_7_159 vpwr vgnd scs8hd_fill_2
XFILLER_19_266 vpwr vgnd scs8hd_fill_2
XFILLER_19_255 vpwr vgnd scs8hd_fill_2
Xmux_right_track_2.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_97 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_206 vgnd vpwr scs8hd_decap_8
XFILLER_25_236 vpwr vgnd scs8hd_fill_2
XFILLER_4_107 vpwr vgnd scs8hd_fill_2
XFILLER_17_95 vpwr vgnd scs8hd_fill_2
XFILLER_17_62 vgnd vpwr scs8hd_decap_8
XFILLER_17_51 vgnd vpwr scs8hd_decap_8
XFILLER_16_236 vpwr vgnd scs8hd_fill_2
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__104__A _103_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_239 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_217 vpwr vgnd scs8hd_fill_2
XFILLER_0_165 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_top_track_0.LATCH_3_.latch data_in mem_top_track_0.LATCH_3_.latch/Q _092_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_272 vgnd vpwr scs8hd_decap_3
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
XFILLER_8_232 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_9.LATCH_0_.latch data_in mem_bottom_track_9.LATCH_0_.latch/Q _144_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_39_114 vgnd vpwr scs8hd_decap_8
XFILLER_5_76 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_52 vgnd vpwr scs8hd_fill_1
XFILLER_39_60 vgnd vpwr scs8hd_fill_1
XANTENNA__101__B _113_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_117 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.INVTX1_2_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_6.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__202__A _202_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_1_.scs8hd_inv_1 top_left_grid_pin_9_ mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_40 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_26_150 vgnd vpwr scs8hd_decap_3
XFILLER_25_62 vpwr vgnd scs8hd_fill_2
XFILLER_25_51 vgnd vpwr scs8hd_decap_8
X_195_ _195_/HI _195_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__112__A _098_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_88 vpwr vgnd scs8hd_fill_2
XFILLER_32_197 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB _123_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_0_.latch data_in mem_top_track_16.LATCH_0_.latch/Q _124_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_175 vpwr vgnd scs8hd_fill_2
XFILLER_11_53 vgnd vpwr scs8hd_decap_4
XANTENNA__107__A _106_/X vgnd vpwr scs8hd_diode_2
X_178_ _178_/A _178_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_245 vgnd vpwr scs8hd_decap_8
XFILLER_28_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_5_.latch data_in mem_bottom_track_1.LATCH_5_.latch/Q _129_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_145 vpwr vgnd scs8hd_fill_2
XFILLER_9_190 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_201 vpwr vgnd scs8hd_fill_2
X_101_ _085_/B _113_/A _101_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_156 vpwr vgnd scs8hd_fill_2
XFILLER_11_123 vgnd vpwr scs8hd_decap_4
XFILLER_7_138 vpwr vgnd scs8hd_fill_2
XFILLER_7_116 vpwr vgnd scs8hd_fill_2
XFILLER_22_96 vpwr vgnd scs8hd_fill_2
XFILLER_19_245 vgnd vpwr scs8hd_fill_1
XFILLER_19_223 vpwr vgnd scs8hd_fill_2
XFILLER_8_65 vgnd vpwr scs8hd_decap_4
XFILLER_8_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_182 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_215 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB _092_/Y vgnd vpwr scs8hd_diode_2
XFILLER_25_259 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.INVTX1_7_.scs8hd_inv_1 bottom_left_grid_pin_13_ mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__210__A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _183_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_31_218 vpwr vgnd scs8hd_fill_2
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_51 vgnd vpwr scs8hd_decap_8
XFILLER_33_62 vgnd vpwr scs8hd_decap_12
XANTENNA__104__B address[4] vgnd vpwr scs8hd_diode_2
XFILLER_3_174 vpwr vgnd scs8hd_fill_2
XANTENNA__120__A _109_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB _153_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_273 vgnd vpwr scs8hd_decap_4
XANTENNA__205__A _205_/A vgnd vpwr scs8hd_diode_2
XANTENNA__115__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_8_255 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_126 vpwr vgnd scs8hd_fill_2
XFILLER_10_3 vgnd vpwr scs8hd_decap_12
XFILLER_5_99 vgnd vpwr scs8hd_decap_4
Xmem_bottom_track_17.LATCH_0_.latch data_in mem_bottom_track_17.LATCH_0_.latch/Q _153_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_top_track_8.LATCH_4_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_14_97 vgnd vpwr scs8hd_fill_1
XFILLER_5_269 vgnd vpwr scs8hd_decap_8
XFILLER_5_258 vpwr vgnd scs8hd_fill_2
XFILLER_5_236 vpwr vgnd scs8hd_fill_2
XFILLER_36_129 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_3_ vgnd vpwr scs8hd_diode_2
XFILLER_27_118 vpwr vgnd scs8hd_fill_2
XFILLER_35_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_228 vgnd vpwr scs8hd_fill_1
XFILLER_2_206 vgnd vpwr scs8hd_decap_8
Xmux_top_track_0.INVTX1_4_.scs8hd_inv_1 chanx_right_in[4] mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_41 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_10.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr
+ scs8hd_diode_2
XFILLER_41_110 vgnd vpwr scs8hd_decap_12
XFILLER_26_184 vpwr vgnd scs8hd_fill_2
X_194_ _194_/HI _194_/LO vgnd vpwr scs8hd_conb_1
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
XANTENNA__112__B _110_/B vgnd vpwr scs8hd_diode_2
XFILLER_2_67 vpwr vgnd scs8hd_fill_2
XFILLER_2_23 vgnd vpwr scs8hd_decap_8
XFILLER_32_154 vgnd vpwr scs8hd_decap_8
XFILLER_32_165 vgnd vpwr scs8hd_decap_12
XFILLER_17_140 vgnd vpwr scs8hd_decap_4
XFILLER_23_198 vpwr vgnd scs8hd_fill_2
XFILLER_23_110 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_11_76 vpwr vgnd scs8hd_fill_2
XANTENNA__213__A _213_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_154 vpwr vgnd scs8hd_fill_2
XFILLER_14_143 vgnd vpwr scs8hd_decap_4
X_177_ _177_/A _177_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__123__A _098_/B vgnd vpwr scs8hd_diode_2
XFILLER_20_113 vgnd vpwr scs8hd_decap_8
XFILLER_20_102 vgnd vpwr scs8hd_decap_3
XFILLER_9_180 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1_A bottom_left_grid_pin_1_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_28_213 vgnd vpwr scs8hd_fill_1
X_100_ _099_/X _113_/A vgnd vpwr scs8hd_buf_1
XANTENNA__208__A right_top_grid_pin_10_ vgnd vpwr scs8hd_diode_2
XFILLER_22_64 vgnd vpwr scs8hd_decap_3
XFILLER_11_146 vgnd vpwr scs8hd_decap_4
XANTENNA__118__A _117_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_88 vgnd vpwr scs8hd_decap_4
XFILLER_8_44 vgnd vpwr scs8hd_fill_1
XFILLER_40_3 vgnd vpwr scs8hd_decap_12
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_249 vpwr vgnd scs8hd_fill_2
XFILLER_33_74 vgnd vpwr scs8hd_decap_12
XANTENNA__104__C _081_/C vgnd vpwr scs8hd_diode_2
XFILLER_3_197 vgnd vpwr scs8hd_decap_4
XFILLER_3_142 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA__120__B _119_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_274 vgnd vpwr scs8hd_fill_1
XFILLER_22_219 vgnd vpwr scs8hd_decap_3
XFILLER_22_208 vpwr vgnd scs8hd_fill_2
XFILLER_15_260 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.INVTX1_1_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_2_.latch/Q mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__221__A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_0_178 vpwr vgnd scs8hd_fill_2
XFILLER_0_134 vpwr vgnd scs8hd_fill_2
Xmem_top_track_8.LATCH_4_.latch data_in mem_top_track_8.LATCH_4_.latch/Q _109_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__115__B _115_/B vgnd vpwr scs8hd_diode_2
XANTENNA__131__A _110_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_105 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_32 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ mem_top_track_16.LATCH_5_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA__216__A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_39_62 vgnd vpwr scs8hd_decap_4
XFILLER_29_193 vgnd vpwr scs8hd_decap_4
XANTENNA__126__A _125_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XPHY_64 vgnd vpwr scs8hd_decap_3
X_193_ _193_/HI _193_/LO vgnd vpwr scs8hd_conb_1
XPHY_75 vgnd vpwr scs8hd_decap_3
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_74 vgnd vpwr scs8hd_decap_12
XFILLER_1_251 vpwr vgnd scs8hd_fill_2
XFILLER_1_240 vpwr vgnd scs8hd_fill_2
XFILLER_32_177 vgnd vpwr scs8hd_decap_12
XFILLER_17_174 vpwr vgnd scs8hd_fill_2
XFILLER_17_163 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_99 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_track_1.LATCH_3_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_188 vgnd vpwr scs8hd_decap_4
X_176_ _176_/A _176_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__123__B _119_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_258 vpwr vgnd scs8hd_fill_2
XFILLER_20_136 vpwr vgnd scs8hd_fill_2
XFILLER_28_247 vpwr vgnd scs8hd_fill_2
XFILLER_11_114 vpwr vgnd scs8hd_fill_2
XANTENNA__224__A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_4.LATCH_0_.latch_SLEEPB _162_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_76 vpwr vgnd scs8hd_fill_2
XFILLER_22_32 vgnd vpwr scs8hd_decap_12
XFILLER_0_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_236 vpwr vgnd scs8hd_fill_2
XFILLER_19_214 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_261 vgnd vpwr scs8hd_decap_12
X_159_ _157_/A _155_/X _136_/X _162_/D _159_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__134__A _113_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_162 vgnd vpwr scs8hd_decap_4
XFILLER_33_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_206 vgnd vpwr scs8hd_decap_6
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__219__A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_33_86 vgnd vpwr scs8hd_decap_12
XFILLER_17_76 vpwr vgnd scs8hd_fill_2
XFILLER_3_132 vpwr vgnd scs8hd_fill_2
XANTENNA__129__A _085_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_231 vpwr vgnd scs8hd_fill_2
XFILLER_21_220 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_146 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_264 vgnd vpwr scs8hd_decap_8
XFILLER_12_253 vpwr vgnd scs8hd_fill_2
XFILLER_8_213 vgnd vpwr scs8hd_fill_1
XANTENNA__131__B _128_/X vgnd vpwr scs8hd_diode_2
XANTENNA__115__C _081_/C vgnd vpwr scs8hd_diode_2
XFILLER_5_57 vpwr vgnd scs8hd_fill_2
XFILLER_5_46 vpwr vgnd scs8hd_fill_2
XFILLER_14_44 vgnd vpwr scs8hd_decap_8
XFILLER_30_32 vgnd vpwr scs8hd_decap_12
XFILLER_5_205 vpwr vgnd scs8hd_fill_2
XFILLER_39_74 vpwr vgnd scs8hd_fill_2
XFILLER_39_85 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_2.LATCH_1_.latch_SLEEPB _157_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__142__A _095_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ mem_bottom_track_9.LATCH_5_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_16.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_5_.scs8hd_inv_1 bottom_left_grid_pin_3_ mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_123 vgnd vpwr scs8hd_decap_12
XFILLER_26_142 vgnd vpwr scs8hd_decap_8
XFILLER_25_87 vpwr vgnd scs8hd_fill_2
X_192_ _192_/HI _192_/LO vgnd vpwr scs8hd_conb_1
XFILLER_41_86 vgnd vpwr scs8hd_decap_12
Xmux_right_track_14.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[3] mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB _144_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__137__A _106_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_189 vgnd vpwr scs8hd_decap_4
XFILLER_23_145 vpwr vgnd scs8hd_fill_2
XFILLER_23_123 vpwr vgnd scs8hd_fill_2
XFILLER_11_45 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_167 vgnd vpwr scs8hd_decap_6
X_175_ _175_/A _175_/Y vgnd vpwr scs8hd_inv_8
XFILLER_28_259 vgnd vpwr scs8hd_decap_12
XFILLER_28_215 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_44 vgnd vpwr scs8hd_decap_12
XFILLER_7_108 vpwr vgnd scs8hd_fill_2
Xmux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_2_.scs8hd_inv_1/Y
+ _178_/A mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_34_218 vgnd vpwr scs8hd_decap_12
XFILLER_19_259 vgnd vpwr scs8hd_decap_4
XFILLER_42_273 vgnd vpwr scs8hd_decap_4
X_089_ address[1] _090_/A vgnd vpwr scs8hd_inv_8
X_158_ address[0] _162_/D vgnd vpwr scs8hd_buf_1
XANTENNA__134__B _128_/X vgnd vpwr scs8hd_diode_2
XFILLER_10_181 vpwr vgnd scs8hd_fill_2
XFILLER_6_185 vpwr vgnd scs8hd_fill_2
XANTENNA__150__A _110_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_98 vgnd vpwr scs8hd_decap_12
XFILLER_24_251 vpwr vgnd scs8hd_fill_2
XANTENNA__129__B _128_/X vgnd vpwr scs8hd_diode_2
XANTENNA__145__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_30_243 vgnd vpwr scs8hd_decap_8
XFILLER_30_254 vgnd vpwr scs8hd_decap_12
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XFILLER_21_265 vpwr vgnd scs8hd_fill_2
XFILLER_21_254 vpwr vgnd scs8hd_fill_2
XFILLER_21_243 vgnd vpwr scs8hd_fill_1
XFILLER_0_103 vpwr vgnd scs8hd_fill_2
XFILLER_28_32 vgnd vpwr scs8hd_decap_12
XFILLER_0_169 vpwr vgnd scs8hd_fill_2
XFILLER_12_210 vpwr vgnd scs8hd_fill_2
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
XFILLER_8_236 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_4_.latch_SLEEPB _109_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_25 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_67 vgnd vpwr scs8hd_decap_6
XFILLER_14_56 vgnd vpwr scs8hd_decap_8
XFILLER_30_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_151 vpwr vgnd scs8hd_fill_2
XFILLER_39_97 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__142__B _138_/X vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _197_/HI mem_top_track_0.LATCH_2_.latch/Q
+ mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_35_110 vgnd vpwr scs8hd_decap_12
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_135 vgnd vpwr scs8hd_decap_12
XFILLER_26_165 vgnd vpwr scs8hd_decap_6
XFILLER_26_154 vpwr vgnd scs8hd_fill_2
XFILLER_25_66 vpwr vgnd scs8hd_fill_2
X_191_ _191_/HI _191_/LO vgnd vpwr scs8hd_conb_1
XFILLER_41_98 vgnd vpwr scs8hd_decap_12
XFILLER_2_15 vgnd vpwr scs8hd_decap_4
XFILLER_1_275 vpwr vgnd scs8hd_fill_2
XFILLER_17_110 vgnd vpwr scs8hd_decap_8
XANTENNA__137__B _167_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_190 vgnd vpwr scs8hd_decap_12
XANTENNA__153__A _113_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_179 vpwr vgnd scs8hd_fill_2
XFILLER_11_57 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_1.LATCH_0_.latch data_in mem_bottom_track_1.LATCH_0_.latch/Q _134_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_36_32 vgnd vpwr scs8hd_decap_12
X_174_ _174_/A _174_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__148__A _085_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_12.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[1] mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_149 vgnd vpwr scs8hd_decap_4
XFILLER_9_172 vpwr vgnd scs8hd_fill_2
XFILLER_9_161 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_205 vpwr vgnd scs8hd_fill_2
XFILLER_3_91 vpwr vgnd scs8hd_fill_2
XFILLER_22_56 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB _101_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_4_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
X_157_ _157_/A _155_/X _136_/X _163_/D _157_/Y vgnd vpwr scs8hd_nor4_4
X_226_ _226_/A chany_top_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_8_69 vgnd vpwr scs8hd_fill_1
X_088_ _085_/B _109_/A _088_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__150__B _149_/B vgnd vpwr scs8hd_diode_2
XFILLER_25_219 vpwr vgnd scs8hd_fill_2
XFILLER_19_3 vgnd vpwr scs8hd_decap_12
XFILLER_33_241 vgnd vpwr scs8hd_decap_3
XFILLER_33_263 vgnd vpwr scs8hd_decap_12
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_263 vgnd vpwr scs8hd_decap_12
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.INVTX1_5_.scs8hd_inv_1 chanx_right_in[6] mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_178 vgnd vpwr scs8hd_decap_3
X_209_ _209_/A chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA__161__A _163_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_266 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_5_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_44 vgnd vpwr scs8hd_decap_12
XFILLER_8_204 vpwr vgnd scs8hd_fill_2
XFILLER_5_37 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_10.tap_buf4_0_.scs8hd_inv_1 mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ _203_/A vgnd vpwr scs8hd_inv_1
XANTENNA__156__A _156_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_141 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_56 vgnd vpwr scs8hd_decap_12
XFILLER_5_218 vpwr vgnd scs8hd_fill_2
XFILLER_39_10 vgnd vpwr scs8hd_decap_4
XFILLER_39_21 vgnd vpwr scs8hd_decap_4
XFILLER_39_32 vgnd vpwr scs8hd_decap_12
XFILLER_29_130 vgnd vpwr scs8hd_decap_12
XFILLER_4_240 vgnd vpwr scs8hd_decap_4
Xmux_top_track_0.INVTX1_1_.scs8hd_inv_1 top_left_grid_pin_7_ mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_12 vgnd vpwr scs8hd_decap_3
X_190_ _190_/HI _190_/LO vgnd vpwr scs8hd_conb_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_147 vgnd vpwr scs8hd_decap_12
XFILLER_26_188 vpwr vgnd scs8hd_fill_2
XFILLER_1_232 vpwr vgnd scs8hd_fill_2
XFILLER_1_221 vpwr vgnd scs8hd_fill_2
XFILLER_17_199 vpwr vgnd scs8hd_fill_2
XANTENNA__137__C _136_/X vgnd vpwr scs8hd_diode_2
XANTENNA__153__B _149_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _174_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_158 vpwr vgnd scs8hd_fill_2
XFILLER_23_114 vgnd vpwr scs8hd_decap_8
XFILLER_36_44 vgnd vpwr scs8hd_decap_12
X_173_ _173_/A _173_/Y vgnd vpwr scs8hd_inv_8
XFILLER_22_180 vpwr vgnd scs8hd_fill_2
XFILLER_14_147 vgnd vpwr scs8hd_fill_1
XANTENNA__148__B _149_/B vgnd vpwr scs8hd_diode_2
XANTENNA__164__A _163_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_4_.latch_SLEEPB _130_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_184 vgnd vpwr scs8hd_decap_4
XFILLER_9_140 vpwr vgnd scs8hd_fill_2
XFILLER_42_242 vgnd vpwr scs8hd_decap_6
XFILLER_27_261 vgnd vpwr scs8hd_decap_4
XFILLER_8_15 vgnd vpwr scs8hd_decap_12
X_087_ _086_/X _109_/A vgnd vpwr scs8hd_buf_1
X_156_ _156_/A _163_/D vgnd vpwr scs8hd_buf_1
X_225_ chany_bottom_in[0] chany_top_out[1] vgnd vpwr scs8hd_buf_2
Xmux_bottom_track_1.INVTX1_7_.scs8hd_inv_1 bottom_left_grid_pin_11_ mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_48 vgnd vpwr scs8hd_decap_8
XFILLER_6_198 vpwr vgnd scs8hd_fill_2
XANTENNA__159__A _157_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_250 vpwr vgnd scs8hd_fill_2
XFILLER_33_253 vpwr vgnd scs8hd_fill_2
XFILLER_33_275 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[1] mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_10.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[2] mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_157 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_264 vgnd vpwr scs8hd_decap_12
XFILLER_15_242 vpwr vgnd scs8hd_fill_2
X_139_ _085_/A _138_/X _139_/Y vgnd vpwr scs8hd_nor2_4
X_208_ right_top_grid_pin_10_ chanx_right_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA__161__B _155_/X vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.tap_buf4_0_.scs8hd_inv_1 mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ _206_/A vgnd vpwr scs8hd_inv_1
XFILLER_31_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_190 vpwr vgnd scs8hd_fill_2
XFILLER_21_245 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_10.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_138 vpwr vgnd scs8hd_fill_2
XFILLER_0_116 vpwr vgnd scs8hd_fill_2
XFILLER_28_56 vgnd vpwr scs8hd_decap_12
XFILLER_12_234 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__172__A _157_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__082__A _081_/X vgnd vpwr scs8hd_diode_2
XFILLER_30_68 vgnd vpwr scs8hd_decap_12
XFILLER_39_44 vgnd vpwr scs8hd_decap_12
XFILLER_39_66 vgnd vpwr scs8hd_fill_1
XFILLER_29_142 vpwr vgnd scs8hd_fill_2
XFILLER_29_164 vpwr vgnd scs8hd_fill_2
XFILLER_29_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__167__A _157_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_123 vgnd vpwr scs8hd_decap_12
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XANTENNA__077__A address[1] vgnd vpwr scs8hd_diode_2
XPHY_57 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_79 vgnd vpwr scs8hd_decap_3
XFILLER_41_159 vgnd vpwr scs8hd_decap_12
XFILLER_9_3 vgnd vpwr scs8hd_decap_12
XFILLER_1_200 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_8.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_2_39 vgnd vpwr scs8hd_decap_8
XFILLER_17_178 vpwr vgnd scs8hd_fill_2
XFILLER_17_123 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_17.LATCH_5_.latch_SLEEPB _148_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_track_0.LATCH_4_.latch data_in mem_top_track_0.LATCH_4_.latch/Q _088_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_31_170 vpwr vgnd scs8hd_fill_2
XFILLER_11_15 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_9.LATCH_1_.latch data_in mem_bottom_track_9.LATCH_1_.latch/Q _143_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _183_/A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_36_56 vgnd vpwr scs8hd_decap_12
XFILLER_14_126 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_172_ _157_/A _167_/B _163_/C address[0] _172_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__164__B _155_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _193_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_107 vgnd vpwr scs8hd_decap_3
XANTENNA__180__A _180_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_251 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[5] mux_right_track_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_22_69 vgnd vpwr scs8hd_decap_4
XFILLER_11_129 vpwr vgnd scs8hd_fill_2
XFILLER_11_118 vpwr vgnd scs8hd_fill_2
XANTENNA__090__A _090_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_240 vpwr vgnd scs8hd_fill_2
XFILLER_19_218 vgnd vpwr scs8hd_decap_3
X_224_ chany_bottom_in[1] chany_top_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_8_27 vgnd vpwr scs8hd_decap_4
X_086_ address[1] _075_/Y address[0] _086_/X vgnd vpwr scs8hd_or3_4
X_155_ _155_/A _155_/X vgnd vpwr scs8hd_buf_1
XANTENNA__159__B _155_/X vgnd vpwr scs8hd_diode_2
XANTENNA__175__A _175_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_2_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__085__A _085_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
XFILLER_24_232 vgnd vpwr scs8hd_decap_8
XFILLER_24_210 vpwr vgnd scs8hd_fill_2
XFILLER_3_114 vpwr vgnd scs8hd_fill_2
XFILLER_3_136 vgnd vpwr scs8hd_decap_4
Xmem_top_track_16.LATCH_1_.latch data_in mem_top_track_16.LATCH_1_.latch/Q _123_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_221 vpwr vgnd scs8hd_fill_2
X_207_ _207_/A chanx_right_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_30_224 vpwr vgnd scs8hd_fill_2
XFILLER_15_276 vgnd vpwr scs8hd_fill_1
X_138_ _137_/X _138_/X vgnd vpwr scs8hd_buf_1
XANTENNA__161__C _162_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_24_3 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_2_.scs8hd_inv_1/Y
+ _176_/A mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_16.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_21_235 vpwr vgnd scs8hd_fill_2
XFILLER_21_224 vpwr vgnd scs8hd_fill_2
XFILLER_0_72 vpwr vgnd scs8hd_fill_2
XFILLER_9_92 vgnd vpwr scs8hd_fill_1
XFILLER_28_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_12.LATCH_0_.latch_SLEEPB _168_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_257 vgnd vpwr scs8hd_decap_4
Xmem_right_track_12.LATCH_0_.latch data_in _182_/A _168_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__172__B _167_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_261 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_154 vgnd vpwr scs8hd_decap_12
XFILLER_14_15 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_56 vgnd vpwr scs8hd_decap_4
XFILLER_29_110 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_2_.scs8hd_inv_1 chanx_right_in[2] mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_135 vgnd vpwr scs8hd_decap_12
XANTENNA__167__B _167_/B vgnd vpwr scs8hd_diode_2
XANTENNA__183__A _183_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_0.LATCH_3_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_6_71 vgnd vpwr scs8hd_decap_4
XFILLER_6_60 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.tap_buf4_0_.scs8hd_inv_1 mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _226_/A vgnd vpwr scs8hd_inv_1
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XPHY_69 vgnd vpwr scs8hd_decap_3
XANTENNA__077__B _075_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__093__A _090_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_190 vgnd vpwr scs8hd_decap_12
XFILLER_1_245 vgnd vpwr scs8hd_decap_4
XFILLER_17_146 vpwr vgnd scs8hd_fill_2
XFILLER_32_105 vgnd vpwr scs8hd_decap_12
XFILLER_25_190 vpwr vgnd scs8hd_fill_2
XANTENNA__178__A _178_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_127 vgnd vpwr scs8hd_decap_3
XFILLER_31_182 vgnd vpwr scs8hd_fill_1
XFILLER_11_49 vgnd vpwr scs8hd_fill_1
XFILLER_11_27 vgnd vpwr scs8hd_decap_12
XANTENNA__088__A _085_/B vgnd vpwr scs8hd_diode_2
XFILLER_36_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_171_ _157_/A _167_/B _163_/C _156_/A _171_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_22_193 vgnd vpwr scs8hd_decap_4
Xmem_bottom_track_17.LATCH_1_.latch data_in mem_bottom_track_17.LATCH_1_.latch/Q _152_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_10.LATCH_1_.latch_SLEEPB _165_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_208 vgnd vpwr scs8hd_decap_12
XANTENNA__164__C _163_/C vgnd vpwr scs8hd_diode_2
XFILLER_13_193 vpwr vgnd scs8hd_fill_2
XFILLER_13_171 vgnd vpwr scs8hd_decap_4
XFILLER_9_153 vpwr vgnd scs8hd_fill_2
XFILLER_28_219 vpwr vgnd scs8hd_fill_2
XFILLER_3_72 vpwr vgnd scs8hd_fill_2
XFILLER_36_263 vgnd vpwr scs8hd_decap_12
XFILLER_22_15 vgnd vpwr scs8hd_decap_12
XANTENNA__090__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_0_8 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_2_.scs8hd_inv_1/Y
+ _182_/A mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_42_211 vgnd vpwr scs8hd_decap_6
XFILLER_27_230 vpwr vgnd scs8hd_fill_2
X_223_ chany_bottom_in[2] chany_top_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_10_152 vgnd vpwr scs8hd_fill_1
X_085_ _085_/A _085_/B _085_/Y vgnd vpwr scs8hd_nor2_4
X_154_ _106_/A _157_/A vgnd vpwr scs8hd_buf_1
XFILLER_10_185 vgnd vpwr scs8hd_decap_4
XFILLER_6_178 vgnd vpwr scs8hd_decap_4
XFILLER_6_145 vgnd vpwr scs8hd_decap_8
Xmux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__159__C _136_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_59 vpwr vgnd scs8hd_fill_2
XFILLER_17_15 vgnd vpwr scs8hd_decap_12
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__085__B _085_/B vgnd vpwr scs8hd_diode_2
XFILLER_24_255 vpwr vgnd scs8hd_fill_2
Xmem_right_track_8.LATCH_0_.latch data_in _184_/A _170_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_4.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[6] mux_right_track_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_137_ _106_/A _167_/B _136_/X _137_/X vgnd vpwr scs8hd_or3_4
X_206_ _206_/A chanx_right_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_23_80 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_2_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__161__D _163_/D vgnd vpwr scs8hd_diode_2
XFILLER_17_3 vgnd vpwr scs8hd_decap_12
XANTENNA__186__A _186_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_269 vpwr vgnd scs8hd_fill_2
XFILLER_21_258 vgnd vpwr scs8hd_decap_4
XFILLER_21_214 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_107 vgnd vpwr scs8hd_decap_3
XANTENNA__096__A address[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _180_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_track_8.LATCH_5_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_5_29 vgnd vpwr scs8hd_decap_8
Xmux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__172__C _163_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A top_left_grid_pin_9_ vgnd vpwr scs8hd_diode_2
XFILLER_38_166 vgnd vpwr scs8hd_decap_12
XFILLER_14_27 vgnd vpwr scs8hd_decap_4
XFILLER_30_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_10.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_199 vgnd vpwr scs8hd_decap_4
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XANTENNA__167__C _162_/C vgnd vpwr scs8hd_diode_2
XFILLER_35_147 vgnd vpwr scs8hd_decap_12
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_59 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA__077__C _156_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_59 vpwr vgnd scs8hd_fill_2
XFILLER_25_15 vgnd vpwr scs8hd_decap_12
XANTENNA__093__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_19 vgnd vpwr scs8hd_fill_1
XFILLER_32_117 vgnd vpwr scs8hd_decap_12
Xmem_top_track_8.LATCH_5_.latch data_in mem_top_track_8.LATCH_5_.latch/Q _108_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_39 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1_A bottom_left_grid_pin_7_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA__088__B _109_/A vgnd vpwr scs8hd_diode_2
X_170_ _160_/A _155_/A _169_/C _162_/D _170_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__164__D _162_/D vgnd vpwr scs8hd_diode_2
XFILLER_13_150 vpwr vgnd scs8hd_fill_2
XFILLER_9_176 vgnd vpwr scs8hd_decap_4
XFILLER_9_132 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.INVTX1_1_.scs8hd_inv_1 chany_top_in[5] mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_28_209 vgnd vpwr scs8hd_decap_4
XFILLER_3_95 vpwr vgnd scs8hd_fill_2
XFILLER_3_62 vgnd vpwr scs8hd_fill_1
XANTENNA__090__C _156_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_27 vgnd vpwr scs8hd_decap_4
XANTENNA__099__A address[1] vgnd vpwr scs8hd_diode_2
X_153_ _113_/A _149_/B _153_/Y vgnd vpwr scs8hd_nor2_4
X_222_ _222_/A chany_top_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_10_164 vpwr vgnd scs8hd_fill_2
XFILLER_10_142 vpwr vgnd scs8hd_fill_2
XFILLER_6_124 vpwr vgnd scs8hd_fill_2
XFILLER_6_102 vpwr vgnd scs8hd_fill_2
X_084_ _084_/A _085_/B vgnd vpwr scs8hd_buf_1
XFILLER_12_71 vgnd vpwr scs8hd_decap_4
XFILLER_6_168 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_2.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA__159__D _162_/D vgnd vpwr scs8hd_diode_2
XFILLER_18_231 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.INVTX1_2_.scs8hd_inv_1 top_right_grid_pin_11_ mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_245 vgnd vpwr scs8hd_decap_8
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_6.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_17_27 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_15 vgnd vpwr scs8hd_decap_12
XFILLER_33_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_5_.latch_SLEEPB _139_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_245 vgnd vpwr scs8hd_decap_4
XFILLER_15_212 vgnd vpwr scs8hd_decap_3
X_136_ _135_/X _136_/X vgnd vpwr scs8hd_buf_1
X_205_ _205_/A chanx_right_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_85 vpwr vgnd scs8hd_fill_2
XFILLER_0_63 vgnd vpwr scs8hd_fill_1
XFILLER_28_15 vgnd vpwr scs8hd_decap_12
XANTENNA__096__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_12_215 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _197_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_208 vgnd vpwr scs8hd_decap_3
XFILLER_5_19 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _173_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_34_80 vgnd vpwr scs8hd_decap_12
X_119_ _085_/A _119_/B _119_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__172__D address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_12.INVTX1_0_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
Xmux_right_track_2.INVTX1_2_.scs8hd_inv_1 right_bottom_grid_pin_12_ mux_right_track_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_38_178 vgnd vpwr scs8hd_decap_12
XFILLER_30_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_244 vgnd vpwr scs8hd_fill_1
XFILLER_4_211 vgnd vpwr scs8hd_decap_3
XANTENNA__167__D _163_/D vgnd vpwr scs8hd_diode_2
XFILLER_35_159 vgnd vpwr scs8hd_decap_12
XFILLER_6_84 vpwr vgnd scs8hd_fill_2
XFILLER_6_40 vpwr vgnd scs8hd_fill_2
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XPHY_49 vgnd vpwr scs8hd_decap_3
XFILLER_25_27 vgnd vpwr scs8hd_decap_12
XANTENNA__093__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_track_1.LATCH_4_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_1_236 vpwr vgnd scs8hd_fill_2
XFILLER_1_225 vpwr vgnd scs8hd_fill_2
XFILLER_32_129 vgnd vpwr scs8hd_decap_12
XFILLER_17_159 vpwr vgnd scs8hd_fill_2
XFILLER_15_71 vpwr vgnd scs8hd_fill_2
XFILLER_31_184 vgnd vpwr scs8hd_decap_3
XFILLER_36_15 vgnd vpwr scs8hd_decap_12
XFILLER_39_240 vpwr vgnd scs8hd_fill_2
XFILLER_14_107 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_151 vpwr vgnd scs8hd_fill_2
XFILLER_7_3 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.INVTX1_4_.scs8hd_inv_1 chanx_right_in[7] mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
XANTENNA__099__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_27_276 vgnd vpwr scs8hd_fill_1
X_083_ _106_/A address[6] _162_/C _084_/A vgnd vpwr scs8hd_or3_4
X_152_ _098_/B _149_/B _152_/Y vgnd vpwr scs8hd_nor2_4
X_221_ chany_bottom_in[4] chany_top_out[5] vgnd vpwr scs8hd_buf_2
Xmux_top_track_8.INVTX1_3_.scs8hd_inv_1 chanx_right_in[2] mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_12_50 vgnd vpwr scs8hd_decap_8
XFILLER_10_198 vpwr vgnd scs8hd_fill_2
XFILLER_10_154 vgnd vpwr scs8hd_fill_1
XFILLER_10_121 vpwr vgnd scs8hd_fill_2
XFILLER_6_158 vpwr vgnd scs8hd_fill_2
XFILLER_6_114 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
Xmux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _177_/A mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_33_202 vpwr vgnd scs8hd_fill_2
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
XFILLER_18_254 vpwr vgnd scs8hd_fill_2
XFILLER_33_213 vpwr vgnd scs8hd_fill_2
XFILLER_5_191 vgnd vpwr scs8hd_fill_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB _121_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_39 vgnd vpwr scs8hd_decap_12
XFILLER_33_27 vgnd vpwr scs8hd_decap_12
X_204_ _204_/A chanx_right_out[4] vgnd vpwr scs8hd_buf_2
X_135_ _103_/Y _115_/B _081_/C _135_/X vgnd vpwr scs8hd_or3_4
XANTENNA_mem_top_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_93 vpwr vgnd scs8hd_fill_2
XFILLER_2_194 vgnd vpwr scs8hd_decap_4
XFILLER_21_249 vpwr vgnd scs8hd_fill_2
XFILLER_9_95 vpwr vgnd scs8hd_fill_2
XFILLER_9_73 vpwr vgnd scs8hd_fill_2
XFILLER_9_62 vgnd vpwr scs8hd_decap_4
XFILLER_28_27 vgnd vpwr scs8hd_decap_4
XANTENNA__096__C _156_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_205 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
X_118_ _117_/X _119_/B vgnd vpwr scs8hd_buf_1
XFILLER_7_242 vpwr vgnd scs8hd_fill_2
Xmem_right_track_4.LATCH_0_.latch data_in _176_/A _162_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_3 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_2_.latch/Q mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_2_.scs8hd_inv_1/Y
+ _174_/A mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB _085_/Y vgnd vpwr scs8hd_diode_2
XFILLER_29_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_4_223 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_9.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_30 vgnd vpwr scs8hd_fill_1
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_26_138 vpwr vgnd scs8hd_fill_2
XFILLER_26_105 vgnd vpwr scs8hd_decap_3
XPHY_39 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_17.LATCH_2_.latch_SLEEPB _151_/Y vgnd vpwr scs8hd_diode_2
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XFILLER_25_39 vgnd vpwr scs8hd_decap_12
XFILLER_1_204 vpwr vgnd scs8hd_fill_2
XFILLER_1_259 vpwr vgnd scs8hd_fill_2
XFILLER_40_141 vgnd vpwr scs8hd_decap_12
XFILLER_31_174 vgnd vpwr scs8hd_decap_8
XFILLER_16_193 vpwr vgnd scs8hd_fill_2
XFILLER_31_196 vpwr vgnd scs8hd_fill_2
Xmux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _185_/A mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_36_27 vgnd vpwr scs8hd_decap_4
XFILLER_39_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _195_/HI _178_/Y mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_26_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_53 vpwr vgnd scs8hd_fill_2
XFILLER_3_42 vgnd vpwr scs8hd_decap_4
XFILLER_3_31 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _194_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__099__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_27_211 vpwr vgnd scs8hd_fill_2
X_220_ chany_bottom_in[5] chany_top_out[6] vgnd vpwr scs8hd_buf_2
X_082_ _081_/X _162_/C vgnd vpwr scs8hd_buf_1
X_151_ _095_/B _149_/B _151_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_12_84 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[0] mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _198_/HI vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_8.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_118 vpwr vgnd scs8hd_fill_2
XFILLER_15_225 vpwr vgnd scs8hd_fill_2
X_203_ _203_/A chanx_right_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_206 vgnd vpwr scs8hd_decap_8
XFILLER_30_228 vgnd vpwr scs8hd_decap_12
XFILLER_15_236 vgnd vpwr scs8hd_decap_4
X_134_ _113_/A _128_/X _134_/Y vgnd vpwr scs8hd_nor2_4
Xmem_bottom_track_1.LATCH_1_.latch data_in mem_bottom_track_1.LATCH_1_.latch/Q _133_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_2_.scs8hd_inv_1/Y
+ _180_/A mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_0_54 vpwr vgnd scs8hd_fill_2
XFILLER_0_43 vpwr vgnd scs8hd_fill_2
XFILLER_0_32 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB _170_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_239 vgnd vpwr scs8hd_decap_4
XFILLER_18_72 vgnd vpwr scs8hd_decap_3
X_117_ _106_/A address[6] _169_/C _117_/X vgnd vpwr scs8hd_or3_4
XFILLER_34_93 vgnd vpwr scs8hd_decap_12
XFILLER_7_265 vpwr vgnd scs8hd_fill_2
XFILLER_7_254 vgnd vpwr scs8hd_decap_4
XFILLER_7_221 vgnd vpwr scs8hd_decap_4
XFILLER_15_3 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ _184_/A mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_29_147 vpwr vgnd scs8hd_fill_2
XFILLER_29_158 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_84 vgnd vpwr scs8hd_decap_8
XFILLER_4_257 vgnd vpwr scs8hd_decap_12
XFILLER_4_202 vpwr vgnd scs8hd_fill_2
XFILLER_28_180 vpwr vgnd scs8hd_fill_2
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_26_117 vgnd vpwr scs8hd_decap_12
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XFILLER_25_194 vpwr vgnd scs8hd_fill_2
XFILLER_15_84 vpwr vgnd scs8hd_fill_2
XFILLER_15_62 vpwr vgnd scs8hd_fill_2
XFILLER_15_51 vgnd vpwr scs8hd_decap_8
XFILLER_40_186 vgnd vpwr scs8hd_fill_1
XANTENNA__102__A address[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_275 vpwr vgnd scs8hd_fill_2
XFILLER_39_253 vpwr vgnd scs8hd_fill_2
XFILLER_39_220 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_6.LATCH_1_.latch_SLEEPB _163_/Y vgnd vpwr scs8hd_diode_2
XFILLER_13_197 vpwr vgnd scs8hd_fill_2
XFILLER_13_142 vgnd vpwr scs8hd_decap_4
XFILLER_9_157 vpwr vgnd scs8hd_fill_2
XFILLER_3_76 vpwr vgnd scs8hd_fill_2
XFILLER_8_190 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _179_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_27_245 vgnd vpwr scs8hd_decap_3
XFILLER_27_234 vgnd vpwr scs8hd_decap_4
XFILLER_27_201 vpwr vgnd scs8hd_fill_2
X_150_ _110_/A _149_/B _150_/Y vgnd vpwr scs8hd_nor2_4
X_081_ address[3] address[4] _081_/C _081_/X vgnd vpwr scs8hd_or3_4
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_259 vpwr vgnd scs8hd_fill_2
XFILLER_18_267 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A top_left_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _174_/Y vgnd vpwr
+ scs8hd_diode_2
X_133_ _098_/B _128_/X _133_/Y vgnd vpwr scs8hd_nor2_4
X_202_ _202_/A chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_23_62 vgnd vpwr scs8hd_decap_3
XFILLER_23_51 vgnd vpwr scs8hd_decap_8
XANTENNA__110__A _110_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_84 vpwr vgnd scs8hd_fill_2
X_116_ _116_/A _169_/C vgnd vpwr scs8hd_buf_1
XANTENNA__105__A _104_/X vgnd vpwr scs8hd_diode_2
XFILLER_11_240 vpwr vgnd scs8hd_fill_2
XFILLER_39_17 vpwr vgnd scs8hd_fill_2
XFILLER_39_28 vpwr vgnd scs8hd_fill_2
XFILLER_29_126 vpwr vgnd scs8hd_fill_2
XFILLER_20_74 vgnd vpwr scs8hd_fill_1
XFILLER_4_269 vgnd vpwr scs8hd_decap_6
XFILLER_4_247 vgnd vpwr scs8hd_fill_1
XFILLER_6_32 vgnd vpwr scs8hd_decap_8
XPHY_19 vgnd vpwr scs8hd_decap_3
Xmem_top_track_8.LATCH_0_.latch data_in mem_top_track_8.LATCH_0_.latch/Q _113_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_118 vpwr vgnd scs8hd_fill_2
XFILLER_40_154 vgnd vpwr scs8hd_decap_12
XFILLER_25_184 vgnd vpwr scs8hd_decap_3
XFILLER_31_51 vgnd vpwr scs8hd_decap_8
XFILLER_31_62 vgnd vpwr scs8hd_decap_12
XFILLER_31_110 vgnd vpwr scs8hd_decap_12
XFILLER_16_173 vgnd vpwr scs8hd_fill_1
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_176 vpwr vgnd scs8hd_fill_2
XFILLER_22_165 vpwr vgnd scs8hd_fill_2
XFILLER_22_132 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _176_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__203__A _203_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_84 vgnd vpwr scs8hd_decap_8
XFILLER_42_94 vgnd vpwr scs8hd_decap_12
XFILLER_13_154 vpwr vgnd scs8hd_fill_2
XFILLER_9_136 vpwr vgnd scs8hd_fill_2
XFILLER_9_114 vpwr vgnd scs8hd_fill_2
XANTENNA__113__A _113_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_202 vgnd vpwr scs8hd_decap_12
XFILLER_3_99 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_2_.latch/Q mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_268 vgnd vpwr scs8hd_decap_8
XFILLER_27_257 vpwr vgnd scs8hd_fill_2
X_080_ enable _081_/C vgnd vpwr scs8hd_inv_8
XFILLER_42_249 vgnd vpwr scs8hd_decap_12
XFILLER_10_168 vpwr vgnd scs8hd_fill_2
XFILLER_10_146 vgnd vpwr scs8hd_decap_6
XFILLER_10_102 vpwr vgnd scs8hd_fill_2
XFILLER_6_106 vgnd vpwr scs8hd_decap_6
Xmux_bottom_track_17.INVTX1_7_.scs8hd_inv_1 bottom_left_grid_pin_15_ mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_128 vgnd vpwr scs8hd_decap_8
XFILLER_5_3 vpwr vgnd scs8hd_fill_2
XFILLER_41_260 vgnd vpwr scs8hd_decap_12
XFILLER_18_235 vpwr vgnd scs8hd_fill_2
XANTENNA__108__A _085_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_2_.latch_SLEEPB _142_/Y vgnd vpwr scs8hd_diode_2
XFILLER_38_3 vgnd vpwr scs8hd_decap_12
XFILLER_32_271 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_12.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_132_ _095_/B _128_/X _132_/Y vgnd vpwr scs8hd_nor2_4
X_201_ _201_/A chanx_right_out[7] vgnd vpwr scs8hd_buf_2
Xmem_top_track_0.LATCH_5_.latch data_in mem_top_track_0.LATCH_5_.latch/Q _085_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_271 vgnd vpwr scs8hd_decap_6
Xmem_bottom_track_9.LATCH_2_.latch data_in mem_bottom_track_9.LATCH_2_.latch/Q _142_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__110__B _110_/B vgnd vpwr scs8hd_diode_2
XFILLER_0_23 vpwr vgnd scs8hd_fill_2
XFILLER_0_12 vgnd vpwr scs8hd_decap_8
XFILLER_0_89 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _175_/A mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _174_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_274 vgnd vpwr scs8hd_fill_1
XANTENNA__211__A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
X_115_ address[3] _115_/B _081_/C _116_/A vgnd vpwr scs8hd_or3_4
XANTENNA__121__A _110_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_105 vgnd vpwr scs8hd_decap_12
XFILLER_37_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__206__A _206_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_7_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_29_62 vgnd vpwr scs8hd_decap_12
XFILLER_29_51 vgnd vpwr scs8hd_decap_8
XANTENNA__116__A _116_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_88 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_2_.latch data_in mem_top_track_16.LATCH_2_.latch/Q _122_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_3 vgnd vpwr scs8hd_decap_12
XFILLER_34_141 vgnd vpwr scs8hd_decap_12
XFILLER_19_193 vpwr vgnd scs8hd_fill_2
XFILLER_19_171 vgnd vpwr scs8hd_decap_6
XFILLER_19_160 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _196_/HI _183_/Y mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_166 vgnd vpwr scs8hd_decap_12
XFILLER_25_152 vpwr vgnd scs8hd_fill_2
XFILLER_31_74 vgnd vpwr scs8hd_decap_12
XFILLER_0_273 vgnd vpwr scs8hd_decap_4
XFILLER_16_163 vpwr vgnd scs8hd_fill_2
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_166 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _189_/HI vgnd vpwr
+ scs8hd_diode_2
.ends

