* NGSPICE file created from sb_2__2_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_dfxbp_1 abstract view
.subckt scs8hd_dfxbp_1 CLK D Q QN vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_mux2_1 abstract view
.subckt scs8hd_mux2_1 A0 A1 S X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

.subckt sb_2__2_ bottom_left_grid_pin_34_ bottom_left_grid_pin_35_ bottom_left_grid_pin_36_
+ bottom_left_grid_pin_37_ bottom_left_grid_pin_38_ bottom_left_grid_pin_39_ bottom_left_grid_pin_40_
+ bottom_left_grid_pin_41_ bottom_right_grid_pin_1_ ccff_head ccff_tail chanx_left_in[0]
+ chanx_left_in[10] chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14]
+ chanx_left_in[15] chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19]
+ chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5]
+ chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0]
+ chanx_left_out[10] chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14]
+ chanx_left_out[15] chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19]
+ chanx_left_out[1] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5]
+ chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chany_bottom_in[0]
+ chany_bottom_in[10] chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13]
+ chany_bottom_in[14] chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17]
+ chany_bottom_in[18] chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4]
+ chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8]
+ chany_bottom_out[9] left_top_grid_pin_1_ prog_clk vpwr vgnd
XFILLER_36_19 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_39.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_39.mux_l1_in_0_/S
+ mux_bottom_track_39.mux_l2_in_0_/S mem_bottom_track_39.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_22_166 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_25.scs8hd_buf_4_0_ mux_bottom_track_25.mux_l2_in_0_/X _75_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_9_104 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_3.mux_l1_in_1_ bottom_left_grid_pin_40_ bottom_left_grid_pin_38_
+ mux_bottom_track_3.mux_l1_in_1_/S mux_bottom_track_3.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
X_83_ _83_/A chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_11.mux_l1_in_0__A0 chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_27_269 vgnd vpwr scs8hd_decap_8
XFILLER_6_129 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_19.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_37_62 vgnd vpwr scs8hd_decap_12
XFILLER_37_51 vgnd vpwr scs8hd_decap_8
XFILLER_5_173 vpwr vgnd scs8hd_fill_2
X_66_ chany_bottom_in[0] chanx_left_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_24_239 vgnd vpwr scs8hd_decap_12
XFILLER_23_42 vgnd vpwr scs8hd_decap_6
XFILLER_2_110 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l3_in_0__S mux_bottom_track_1.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_23.scs8hd_dfxbp_1_0__D mux_bottom_track_21.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
X_49_ chany_bottom_in[17] chanx_left_out[18] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_2__D mux_bottom_track_5.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_7.mux_l2_in_1__S mux_bottom_track_7.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_75 vgnd vpwr scs8hd_decap_12
XFILLER_11_220 vgnd vpwr scs8hd_decap_3
XFILLER_11_242 vpwr vgnd scs8hd_fill_2
XFILLER_7_235 vgnd vpwr scs8hd_decap_8
XFILLER_38_117 vgnd vpwr scs8hd_decap_12
XFILLER_22_7 vgnd vpwr scs8hd_decap_12
XFILLER_39_19 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_0_ chanx_left_in[9] bottom_left_grid_pin_37_ mux_bottom_track_17.mux_l1_in_0_/S
+ mux_bottom_track_17.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_29_74 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_29.mux_l2_in_0_ _45_/HI mux_bottom_track_29.mux_l1_in_0_/X mux_bottom_track_29.mux_l2_in_0_/S
+ mux_bottom_track_29.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_6_23 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_13.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_11.mux_l2_in_0_/S
+ mux_bottom_track_13.mux_l1_in_0_/S mem_bottom_track_13.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_6_45 vgnd vpwr scs8hd_fill_1
XFILLER_6_56 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_19.mux_l2_in_0__S mux_bottom_track_19.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_3 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_31.mux_l2_in_0_ _47_/HI mux_bottom_track_31.mux_l1_in_0_/X mux_bottom_track_31.mux_l2_in_0_/S
+ mux_bottom_track_31.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_bottom_track_33.scs8hd_buf_4_0_ mux_bottom_track_33.mux_l2_in_0_/X _71_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_40_178 vgnd vpwr scs8hd_decap_12
XFILLER_31_31 vgnd vpwr scs8hd_decap_12
XFILLER_15_87 vgnd vpwr scs8hd_decap_12
XFILLER_0_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_3.mux_l1_in_1__A0 bottom_left_grid_pin_40_ vgnd vpwr scs8hd_diode_2
XFILLER_31_123 vgnd vpwr scs8hd_decap_12
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_245 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_39.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_37.mux_l2_in_0_/S
+ mux_bottom_track_39.mux_l1_in_0_/S mem_bottom_track_39.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_22_178 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_21.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_27.scs8hd_buf_4_0__A mux_bottom_track_27.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_112 vpwr vgnd scs8hd_fill_2
XFILLER_13_123 vgnd vpwr scs8hd_decap_6
XFILLER_42_63 vgnd vpwr scs8hd_decap_12
XFILLER_9_138 vgnd vpwr scs8hd_decap_4
XFILLER_13_178 vgnd vpwr scs8hd_decap_4
XFILLER_3_79 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_3.mux_l1_in_0_ bottom_left_grid_pin_36_ bottom_left_grid_pin_34_
+ mux_bottom_track_3.mux_l1_in_1_/S mux_bottom_track_3.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_36_215 vgnd vpwr scs8hd_decap_12
X_82_ _82_/A chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_11.mux_l1_in_0__A1 bottom_left_grid_pin_34_ vgnd vpwr scs8hd_diode_2
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_39.mux_l2_in_0__A0 _27_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0__A0 mux_bottom_track_3.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_12_55 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_1__D mux_bottom_track_7.mux_l1_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_74 vgnd vpwr scs8hd_decap_12
XFILLER_18_215 vgnd vpwr scs8hd_decap_12
XFILLER_5_152 vpwr vgnd scs8hd_fill_2
X_65_ _65_/A chanx_left_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_32_251 vgnd vpwr scs8hd_decap_12
XFILLER_23_21 vgnd vpwr scs8hd_decap_6
XFILLER_2_133 vpwr vgnd scs8hd_fill_2
XFILLER_0_58 vpwr vgnd scs8hd_fill_2
XFILLER_9_56 vgnd vpwr scs8hd_decap_3
XFILLER_14_251 vgnd vpwr scs8hd_decap_12
X_48_ chany_bottom_in[18] chanx_left_out[19] vgnd vpwr scs8hd_buf_2
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
Xmem_left_track_1.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_1.mux_l1_in_0_/S mux_left_track_1.mux_l2_in_0_/S
+ mem_left_track_1.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_18_87 vgnd vpwr scs8hd_decap_4
XFILLER_38_129 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_3.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_track_3.mux_l2_in_0_/S mux_bottom_track_3.mux_l3_in_0_/S
+ mem_bottom_track_3.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_37_184 vgnd vpwr scs8hd_decap_12
XFILLER_20_11 vgnd vpwr scs8hd_fill_1
XFILLER_20_55 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_bottom_track_35.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_19_184 vgnd vpwr scs8hd_decap_12
XFILLER_34_154 vgnd vpwr scs8hd_decap_12
XFILLER_15_11 vgnd vpwr scs8hd_decap_3
XFILLER_15_22 vgnd vpwr scs8hd_fill_1
XFILLER_25_121 vgnd vpwr scs8hd_fill_1
XFILLER_31_43 vgnd vpwr scs8hd_decap_12
XFILLER_15_99 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__D mux_bottom_track_7.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_275 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_1__A1 bottom_left_grid_pin_38_ vgnd vpwr scs8hd_diode_2
XFILLER_31_135 vgnd vpwr scs8hd_decap_12
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_154 vgnd vpwr scs8hd_decap_12
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_257 vgnd vpwr scs8hd_decap_12
XFILLER_30_190 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_29.mux_l1_in_0_ chanx_left_in[15] bottom_left_grid_pin_35_ mux_bottom_track_29.mux_l1_in_0_/S
+ mux_bottom_track_29.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_26_32 vgnd vpwr scs8hd_decap_12
XFILLER_42_75 vgnd vpwr scs8hd_decap_12
X_81_ _81_/A chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_3_58 vgnd vpwr scs8hd_fill_1
XFILLER_36_227 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_31.mux_l1_in_0_ chanx_left_in[16] bottom_left_grid_pin_36_ mux_bottom_track_31.mux_l1_in_0_/S
+ mux_bottom_track_31.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_8_150 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_23.mux_l1_in_0__S mux_bottom_track_23.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_39.mux_l2_in_0__A1 mux_bottom_track_39.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0__A1 mux_bottom_track_3.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_10_127 vpwr vgnd scs8hd_fill_2
XFILLER_10_149 vpwr vgnd scs8hd_fill_2
XFILLER_12_23 vpwr vgnd scs8hd_fill_2
XFILLER_37_86 vgnd vpwr scs8hd_decap_12
XFILLER_33_208 vgnd vpwr scs8hd_decap_12
XFILLER_18_227 vgnd vpwr scs8hd_decap_12
X_64_ chany_bottom_in[2] chanx_left_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_32_263 vgnd vpwr scs8hd_decap_12
XFILLER_15_208 vgnd vpwr scs8hd_decap_12
XFILLER_23_55 vpwr vgnd scs8hd_fill_2
XFILLER_2_145 vpwr vgnd scs8hd_fill_2
XFILLER_2_167 vpwr vgnd scs8hd_fill_2
XFILLER_9_35 vpwr vgnd scs8hd_fill_2
XFILLER_14_263 vgnd vpwr scs8hd_decap_12
XFILLER_9_68 vpwr vgnd scs8hd_fill_2
X_47_ _47_/HI _47_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mem_bottom_track_27.scs8hd_dfxbp_1_1__D mux_bottom_track_27.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_11 vgnd vpwr scs8hd_fill_1
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
Xmem_left_track_1.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_39.mux_l2_in_0_/S mux_left_track_1.mux_l1_in_0_/S
+ mem_left_track_1.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
Xmem_bottom_track_3.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_3.mux_l1_in_1_/S mux_bottom_track_3.mux_l2_in_0_/S
+ mem_bottom_track_3.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_37_196 vgnd vpwr scs8hd_decap_12
XFILLER_4_218 vgnd vpwr scs8hd_decap_8
XFILLER_4_229 vgnd vpwr scs8hd_decap_12
XFILLER_28_141 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_3.mux_l2_in_1__S mux_bottom_track_3.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_34_166 vgnd vpwr scs8hd_decap_12
XFILLER_19_196 vgnd vpwr scs8hd_decap_12
XFILLER_31_55 vgnd vpwr scs8hd_decap_6
XFILLER_0_221 vgnd vpwr scs8hd_decap_12
XFILLER_16_166 vgnd vpwr scs8hd_decap_12
XFILLER_31_147 vgnd vpwr scs8hd_decap_12
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_15.mux_l2_in_0__S mux_bottom_track_15.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_15.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_26_44 vgnd vpwr scs8hd_decap_6
XFILLER_42_87 vgnd vpwr scs8hd_decap_6
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XFILLER_9_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_13.mux_l2_in_0__A0 _37_/HI vgnd vpwr scs8hd_diode_2
X_80_ _80_/A chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_3_37 vpwr vgnd scs8hd_fill_2
XFILLER_3_26 vpwr vgnd scs8hd_fill_2
XFILLER_36_239 vgnd vpwr scs8hd_decap_12
XFILLER_8_140 vgnd vpwr scs8hd_decap_4
XFILLER_8_173 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_5.scs8hd_buf_4_0_ mux_bottom_track_5.mux_l3_in_0_/X _85_/A vgnd
+ vpwr scs8hd_buf_1
Xmem_bottom_track_21.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_21.mux_l1_in_0_/S
+ mux_bottom_track_21.mux_l2_in_0_/S mem_bottom_track_21.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XANTENNA_mem_bottom_track_29.scs8hd_dfxbp_1_0__D mux_bottom_track_27.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_220 vgnd vpwr scs8hd_decap_12
XFILLER_37_98 vgnd vpwr scs8hd_decap_12
XFILLER_18_239 vgnd vpwr scs8hd_decap_12
XFILLER_5_110 vgnd vpwr scs8hd_fill_1
XFILLER_38_7 vgnd vpwr scs8hd_decap_12
XFILLER_5_198 vgnd vpwr scs8hd_decap_6
X_63_ _63_/A chanx_left_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_23_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_7.mux_l1_in_0__A0 bottom_left_grid_pin_36_ vgnd vpwr scs8hd_diode_2
XFILLER_0_27 vpwr vgnd scs8hd_fill_2
X_46_ _46_/HI _46_/LO vgnd vpwr scs8hd_conb_1
Xmem_left_track_9.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_9.mux_l1_in_0_/S mux_left_track_9.mux_l2_in_0_/S
+ mem_left_track_9.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_18_23 vgnd vpwr scs8hd_decap_6
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_2__A0 chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_7_227 vpwr vgnd scs8hd_fill_2
XFILLER_11_234 vgnd vpwr scs8hd_decap_8
XFILLER_11_245 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_3.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_1.mux_l3_in_0_/S mux_bottom_track_3.mux_l1_in_1_/S
+ mem_bottom_track_3.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
X_29_ _29_/HI _29_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_70 vpwr vgnd scs8hd_fill_2
XFILLER_29_11 vgnd vpwr scs8hd_decap_12
XFILLER_20_68 vgnd vpwr scs8hd_decap_12
XFILLER_6_48 vpwr vgnd scs8hd_fill_2
XFILLER_20_7 vgnd vpwr scs8hd_decap_4
XFILLER_34_178 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l2_in_1__A0 _28_/HI vgnd vpwr scs8hd_diode_2
XFILLER_25_123 vgnd vpwr scs8hd_decap_12
XFILLER_15_46 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_21.mux_l2_in_0__A0 _41_/HI vgnd vpwr scs8hd_diode_2
XFILLER_0_244 vgnd vpwr scs8hd_decap_4
XFILLER_0_233 vgnd vpwr scs8hd_decap_4
XFILLER_0_200 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__D mux_left_track_25.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_16_178 vgnd vpwr scs8hd_decap_12
XFILLER_31_159 vgnd vpwr scs8hd_decap_12
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_91 vpwr vgnd scs8hd_fill_2
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XFILLER_9_108 vgnd vpwr scs8hd_decap_3
Xmux_left_track_9.scs8hd_buf_4_0_ mux_left_track_9.mux_l2_in_0_/X _63_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mux_bottom_track_13.mux_l2_in_0__A1 mux_bottom_track_13.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l3_in_0__A0 mux_bottom_track_5.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_196 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_21.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_19.mux_l2_in_0_/S
+ mux_bottom_track_21.mux_l1_in_0_/S mem_bottom_track_21.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_12_14 vpwr vgnd scs8hd_fill_2
XFILLER_37_11 vpwr vgnd scs8hd_fill_2
XFILLER_41_232 vgnd vpwr scs8hd_decap_12
XFILLER_26_251 vgnd vpwr scs8hd_decap_12
XFILLER_5_177 vgnd vpwr scs8hd_decap_4
X_62_ chany_bottom_in[4] chanx_left_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.mux_l2_in_0__A0 _31_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_7.mux_l1_in_0__A1 bottom_left_grid_pin_34_ vgnd vpwr scs8hd_diode_2
XFILLER_23_232 vgnd vpwr scs8hd_decap_12
XFILLER_23_13 vgnd vpwr scs8hd_fill_1
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_35.scs8hd_buf_4_0__A mux_bottom_track_35.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
X_45_ _45_/HI _45_/LO vgnd vpwr scs8hd_conb_1
Xmem_left_track_9.scs8hd_dfxbp_1_0_ prog_clk mux_left_track_5.mux_l2_in_0_/S mux_left_track_9.mux_l1_in_0_/S
+ mem_left_track_9.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_20_202 vgnd vpwr scs8hd_decap_12
XFILLER_34_56 vgnd vpwr scs8hd_decap_12
XFILLER_11_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l1_in_2__A1 bottom_left_grid_pin_41_ vgnd vpwr scs8hd_diode_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_110 vgnd vpwr scs8hd_decap_12
X_28_ _28_/HI _28_/LO vgnd vpwr scs8hd_conb_1
XFILLER_20_14 vgnd vpwr scs8hd_fill_1
XFILLER_29_78 vgnd vpwr scs8hd_decap_12
XFILLER_29_23 vgnd vpwr scs8hd_decap_12
XFILLER_28_154 vgnd vpwr scs8hd_decap_12
XFILLER_6_27 vpwr vgnd scs8hd_fill_2
XFILLER_13_7 vpwr vgnd scs8hd_fill_2
XFILLER_19_110 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l2_in_1__A1 mux_bottom_track_5.mux_l1_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_25_135 vgnd vpwr scs8hd_decap_12
XFILLER_40_105 vgnd vpwr scs8hd_decap_12
XFILLER_15_25 vpwr vgnd scs8hd_fill_2
XFILLER_15_58 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_21.mux_l2_in_0__A1 mux_bottom_track_21.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_0_212 vpwr vgnd scs8hd_fill_2
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_190 vgnd vpwr scs8hd_decap_12
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_105 vgnd vpwr scs8hd_decap_12
XFILLER_13_116 vgnd vpwr scs8hd_decap_6
XFILLER_42_56 vgnd vpwr scs8hd_decap_6
XFILLER_21_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_2__S mux_bottom_track_5.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_bottom_track_29.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_29.mux_l1_in_0_/S
+ mux_bottom_track_29.mux_l2_in_0_/S mem_bottom_track_29.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_5.mux_l3_in_0__A1 mux_bottom_track_5.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_27_208 vgnd vpwr scs8hd_decap_12
XFILLER_12_59 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.mux_l2_in_0__S mux_bottom_track_9.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_11.mux_l2_in_0__S mux_bottom_track_11.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_26_263 vgnd vpwr scs8hd_decap_12
XFILLER_5_123 vgnd vpwr scs8hd_decap_4
XFILLER_5_156 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0__A0 chanx_left_in[9] vgnd vpwr scs8hd_diode_2
X_61_ chany_bottom_in[5] chanx_left_out[6] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_track_1.mux_l2_in_0__A1 mux_left_track_1.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_71 vpwr vgnd scs8hd_fill_2
XFILLER_2_137 vpwr vgnd scs8hd_fill_2
XFILLER_14_211 vgnd vpwr scs8hd_decap_3
XFILLER_9_16 vpwr vgnd scs8hd_fill_2
X_44_ _44_/HI _44_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_11.scs8hd_dfxbp_1_0__D mux_bottom_track_9.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_14 vpwr vgnd scs8hd_fill_2
XFILLER_34_68 vgnd vpwr scs8hd_decap_12
XFILLER_11_269 vgnd vpwr scs8hd_decap_8
XFILLER_1_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_31.scs8hd_dfxbp_1_0__D mux_bottom_track_29.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_90 vpwr vgnd scs8hd_fill_2
X_27_ _27_/HI _27_/LO vgnd vpwr scs8hd_conb_1
XFILLER_20_26 vgnd vpwr scs8hd_decap_3
XFILLER_29_35 vgnd vpwr scs8hd_decap_12
XFILLER_28_166 vgnd vpwr scs8hd_decap_12
XFILLER_3_243 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_13.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_42_180 vgnd vpwr scs8hd_decap_6
XFILLER_40_117 vgnd vpwr scs8hd_decap_12
XFILLER_25_147 vgnd vpwr scs8hd_decap_12
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_39.scs8hd_buf_4_0_ mux_bottom_track_39.mux_l2_in_0_/X _68_/A vgnd
+ vpwr scs8hd_buf_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_0 vgnd vpwr scs8hd_decap_3
XFILLER_22_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_1__A0 _30_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_25.mux_l1_in_0__A0 bottom_left_grid_pin_41_ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_13.mux_l2_in_0_ _37_/HI mux_bottom_track_13.mux_l1_in_0_/X mux_bottom_track_13.mux_l2_in_0_/S
+ mux_bottom_track_13.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmem_bottom_track_29.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_27.mux_l2_in_0_/S
+ mux_bottom_track_29.mux_l1_in_0_/S mem_bottom_track_29.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_8_110 vpwr vgnd scs8hd_fill_2
XFILLER_8_154 vpwr vgnd scs8hd_fill_2
XFILLER_16_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_17.scs8hd_buf_4_0__A mux_bottom_track_17.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_220 vgnd vpwr scs8hd_decap_12
XFILLER_12_27 vpwr vgnd scs8hd_fill_2
XFILLER_41_245 vgnd vpwr scs8hd_decap_12
XFILLER_5_102 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0__A1 bottom_left_grid_pin_37_ vgnd vpwr scs8hd_diode_2
X_60_ chany_bottom_in[6] chanx_left_out[7] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0__A0 mux_bottom_track_9.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_17_220 vgnd vpwr scs8hd_decap_12
XFILLER_23_48 vgnd vpwr scs8hd_fill_1
XFILLER_23_59 vpwr vgnd scs8hd_fill_2
XFILLER_23_245 vgnd vpwr scs8hd_decap_12
XFILLER_2_149 vpwr vgnd scs8hd_fill_2
XFILLER_9_39 vpwr vgnd scs8hd_fill_2
XFILLER_13_81 vpwr vgnd scs8hd_fill_2
XFILLER_36_7 vgnd vpwr scs8hd_decap_12
XFILLER_1_193 vpwr vgnd scs8hd_fill_2
X_43_ _43_/HI _43_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_left_track_5.mux_l1_in_0__A0 left_top_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XFILLER_20_215 vgnd vpwr scs8hd_decap_12
XFILLER_7_208 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_27.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_11_226 vpwr vgnd scs8hd_fill_2
XFILLER_6_274 vgnd vpwr scs8hd_fill_1
XFILLER_37_123 vgnd vpwr scs8hd_decap_12
X_26_ _26_/HI _26_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_51 vpwr vgnd scs8hd_fill_2
XFILLER_1_62 vpwr vgnd scs8hd_fill_2
XFILLER_29_47 vgnd vpwr scs8hd_decap_12
XFILLER_28_178 vgnd vpwr scs8hd_decap_12
XANTENNA__50__A chany_bottom_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_3_200 vpwr vgnd scs8hd_fill_2
XFILLER_19_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_37.mux_l1_in_0__S mux_bottom_track_37.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_40_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_33.mux_l1_in_0__A0 chanx_left_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_15_16 vgnd vpwr scs8hd_decap_6
XFILLER_15_38 vpwr vgnd scs8hd_fill_2
XFILLER_25_159 vgnd vpwr scs8hd_decap_12
XFILLER_0_203 vgnd vpwr scs8hd_fill_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_22_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_1__A1 chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_38_251 vgnd vpwr scs8hd_decap_12
XFILLER_13_129 vgnd vpwr scs8hd_fill_1
XFILLER_26_59 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_25.mux_l1_in_0__A1 bottom_right_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XFILLER_21_184 vgnd vpwr scs8hd_decap_12
XFILLER_32_80 vgnd vpwr scs8hd_decap_12
XFILLER_35_232 vgnd vpwr scs8hd_decap_12
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
XFILLER_41_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.scs8hd_buf_4_0__A mux_bottom_track_5.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_5_114 vpwr vgnd scs8hd_fill_2
XFILLER_32_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_2__S mux_bottom_track_1.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0__A1 mux_bottom_track_9.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_17_232 vgnd vpwr scs8hd_decap_12
XFILLER_4_180 vgnd vpwr scs8hd_decap_4
XFILLER_4_84 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_13.mux_l1_in_0_ chanx_left_in[7] bottom_left_grid_pin_35_ mux_bottom_track_13.mux_l1_in_0_/S
+ mux_bottom_track_13.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_23_257 vgnd vpwr scs8hd_decap_12
XFILLER_2_106 vpwr vgnd scs8hd_fill_2
XANTENNA__53__A chany_bottom_in[13] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0__S mux_bottom_track_5.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_25.mux_l2_in_0_ mux_bottom_track_25.mux_l1_in_1_/X mux_bottom_track_25.mux_l1_in_0_/X
+ mux_bottom_track_25.mux_l2_in_0_/S mux_bottom_track_25.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_mux2_1
XFILLER_29_7 vpwr vgnd scs8hd_fill_2
X_42_ _42_/HI _42_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_left_track_5.mux_l1_in_0__A1 chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_20_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_15.scs8hd_dfxbp_1_1__D mux_bottom_track_15.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA__48__A chany_bottom_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_40_80 vgnd vpwr scs8hd_decap_12
XFILLER_6_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_29.mux_l2_in_0__S mux_bottom_track_29.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_37_135 vgnd vpwr scs8hd_decap_12
XFILLER_1_74 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_35.scs8hd_dfxbp_1_1__D mux_bottom_track_35.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
X_25_ _25_/HI _25_/LO vgnd vpwr scs8hd_conb_1
XFILLER_29_59 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_25.mux_l1_in_1_ _43_/HI chanx_left_in[13] mux_bottom_track_25.mux_l1_in_1_/S
+ mux_bottom_track_25.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_36_190 vgnd vpwr scs8hd_decap_12
XFILLER_3_245 vgnd vpwr scs8hd_decap_12
XFILLER_3_212 vpwr vgnd scs8hd_fill_2
XFILLER_10_83 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l2_in_0_ mux_bottom_track_9.mux_l1_in_1_/X mux_bottom_track_9.mux_l1_in_0_/X
+ mux_bottom_track_9.mux_l2_in_0_/S mux_bottom_track_9.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_34_105 vgnd vpwr scs8hd_decap_12
XFILLER_19_135 vgnd vpwr scs8hd_decap_12
XFILLER_25_105 vgnd vpwr scs8hd_decap_12
XFILLER_33_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_33.mux_l1_in_0__A1 bottom_left_grid_pin_37_ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_13.scs8hd_buf_4_0_ mux_bottom_track_13.mux_l2_in_0_/X _81_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_18_190 vgnd vpwr scs8hd_decap_12
XFILLER_0_259 vpwr vgnd scs8hd_fill_2
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_105 vgnd vpwr scs8hd_decap_12
XFILLER_31_108 vgnd vpwr scs8hd_decap_12
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__61__A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_21_71 vgnd vpwr scs8hd_decap_12
XFILLER_39_208 vgnd vpwr scs8hd_decap_12
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_15_171 vgnd vpwr scs8hd_decap_12
XFILLER_30_141 vgnd vpwr scs8hd_decap_12
XFILLER_7_62 vgnd vpwr scs8hd_decap_3
XFILLER_38_263 vgnd vpwr scs8hd_decap_12
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.mux_l1_in_1_ _30_/HI chanx_left_in[5] mux_bottom_track_9.mux_l1_in_0_/S
+ mux_bottom_track_9.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_21_196 vgnd vpwr scs8hd_decap_12
XANTENNA__56__A chany_bottom_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_16_93 vgnd vpwr scs8hd_decap_12
XFILLER_8_123 vpwr vgnd scs8hd_fill_2
XFILLER_12_152 vgnd vpwr scs8hd_fill_1
XFILLER_12_163 vgnd vpwr scs8hd_decap_12
XFILLER_12_18 vgnd vpwr scs8hd_decap_3
XFILLER_37_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_19.mux_l2_in_0__A0 _40_/HI vgnd vpwr scs8hd_diode_2
XFILLER_37_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_0__D mux_bottom_track_15.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_269 vgnd vpwr scs8hd_decap_8
Xmem_bottom_track_11.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_11.mux_l1_in_0_/S
+ mux_bottom_track_11.mux_l2_in_0_/S mem_bottom_track_11.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_4_192 vgnd vpwr scs8hd_decap_8
XFILLER_4_41 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_37.scs8hd_dfxbp_1_0__D mux_bottom_track_35.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_17 vpwr vgnd scs8hd_fill_2
XFILLER_23_269 vgnd vpwr scs8hd_decap_8
XFILLER_14_203 vgnd vpwr scs8hd_decap_8
X_41_ _41_/HI _41_/LO vgnd vpwr scs8hd_conb_1
XFILLER_38_80 vgnd vpwr scs8hd_decap_12
XFILLER_20_239 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_37.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_37.mux_l1_in_0_/S
+ mux_bottom_track_37.mux_l2_in_0_/S mem_bottom_track_37.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XANTENNA__64__A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_10_250 vgnd vpwr scs8hd_decap_12
XFILLER_24_93 vgnd vpwr scs8hd_decap_12
XFILLER_6_232 vgnd vpwr scs8hd_decap_12
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_9.mux_l2_in_0__S mux_left_track_9.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_147 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_21.scs8hd_buf_4_0_ mux_bottom_track_21.mux_l2_in_0_/X _77_/A vgnd
+ vpwr scs8hd_buf_1
X_24_ _24_/HI _24_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_1_97 vpwr vgnd scs8hd_fill_2
XFILLER_20_18 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_25.mux_l1_in_0_ bottom_left_grid_pin_41_ bottom_right_grid_pin_1_
+ mux_bottom_track_25.mux_l1_in_1_/S mux_bottom_track_25.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_mux2_1
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__D mux_left_track_1.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_257 vgnd vpwr scs8hd_decap_12
XFILLER_3_235 vpwr vgnd scs8hd_fill_2
XFILLER_3_224 vpwr vgnd scs8hd_fill_2
XFILLER_10_62 vpwr vgnd scs8hd_fill_2
XANTENNA__59__A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_19_60 vgnd vpwr scs8hd_fill_1
XFILLER_19_147 vgnd vpwr scs8hd_decap_12
XFILLER_34_117 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_37.mux_l2_in_0_ _26_/HI mux_bottom_track_37.mux_l1_in_0_/X mux_bottom_track_37.mux_l2_in_0_/S
+ mux_bottom_track_37.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_25_117 vgnd vpwr scs8hd_decap_4
XFILLER_0_249 vgnd vpwr scs8hd_decap_6
XFILLER_0_216 vgnd vpwr scs8hd_fill_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_117 vgnd vpwr scs8hd_decap_12
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_83 vgnd vpwr scs8hd_decap_12
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_7_30 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_27.mux_l2_in_0__A0 _44_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_33.mux_l1_in_0__S mux_bottom_track_33.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_9.mux_l1_in_0_ bottom_left_grid_pin_41_ bottom_right_grid_pin_1_
+ mux_bottom_track_9.mux_l1_in_0_/S mux_bottom_track_9.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_29_220 vgnd vpwr scs8hd_decap_12
XANTENNA__72__A _72_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_93 vgnd vpwr scs8hd_decap_12
XFILLER_8_146 vgnd vpwr scs8hd_decap_4
XFILLER_12_175 vgnd vpwr scs8hd_decap_12
XFILLER_35_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_19.mux_l2_in_0__A1 mux_bottom_track_19.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_37_27 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_11.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_9.mux_l2_in_0_/S
+ mux_bottom_track_11.mux_l1_in_0_/S mem_bottom_track_11.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XANTENNA__67__A _67_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_245 vgnd vpwr scs8hd_decap_12
XFILLER_32_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_23_29 vpwr vgnd scs8hd_fill_2
XFILLER_13_51 vpwr vgnd scs8hd_fill_2
XFILLER_14_215 vgnd vpwr scs8hd_decap_12
XFILLER_1_152 vpwr vgnd scs8hd_fill_2
X_40_ _40_/HI _40_/LO vgnd vpwr scs8hd_conb_1
Xmem_bottom_track_37.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_35.mux_l2_in_0_/S
+ mux_bottom_track_37.mux_l1_in_0_/S mem_bottom_track_37.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_18_18 vpwr vgnd scs8hd_fill_2
XFILLER_1_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_25.scs8hd_buf_4_0__A mux_bottom_track_25.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA__80__A _80_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_211 vgnd vpwr scs8hd_decap_3
XFILLER_6_244 vgnd vpwr scs8hd_decap_12
XFILLER_10_262 vgnd vpwr scs8hd_decap_12
XFILLER_40_93 vgnd vpwr scs8hd_decap_12
XFILLER_34_7 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l2_in_0__S mux_bottom_track_1.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_37_159 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_7.mux_l1_in_1__S mux_bottom_track_7.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_269 vgnd vpwr scs8hd_decap_8
XANTENNA__75__A _75_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_159 vgnd vpwr scs8hd_decap_12
XFILLER_34_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_35.mux_l2_in_0__A0 _25_/HI vgnd vpwr scs8hd_diode_2
XFILLER_25_3 vgnd vpwr scs8hd_decap_12
XFILLER_33_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_25.mux_l2_in_0__S mux_bottom_track_25.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_129 vgnd vpwr scs8hd_decap_12
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_25.mux_l2_in_0__A0 _32_/HI vgnd vpwr scs8hd_diode_2
XFILLER_21_95 vgnd vpwr scs8hd_decap_12
XFILLER_30_154 vgnd vpwr scs8hd_decap_12
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_15_184 vgnd vpwr scs8hd_decap_12
XFILLER_7_53 vpwr vgnd scs8hd_fill_2
XFILLER_7_86 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_19.mux_l1_in_0__S mux_bottom_track_19.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_27.mux_l2_in_0__A1 mux_bottom_track_27.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_37.mux_l1_in_0_ chanx_left_in[19] bottom_left_grid_pin_39_ mux_bottom_track_37.mux_l1_in_0_/S
+ mux_bottom_track_37.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_29_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_39.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_12_110 vpwr vgnd scs8hd_fill_2
XFILLER_12_187 vgnd vpwr scs8hd_decap_12
XFILLER_8_158 vpwr vgnd scs8hd_fill_2
XFILLER_8_169 vpwr vgnd scs8hd_fill_2
XFILLER_35_257 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_1.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_track_1.mux_l2_in_0_/S mux_bottom_track_1.mux_l3_in_0_/S
+ mem_bottom_track_1.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
Xmem_bottom_track_19.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_19.mux_l1_in_0_/S
+ mux_bottom_track_19.mux_l2_in_0_/S mem_bottom_track_19.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_37_39 vgnd vpwr scs8hd_decap_12
XFILLER_26_202 vgnd vpwr scs8hd_decap_12
XFILLER_5_106 vpwr vgnd scs8hd_fill_2
XFILLER_32_227 vgnd vpwr scs8hd_decap_12
XANTENNA__83__A _83_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_257 vgnd vpwr scs8hd_decap_12
XFILLER_4_54 vgnd vpwr scs8hd_decap_3
XFILLER_4_32 vpwr vgnd scs8hd_fill_2
XFILLER_4_10 vpwr vgnd scs8hd_fill_2
XFILLER_14_227 vgnd vpwr scs8hd_decap_12
XFILLER_13_30 vpwr vgnd scs8hd_fill_2
XANTENNA__78__A _78_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_142 vgnd vpwr scs8hd_decap_4
XFILLER_13_85 vpwr vgnd scs8hd_fill_2
XFILLER_38_93 vgnd vpwr scs8hd_decap_12
XFILLER_1_197 vpwr vgnd scs8hd_fill_2
XFILLER_1_175 vpwr vgnd scs8hd_fill_2
XFILLER_9_253 vpwr vgnd scs8hd_fill_2
XFILLER_11_208 vgnd vpwr scs8hd_decap_12
XFILLER_6_256 vgnd vpwr scs8hd_decap_12
XFILLER_10_274 vgnd vpwr scs8hd_fill_1
XFILLER_24_62 vpwr vgnd scs8hd_fill_2
XFILLER_27_7 vpwr vgnd scs8hd_fill_2
XFILLER_1_11 vpwr vgnd scs8hd_fill_2
XFILLER_1_55 vgnd vpwr scs8hd_decap_4
XFILLER_1_66 vgnd vpwr scs8hd_fill_1
XFILLER_28_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_2__D mux_bottom_track_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_204 vpwr vgnd scs8hd_fill_2
XFILLER_10_20 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__D mux_left_track_9.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_27_171 vgnd vpwr scs8hd_decap_12
XFILLER_19_62 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_35.mux_l2_in_0__A1 mux_bottom_track_35.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l2_in_0__S mux_left_track_5.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_196 vgnd vpwr scs8hd_decap_12
XFILLER_31_19 vgnd vpwr scs8hd_decap_12
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_141 vgnd vpwr scs8hd_decap_12
XFILLER_21_30 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_25.mux_l2_in_0__A1 mux_left_track_25.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA__86__A _86_/A vgnd vpwr scs8hd_diode_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_30_166 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_15_196 vgnd vpwr scs8hd_decap_12
XFILLER_26_19 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_12_144 vgnd vpwr scs8hd_decap_8
XFILLER_12_199 vgnd vpwr scs8hd_decap_12
XFILLER_35_269 vgnd vpwr scs8hd_decap_8
Xmem_bottom_track_1.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_1.mux_l1_in_0_/S mux_bottom_track_1.mux_l2_in_0_/S
+ mem_bottom_track_1.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
Xmem_bottom_track_19.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_17.mux_l2_in_0_/S
+ mux_bottom_track_19.mux_l1_in_0_/S mem_bottom_track_19.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_5_118 vpwr vgnd scs8hd_fill_2
XFILLER_5_129 vpwr vgnd scs8hd_fill_2
XFILLER_32_239 vgnd vpwr scs8hd_decap_12
XFILLER_17_269 vgnd vpwr scs8hd_decap_8
XFILLER_27_62 vgnd vpwr scs8hd_decap_12
XFILLER_4_88 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_19.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_1__D mux_bottom_track_3.mux_l1_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_239 vgnd vpwr scs8hd_decap_12
XFILLER_9_243 vgnd vpwr scs8hd_fill_1
XFILLER_34_19 vgnd vpwr scs8hd_decap_12
XFILLER_24_52 vgnd vpwr scs8hd_fill_1
XFILLER_6_268 vgnd vpwr scs8hd_decap_6
XFILLER_10_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_1_34 vpwr vgnd scs8hd_fill_2
XFILLER_28_117 vgnd vpwr scs8hd_decap_12
XFILLER_3_216 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.scs8hd_buf_4_0_ mux_bottom_track_1.mux_l3_in_0_/X _87_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_10_87 vgnd vpwr scs8hd_decap_3
XFILLER_19_74 vgnd vpwr scs8hd_decap_12
XFILLER_35_62 vgnd vpwr scs8hd_decap_12
XFILLER_0_208 vpwr vgnd scs8hd_fill_2
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0__A0 bottom_left_grid_pin_36_ vgnd vpwr scs8hd_diode_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_3.mux_l1_in_1__S mux_bottom_track_3.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_39.mux_l1_in_0__A0 chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_30_178 vgnd vpwr scs8hd_decap_12
Xmem_left_track_25.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_25.mux_l1_in_0_/S ccff_tail
+ mem_left_track_25.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_30_3 vgnd vpwr scs8hd_decap_12
XFILLER_21_123 vgnd vpwr scs8hd_decap_12
XFILLER_29_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__D mux_bottom_track_3.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_21.mux_l2_in_0__S mux_bottom_track_21.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_127 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_21.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.scs8hd_dfxbp_1_0_ prog_clk ccff_head mux_bottom_track_1.mux_l1_in_0_/S
+ mem_bottom_track_1.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_1.mux_l1_in_2__A0 chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_7_193 vpwr vgnd scs8hd_fill_2
XFILLER_26_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_15.mux_l1_in_0__S mux_bottom_track_15.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_40_251 vgnd vpwr scs8hd_decap_12
XFILLER_27_74 vgnd vpwr scs8hd_decap_12
XFILLER_4_163 vpwr vgnd scs8hd_fill_2
XFILLER_4_67 vpwr vgnd scs8hd_fill_2
XFILLER_4_23 vpwr vgnd scs8hd_fill_2
XFILLER_22_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l2_in_1__A0 _35_/HI vgnd vpwr scs8hd_diode_2
XFILLER_8_3 vgnd vpwr scs8hd_decap_4
XFILLER_9_222 vgnd vpwr scs8hd_decap_12
XFILLER_10_232 vgnd vpwr scs8hd_decap_3
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
Xmux_left_track_5.scs8hd_buf_4_0_ mux_left_track_5.mux_l2_in_0_/X _65_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mem_bottom_track_23.scs8hd_dfxbp_1_1__D mux_bottom_track_23.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l3_in_0__A0 mux_bottom_track_1.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_239 vgnd vpwr scs8hd_decap_4
XFILLER_3_228 vgnd vpwr scs8hd_decap_4
XFILLER_10_66 vpwr vgnd scs8hd_fill_2
XFILLER_19_42 vgnd vpwr scs8hd_decap_12
XFILLER_35_74 vgnd vpwr scs8hd_decap_12
XFILLER_27_184 vgnd vpwr scs8hd_decap_12
XFILLER_19_86 vgnd vpwr scs8hd_decap_12
XFILLER_42_187 vgnd vpwr scs8hd_decap_12
XFILLER_32_7 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_37.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_33_110 vgnd vpwr scs8hd_decap_12
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_3.mux_l1_in_0__A1 bottom_left_grid_pin_34_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_39.mux_l1_in_0__A1 bottom_left_grid_pin_40_ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_19.scs8hd_buf_4_0_ mux_bottom_track_19.mux_l2_in_0_/X _78_/A vgnd
+ vpwr scs8hd_buf_1
XPHY_7 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_33.scs8hd_buf_4_0__A mux_bottom_track_33.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_25.scs8hd_dfxbp_1_0_ prog_clk mux_left_track_9.mux_l2_in_0_/S mux_left_track_25.mux_l1_in_0_/S
+ mem_left_track_25.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_38_202 vgnd vpwr scs8hd_decap_12
XFILLER_23_3 vpwr vgnd scs8hd_fill_2
XFILLER_21_135 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l2_in_0__S mux_left_track_1.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_257 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_9.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_9.mux_l1_in_0_/S mux_bottom_track_9.mux_l2_in_0_/S
+ mem_bottom_track_9.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_12_102 vpwr vgnd scs8hd_fill_2
XFILLER_16_32 vpwr vgnd scs8hd_fill_2
XFILLER_8_106 vpwr vgnd scs8hd_fill_2
XFILLER_20_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_2__A1 bottom_left_grid_pin_41_ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_5.mux_l3_in_0_ mux_bottom_track_5.mux_l2_in_1_/X mux_bottom_track_5.mux_l2_in_0_/X
+ mux_bottom_track_5.mux_l3_in_0_/S mux_bottom_track_5.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_41_208 vgnd vpwr scs8hd_decap_12
XFILLER_26_227 vgnd vpwr scs8hd_decap_12
XFILLER_27_86 vgnd vpwr scs8hd_decap_12
XFILLER_40_263 vgnd vpwr scs8hd_decap_12
XFILLER_4_186 vpwr vgnd scs8hd_fill_2
XFILLER_23_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__D mux_bottom_track_23.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_11 vgnd vpwr scs8hd_decap_3
XFILLER_22_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_2__D mux_bottom_track_7.mux_l2_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_55 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.mux_l2_in_1__A1 mux_bottom_track_1.mux_l1_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_1_101 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_5.mux_l2_in_1_ _28_/HI mux_bottom_track_5.mux_l1_in_2_/X mux_bottom_track_5.mux_l2_in_0_/S
+ mux_bottom_track_5.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_9_234 vgnd vpwr scs8hd_fill_1
XFILLER_39_171 vgnd vpwr scs8hd_decap_12
XFILLER_6_215 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_27.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_27.mux_l1_in_0_/S
+ mux_bottom_track_27.mux_l2_in_0_/S mem_bottom_track_27.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_24_32 vpwr vgnd scs8hd_fill_2
XFILLER_36_141 vgnd vpwr scs8hd_decap_12
X_79_ _79_/A chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_1.mux_l3_in_0__A1 mux_bottom_track_1.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_5.mux_l1_in_2_ chanx_left_in[3] bottom_left_grid_pin_41_ mux_bottom_track_5.mux_l1_in_1_/S
+ mux_bottom_track_5.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
Xmux_bottom_track_27.scs8hd_buf_4_0_ mux_bottom_track_27.mux_l2_in_0_/X _74_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_10_12 vpwr vgnd scs8hd_fill_2
XFILLER_19_21 vpwr vgnd scs8hd_fill_2
XFILLER_19_54 vgnd vpwr scs8hd_decap_6
XFILLER_19_98 vgnd vpwr scs8hd_decap_12
XFILLER_35_86 vgnd vpwr scs8hd_decap_12
XFILLER_35_31 vgnd vpwr scs8hd_decap_12
XFILLER_27_196 vgnd vpwr scs8hd_decap_12
XFILLER_42_199 vgnd vpwr scs8hd_decap_12
XFILLER_2_240 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_13.mux_l1_in_0__A0 chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_166 vgnd vpwr scs8hd_decap_12
XFILLER_21_11 vpwr vgnd scs8hd_fill_2
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_15_111 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_5.scs8hd_buf_4_0__A mux_left_track_5.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_57 vpwr vgnd scs8hd_fill_2
XFILLER_16_3 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_19.mux_l2_in_0_ _40_/HI mux_bottom_track_19.mux_l1_in_0_/X mux_bottom_track_19.mux_l2_in_0_/S
+ mux_bottom_track_19.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_21_147 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_29_269 vgnd vpwr scs8hd_decap_8
Xmem_bottom_track_9.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_7.mux_l3_in_0_/S mux_bottom_track_9.mux_l1_in_0_/S
+ mem_bottom_track_9.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_12_114 vgnd vpwr scs8hd_decap_6
XFILLER_16_55 vgnd vpwr scs8hd_decap_12
XFILLER_32_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__D mux_bottom_track_9.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_21.mux_l2_in_0_ _41_/HI mux_bottom_track_21.mux_l1_in_0_/X mux_bottom_track_21.mux_l2_in_0_/S
+ mux_bottom_track_21.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_26_239 vgnd vpwr scs8hd_decap_12
XFILLER_27_98 vgnd vpwr scs8hd_decap_12
XFILLER_4_143 vpwr vgnd scs8hd_fill_2
XFILLER_31_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_0__S mux_bottom_track_9.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_34 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_11.mux_l1_in_0__S mux_bottom_track_11.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_89 vpwr vgnd scs8hd_fill_2
XFILLER_1_179 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_5.mux_l2_in_0_ mux_bottom_track_5.mux_l1_in_1_/X mux_bottom_track_5.mux_l1_in_0_/X
+ mux_bottom_track_5.mux_l2_in_0_/S mux_bottom_track_5.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_13_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_39.mux_l2_in_0__S mux_bottom_track_39.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_257 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_35.scs8hd_buf_4_0_ mux_bottom_track_35.mux_l2_in_0_/X _70_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_27.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_25.mux_l2_in_0_/S
+ mux_bottom_track_27.mux_l1_in_0_/S mem_bottom_track_27.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_24_66 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_1__A0 bottom_left_grid_pin_39_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_21.mux_l1_in_0__A0 chanx_left_in[11] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_15.scs8hd_buf_4_0__A mux_bottom_track_15.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
X_78_ _78_/A chany_bottom_out[9] vgnd vpwr scs8hd_buf_2
Xmux_bottom_track_5.mux_l1_in_1_ bottom_left_grid_pin_39_ bottom_left_grid_pin_37_
+ mux_bottom_track_5.mux_l1_in_1_/S mux_bottom_track_5.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_10_24 vpwr vgnd scs8hd_fill_2
XFILLER_10_35 vpwr vgnd scs8hd_fill_2
XFILLER_10_79 vpwr vgnd scs8hd_fill_2
XFILLER_42_156 vgnd vpwr scs8hd_decap_12
XFILLER_35_98 vgnd vpwr scs8hd_decap_12
XFILLER_35_43 vgnd vpwr scs8hd_decap_12
XFILLER_2_274 vgnd vpwr scs8hd_fill_1
XFILLER_33_123 vgnd vpwr scs8hd_decap_12
XFILLER_18_7 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_13.mux_l1_in_0__A1 bottom_left_grid_pin_35_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0__A0 mux_bottom_track_5.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_178 vgnd vpwr scs8hd_decap_12
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_15_123 vgnd vpwr scs8hd_decap_12
XFILLER_38_215 vgnd vpwr scs8hd_decap_12
XFILLER_21_159 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l1_in_0__A0 left_top_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XFILLER_16_23 vgnd vpwr scs8hd_decap_6
XFILLER_32_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_7.mux_l3_in_0__S mux_bottom_track_7.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_16_67 vgnd vpwr scs8hd_decap_12
XFILLER_7_152 vpwr vgnd scs8hd_fill_2
XFILLER_34_251 vgnd vpwr scs8hd_decap_12
XFILLER_27_11 vgnd vpwr scs8hd_decap_4
XFILLER_27_22 vgnd vpwr scs8hd_decap_12
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
XFILLER_4_122 vpwr vgnd scs8hd_fill_2
XFILLER_4_59 vgnd vpwr scs8hd_decap_3
XFILLER_4_37 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_19.mux_l1_in_0_ chanx_left_in[10] bottom_left_grid_pin_38_ mux_bottom_track_19.mux_l1_in_0_/S
+ mux_bottom_track_19.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_31_232 vgnd vpwr scs8hd_decap_12
XFILLER_16_251 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_21.mux_l1_in_0_ chanx_left_in[11] bottom_left_grid_pin_39_ mux_bottom_track_21.mux_l1_in_0_/S
+ mux_bottom_track_21.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_bottom_track_29.scs8hd_dfxbp_1_1__D mux_bottom_track_29.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_1_114 vpwr vgnd scs8hd_fill_2
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XFILLER_9_203 vgnd vpwr scs8hd_decap_8
XFILLER_9_214 vpwr vgnd scs8hd_fill_2
XFILLER_13_232 vgnd vpwr scs8hd_decap_12
XFILLER_9_269 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_33.mux_l2_in_0_ _24_/HI mux_bottom_track_33.mux_l1_in_0_/X mux_bottom_track_33.mux_l2_in_0_/S
+ mux_bottom_track_33.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_39_184 vgnd vpwr scs8hd_decap_12
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_1__A1 bottom_left_grid_pin_37_ vgnd vpwr scs8hd_diode_2
XFILLER_10_213 vgnd vpwr scs8hd_fill_1
XFILLER_24_78 vgnd vpwr scs8hd_decap_12
XFILLER_6_3 vgnd vpwr scs8hd_fill_1
XFILLER_1_38 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_21.mux_l1_in_0__A1 bottom_left_grid_pin_39_ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_36_154 vgnd vpwr scs8hd_decap_12
X_77_ _77_/A chany_bottom_out[10] vgnd vpwr scs8hd_buf_2
Xmux_bottom_track_5.mux_l1_in_0_ bottom_left_grid_pin_35_ bottom_right_grid_pin_1_
+ mux_bottom_track_5.mux_l1_in_1_/S mux_bottom_track_5.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_3.scs8hd_buf_4_0__A mux_bottom_track_3.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_27_110 vgnd vpwr scs8hd_decap_12
XFILLER_42_168 vgnd vpwr scs8hd_decap_12
XFILLER_35_55 vgnd vpwr scs8hd_decap_6
XFILLER_33_135 vgnd vpwr scs8hd_decap_12
XFILLER_18_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l2_in_0__A1 mux_bottom_track_5.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_2_81 vpwr vgnd scs8hd_fill_2
XFILLER_32_190 vgnd vpwr scs8hd_decap_12
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_57 vpwr vgnd scs8hd_fill_2
XFILLER_15_135 vgnd vpwr scs8hd_decap_12
XFILLER_30_105 vgnd vpwr scs8hd_decap_12
XFILLER_7_26 vpwr vgnd scs8hd_fill_2
XFILLER_38_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l1_in_0__A1 chany_bottom_in[19] vgnd vpwr scs8hd_diode_2
XFILLER_32_56 vgnd vpwr scs8hd_decap_12
XFILLER_16_79 vgnd vpwr scs8hd_decap_12
XFILLER_35_208 vgnd vpwr scs8hd_decap_12
XFILLER_7_142 vpwr vgnd scs8hd_fill_2
XFILLER_7_175 vpwr vgnd scs8hd_fill_2
XFILLER_7_197 vpwr vgnd scs8hd_fill_2
XFILLER_11_182 vgnd vpwr scs8hd_fill_1
XFILLER_34_263 vgnd vpwr scs8hd_decap_12
XFILLER_17_208 vgnd vpwr scs8hd_decap_12
XFILLER_27_34 vgnd vpwr scs8hd_decap_12
XFILLER_4_112 vgnd vpwr scs8hd_fill_1
XFILLER_4_167 vpwr vgnd scs8hd_fill_2
XFILLER_4_27 vpwr vgnd scs8hd_fill_2
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_263 vgnd vpwr scs8hd_decap_12
XFILLER_1_148 vpwr vgnd scs8hd_fill_2
XFILLER_38_44 vgnd vpwr scs8hd_decap_12
XFILLER_9_237 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_39_196 vgnd vpwr scs8hd_decap_12
XFILLER_40_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_0__S mux_bottom_track_5.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
X_76_ _76_/A chany_bottom_out[11] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_35.mux_l2_in_0__S mux_bottom_track_35.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_166 vgnd vpwr scs8hd_decap_12
XFILLER_42_125 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_33.mux_l1_in_0_ chanx_left_in[17] bottom_left_grid_pin_37_ mux_bottom_track_33.mux_l1_in_0_/S
+ mux_bottom_track_33.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_15.mux_l2_in_0__A0 _38_/HI vgnd vpwr scs8hd_diode_2
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_147 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_7.scs8hd_buf_4_0_ mux_bottom_track_7.mux_l3_in_0_/X _84_/A vgnd
+ vpwr scs8hd_buf_1
XANTENNA_mux_bottom_track_29.mux_l1_in_0__S mux_bottom_track_29.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_166 vgnd vpwr scs8hd_decap_12
X_59_ chany_bottom_in[7] chanx_left_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_2_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_13.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_117 vgnd vpwr scs8hd_decap_12
XFILLER_15_147 vgnd vpwr scs8hd_decap_12
XFILLER_23_7 vgnd vpwr scs8hd_decap_6
XFILLER_38_239 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_35.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_35.mux_l1_in_0_/S
+ mux_bottom_track_35.mux_l2_in_0_/S mem_bottom_track_35.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_14_191 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A0 bottom_left_grid_pin_41_ vgnd vpwr scs8hd_diode_2
XFILLER_12_106 vpwr vgnd scs8hd_fill_2
XFILLER_32_68 vgnd vpwr scs8hd_decap_12
XFILLER_12_139 vgnd vpwr scs8hd_decap_3
XFILLER_11_161 vpwr vgnd scs8hd_fill_2
XFILLER_22_90 vpwr vgnd scs8hd_fill_2
XFILLER_14_3 vpwr vgnd scs8hd_fill_2
XFILLER_27_46 vgnd vpwr scs8hd_decap_12
XFILLER_25_220 vgnd vpwr scs8hd_decap_12
XFILLER_4_102 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_3.mux_l3_in_0__S mux_bottom_track_3.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_245 vgnd vpwr scs8hd_decap_12
XFILLER_38_56 vgnd vpwr scs8hd_decap_12
XFILLER_9_249 vpwr vgnd scs8hd_fill_2
XFILLER_13_245 vgnd vpwr scs8hd_decap_12
XFILLER_0_182 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_7.mux_l2_in_1__A0 _29_/HI vgnd vpwr scs8hd_diode_2
XFILLER_5_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_23.mux_l2_in_0__A0 _42_/HI vgnd vpwr scs8hd_diode_2
XFILLER_10_215 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_29.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_24_36 vgnd vpwr scs8hd_decap_12
XFILLER_40_68 vgnd vpwr scs8hd_decap_12
XFILLER_36_178 vgnd vpwr scs8hd_decap_12
X_75_ _75_/A chany_bottom_out[12] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_bottom_track_11.scs8hd_dfxbp_1_1__D mux_bottom_track_11.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_16 vpwr vgnd scs8hd_fill_2
XFILLER_19_25 vpwr vgnd scs8hd_fill_2
XFILLER_42_137 vgnd vpwr scs8hd_decap_12
XFILLER_27_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_15.mux_l2_in_0__A1 mux_bottom_track_15.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_2_244 vgnd vpwr scs8hd_decap_12
XFILLER_2_222 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_7.mux_l3_in_0__A0 mux_bottom_track_7.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_33_159 vgnd vpwr scs8hd_decap_12
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_bottom_track_31.scs8hd_dfxbp_1_1__D mux_bottom_track_31.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_178 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0__S mux_left_track_9.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
X_58_ chany_bottom_in[8] chanx_left_out[9] vgnd vpwr scs8hd_buf_2
XFILLER_21_15 vgnd vpwr scs8hd_decap_12
XFILLER_30_129 vgnd vpwr scs8hd_decap_12
XFILLER_15_159 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_35.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_33.mux_l2_in_0_/S
+ mux_bottom_track_35.mux_l1_in_0_/S mem_bottom_track_35.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_21_107 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A1 bottom_right_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_23.scs8hd_buf_4_0__A mux_bottom_track_23.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_15 vgnd vpwr scs8hd_decap_4
XFILLER_28_251 vgnd vpwr scs8hd_decap_12
XFILLER_11_184 vgnd vpwr scs8hd_decap_12
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
Xmux_left_track_9.mux_l2_in_0_ _34_/HI mux_left_track_9.mux_l1_in_0_/X mux_left_track_9.mux_l2_in_0_/S
+ mux_left_track_9.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_8_82 vpwr vgnd scs8hd_fill_2
XFILLER_8_93 vpwr vgnd scs8hd_fill_2
XFILLER_25_232 vgnd vpwr scs8hd_decap_12
XFILLER_27_58 vgnd vpwr scs8hd_decap_3
XFILLER_40_202 vgnd vpwr scs8hd_decap_12
XFILLER_4_147 vgnd vpwr scs8hd_decap_4
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_31.mux_l2_in_0__A0 _47_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_31.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_13_16 vgnd vpwr scs8hd_decap_3
XFILLER_13_38 vpwr vgnd scs8hd_fill_2
XFILLER_22_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_13.scs8hd_dfxbp_1_0__D mux_bottom_track_11.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_68 vgnd vpwr scs8hd_decap_12
XFILLER_8_9 vpwr vgnd scs8hd_fill_2
XFILLER_13_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_0__D mux_bottom_track_31.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_272 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_7.mux_l2_in_1__A1 chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_39_110 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_23.mux_l2_in_0__A1 mux_bottom_track_23.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_24_48 vgnd vpwr scs8hd_decap_4
XFILLER_5_220 vpwr vgnd scs8hd_fill_2
XFILLER_5_231 vpwr vgnd scs8hd_fill_2
XFILLER_30_80 vgnd vpwr scs8hd_decap_12
X_74_ _74_/A chany_bottom_out[13] vgnd vpwr scs8hd_buf_2
Xmem_bottom_track_17.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_17.mux_l1_in_0_/S
+ mux_bottom_track_17.mux_l2_in_0_/S mem_bottom_track_17.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_10_28 vgnd vpwr scs8hd_decap_3
XFILLER_10_39 vpwr vgnd scs8hd_fill_2
XFILLER_27_135 vgnd vpwr scs8hd_decap_12
XFILLER_42_149 vgnd vpwr scs8hd_decap_6
XFILLER_2_256 vgnd vpwr scs8hd_decap_12
XFILLER_2_234 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_7.mux_l3_in_0__A1 mux_bottom_track_7.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_41_171 vgnd vpwr scs8hd_decap_12
XPHY_80 vgnd vpwr scs8hd_decap_3
XFILLER_26_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_0__S mux_bottom_track_1.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_57_ chany_bottom_in[9] chanx_left_out[10] vgnd vpwr scs8hd_buf_2
XFILLER_24_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__D mux_bottom_track_39.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_27 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_31.mux_l2_in_0__S mux_bottom_track_31.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_19.mux_l1_in_0__A0 chanx_left_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_23_171 vgnd vpwr scs8hd_decap_12
XANTENNA__51__A chany_bottom_in[15] vgnd vpwr scs8hd_diode_2
XFILLER_21_119 vgnd vpwr scs8hd_decap_3
XFILLER_29_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_25.mux_l1_in_0__S mux_bottom_track_25.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_20_141 vgnd vpwr scs8hd_decap_12
XFILLER_28_263 vgnd vpwr scs8hd_decap_12
XFILLER_11_174 vpwr vgnd scs8hd_fill_2
XFILLER_11_196 vgnd vpwr scs8hd_decap_12
XFILLER_22_70 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_4_126 vpwr vgnd scs8hd_fill_2
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_269 vgnd vpwr scs8hd_decap_8
XFILLER_3_192 vpwr vgnd scs8hd_fill_2
XFILLER_3_170 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_31.mux_l2_in_0__A1 mux_bottom_track_31.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_1_118 vpwr vgnd scs8hd_fill_2
XFILLER_9_218 vpwr vgnd scs8hd_fill_2
XFILLER_13_269 vgnd vpwr scs8hd_decap_8
XFILLER_0_151 vpwr vgnd scs8hd_fill_2
XFILLER_0_162 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l1_in_0_ left_top_grid_pin_1_ chany_bottom_in[3] mux_left_track_9.mux_l1_in_0_/S
+ mux_left_track_9.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_28_80 vgnd vpwr scs8hd_decap_12
XFILLER_10_239 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_track_11.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA__54__A chany_bottom_in[12] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l2_in_1__S mux_bottom_track_5.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_5_243 vgnd vpwr scs8hd_fill_1
XFILLER_39_7 vpwr vgnd scs8hd_fill_2
X_73_ _73_/A chany_bottom_out[14] vgnd vpwr scs8hd_buf_2
Xmem_bottom_track_17.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_15.mux_l2_in_0_/S
+ mux_bottom_track_17.mux_l1_in_0_/S mem_bottom_track_17.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_27_147 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_27.mux_l1_in_0__A0 chanx_left_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_19_38 vpwr vgnd scs8hd_fill_2
XFILLER_42_106 vgnd vpwr scs8hd_decap_12
XFILLER_2_202 vpwr vgnd scs8hd_fill_2
XANTENNA__49__A chany_bottom_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_2_268 vgnd vpwr scs8hd_decap_6
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_25_81 vgnd vpwr scs8hd_decap_12
X_56_ chany_bottom_in[10] chanx_left_out[11] vgnd vpwr scs8hd_buf_2
Xmux_bottom_track_1.mux_l3_in_0_ mux_bottom_track_1.mux_l2_in_1_/X mux_bottom_track_1.mux_l2_in_0_/X
+ mux_bottom_track_1.mux_l3_in_0_/S mux_bottom_track_1.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_2_85 vpwr vgnd scs8hd_fill_2
XFILLER_2_41 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_17.mux_l2_in_0__S mux_bottom_track_17.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_24_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_19.mux_l1_in_0__A1 bottom_left_grid_pin_38_ vgnd vpwr scs8hd_diode_2
XFILLER_11_50 vgnd vpwr scs8hd_decap_8
XFILLER_36_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_5.mux_l1_in_0__S mux_left_track_5.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_220 vgnd vpwr scs8hd_decap_12
X_39_ _39_/HI _39_/LO vgnd vpwr scs8hd_conb_1
Xmux_bottom_track_1.mux_l2_in_1_ _35_/HI mux_bottom_track_1.mux_l1_in_2_/X mux_bottom_track_1.mux_l2_in_0_/S
+ mux_bottom_track_1.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_7_146 vgnd vpwr scs8hd_decap_4
XFILLER_7_179 vpwr vgnd scs8hd_fill_2
XFILLER_22_82 vgnd vpwr scs8hd_decap_8
XFILLER_22_93 vgnd vpwr scs8hd_decap_12
XANTENNA__62__A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_19_220 vgnd vpwr scs8hd_decap_12
XFILLER_21_7 vpwr vgnd scs8hd_fill_2
XFILLER_8_40 vgnd vpwr scs8hd_decap_3
XFILLER_40_215 vgnd vpwr scs8hd_decap_12
XFILLER_25_245 vgnd vpwr scs8hd_decap_12
XANTENNA__57__A chany_bottom_in[9] vgnd vpwr scs8hd_diode_2
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_60 vgnd vpwr scs8hd_fill_1
XFILLER_3_182 vgnd vpwr scs8hd_fill_1
XFILLER_12_3 vpwr vgnd scs8hd_fill_2
XFILLER_22_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_2_ chanx_left_in[1] bottom_left_grid_pin_41_ mux_bottom_track_1.mux_l1_in_0_/S
+ mux_bottom_track_1.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_1__D mux_bottom_track_17.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_196 vgnd vpwr scs8hd_decap_4
Xmem_left_track_5.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_5.mux_l1_in_0_/S mux_left_track_5.mux_l2_in_0_/S
+ mem_left_track_5.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_8_252 vgnd vpwr scs8hd_decap_12
XFILLER_39_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_37.scs8hd_dfxbp_1_1__D mux_bottom_track_37.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_35.mux_l1_in_0__A0 chanx_left_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_10_207 vgnd vpwr scs8hd_decap_6
Xmem_bottom_track_7.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_track_7.mux_l2_in_1_/S mux_bottom_track_7.mux_l3_in_0_/S
+ mem_bottom_track_7.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA__70__A _70_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_93 vgnd vpwr scs8hd_decap_12
X_72_ _72_/A chany_bottom_out[15] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_track_25.mux_l1_in_0__A0 left_top_grid_pin_1_ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_15.mux_l2_in_0_ _38_/HI mux_bottom_track_15.mux_l1_in_0_/X mux_bottom_track_15.mux_l2_in_0_/S
+ mux_bottom_track_15.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_42_118 vgnd vpwr scs8hd_decap_6
XFILLER_27_159 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_27.mux_l1_in_0__A1 bottom_left_grid_pin_34_ vgnd vpwr scs8hd_diode_2
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_18_137 vgnd vpwr scs8hd_decap_12
XANTENNA__65__A _65_/A vgnd vpwr scs8hd_diode_2
XFILLER_41_184 vgnd vpwr scs8hd_decap_12
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_25_93 vgnd vpwr scs8hd_decap_12
X_55_ _55_/A chanx_left_out[12] vgnd vpwr scs8hd_buf_2
XFILLER_24_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__D mux_left_track_5.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_184 vgnd vpwr scs8hd_decap_12
XFILLER_11_73 vpwr vgnd scs8hd_fill_2
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_232 vgnd vpwr scs8hd_decap_12
X_38_ _38_/HI _38_/LO vgnd vpwr scs8hd_conb_1
XFILLER_20_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_19.scs8hd_dfxbp_1_0__D mux_bottom_track_17.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
XFILLER_11_132 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l2_in_0_ mux_bottom_track_1.mux_l1_in_1_/X mux_bottom_track_1.mux_l1_in_0_/X
+ mux_bottom_track_1.mux_l2_in_0_/S mux_bottom_track_1.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_7_114 vpwr vgnd scs8hd_fill_2
XFILLER_11_165 vpwr vgnd scs8hd_fill_2
XFILLER_34_202 vgnd vpwr scs8hd_decap_12
XFILLER_14_7 vpwr vgnd scs8hd_fill_2
XFILLER_19_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_39.scs8hd_dfxbp_1_0__D mux_bottom_track_37.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.scs8hd_buf_4_0_ mux_left_track_1.mux_l2_in_0_/X _67_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_40_227 vgnd vpwr scs8hd_decap_12
XFILLER_25_257 vgnd vpwr scs8hd_decap_12
XFILLER_4_139 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_21.mux_l1_in_0__S mux_bottom_track_21.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_16_202 vgnd vpwr scs8hd_decap_12
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__73__A _73_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_227 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.mux_l1_in_1_ bottom_left_grid_pin_39_ bottom_left_grid_pin_37_
+ mux_bottom_track_1.mux_l1_in_0_/S mux_bottom_track_1.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA__68__A _68_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_175 vgnd vpwr scs8hd_decap_4
XFILLER_0_120 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_31.scs8hd_buf_4_0__A mux_bottom_track_31.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_93 vgnd vpwr scs8hd_decap_12
Xmem_left_track_5.scs8hd_dfxbp_1_0_ prog_clk mux_left_track_1.mux_l2_in_0_/S mux_left_track_5.mux_l1_in_0_/S
+ mem_left_track_5.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_8_264 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_15.scs8hd_buf_4_0_ mux_bottom_track_15.mux_l2_in_0_/X _80_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_5_53 vgnd vpwr scs8hd_decap_4
XFILLER_5_75 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_35.mux_l1_in_0__A1 bottom_left_grid_pin_38_ vgnd vpwr scs8hd_diode_2
XFILLER_39_135 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_7.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_7.mux_l1_in_1_/S mux_bottom_track_7.mux_l2_in_1_/S
+ mem_bottom_track_7.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_38_190 vgnd vpwr scs8hd_decap_12
XFILLER_14_40 vpwr vgnd scs8hd_fill_2
XFILLER_5_245 vgnd vpwr scs8hd_decap_12
XFILLER_36_105 vgnd vpwr scs8hd_decap_12
X_71_ _71_/A chany_bottom_out[16] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_track_25.mux_l1_in_0__A1 chany_bottom_in[11] vgnd vpwr scs8hd_diode_2
XFILLER_35_171 vgnd vpwr scs8hd_decap_12
XFILLER_4_6 vpwr vgnd scs8hd_fill_2
XFILLER_18_105 vgnd vpwr scs8hd_decap_12
XFILLER_18_149 vgnd vpwr scs8hd_decap_4
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XANTENNA__81__A _81_/A vgnd vpwr scs8hd_diode_2
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_50 vgnd vpwr scs8hd_decap_3
XFILLER_41_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l2_in_1__S mux_bottom_track_1.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_2_32 vpwr vgnd scs8hd_fill_2
X_54_ chany_bottom_in[12] chanx_left_out[13] vgnd vpwr scs8hd_buf_2
XFILLER_2_54 vpwr vgnd scs8hd_fill_2
XFILLER_32_141 vgnd vpwr scs8hd_decap_12
XFILLER_15_119 vgnd vpwr scs8hd_decap_3
XFILLER_23_196 vgnd vpwr scs8hd_decap_12
XFILLER_2_3 vgnd vpwr scs8hd_fill_1
XFILLER_11_96 vpwr vgnd scs8hd_fill_2
XANTENNA__76__A _76_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_93 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_15.mux_l1_in_0_ chanx_left_in[8] bottom_left_grid_pin_36_ mux_bottom_track_15.mux_l1_in_0_/S
+ mux_bottom_track_15.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_14_141 vgnd vpwr scs8hd_decap_12
XFILLER_35_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
X_37_ _37_/HI _37_/LO vgnd vpwr scs8hd_conb_1
XFILLER_16_19 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_27.mux_l2_in_0_ _44_/HI mux_bottom_track_27.mux_l1_in_0_/X mux_bottom_track_27.mux_l2_in_0_/S
+ mux_bottom_track_27.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_20_166 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_13.mux_l2_in_0__S mux_bottom_track_13.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_bottom_track_25.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_25.mux_l1_in_1_/S
+ mux_bottom_track_25.mux_l2_in_0_/S mem_bottom_track_25.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_11_100 vpwr vgnd scs8hd_fill_2
XFILLER_8_86 vgnd vpwr scs8hd_decap_4
XFILLER_6_192 vgnd vpwr scs8hd_decap_4
XFILLER_27_18 vpwr vgnd scs8hd_fill_2
XFILLER_40_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l1_in_0__S mux_left_track_1.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__D ccff_head vgnd vpwr scs8hd_diode_2
XFILLER_25_269 vgnd vpwr scs8hd_decap_8
XFILLER_17_62 vgnd vpwr scs8hd_decap_12
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_23.scs8hd_buf_4_0_ mux_bottom_track_23.mux_l2_in_0_/X _76_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_22_239 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.mux_l1_in_0_ bottom_left_grid_pin_35_ bottom_right_grid_pin_1_
+ mux_bottom_track_1.mux_l1_in_0_/S mux_bottom_track_1.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA__84__A _84_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
XFILLER_5_43 vpwr vgnd scs8hd_fill_2
XFILLER_5_98 vpwr vgnd scs8hd_fill_2
XFILLER_39_147 vgnd vpwr scs8hd_decap_12
XFILLER_24_19 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_7.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_5.mux_l3_in_0_/S mux_bottom_track_7.mux_l1_in_1_/S
+ mem_bottom_track_7.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_5_213 vpwr vgnd scs8hd_fill_2
XFILLER_5_224 vgnd vpwr scs8hd_decap_4
XFILLER_5_235 vgnd vpwr scs8hd_decap_8
XFILLER_14_96 vgnd vpwr scs8hd_decap_8
XANTENNA__79__A _79_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_257 vgnd vpwr scs8hd_decap_12
XFILLER_36_117 vgnd vpwr scs8hd_decap_12
X_70_ _70_/A chany_bottom_out[17] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_29.mux_l2_in_0__A0 _45_/HI vgnd vpwr scs8hd_diode_2
XFILLER_18_117 vgnd vpwr scs8hd_fill_1
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_37_7 vpwr vgnd scs8hd_fill_2
X_53_ chany_bottom_in[13] chanx_left_out[14] vgnd vpwr scs8hd_buf_2
XFILLER_2_44 vgnd vpwr scs8hd_fill_1
XFILLER_11_20 vgnd vpwr scs8hd_decap_4
XFILLER_37_245 vgnd vpwr scs8hd_decap_12
X_36_ _36_/HI _36_/LO vgnd vpwr scs8hd_conb_1
XFILLER_32_19 vgnd vpwr scs8hd_decap_12
XFILLER_20_178 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l2_in_0__A0 _34_/HI vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_25.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_23.mux_l2_in_0_/S
+ mux_bottom_track_25.mux_l1_in_1_/S mem_bottom_track_25.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
Xmux_bottom_track_31.scs8hd_buf_4_0_ mux_bottom_track_31.mux_l2_in_0_/X _72_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_11_178 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_23.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA__87__A _87_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_245 vgnd vpwr scs8hd_decap_12
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_13.scs8hd_buf_4_0__A mux_bottom_track_13.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1__A0 bottom_left_grid_pin_39_ vgnd vpwr scs8hd_diode_2
XFILLER_8_32 vpwr vgnd scs8hd_fill_2
XFILLER_8_65 vpwr vgnd scs8hd_fill_2
XFILLER_4_108 vpwr vgnd scs8hd_fill_2
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_215 vgnd vpwr scs8hd_decap_12
XFILLER_17_74 vgnd vpwr scs8hd_decap_12
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_62 vgnd vpwr scs8hd_decap_12
XFILLER_3_174 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_27.mux_l1_in_0_ chanx_left_in[14] bottom_left_grid_pin_34_ mux_bottom_track_27.mux_l1_in_0_/S
+ mux_bottom_track_27.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_30_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_39.scs8hd_buf_4_0__A mux_bottom_track_39.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_39.mux_l2_in_0_ _27_/HI mux_bottom_track_39.mux_l1_in_0_/X mux_bottom_track_39.mux_l2_in_0_/S
+ mux_bottom_track_39.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_37.mux_l2_in_0__A0 _26_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0__A0 mux_bottom_track_1.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_233 vgnd vpwr scs8hd_decap_12
XFILLER_39_159 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_21.scs8hd_dfxbp_1_0__D mux_bottom_track_19.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_19 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_2__D mux_bottom_track_3.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_269 vgnd vpwr scs8hd_decap_8
XFILLER_14_64 vpwr vgnd scs8hd_fill_2
XFILLER_36_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_39.mux_l1_in_0__S mux_bottom_track_39.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_29.mux_l2_in_0__A1 mux_bottom_track_29.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_35_184 vgnd vpwr scs8hd_decap_12
XFILLER_35_19 vgnd vpwr scs8hd_decap_12
XFILLER_2_206 vgnd vpwr scs8hd_decap_8
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_110 vgnd vpwr scs8hd_decap_12
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_41 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
X_52_ chany_bottom_in[14] chanx_left_out[15] vgnd vpwr scs8hd_buf_2
XFILLER_2_89 vgnd vpwr scs8hd_decap_3
XFILLER_2_23 vpwr vgnd scs8hd_fill_2
XFILLER_1_261 vgnd vpwr scs8hd_decap_12
XFILLER_32_154 vgnd vpwr scs8hd_decap_12
XFILLER_17_151 vgnd vpwr scs8hd_decap_12
XFILLER_17_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_37.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_23_121 vgnd vpwr scs8hd_fill_1
XFILLER_11_65 vpwr vgnd scs8hd_fill_2
XFILLER_14_154 vgnd vpwr scs8hd_decap_12
XFILLER_37_257 vgnd vpwr scs8hd_decap_12
X_35_ _35_/HI _35_/LO vgnd vpwr scs8hd_conb_1
XFILLER_28_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l2_in_0__A1 mux_left_track_9.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_113 vgnd vpwr scs8hd_decap_3
XFILLER_19_257 vgnd vpwr scs8hd_decap_12
XFILLER_34_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_1__A1 bottom_left_grid_pin_37_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.scs8hd_buf_4_0__A mux_bottom_track_1.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__D mux_bottom_track_5.mux_l1_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_7.mux_l2_in_0__S mux_bottom_track_7.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_208 vgnd vpwr scs8hd_decap_12
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_227 vgnd vpwr scs8hd_decap_12
XFILLER_17_86 vgnd vpwr scs8hd_decap_12
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_74 vgnd vpwr scs8hd_decap_12
XFILLER_30_263 vgnd vpwr scs8hd_decap_12
XFILLER_38_19 vgnd vpwr scs8hd_decap_12
XFILLER_13_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l2_in_0__A1 mux_bottom_track_1.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_0_156 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_37.mux_l2_in_0__A1 mux_bottom_track_37.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_245 vgnd vpwr scs8hd_decap_3
XFILLER_12_274 vgnd vpwr scs8hd_fill_1
XFILLER_5_12 vpwr vgnd scs8hd_fill_2
XFILLER_14_32 vgnd vpwr scs8hd_decap_8
XFILLER_5_204 vgnd vpwr scs8hd_fill_1
XFILLER_39_62 vgnd vpwr scs8hd_decap_12
XFILLER_29_171 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_39.mux_l1_in_0_ chanx_left_in[0] bottom_left_grid_pin_40_ mux_bottom_track_39.mux_l1_in_0_/S
+ mux_bottom_track_39.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_35_196 vgnd vpwr scs8hd_decap_12
XFILLER_2_218 vpwr vgnd scs8hd_fill_2
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_26_141 vgnd vpwr scs8hd_decap_12
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XFILLER_25_53 vpwr vgnd scs8hd_fill_2
XFILLER_41_74 vgnd vpwr scs8hd_decap_12
XPHY_75 vgnd vpwr scs8hd_decap_3
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_1_240 vgnd vpwr scs8hd_fill_1
X_51_ chany_bottom_in[15] chanx_left_out[16] vgnd vpwr scs8hd_buf_2
XFILLER_1_273 vgnd vpwr scs8hd_decap_4
XFILLER_32_166 vgnd vpwr scs8hd_decap_12
XFILLER_17_163 vgnd vpwr scs8hd_decap_12
XFILLER_17_196 vgnd vpwr scs8hd_decap_12
Xmux_left_track_5.mux_l2_in_0_ _33_/HI mux_left_track_5.mux_l1_in_0_/X mux_left_track_5.mux_l2_in_0_/S
+ mux_left_track_5.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_0__D mux_bottom_track_5.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_166 vgnd vpwr scs8hd_decap_6
XFILLER_37_269 vgnd vpwr scs8hd_decap_8
X_34_ _34_/HI _34_/LO vgnd vpwr scs8hd_conb_1
XFILLER_7_118 vpwr vgnd scs8hd_fill_2
XFILLER_11_136 vgnd vpwr scs8hd_decap_4
XFILLER_11_169 vpwr vgnd scs8hd_fill_2
XFILLER_22_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_34_239 vgnd vpwr scs8hd_decap_12
XFILLER_19_269 vgnd vpwr scs8hd_decap_8
XFILLER_42_261 vgnd vpwr scs8hd_decap_12
XFILLER_8_23 vgnd vpwr scs8hd_decap_3
XFILLER_8_45 vgnd vpwr scs8hd_fill_1
XFILLER_10_180 vgnd vpwr scs8hd_decap_4
XFILLER_10_191 vpwr vgnd scs8hd_fill_2
XFILLER_33_3 vpwr vgnd scs8hd_fill_2
XFILLER_16_239 vgnd vpwr scs8hd_decap_12
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_86 vgnd vpwr scs8hd_decap_12
XFILLER_33_31 vgnd vpwr scs8hd_decap_12
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_98 vgnd vpwr scs8hd_decap_12
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_143 vpwr vgnd scs8hd_fill_2
XFILLER_3_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_11.mux_l2_in_0__A0 _36_/HI vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_3.scs8hd_buf_4_0_ mux_bottom_track_3.mux_l3_in_0_/X _86_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_21_220 vgnd vpwr scs8hd_decap_12
XFILLER_0_179 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_33.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_33.mux_l1_in_0_/S
+ mux_bottom_track_33.mux_l2_in_0_/S mem_bottom_track_33.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__D mux_bottom_track_25.mux_l1_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_11 vgnd vpwr scs8hd_decap_3
XFILLER_14_44 vgnd vpwr scs8hd_decap_6
XFILLER_14_77 vgnd vpwr scs8hd_decap_12
XFILLER_30_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A0 bottom_left_grid_pin_35_ vgnd vpwr scs8hd_diode_2
XFILLER_39_74 vgnd vpwr scs8hd_decap_12
XFILLER_41_123 vgnd vpwr scs8hd_decap_12
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XFILLER_25_65 vpwr vgnd scs8hd_fill_2
XPHY_54 vgnd vpwr scs8hd_decap_3
XFILLER_41_86 vgnd vpwr scs8hd_decap_12
X_50_ chany_bottom_in[16] chanx_left_out[17] vgnd vpwr scs8hd_buf_2
XFILLER_2_58 vpwr vgnd scs8hd_fill_2
XFILLER_17_120 vpwr vgnd scs8hd_fill_2
XFILLER_32_178 vgnd vpwr scs8hd_decap_12
XFILLER_17_175 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_35.mux_l1_in_0__S mux_bottom_track_35.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_123 vgnd vpwr scs8hd_decap_12
Xmux_left_track_25.mux_l2_in_0_ _32_/HI mux_left_track_25.mux_l1_in_0_/X ccff_tail
+ mux_left_track_25.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_11_12 vpwr vgnd scs8hd_fill_2
XFILLER_14_134 vgnd vpwr scs8hd_decap_4
XFILLER_35_7 vgnd vpwr scs8hd_decap_12
X_33_ _33_/HI _33_/LO vgnd vpwr scs8hd_conb_1
XFILLER_9_182 vgnd vpwr scs8hd_fill_1
XFILLER_28_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_3.mux_l2_in_1__A0 _46_/HI vgnd vpwr scs8hd_diode_2
XFILLER_22_66 vpwr vgnd scs8hd_fill_2
Xmux_left_track_5.mux_l1_in_0_ left_top_grid_pin_1_ chany_bottom_in[1] mux_left_track_5.mux_l1_in_0_/S
+ mux_left_track_5.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_42_273 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.scs8hd_buf_4_0__A mux_bottom_track_9.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_13 vgnd vpwr scs8hd_fill_1
XFILLER_6_163 vpwr vgnd scs8hd_fill_2
XFILLER_26_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_27.scs8hd_dfxbp_1_0__D mux_bottom_track_25.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_22 vgnd vpwr scs8hd_fill_1
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_98 vgnd vpwr scs8hd_decap_12
XFILLER_33_43 vgnd vpwr scs8hd_decap_12
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_251 vgnd vpwr scs8hd_decap_12
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_188 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_11.mux_l2_in_0__A1 mux_bottom_track_11.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_3.mux_l3_in_0__A0 mux_bottom_track_3.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_232 vgnd vpwr scs8hd_decap_12
XFILLER_0_103 vpwr vgnd scs8hd_fill_2
XFILLER_28_32 vgnd vpwr scs8hd_decap_12
XFILLER_0_125 vgnd vpwr scs8hd_decap_3
XFILLER_0_147 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0__S mux_bottom_track_3.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_12_232 vgnd vpwr scs8hd_decap_12
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
XFILLER_5_47 vgnd vpwr scs8hd_decap_3
Xmem_bottom_track_33.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_31.mux_l2_in_0_/S
+ mux_bottom_track_33.mux_l1_in_0_/S mem_bottom_track_33.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_21.scs8hd_buf_4_0__A mux_bottom_track_21.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1__S mux_bottom_track_9.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_14_23 vgnd vpwr scs8hd_decap_6
XFILLER_14_89 vgnd vpwr scs8hd_decap_3
XFILLER_30_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A1 bottom_right_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_25.mux_l2_in_0__S ccff_tail vgnd vpwr scs8hd_diode_2
XFILLER_39_86 vgnd vpwr scs8hd_decap_12
XFILLER_29_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_35.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_35_110 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_27.mux_l2_in_0__S mux_bottom_track_27.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_41_135 vgnd vpwr scs8hd_decap_12
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_154 vgnd vpwr scs8hd_decap_12
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XFILLER_41_98 vgnd vpwr scs8hd_decap_12
XFILLER_2_37 vgnd vpwr scs8hd_decap_4
XFILLER_17_110 vgnd vpwr scs8hd_decap_8
XFILLER_40_190 vgnd vpwr scs8hd_decap_12
XFILLER_23_135 vgnd vpwr scs8hd_decap_12
XFILLER_11_24 vgnd vpwr scs8hd_fill_1
XFILLER_36_32 vgnd vpwr scs8hd_decap_12
XFILLER_22_190 vgnd vpwr scs8hd_decap_12
XFILLER_28_7 vgnd vpwr scs8hd_decap_12
X_32_ _32_/HI _32_/LO vgnd vpwr scs8hd_conb_1
XFILLER_20_105 vgnd vpwr scs8hd_decap_12
XFILLER_28_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_3.mux_l2_in_1__A1 chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_22_45 vpwr vgnd scs8hd_fill_2
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
XFILLER_8_36 vpwr vgnd scs8hd_fill_2
XFILLER_8_69 vpwr vgnd scs8hd_fill_2
Xmux_left_track_25.mux_l1_in_0_ left_top_grid_pin_1_ chany_bottom_in[11] mux_left_track_25.mux_l1_in_0_/S
+ mux_left_track_25.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmem_bottom_track_15.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_15.mux_l1_in_0_/S
+ mux_bottom_track_15.mux_l2_in_0_/S mem_bottom_track_15.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_19_3 vpwr vgnd scs8hd_fill_2
XFILLER_25_208 vgnd vpwr scs8hd_decap_12
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_12 vpwr vgnd scs8hd_fill_2
XFILLER_24_263 vgnd vpwr scs8hd_decap_12
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_55 vgnd vpwr scs8hd_decap_6
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_178 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l3_in_0__A1 mux_bottom_track_3.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_11.mux_l2_in_0_ _36_/HI mux_bottom_track_11.mux_l1_in_0_/X mux_bottom_track_11.mux_l2_in_0_/S
+ mux_bottom_track_11.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_bottom_track_29.scs8hd_buf_4_0_ mux_bottom_track_29.mux_l2_in_0_/X _73_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_28_44 vgnd vpwr scs8hd_decap_12
XFILLER_12_211 vgnd vpwr scs8hd_decap_3
XFILLER_12_244 vgnd vpwr scs8hd_decap_12
XFILLER_8_215 vgnd vpwr scs8hd_decap_12
XFILLER_5_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_15.mux_l1_in_0__A0 chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_38_141 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_30_56 vgnd vpwr scs8hd_decap_12
XFILLER_39_98 vgnd vpwr scs8hd_decap_12
XFILLER_29_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__D mux_left_track_9.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_4_273 vpwr vgnd scs8hd_fill_2
XFILLER_6_80 vpwr vgnd scs8hd_fill_2
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_41_147 vgnd vpwr scs8hd_decap_12
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XFILLER_26_166 vgnd vpwr scs8hd_decap_12
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_7.mux_l3_in_0_ mux_bottom_track_7.mux_l2_in_1_/X mux_bottom_track_7.mux_l2_in_0_/X
+ mux_bottom_track_7.mux_l3_in_0_/S mux_bottom_track_7.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XFILLER_1_210 vpwr vgnd scs8hd_fill_2
XFILLER_2_27 vpwr vgnd scs8hd_fill_2
XFILLER_1_243 vgnd vpwr scs8hd_fill_1
XFILLER_1_232 vpwr vgnd scs8hd_fill_2
XFILLER_1_221 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_15.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_23_147 vgnd vpwr scs8hd_decap_12
XFILLER_11_58 vgnd vpwr scs8hd_decap_3
XFILLER_11_69 vpwr vgnd scs8hd_fill_2
XFILLER_36_44 vgnd vpwr scs8hd_decap_12
X_31_ _31_/HI _31_/LO vgnd vpwr scs8hd_conb_1
XFILLER_20_117 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_7.mux_l2_in_1_ _29_/HI chanx_left_in[4] mux_bottom_track_7.mux_l2_in_1_/S
+ mux_bottom_track_7.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_28_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_31.mux_l1_in_0__S mux_bottom_track_31.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_0_6 vpwr vgnd scs8hd_fill_2
XFILLER_42_242 vgnd vpwr scs8hd_decap_6
XFILLER_6_154 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_40_7 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_15.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_13.mux_l2_in_0_/S
+ mux_bottom_track_15.mux_l1_in_0_/S mem_bottom_track_15.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_33_220 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_37.scs8hd_buf_4_0_ mux_bottom_track_37.mux_l2_in_0_/X _69_/A vgnd
+ vpwr scs8hd_buf_1
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_7.mux_l1_in_1__A0 bottom_left_grid_pin_40_ vgnd vpwr scs8hd_diode_2
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_102 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_23.mux_l1_in_0__A0 chanx_left_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_15_220 vgnd vpwr scs8hd_decap_12
XFILLER_31_3 vpwr vgnd scs8hd_fill_2
XFILLER_2_190 vpwr vgnd scs8hd_fill_2
XFILLER_0_82 vgnd vpwr scs8hd_decap_4
XFILLER_21_245 vgnd vpwr scs8hd_decap_12
XFILLER_0_116 vpwr vgnd scs8hd_fill_2
XFILLER_28_56 vgnd vpwr scs8hd_decap_12
XFILLER_8_227 vpwr vgnd scs8hd_fill_2
XFILLER_12_256 vgnd vpwr scs8hd_decap_12
XFILLER_5_16 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_29.scs8hd_buf_4_0__A mux_bottom_track_29.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_15.mux_l1_in_0__A1 bottom_left_grid_pin_36_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_7.mux_l2_in_0__A0 mux_bottom_track_7.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_30_68 vgnd vpwr scs8hd_decap_12
XFILLER_39_11 vpwr vgnd scs8hd_fill_2
Xmux_left_track_25.scs8hd_buf_4_0_ mux_left_track_25.mux_l2_in_0_/X _55_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mem_bottom_track_29.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_4_241 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_11.mux_l1_in_0_ chanx_left_in[6] bottom_left_grid_pin_34_ mux_bottom_track_11.mux_l1_in_0_/S
+ mux_bottom_track_11.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_35_123 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_23.mux_l2_in_0_ _42_/HI mux_bottom_track_23.mux_l1_in_0_/X mux_bottom_track_23.mux_l2_in_0_/S
+ mux_bottom_track_23.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_26_178 vgnd vpwr scs8hd_decap_12
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XFILLER_41_159 vgnd vpwr scs8hd_decap_12
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_25_57 vpwr vgnd scs8hd_fill_2
XFILLER_9_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l1_in_1__S mux_bottom_track_5.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_17_123 vpwr vgnd scs8hd_fill_2
XFILLER_23_159 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_23.mux_l2_in_0__S mux_bottom_track_23.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_56 vgnd vpwr scs8hd_decap_12
XFILLER_14_104 vgnd vpwr scs8hd_decap_3
XFILLER_14_126 vgnd vpwr scs8hd_decap_6
X_30_ _30_/HI _30_/LO vgnd vpwr scs8hd_conb_1
XFILLER_20_129 vgnd vpwr scs8hd_decap_12
XFILLER_9_163 vpwr vgnd scs8hd_fill_2
XFILLER_9_174 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0__S mux_bottom_track_17.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_7.mux_l2_in_0_ mux_bottom_track_7.mux_l1_in_1_/X mux_bottom_track_7.mux_l1_in_0_/X
+ mux_bottom_track_7.mux_l2_in_1_/S mux_bottom_track_7.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_36_251 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_5.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_track_5.mux_l2_in_0_/S mux_bottom_track_5.mux_l3_in_0_/S
+ mem_bottom_track_5.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_11_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_31.mux_l1_in_0__A0 chanx_left_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_6_133 vpwr vgnd scs8hd_fill_2
XFILLER_6_188 vpwr vgnd scs8hd_fill_2
XFILLER_6_199 vgnd vpwr scs8hd_decap_12
XFILLER_10_195 vgnd vpwr scs8hd_decap_12
XFILLER_33_7 vgnd vpwr scs8hd_decap_12
XFILLER_33_232 vgnd vpwr scs8hd_decap_12
XFILLER_18_251 vgnd vpwr scs8hd_decap_12
XFILLER_17_25 vpwr vgnd scs8hd_fill_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_7.mux_l1_in_1__A1 bottom_left_grid_pin_38_ vgnd vpwr scs8hd_diode_2
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_114 vpwr vgnd scs8hd_fill_2
XFILLER_3_147 vpwr vgnd scs8hd_fill_2
XFILLER_3_136 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_23.mux_l1_in_0__A1 bottom_left_grid_pin_40_ vgnd vpwr scs8hd_diode_2
XFILLER_15_232 vgnd vpwr scs8hd_decap_12
XFILLER_30_202 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_7.mux_l1_in_1_ bottom_left_grid_pin_40_ bottom_left_grid_pin_38_
+ mux_bottom_track_7.mux_l1_in_1_/S mux_bottom_track_7.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_0_94 vgnd vpwr scs8hd_fill_1
XFILLER_21_257 vgnd vpwr scs8hd_decap_12
XFILLER_28_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_31.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_12_268 vgnd vpwr scs8hd_decap_6
XFILLER_5_39 vpwr vgnd scs8hd_fill_2
XFILLER_7_250 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_7.mux_l2_in_0__A1 mux_bottom_track_7.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_38_154 vgnd vpwr scs8hd_decap_12
XFILLER_14_59 vgnd vpwr scs8hd_decap_3
XFILLER_5_209 vpwr vgnd scs8hd_fill_2
XFILLER_39_23 vgnd vpwr scs8hd_decap_12
XFILLER_4_253 vgnd vpwr scs8hd_decap_12
XFILLER_20_80 vgnd vpwr scs8hd_decap_12
XFILLER_35_135 vgnd vpwr scs8hd_decap_12
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XFILLER_25_69 vgnd vpwr scs8hd_decap_12
XFILLER_34_190 vgnd vpwr scs8hd_decap_12
XFILLER_1_245 vgnd vpwr scs8hd_decap_8
XFILLER_32_105 vgnd vpwr scs8hd_decap_12
XFILLER_23_105 vgnd vpwr scs8hd_decap_12
XFILLER_31_171 vgnd vpwr scs8hd_decap_12
XFILLER_16_190 vgnd vpwr scs8hd_decap_12
XFILLER_11_16 vpwr vgnd scs8hd_fill_2
XFILLER_11_27 vpwr vgnd scs8hd_fill_2
XFILLER_36_68 vgnd vpwr scs8hd_decap_12
XFILLER_37_208 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_23.mux_l1_in_0_ chanx_left_in[12] bottom_left_grid_pin_40_ mux_bottom_track_23.mux_l1_in_0_/S
+ mux_bottom_track_23.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_13_171 vgnd vpwr scs8hd_fill_1
XFILLER_13_182 vgnd vpwr scs8hd_fill_1
XFILLER_3_50 vpwr vgnd scs8hd_fill_2
XFILLER_36_263 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_5.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_5.mux_l1_in_1_/S mux_bottom_track_5.mux_l2_in_0_/S
+ mem_bottom_track_5.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_bottom_track_35.mux_l2_in_0_ _25_/HI mux_bottom_track_35.mux_l1_in_0_/X mux_bottom_track_35.mux_l2_in_0_/S
+ mux_bottom_track_35.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_bottom_track_11.scs8hd_buf_4_0_ mux_bottom_track_11.mux_l2_in_0_/X _82_/A vgnd
+ vpwr scs8hd_buf_1
XANTENNA_mux_bottom_track_31.mux_l1_in_0__A1 bottom_left_grid_pin_36_ vgnd vpwr scs8hd_diode_2
XFILLER_22_37 vgnd vpwr scs8hd_decap_8
XFILLER_42_211 vgnd vpwr scs8hd_decap_6
XFILLER_19_208 vgnd vpwr scs8hd_decap_12
XFILLER_8_28 vgnd vpwr scs8hd_decap_3
XFILLER_6_145 vpwr vgnd scs8hd_fill_2
XFILLER_6_167 vpwr vgnd scs8hd_fill_2
XFILLER_10_163 vgnd vpwr scs8hd_decap_8
XFILLER_26_7 vgnd vpwr scs8hd_decap_12
XFILLER_18_263 vgnd vpwr scs8hd_decap_12
XFILLER_17_48 vgnd vpwr scs8hd_decap_12
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_7.mux_l1_in_0_ bottom_left_grid_pin_36_ bottom_left_grid_pin_34_
+ mux_bottom_track_7.mux_l1_in_1_/S mux_bottom_track_7.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_17_3 vpwr vgnd scs8hd_fill_2
XFILLER_21_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_17.mux_l2_in_0__A0 _39_/HI vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.scs8hd_buf_4_0_ mux_bottom_track_9.mux_l2_in_0_/X _83_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_18_91 vgnd vpwr scs8hd_fill_1
XFILLER_7_262 vgnd vpwr scs8hd_decap_12
XFILLER_38_166 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_13.scs8hd_dfxbp_1_1__D mux_bottom_track_13.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_15 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_23.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_23.mux_l1_in_0_/S
+ mux_bottom_track_23.mux_l2_in_0_/S mem_bottom_track_23.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_39_35 vgnd vpwr scs8hd_decap_12
XFILLER_4_265 vgnd vpwr scs8hd_decap_8
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XFILLER_35_147 vgnd vpwr scs8hd_decap_12
XFILLER_29_90 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_11.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_1__D mux_bottom_track_33.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XPHY_59 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XFILLER_25_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_257 vpwr vgnd scs8hd_fill_2
XFILLER_32_117 vgnd vpwr scs8hd_decap_12
XFILLER_31_80 vpwr vgnd scs8hd_fill_2
XFILLER_23_117 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.scs8hd_buf_4_0__A mux_left_track_1.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_25.mux_l1_in_1__A0 _43_/HI vgnd vpwr scs8hd_diode_2
XFILLER_26_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_1.mux_l1_in_1__S mux_bottom_track_1.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_62 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_5.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_3.mux_l3_in_0_/S mux_bottom_track_5.mux_l1_in_1_/S
+ mem_bottom_track_5.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__D mux_left_track_1.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_27_220 vgnd vpwr scs8hd_decap_12
XANTENNA__52__A chany_bottom_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_6_102 vpwr vgnd scs8hd_fill_2
XFILLER_10_131 vgnd vpwr scs8hd_decap_3
XFILLER_10_186 vpwr vgnd scs8hd_fill_2
XFILLER_19_7 vgnd vpwr scs8hd_decap_3
XFILLER_33_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_25.mux_l2_in_0__A0 mux_bottom_track_25.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_25.mux_l1_in_1__S mux_bottom_track_25.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_17_16 vgnd vpwr scs8hd_decap_6
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_bottom_track_15.scs8hd_dfxbp_1_0__D mux_bottom_track_13.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_13.mux_l1_in_0__S mux_bottom_track_13.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_30_215 vgnd vpwr scs8hd_decap_12
XFILLER_15_245 vgnd vpwr scs8hd_decap_12
XFILLER_23_81 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_35.mux_l1_in_0_ chanx_left_in[18] bottom_left_grid_pin_38_ mux_bottom_track_35.mux_l1_in_0_/S
+ mux_bottom_track_35.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_bottom_track_35.scs8hd_dfxbp_1_0__D mux_bottom_track_33.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_72 vpwr vgnd scs8hd_fill_2
XFILLER_9_83 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_27.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0__A1 mux_bottom_track_17.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_12_215 vgnd vpwr scs8hd_decap_12
XFILLER_8_208 vgnd vpwr scs8hd_decap_6
XFILLER_34_80 vgnd vpwr scs8hd_decap_12
XFILLER_7_274 vgnd vpwr scs8hd_decap_3
Xmux_left_track_1.mux_l2_in_0_ _31_/HI mux_left_track_1.mux_l1_in_0_/X mux_left_track_1.mux_l2_in_0_/S
+ mux_left_track_1.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_38_178 vgnd vpwr scs8hd_decap_12
XFILLER_30_27 vgnd vpwr scs8hd_decap_4
Xmem_bottom_track_23.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_21.mux_l2_in_0_/S
+ mux_bottom_track_23.mux_l1_in_0_/S mem_bottom_track_23.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_39_47 vgnd vpwr scs8hd_decap_12
XFILLER_29_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_11.scs8hd_buf_4_0__A mux_bottom_track_11.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l2_in_0__A0 _33_/HI vgnd vpwr scs8hd_diode_2
XANTENNA__60__A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_20_93 vgnd vpwr scs8hd_decap_12
XFILLER_35_159 vgnd vpwr scs8hd_decap_12
XFILLER_6_84 vpwr vgnd scs8hd_fill_2
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XPHY_49 vgnd vpwr scs8hd_decap_3
XFILLER_25_27 vgnd vpwr scs8hd_decap_12
XFILLER_25_49 vpwr vgnd scs8hd_fill_2
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_236 vgnd vpwr scs8hd_decap_4
XFILLER_1_225 vgnd vpwr scs8hd_decap_4
XFILLER_1_214 vgnd vpwr scs8hd_decap_4
XFILLER_32_129 vgnd vpwr scs8hd_decap_12
XANTENNA__55__A _55_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_82 vpwr vgnd scs8hd_fill_2
XFILLER_31_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_37.scs8hd_buf_4_0__A mux_bottom_track_37.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_25.mux_l1_in_1__A1 chanx_left_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_7_3 vpwr vgnd scs8hd_fill_2
XFILLER_9_100 vpwr vgnd scs8hd_fill_2
XFILLER_13_151 vgnd vpwr scs8hd_decap_12
XFILLER_9_133 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_33.mux_l2_in_0__A0 _24_/HI vgnd vpwr scs8hd_diode_2
XFILLER_13_184 vgnd vpwr scs8hd_decap_12
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
X_87_ _87_/A chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_27_232 vgnd vpwr scs8hd_decap_12
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_25.mux_l2_in_0__A1 mux_bottom_track_25.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_202 vgnd vpwr scs8hd_decap_12
XFILLER_3_106 vgnd vpwr scs8hd_decap_3
XFILLER_30_227 vgnd vpwr scs8hd_decap_12
XFILLER_15_257 vgnd vpwr scs8hd_decap_12
XANTENNA__63__A _63_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_93 vgnd vpwr scs8hd_decap_12
XFILLER_31_7 vgnd vpwr scs8hd_decap_12
XFILLER_2_194 vgnd vpwr scs8hd_decap_4
XFILLER_0_86 vgnd vpwr scs8hd_fill_1
XFILLER_9_62 vgnd vpwr scs8hd_decap_4
XFILLER_12_227 vpwr vgnd scs8hd_fill_2
XANTENNA__58__A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_18_93 vgnd vpwr scs8hd_decap_12
XFILLER_7_220 vgnd vpwr scs8hd_decap_3
XFILLER_7_231 vpwr vgnd scs8hd_fill_2
XFILLER_39_59 vpwr vgnd scs8hd_fill_2
XFILLER_29_102 vgnd vpwr scs8hd_decap_12
XFILLER_29_135 vgnd vpwr scs8hd_decap_12
XFILLER_4_212 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l2_in_0__A1 mux_left_track_5.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_61 vgnd vpwr scs8hd_fill_1
XFILLER_28_190 vgnd vpwr scs8hd_decap_12
XFILLER_6_41 vgnd vpwr scs8hd_decap_4
XFILLER_6_52 vpwr vgnd scs8hd_fill_2
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_26_105 vgnd vpwr scs8hd_decap_12
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_25_39 vgnd vpwr scs8hd_decap_4
XFILLER_17_127 vgnd vpwr scs8hd_decap_12
XFILLER_25_171 vgnd vpwr scs8hd_decap_12
XFILLER_40_141 vgnd vpwr scs8hd_decap_12
XANTENNA__71__A _71_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_0_ left_top_grid_pin_1_ chany_bottom_in[19] mux_left_track_1.mux_l1_in_0_/S
+ mux_left_track_1.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_9.scs8hd_buf_4_0__A mux_left_track_9.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_31_196 vgnd vpwr scs8hd_decap_12
XFILLER_22_141 vgnd vpwr scs8hd_decap_12
XANTENNA__66__A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_9_123 vgnd vpwr scs8hd_fill_1
XFILLER_13_163 vgnd vpwr scs8hd_decap_8
XFILLER_13_174 vpwr vgnd scs8hd_fill_2
XFILLER_26_71 vgnd vpwr scs8hd_decap_12
XFILLER_26_93 vgnd vpwr scs8hd_decap_12
XFILLER_9_167 vpwr vgnd scs8hd_fill_2
XFILLER_9_178 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_33.mux_l2_in_0__A1 mux_bottom_track_33.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_196 vgnd vpwr scs8hd_decap_12
XFILLER_3_75 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
X_86_ _86_/A chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_6_137 vgnd vpwr scs8hd_decap_3
XFILLER_6_159 vpwr vgnd scs8hd_fill_2
XFILLER_12_51 vpwr vgnd scs8hd_fill_2
XFILLER_12_84 vgnd vpwr scs8hd_decap_6
XFILLER_33_269 vgnd vpwr scs8hd_decap_8
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_69_ _69_/A chany_bottom_out[18] vgnd vpwr scs8hd_buf_2
XFILLER_3_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_19.scs8hd_dfxbp_1_1__D mux_bottom_track_19.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_239 vgnd vpwr scs8hd_decap_12
XFILLER_15_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_25.scs8hd_buf_4_0__A mux_left_track_25.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_0_10 vpwr vgnd scs8hd_fill_2
XFILLER_24_7 vgnd vpwr scs8hd_decap_12
XFILLER_0_32 vgnd vpwr scs8hd_decap_3
XFILLER_0_54 vpwr vgnd scs8hd_fill_2
XFILLER_9_52 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_39.scs8hd_dfxbp_1_1__D mux_bottom_track_39.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_29.mux_l1_in_0__A0 chanx_left_in[15] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_7.mux_l1_in_0__S mux_bottom_track_7.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA__74__A _74_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_34_93 vgnd vpwr scs8hd_decap_12
XFILLER_7_243 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_37.mux_l2_in_0__S mux_bottom_track_37.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_15_3 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_19.scs8hd_buf_4_0__A mux_bottom_track_19.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_114 vgnd vpwr scs8hd_decap_8
XFILLER_29_147 vgnd vpwr scs8hd_decap_12
XANTENNA__69__A _69_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_51 vpwr vgnd scs8hd_fill_2
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_26_117 vgnd vpwr scs8hd_decap_12
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XFILLER_15_62 vgnd vpwr scs8hd_decap_12
XFILLER_17_139 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0__A0 left_top_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XFILLER_31_120 vpwr vgnd scs8hd_fill_2
XFILLER_39_220 vgnd vpwr scs8hd_decap_12
XANTENNA__82__A _82_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_31.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_31.mux_l1_in_0_/S
+ mux_bottom_track_31.mux_l2_in_0_/S mem_bottom_track_31.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_26_83 vgnd vpwr scs8hd_decap_8
XFILLER_3_54 vgnd vpwr scs8hd_decap_4
X_85_ _85_/A chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_22_19 vgnd vpwr scs8hd_decap_12
XFILLER_27_245 vgnd vpwr scs8hd_decap_12
XFILLER_10_112 vgnd vpwr scs8hd_decap_8
XFILLER_10_123 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l3_in_0__S mux_bottom_track_5.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_6_149 vpwr vgnd scs8hd_fill_2
XFILLER_10_145 vpwr vgnd scs8hd_fill_2
XANTENNA__77__A _77_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_37.mux_l1_in_0__A0 chanx_left_in[19] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A0 bottom_left_grid_pin_35_ vgnd vpwr scs8hd_diode_2
XFILLER_5_160 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_23.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_5_193 vgnd vpwr scs8hd_decap_3
X_68_ _68_/A chany_bottom_out[19] vgnd vpwr scs8hd_buf_2
XFILLER_24_215 vgnd vpwr scs8hd_decap_12
XFILLER_23_51 vpwr vgnd scs8hd_fill_2
XFILLER_2_163 vpwr vgnd scs8hd_fill_2
XFILLER_17_7 vpwr vgnd scs8hd_fill_2
XFILLER_0_99 vpwr vgnd scs8hd_fill_2
XFILLER_9_20 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_29.mux_l1_in_0__A1 bottom_left_grid_pin_35_ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__D mux_bottom_track_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_251 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_3.mux_l3_in_0_ mux_bottom_track_3.mux_l2_in_1_/X mux_bottom_track_3.mux_l2_in_0_/X
+ mux_bottom_track_3.mux_l3_in_0_/S mux_bottom_track_3.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__D mux_left_track_5.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_51 vgnd vpwr scs8hd_decap_12
XFILLER_29_159 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_7.scs8hd_buf_4_0__A mux_bottom_track_7.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA__85__A _85_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_76 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_3.mux_l2_in_1_ _46_/HI chanx_left_in[2] mux_bottom_track_3.mux_l2_in_0_/S
+ mux_bottom_track_3.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XPHY_19 vgnd vpwr scs8hd_decap_3
XFILLER_26_129 vgnd vpwr scs8hd_decap_12
XFILLER_40_154 vgnd vpwr scs8hd_decap_12
XFILLER_15_74 vgnd vpwr scs8hd_decap_8
XFILLER_25_184 vgnd vpwr scs8hd_decap_12
XFILLER_31_84 vgnd vpwr scs8hd_decap_12
XFILLER_31_62 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0__A1 chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_39.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_22_154 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_31.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_29.mux_l2_in_0_/S
+ mux_bottom_track_31.mux_l1_in_0_/S mem_bottom_track_31.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_42_94 vgnd vpwr scs8hd_decap_12
XFILLER_9_114 vpwr vgnd scs8hd_fill_2
XFILLER_3_22 vpwr vgnd scs8hd_fill_2
XFILLER_36_202 vgnd vpwr scs8hd_decap_12
X_84_ _84_/A chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_3_33 vpwr vgnd scs8hd_fill_2
XFILLER_27_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_0__D mux_bottom_track_1.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_249 vgnd vpwr scs8hd_decap_12
XFILLER_6_106 vpwr vgnd scs8hd_fill_2
XFILLER_12_64 vgnd vpwr scs8hd_fill_1
XFILLER_18_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_37.mux_l1_in_0__A1 bottom_left_grid_pin_39_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A1 bottom_right_grid_pin_1_ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.scs8hd_buf_4_0_ mux_bottom_track_17.mux_l2_in_0_/X _79_/A vgnd
+ vpwr scs8hd_buf_1
X_67_ _67_/A chanx_left_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_24_227 vgnd vpwr scs8hd_decap_12
XFILLER_33_19 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l2_in_0_ _39_/HI mux_bottom_track_17.mux_l1_in_0_/X mux_bottom_track_17.mux_l2_in_0_/S
+ mux_bottom_track_17.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_0_23 vpwr vgnd scs8hd_fill_2
XFILLER_0_89 vpwr vgnd scs8hd_fill_2
XFILLER_9_87 vpwr vgnd scs8hd_fill_2
XFILLER_21_208 vgnd vpwr scs8hd_decap_12
XFILLER_28_19 vgnd vpwr scs8hd_decap_12
XFILLER_20_263 vgnd vpwr scs8hd_decap_12
XFILLER_18_63 vgnd vpwr scs8hd_decap_12
XFILLER_11_230 vpwr vgnd scs8hd_fill_2
XFILLER_7_201 vgnd vpwr scs8hd_decap_4
XFILLER_7_212 vgnd vpwr scs8hd_decap_8
XFILLER_7_245 vgnd vpwr scs8hd_decap_3
XFILLER_38_105 vgnd vpwr scs8hd_decap_12
XFILLER_37_171 vgnd vpwr scs8hd_decap_12
XFILLER_4_204 vgnd vpwr scs8hd_decap_8
XFILLER_29_62 vgnd vpwr scs8hd_decap_8
XFILLER_20_64 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0__S mux_bottom_track_3.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_bottom_track_13.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_13.mux_l1_in_0_/S
+ mux_bottom_track_13.mux_l2_in_0_/S mem_bottom_track_13.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_6_88 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_21.scs8hd_dfxbp_1_1__D mux_bottom_track_21.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_141 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_3.mux_l2_in_0_ mux_bottom_track_3.mux_l1_in_1_/X mux_bottom_track_3.mux_l1_in_0_/X
+ mux_bottom_track_3.mux_l2_in_0_/S mux_bottom_track_3.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_19_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_33.mux_l2_in_0__S mux_bottom_track_33.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_40_166 vgnd vpwr scs8hd_decap_12
XFILLER_15_42 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_25.mux_l1_in_0__S mux_left_track_25.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_25_196 vgnd vpwr scs8hd_decap_12
XFILLER_31_96 vgnd vpwr scs8hd_decap_12
XFILLER_31_74 vpwr vgnd scs8hd_fill_2
XFILLER_0_240 vpwr vgnd scs8hd_fill_2
XFILLER_16_141 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_27.mux_l1_in_0__S mux_bottom_track_27.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
.ends

