VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cby_1__1_
  CLASS BLOCK ;
  FOREIGN cby_1__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 85.000 BY 100.000 ;
  PIN Test_en_E_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 82.600 83.000 85.000 83.600 ;
    END
  END Test_en_E_in
  PIN Test_en_E_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 82.600 49.680 85.000 50.280 ;
    END
  END Test_en_E_out
  PIN Test_en_N_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 15.730 97.600 16.010 100.000 ;
    END
  END Test_en_N_out
  PIN Test_en_S_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 2.400 ;
    END
  END Test_en_S_in
  PIN Test_en_W_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 2.400 87.000 ;
    END
  END Test_en_W_in
  PIN Test_en_W_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 2.400 92.440 ;
    END
  END Test_en_W_out
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 2.400 2.680 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 82.600 16.360 85.000 16.960 ;
    END
  END ccff_tail
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 2.400 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 2.400 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 2.400 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 2.400 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 2.400 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 2.400 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 2.400 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 2.400 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 2.400 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 2.400 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 2.400 ;
    END
  END chany_bottom_in[19]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 2.400 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 2.400 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 2.400 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 2.400 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 2.400 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.710 0.000 44.990 2.400 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 2.400 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 2.400 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 2.400 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 0.550 0.000 0.830 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 2.400 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 2.400 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 2.400 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 2.400 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 2.400 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 2.400 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 2.400 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 2.400 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 2.400 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 2.400 ;
    END
  END chany_bottom_out[19]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 2.400 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 2.400 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 2.400 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 2.400 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 2.400 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 10.670 0.000 10.950 2.400 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 2.400 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 2.400 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 2.400 ;
    END
  END chany_bottom_out[9]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 51.610 97.600 51.890 100.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.630 97.600 68.910 100.000 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.010 97.600 70.290 100.000 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 71.850 97.600 72.130 100.000 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 73.690 97.600 73.970 100.000 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.070 97.600 75.350 100.000 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 76.910 97.600 77.190 100.000 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.750 97.600 79.030 100.000 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.130 97.600 80.410 100.000 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 81.970 97.600 82.250 100.000 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 83.810 97.600 84.090 100.000 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.990 97.600 53.270 100.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 54.830 97.600 55.110 100.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.670 97.600 56.950 100.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.050 97.600 58.330 100.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.890 97.600 60.170 100.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.730 97.600 62.010 100.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.110 97.600 63.390 100.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.950 97.600 65.230 100.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 66.790 97.600 67.070 100.000 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 17.570 97.600 17.850 100.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 34.590 97.600 34.870 100.000 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 35.970 97.600 36.250 100.000 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 37.810 97.600 38.090 100.000 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 39.650 97.600 39.930 100.000 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 41.030 97.600 41.310 100.000 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 42.870 97.600 43.150 100.000 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 44.710 97.600 44.990 100.000 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 46.090 97.600 46.370 100.000 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 47.930 97.600 48.210 100.000 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 49.770 97.600 50.050 100.000 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 18.950 97.600 19.230 100.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 20.790 97.600 21.070 100.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 22.630 97.600 22.910 100.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.010 97.600 24.290 100.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 25.850 97.600 26.130 100.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 27.690 97.600 27.970 100.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 29.070 97.600 29.350 100.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 30.910 97.600 31.190 100.000 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 32.750 97.600 33.030 100.000 ;
    END
  END chany_top_out[9]
  PIN clk_2_N_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 0.550 97.600 0.830 100.000 ;
    END
  END clk_2_N_in
  PIN clk_2_N_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 6.990 97.600 7.270 100.000 ;
    END
  END clk_2_N_out
  PIN clk_2_S_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 2.400 ;
    END
  END clk_2_S_in
  PIN clk_2_S_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 2.400 ;
    END
  END clk_2_S_out
  PIN clk_3_N_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.930 97.600 2.210 100.000 ;
    END
  END clk_3_N_in
  PIN clk_3_N_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 8.830 97.600 9.110 100.000 ;
    END
  END clk_3_N_out
  PIN clk_3_S_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 2.400 ;
    END
  END clk_3_S_in
  PIN clk_3_S_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 2.400 ;
    END
  END clk_3_S_out
  PIN left_grid_pin_16_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 2.400 7.440 ;
    END
  END left_grid_pin_16_
  PIN left_grid_pin_17_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.600 2.400 12.200 ;
    END
  END left_grid_pin_17_
  PIN left_grid_pin_18_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 2.400 17.640 ;
    END
  END left_grid_pin_18_
  PIN left_grid_pin_19_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 2.400 22.400 ;
    END
  END left_grid_pin_19_
  PIN left_grid_pin_20_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 2.400 27.160 ;
    END
  END left_grid_pin_20_
  PIN left_grid_pin_21_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.000 2.400 32.600 ;
    END
  END left_grid_pin_21_
  PIN left_grid_pin_22_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 2.400 37.360 ;
    END
  END left_grid_pin_22_
  PIN left_grid_pin_23_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.520 2.400 42.120 ;
    END
  END left_grid_pin_23_
  PIN left_grid_pin_24_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.960 2.400 47.560 ;
    END
  END left_grid_pin_24_
  PIN left_grid_pin_25_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 2.400 52.320 ;
    END
  END left_grid_pin_25_
  PIN left_grid_pin_26_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 2.400 57.080 ;
    END
  END left_grid_pin_26_
  PIN left_grid_pin_27_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.920 2.400 62.520 ;
    END
  END left_grid_pin_27_
  PIN left_grid_pin_28_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 2.400 67.280 ;
    END
  END left_grid_pin_28_
  PIN left_grid_pin_29_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 2.400 72.040 ;
    END
  END left_grid_pin_29_
  PIN left_grid_pin_30_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 2.400 77.480 ;
    END
  END left_grid_pin_30_
  PIN left_grid_pin_31_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 2.400 82.240 ;
    END
  END left_grid_pin_31_
  PIN prog_clk_0_N_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 10.670 97.600 10.950 100.000 ;
    END
  END prog_clk_0_N_out
  PIN prog_clk_0_S_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 2.400 ;
    END
  END prog_clk_0_S_out
  PIN prog_clk_0_W_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 2.400 97.200 ;
    END
  END prog_clk_0_W_in
  PIN prog_clk_2_N_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.770 97.600 4.050 100.000 ;
    END
  END prog_clk_2_N_in
  PIN prog_clk_2_N_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 12.050 97.600 12.330 100.000 ;
    END
  END prog_clk_2_N_out
  PIN prog_clk_2_S_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 2.400 ;
    END
  END prog_clk_2_S_in
  PIN prog_clk_2_S_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 2.400 ;
    END
  END prog_clk_2_S_out
  PIN prog_clk_3_N_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.610 97.600 5.890 100.000 ;
    END
  END prog_clk_3_N_in
  PIN prog_clk_3_N_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 13.890 97.600 14.170 100.000 ;
    END
  END prog_clk_3_N_out
  PIN prog_clk_3_S_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 2.400 ;
    END
  END prog_clk_3_S_in
  PIN prog_clk_3_S_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 2.400 ;
    END
  END prog_clk_3_S_out
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 17.045 10.640 18.645 87.280 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 29.375 10.640 30.975 87.280 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 4.745 9.945 79.120 89.675 ;
      LAYER met1 ;
        RECT 0.530 6.160 84.110 90.400 ;
      LAYER met2 ;
        RECT 1.110 97.320 1.650 97.600 ;
        RECT 2.490 97.320 3.490 97.600 ;
        RECT 4.330 97.320 5.330 97.600 ;
        RECT 6.170 97.320 6.710 97.600 ;
        RECT 7.550 97.320 8.550 97.600 ;
        RECT 9.390 97.320 10.390 97.600 ;
        RECT 11.230 97.320 11.770 97.600 ;
        RECT 12.610 97.320 13.610 97.600 ;
        RECT 14.450 97.320 15.450 97.600 ;
        RECT 16.290 97.320 17.290 97.600 ;
        RECT 18.130 97.320 18.670 97.600 ;
        RECT 19.510 97.320 20.510 97.600 ;
        RECT 21.350 97.320 22.350 97.600 ;
        RECT 23.190 97.320 23.730 97.600 ;
        RECT 24.570 97.320 25.570 97.600 ;
        RECT 26.410 97.320 27.410 97.600 ;
        RECT 28.250 97.320 28.790 97.600 ;
        RECT 29.630 97.320 30.630 97.600 ;
        RECT 31.470 97.320 32.470 97.600 ;
        RECT 33.310 97.320 34.310 97.600 ;
        RECT 35.150 97.320 35.690 97.600 ;
        RECT 36.530 97.320 37.530 97.600 ;
        RECT 38.370 97.320 39.370 97.600 ;
        RECT 40.210 97.320 40.750 97.600 ;
        RECT 41.590 97.320 42.590 97.600 ;
        RECT 43.430 97.320 44.430 97.600 ;
        RECT 45.270 97.320 45.810 97.600 ;
        RECT 46.650 97.320 47.650 97.600 ;
        RECT 48.490 97.320 49.490 97.600 ;
        RECT 50.330 97.320 51.330 97.600 ;
        RECT 52.170 97.320 52.710 97.600 ;
        RECT 53.550 97.320 54.550 97.600 ;
        RECT 55.390 97.320 56.390 97.600 ;
        RECT 57.230 97.320 57.770 97.600 ;
        RECT 58.610 97.320 59.610 97.600 ;
        RECT 60.450 97.320 61.450 97.600 ;
        RECT 62.290 97.320 62.830 97.600 ;
        RECT 63.670 97.320 64.670 97.600 ;
        RECT 65.510 97.320 66.510 97.600 ;
        RECT 67.350 97.320 68.350 97.600 ;
        RECT 69.190 97.320 69.730 97.600 ;
        RECT 70.570 97.320 71.570 97.600 ;
        RECT 72.410 97.320 73.410 97.600 ;
        RECT 74.250 97.320 74.790 97.600 ;
        RECT 75.630 97.320 76.630 97.600 ;
        RECT 77.470 97.320 78.470 97.600 ;
        RECT 79.310 97.320 79.850 97.600 ;
        RECT 80.690 97.320 81.690 97.600 ;
        RECT 82.530 97.320 83.530 97.600 ;
        RECT 0.560 2.680 84.090 97.320 ;
        RECT 1.110 2.195 1.650 2.680 ;
        RECT 2.490 2.195 3.490 2.680 ;
        RECT 4.330 2.195 5.330 2.680 ;
        RECT 6.170 2.195 6.710 2.680 ;
        RECT 7.550 2.195 8.550 2.680 ;
        RECT 9.390 2.195 10.390 2.680 ;
        RECT 11.230 2.195 11.770 2.680 ;
        RECT 12.610 2.195 13.610 2.680 ;
        RECT 14.450 2.195 15.450 2.680 ;
        RECT 16.290 2.195 17.290 2.680 ;
        RECT 18.130 2.195 18.670 2.680 ;
        RECT 19.510 2.195 20.510 2.680 ;
        RECT 21.350 2.195 22.350 2.680 ;
        RECT 23.190 2.195 23.730 2.680 ;
        RECT 24.570 2.195 25.570 2.680 ;
        RECT 26.410 2.195 27.410 2.680 ;
        RECT 28.250 2.195 28.790 2.680 ;
        RECT 29.630 2.195 30.630 2.680 ;
        RECT 31.470 2.195 32.470 2.680 ;
        RECT 33.310 2.195 34.310 2.680 ;
        RECT 35.150 2.195 35.690 2.680 ;
        RECT 36.530 2.195 37.530 2.680 ;
        RECT 38.370 2.195 39.370 2.680 ;
        RECT 40.210 2.195 40.750 2.680 ;
        RECT 41.590 2.195 42.590 2.680 ;
        RECT 43.430 2.195 44.430 2.680 ;
        RECT 45.270 2.195 45.810 2.680 ;
        RECT 46.650 2.195 47.650 2.680 ;
        RECT 48.490 2.195 49.490 2.680 ;
        RECT 50.330 2.195 51.330 2.680 ;
        RECT 52.170 2.195 52.710 2.680 ;
        RECT 53.550 2.195 54.550 2.680 ;
        RECT 55.390 2.195 56.390 2.680 ;
        RECT 57.230 2.195 57.770 2.680 ;
        RECT 58.610 2.195 59.610 2.680 ;
        RECT 60.450 2.195 61.450 2.680 ;
        RECT 62.290 2.195 62.830 2.680 ;
        RECT 63.670 2.195 64.670 2.680 ;
        RECT 65.510 2.195 66.510 2.680 ;
        RECT 67.350 2.195 68.350 2.680 ;
        RECT 69.190 2.195 69.730 2.680 ;
        RECT 70.570 2.195 71.570 2.680 ;
        RECT 72.410 2.195 73.410 2.680 ;
        RECT 74.250 2.195 74.790 2.680 ;
        RECT 75.630 2.195 76.630 2.680 ;
        RECT 77.470 2.195 78.470 2.680 ;
        RECT 79.310 2.195 79.850 2.680 ;
        RECT 80.690 2.195 81.690 2.680 ;
        RECT 82.530 2.195 83.530 2.680 ;
      LAYER met3 ;
        RECT 2.800 96.200 84.115 97.065 ;
        RECT 2.400 92.840 84.115 96.200 ;
        RECT 2.800 91.440 84.115 92.840 ;
        RECT 2.400 87.400 84.115 91.440 ;
        RECT 2.800 86.000 84.115 87.400 ;
        RECT 2.400 84.000 84.115 86.000 ;
        RECT 2.400 82.640 82.200 84.000 ;
        RECT 2.800 82.600 82.200 82.640 ;
        RECT 2.800 81.240 84.115 82.600 ;
        RECT 2.400 77.880 84.115 81.240 ;
        RECT 2.800 76.480 84.115 77.880 ;
        RECT 2.400 72.440 84.115 76.480 ;
        RECT 2.800 71.040 84.115 72.440 ;
        RECT 2.400 67.680 84.115 71.040 ;
        RECT 2.800 66.280 84.115 67.680 ;
        RECT 2.400 62.920 84.115 66.280 ;
        RECT 2.800 61.520 84.115 62.920 ;
        RECT 2.400 57.480 84.115 61.520 ;
        RECT 2.800 56.080 84.115 57.480 ;
        RECT 2.400 52.720 84.115 56.080 ;
        RECT 2.800 51.320 84.115 52.720 ;
        RECT 2.400 50.680 84.115 51.320 ;
        RECT 2.400 49.280 82.200 50.680 ;
        RECT 2.400 47.960 84.115 49.280 ;
        RECT 2.800 46.560 84.115 47.960 ;
        RECT 2.400 42.520 84.115 46.560 ;
        RECT 2.800 41.120 84.115 42.520 ;
        RECT 2.400 37.760 84.115 41.120 ;
        RECT 2.800 36.360 84.115 37.760 ;
        RECT 2.400 33.000 84.115 36.360 ;
        RECT 2.800 31.600 84.115 33.000 ;
        RECT 2.400 27.560 84.115 31.600 ;
        RECT 2.800 26.160 84.115 27.560 ;
        RECT 2.400 22.800 84.115 26.160 ;
        RECT 2.800 21.400 84.115 22.800 ;
        RECT 2.400 18.040 84.115 21.400 ;
        RECT 2.800 17.360 84.115 18.040 ;
        RECT 2.800 16.640 82.200 17.360 ;
        RECT 2.400 15.960 82.200 16.640 ;
        RECT 2.400 12.600 84.115 15.960 ;
        RECT 2.800 11.200 84.115 12.600 ;
        RECT 2.400 7.840 84.115 11.200 ;
        RECT 2.800 6.440 84.115 7.840 ;
        RECT 2.400 3.080 84.115 6.440 ;
        RECT 2.800 2.215 84.115 3.080 ;
      LAYER met4 ;
        RECT 12.255 10.640 16.645 87.280 ;
        RECT 19.045 10.640 28.975 87.280 ;
        RECT 31.375 10.640 72.385 87.280 ;
  END
END cby_1__1_
END LIBRARY

