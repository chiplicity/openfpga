magic
tech sky130A
magscale 1 2
timestamp 1605004454
<< locali >>
rect 15301 22083 15335 22185
rect 8953 20247 8987 20553
rect 12449 20315 12483 20417
rect 13461 16439 13495 16609
rect 6101 15895 6135 15997
rect 8309 15963 8343 16201
rect 13277 12087 13311 12189
rect 4997 9367 5031 9469
rect 13461 8415 13495 8517
rect 11069 7735 11103 8041
rect 14933 7803 14967 7973
rect 10517 7191 10551 7293
rect 16129 3995 16163 4097
rect 17693 3995 17727 4097
<< viali >>
rect 1593 25449 1627 25483
rect 7113 25449 7147 25483
rect 8217 25449 8251 25483
rect 1409 25313 1443 25347
rect 2513 25313 2547 25347
rect 4077 25313 4111 25347
rect 5181 25313 5215 25347
rect 6929 25313 6963 25347
rect 8033 25313 8067 25347
rect 9781 25313 9815 25347
rect 15485 25313 15519 25347
rect 5825 25245 5859 25279
rect 2697 25177 2731 25211
rect 5365 25177 5399 25211
rect 9965 25177 9999 25211
rect 2053 25109 2087 25143
rect 4261 25109 4295 25143
rect 15669 25109 15703 25143
rect 7021 24905 7055 24939
rect 8125 24905 8159 24939
rect 7757 24837 7791 24871
rect 5825 24769 5859 24803
rect 7481 24769 7515 24803
rect 9781 24769 9815 24803
rect 12633 24769 12667 24803
rect 1501 24701 1535 24735
rect 2329 24701 2363 24735
rect 2789 24701 2823 24735
rect 3341 24701 3375 24735
rect 3893 24701 3927 24735
rect 6837 24701 6871 24735
rect 7941 24701 7975 24735
rect 8493 24701 8527 24735
rect 9505 24701 9539 24735
rect 9597 24701 9631 24735
rect 10333 24701 10367 24735
rect 12449 24701 12483 24735
rect 15117 24701 15151 24735
rect 16221 24701 16255 24735
rect 16773 24701 16807 24735
rect 18061 24701 18095 24735
rect 18613 24701 18647 24735
rect 1777 24633 1811 24667
rect 3709 24633 3743 24667
rect 5089 24633 5123 24667
rect 5641 24633 5675 24667
rect 15025 24633 15059 24667
rect 2605 24565 2639 24599
rect 2973 24565 3007 24599
rect 4077 24565 4111 24599
rect 4445 24565 4479 24599
rect 5181 24565 5215 24599
rect 5549 24565 5583 24599
rect 6285 24565 6319 24599
rect 6653 24565 6687 24599
rect 8861 24565 8895 24599
rect 13185 24565 13219 24599
rect 13645 24565 13679 24599
rect 15301 24565 15335 24599
rect 15669 24565 15703 24599
rect 16405 24565 16439 24599
rect 18245 24565 18279 24599
rect 8401 24361 8435 24395
rect 9505 24361 9539 24395
rect 10425 24361 10459 24395
rect 11529 24361 11563 24395
rect 11989 24361 12023 24395
rect 13093 24361 13127 24395
rect 15485 24361 15519 24395
rect 17693 24361 17727 24395
rect 18797 24361 18831 24395
rect 22201 24361 22235 24395
rect 23305 24361 23339 24395
rect 1961 24293 1995 24327
rect 1685 24225 1719 24259
rect 4077 24225 4111 24259
rect 4629 24225 4663 24259
rect 5540 24225 5574 24259
rect 8493 24225 8527 24259
rect 10333 24225 10367 24259
rect 11897 24225 11931 24259
rect 13461 24225 13495 24259
rect 15301 24225 15335 24259
rect 16405 24225 16439 24259
rect 17509 24225 17543 24259
rect 18613 24225 18647 24259
rect 20913 24225 20947 24259
rect 22017 24225 22051 24259
rect 23121 24225 23155 24259
rect 3249 24157 3283 24191
rect 5273 24157 5307 24191
rect 7941 24157 7975 24191
rect 8677 24157 8711 24191
rect 10517 24157 10551 24191
rect 12173 24157 12207 24191
rect 13553 24157 13587 24191
rect 13737 24157 13771 24191
rect 9965 24089 9999 24123
rect 13001 24089 13035 24123
rect 16589 24089 16623 24123
rect 21097 24089 21131 24123
rect 4261 24021 4295 24055
rect 6653 24021 6687 24055
rect 7205 24021 7239 24055
rect 8033 24021 8067 24055
rect 14105 24021 14139 24055
rect 2329 23817 2363 23851
rect 5365 23817 5399 23851
rect 8401 23817 8435 23851
rect 9045 23817 9079 23851
rect 9321 23817 9355 23851
rect 11253 23817 11287 23851
rect 11897 23817 11931 23851
rect 14933 23817 14967 23851
rect 16773 23817 16807 23851
rect 18245 23817 18279 23851
rect 19349 23817 19383 23851
rect 20453 23817 20487 23851
rect 21557 23817 21591 23851
rect 22661 23817 22695 23851
rect 23857 23817 23891 23851
rect 12633 23749 12667 23783
rect 1777 23681 1811 23715
rect 3157 23681 3191 23715
rect 7021 23681 7055 23715
rect 16221 23681 16255 23715
rect 18613 23681 18647 23715
rect 1501 23613 1535 23647
rect 5641 23613 5675 23647
rect 9873 23613 9907 23647
rect 12449 23613 12483 23647
rect 13001 23613 13035 23647
rect 13553 23613 13587 23647
rect 16037 23613 16071 23647
rect 18061 23613 18095 23647
rect 19165 23613 19199 23647
rect 19717 23613 19751 23647
rect 20269 23613 20303 23647
rect 21373 23613 21407 23647
rect 21925 23613 21959 23647
rect 22477 23613 22511 23647
rect 23029 23613 23063 23647
rect 23673 23613 23707 23647
rect 24225 23613 24259 23647
rect 3065 23545 3099 23579
rect 3424 23545 3458 23579
rect 6653 23545 6687 23579
rect 7266 23545 7300 23579
rect 10140 23545 10174 23579
rect 13820 23545 13854 23579
rect 15853 23545 15887 23579
rect 18981 23545 19015 23579
rect 2697 23477 2731 23511
rect 4537 23477 4571 23511
rect 5825 23477 5859 23511
rect 6193 23477 6227 23511
rect 9781 23477 9815 23511
rect 12265 23477 12299 23511
rect 13369 23477 13403 23511
rect 15485 23477 15519 23511
rect 17509 23477 17543 23511
rect 20085 23477 20119 23511
rect 20913 23477 20947 23511
rect 22293 23477 22327 23511
rect 23397 23477 23431 23511
rect 1869 23273 1903 23307
rect 2421 23273 2455 23307
rect 7021 23273 7055 23307
rect 8493 23273 8527 23307
rect 9505 23273 9539 23307
rect 10057 23273 10091 23307
rect 11621 23273 11655 23307
rect 14105 23273 14139 23307
rect 15761 23273 15795 23307
rect 19625 23273 19659 23307
rect 10508 23205 10542 23239
rect 12265 23205 12299 23239
rect 12633 23205 12667 23239
rect 17141 23205 17175 23239
rect 21189 23205 21223 23239
rect 22753 23205 22787 23239
rect 1409 23137 1443 23171
rect 2789 23137 2823 23171
rect 4333 23137 4367 23171
rect 6101 23137 6135 23171
rect 7113 23137 7147 23171
rect 7380 23137 7414 23171
rect 12992 23137 13026 23171
rect 15669 23137 15703 23171
rect 16865 23137 16899 23171
rect 18153 23137 18187 23171
rect 18429 23137 18463 23171
rect 19441 23137 19475 23171
rect 20913 23137 20947 23171
rect 22477 23137 22511 23171
rect 2329 23069 2363 23103
rect 2881 23069 2915 23103
rect 2973 23069 3007 23103
rect 4077 23069 4111 23103
rect 9137 23069 9171 23103
rect 10241 23069 10275 23103
rect 12725 23069 12759 23103
rect 15945 23069 15979 23103
rect 3525 22933 3559 22967
rect 5457 22933 5491 22967
rect 15301 22933 15335 22967
rect 16313 22933 16347 22967
rect 2421 22729 2455 22763
rect 2973 22729 3007 22763
rect 5641 22729 5675 22763
rect 7021 22729 7055 22763
rect 8493 22729 8527 22763
rect 10517 22729 10551 22763
rect 12817 22729 12851 22763
rect 13277 22729 13311 22763
rect 14933 22729 14967 22763
rect 19441 22729 19475 22763
rect 20913 22729 20947 22763
rect 2789 22661 2823 22695
rect 4537 22661 4571 22695
rect 16865 22661 16899 22695
rect 1961 22593 1995 22627
rect 3617 22593 3651 22627
rect 5181 22593 5215 22627
rect 7573 22593 7607 22627
rect 8033 22593 8067 22627
rect 13185 22593 13219 22627
rect 13737 22593 13771 22627
rect 13921 22593 13955 22627
rect 15485 22593 15519 22627
rect 1685 22525 1719 22559
rect 3985 22525 4019 22559
rect 4997 22525 5031 22559
rect 6285 22525 6319 22559
rect 8585 22525 8619 22559
rect 8841 22525 8875 22559
rect 13645 22525 13679 22559
rect 22477 22525 22511 22559
rect 4445 22457 4479 22491
rect 6653 22457 6687 22491
rect 10977 22457 11011 22491
rect 14657 22457 14691 22491
rect 15730 22457 15764 22491
rect 17417 22457 17451 22491
rect 3341 22389 3375 22423
rect 3433 22389 3467 22423
rect 4905 22389 4939 22423
rect 7389 22389 7423 22423
rect 7481 22389 7515 22423
rect 9965 22389 9999 22423
rect 11069 22389 11103 22423
rect 12265 22389 12299 22423
rect 15301 22389 15335 22423
rect 18245 22389 18279 22423
rect 11345 22185 11379 22219
rect 12633 22185 12667 22219
rect 13737 22185 13771 22219
rect 15301 22185 15335 22219
rect 3433 22117 3467 22151
rect 5172 22117 5206 22151
rect 8033 22117 8067 22151
rect 1593 22049 1627 22083
rect 1869 22049 1903 22083
rect 2513 22049 2547 22083
rect 2881 22049 2915 22083
rect 10149 22049 10183 22083
rect 13829 22049 13863 22083
rect 14105 22049 14139 22083
rect 15301 22049 15335 22083
rect 15393 22049 15427 22083
rect 15660 22049 15694 22083
rect 4905 21981 4939 22015
rect 8125 21981 8159 22015
rect 8309 21981 8343 22015
rect 10241 21981 10275 22015
rect 10425 21981 10459 22015
rect 15117 21981 15151 22015
rect 6285 21913 6319 21947
rect 7573 21913 7607 21947
rect 9781 21913 9815 21947
rect 3065 21845 3099 21879
rect 3893 21845 3927 21879
rect 4537 21845 4571 21879
rect 7113 21845 7147 21879
rect 7665 21845 7699 21879
rect 8769 21845 8803 21879
rect 9045 21845 9079 21879
rect 10793 21845 10827 21879
rect 12541 21845 12575 21879
rect 13277 21845 13311 21879
rect 16773 21845 16807 21879
rect 2881 21641 2915 21675
rect 4169 21641 4203 21675
rect 5273 21641 5307 21675
rect 6653 21641 6687 21675
rect 7389 21641 7423 21675
rect 11345 21641 11379 21675
rect 12173 21573 12207 21607
rect 2145 21505 2179 21539
rect 3157 21505 3191 21539
rect 4813 21505 4847 21539
rect 5733 21505 5767 21539
rect 10609 21505 10643 21539
rect 13001 21505 13035 21539
rect 14013 21505 14047 21539
rect 1869 21437 1903 21471
rect 4077 21437 4111 21471
rect 4629 21437 4663 21471
rect 7481 21437 7515 21471
rect 10425 21437 10459 21471
rect 7748 21369 7782 21403
rect 9413 21369 9447 21403
rect 10333 21369 10367 21403
rect 10977 21369 11011 21403
rect 12909 21369 12943 21403
rect 14258 21369 14292 21403
rect 1777 21301 1811 21335
rect 3617 21301 3651 21335
rect 4537 21301 4571 21335
rect 5641 21301 5675 21335
rect 6193 21301 6227 21335
rect 8861 21301 8895 21335
rect 9781 21301 9815 21335
rect 9965 21301 9999 21335
rect 11897 21301 11931 21335
rect 12449 21301 12483 21335
rect 12817 21301 12851 21335
rect 13461 21301 13495 21335
rect 13829 21301 13863 21335
rect 15393 21301 15427 21335
rect 15945 21301 15979 21335
rect 16405 21301 16439 21335
rect 1593 21097 1627 21131
rect 4353 21097 4387 21131
rect 8401 21097 8435 21131
rect 12081 21097 12115 21131
rect 12909 21097 12943 21131
rect 14013 21097 14047 21131
rect 15761 21097 15795 21131
rect 2237 21029 2271 21063
rect 5150 21029 5184 21063
rect 9965 21029 9999 21063
rect 1961 20961 1995 20995
rect 2789 20961 2823 20995
rect 3157 20961 3191 20995
rect 4813 20961 4847 20995
rect 4905 20961 4939 20995
rect 7757 20961 7791 20995
rect 10324 20961 10358 20995
rect 15669 20961 15703 20995
rect 7849 20893 7883 20927
rect 8033 20893 8067 20927
rect 10057 20893 10091 20927
rect 12449 20893 12483 20927
rect 13001 20893 13035 20927
rect 13093 20893 13127 20927
rect 14197 20893 14231 20927
rect 15853 20893 15887 20927
rect 7297 20825 7331 20859
rect 12541 20825 12575 20859
rect 15301 20825 15335 20859
rect 6285 20757 6319 20791
rect 6837 20757 6871 20791
rect 7389 20757 7423 20791
rect 9045 20757 9079 20791
rect 9413 20757 9447 20791
rect 11437 20757 11471 20791
rect 13553 20757 13587 20791
rect 1685 20553 1719 20587
rect 2513 20553 2547 20587
rect 8953 20553 8987 20587
rect 11897 20553 11931 20587
rect 12265 20553 12299 20587
rect 14013 20553 14047 20587
rect 14565 20553 14599 20587
rect 16129 20553 16163 20587
rect 4353 20485 4387 20519
rect 8769 20485 8803 20519
rect 2053 20417 2087 20451
rect 4721 20417 4755 20451
rect 5365 20417 5399 20451
rect 1777 20349 1811 20383
rect 3065 20349 3099 20383
rect 3985 20349 4019 20383
rect 5273 20349 5307 20383
rect 6285 20349 6319 20383
rect 6561 20349 6595 20383
rect 6837 20349 6871 20383
rect 7093 20349 7127 20383
rect 5181 20281 5215 20315
rect 5825 20281 5859 20315
rect 15117 20485 15151 20519
rect 12449 20417 12483 20451
rect 15761 20417 15795 20451
rect 16497 20417 16531 20451
rect 16681 20417 16715 20451
rect 9321 20349 9355 20383
rect 12633 20349 12667 20383
rect 15485 20349 15519 20383
rect 9566 20281 9600 20315
rect 12449 20281 12483 20315
rect 12878 20281 12912 20315
rect 2881 20213 2915 20247
rect 3249 20213 3283 20247
rect 4813 20213 4847 20247
rect 6377 20213 6411 20247
rect 8217 20213 8251 20247
rect 8953 20213 8987 20247
rect 9229 20213 9263 20247
rect 10701 20213 10735 20247
rect 11253 20213 11287 20247
rect 15025 20213 15059 20247
rect 15577 20213 15611 20247
rect 3893 20009 3927 20043
rect 4353 20009 4387 20043
rect 5917 20009 5951 20043
rect 6285 20009 6319 20043
rect 7849 20009 7883 20043
rect 8861 20009 8895 20043
rect 10149 20009 10183 20043
rect 12725 20009 12759 20043
rect 13277 20009 13311 20043
rect 15117 20009 15151 20043
rect 16037 20009 16071 20043
rect 16773 20009 16807 20043
rect 1685 19941 1719 19975
rect 2973 19941 3007 19975
rect 6929 19941 6963 19975
rect 14105 19941 14139 19975
rect 1409 19873 1443 19907
rect 2697 19873 2731 19907
rect 4721 19873 4755 19907
rect 4813 19873 4847 19907
rect 6377 19873 6411 19907
rect 7941 19873 7975 19907
rect 9229 19873 9263 19907
rect 11601 19873 11635 19907
rect 13829 19873 13863 19907
rect 15301 19873 15335 19907
rect 15577 19873 15611 19907
rect 16589 19873 16623 19907
rect 2237 19805 2271 19839
rect 4997 19805 5031 19839
rect 6561 19805 6595 19839
rect 8033 19805 8067 19839
rect 10241 19805 10275 19839
rect 10333 19805 10367 19839
rect 11345 19805 11379 19839
rect 5825 19737 5859 19771
rect 7481 19737 7515 19771
rect 9781 19737 9815 19771
rect 2513 19669 2547 19703
rect 3433 19669 3467 19703
rect 5365 19669 5399 19703
rect 7389 19669 7423 19703
rect 8585 19669 8619 19703
rect 9045 19669 9079 19703
rect 10885 19669 10919 19703
rect 11253 19669 11287 19703
rect 6561 19465 6595 19499
rect 9873 19465 9907 19499
rect 11805 19465 11839 19499
rect 13001 19465 13035 19499
rect 17325 19465 17359 19499
rect 10793 19397 10827 19431
rect 2145 19329 2179 19363
rect 7297 19329 7331 19363
rect 7481 19329 7515 19363
rect 8953 19329 8987 19363
rect 10333 19329 10367 19363
rect 11345 19329 11379 19363
rect 13553 19329 13587 19363
rect 1869 19261 1903 19295
rect 3065 19261 3099 19295
rect 5549 19261 5583 19295
rect 6193 19261 6227 19295
rect 8309 19261 8343 19295
rect 8769 19261 8803 19295
rect 9505 19261 9539 19295
rect 11253 19261 11287 19295
rect 14841 19261 14875 19295
rect 15393 19261 15427 19295
rect 3310 19193 3344 19227
rect 7941 19193 7975 19227
rect 10701 19193 10735 19227
rect 11161 19193 11195 19227
rect 12173 19193 12207 19227
rect 12909 19193 12943 19227
rect 13369 19193 13403 19227
rect 15301 19193 15335 19227
rect 15660 19193 15694 19227
rect 1501 19125 1535 19159
rect 1961 19125 1995 19159
rect 2605 19125 2639 19159
rect 2973 19125 3007 19159
rect 4445 19125 4479 19159
rect 4997 19125 5031 19159
rect 5365 19125 5399 19159
rect 5733 19125 5767 19159
rect 6837 19125 6871 19159
rect 7205 19125 7239 19159
rect 8401 19125 8435 19159
rect 8861 19125 8895 19159
rect 13461 19125 13495 19159
rect 14013 19125 14047 19159
rect 14565 19125 14599 19159
rect 16773 19125 16807 19159
rect 1409 18921 1443 18955
rect 2789 18921 2823 18955
rect 2973 18921 3007 18955
rect 7757 18921 7791 18955
rect 8125 18921 8159 18955
rect 8769 18921 8803 18955
rect 9229 18921 9263 18955
rect 9965 18921 9999 18955
rect 10517 18921 10551 18955
rect 11621 18921 11655 18955
rect 13645 18921 13679 18955
rect 16681 18921 16715 18955
rect 3433 18853 3467 18887
rect 4629 18853 4663 18887
rect 5181 18853 5215 18887
rect 6000 18853 6034 18887
rect 11437 18853 11471 18887
rect 12081 18853 12115 18887
rect 1777 18785 1811 18819
rect 3801 18785 3835 18819
rect 4537 18785 4571 18819
rect 5733 18785 5767 18819
rect 8217 18785 8251 18819
rect 10425 18785 10459 18819
rect 11989 18785 12023 18819
rect 13553 18785 13587 18819
rect 14013 18785 14047 18819
rect 14105 18785 14139 18819
rect 15025 18785 15059 18819
rect 15568 18785 15602 18819
rect 1869 18717 1903 18751
rect 2053 18717 2087 18751
rect 4721 18717 4755 18751
rect 10609 18717 10643 18751
rect 12173 18717 12207 18751
rect 14289 18717 14323 18751
rect 15301 18717 15335 18751
rect 8401 18649 8435 18683
rect 2513 18581 2547 18615
rect 4169 18581 4203 18615
rect 5549 18581 5583 18615
rect 7113 18581 7147 18615
rect 10057 18581 10091 18615
rect 11161 18581 11195 18615
rect 12633 18581 12667 18615
rect 13093 18581 13127 18615
rect 4169 18377 4203 18411
rect 4537 18377 4571 18411
rect 5181 18377 5215 18411
rect 8493 18377 8527 18411
rect 9597 18377 9631 18411
rect 11897 18377 11931 18411
rect 14933 18377 14967 18411
rect 14381 18309 14415 18343
rect 14749 18309 14783 18343
rect 5089 18241 5123 18275
rect 5733 18241 5767 18275
rect 6561 18241 6595 18275
rect 9689 18241 9723 18275
rect 11345 18241 11379 18275
rect 12173 18241 12207 18275
rect 15393 18241 15427 18275
rect 15577 18241 15611 18275
rect 2053 18173 2087 18207
rect 5641 18173 5675 18207
rect 7113 18173 7147 18207
rect 7369 18173 7403 18207
rect 11161 18173 11195 18207
rect 12449 18173 12483 18207
rect 12705 18173 12739 18207
rect 1961 18105 1995 18139
rect 2320 18105 2354 18139
rect 10241 18105 10275 18139
rect 10609 18105 10643 18139
rect 15301 18105 15335 18139
rect 16497 18105 16531 18139
rect 3433 18037 3467 18071
rect 5549 18037 5583 18071
rect 6193 18037 6227 18071
rect 9137 18037 9171 18071
rect 10793 18037 10827 18071
rect 11253 18037 11287 18071
rect 13829 18037 13863 18071
rect 15945 18037 15979 18071
rect 16405 18037 16439 18071
rect 2789 17833 2823 17867
rect 6929 17833 6963 17867
rect 9689 17833 9723 17867
rect 10701 17833 10735 17867
rect 12173 17833 12207 17867
rect 12725 17833 12759 17867
rect 13737 17833 13771 17867
rect 15025 17833 15059 17867
rect 4690 17765 4724 17799
rect 11060 17765 11094 17799
rect 15669 17765 15703 17799
rect 2881 17697 2915 17731
rect 4445 17697 4479 17731
rect 7297 17697 7331 17731
rect 13645 17697 13679 17731
rect 16313 17697 16347 17731
rect 17233 17697 17267 17731
rect 1685 17629 1719 17663
rect 3065 17629 3099 17663
rect 7389 17629 7423 17663
rect 7481 17629 7515 17663
rect 8493 17629 8527 17663
rect 10793 17629 10827 17663
rect 13185 17629 13219 17663
rect 13829 17629 13863 17663
rect 15761 17629 15795 17663
rect 15945 17629 15979 17663
rect 17325 17629 17359 17663
rect 17509 17629 17543 17663
rect 3433 17561 3467 17595
rect 6745 17561 6779 17595
rect 9321 17561 9355 17595
rect 13277 17561 13311 17595
rect 1961 17493 1995 17527
rect 2421 17493 2455 17527
rect 3893 17493 3927 17527
rect 4353 17493 4387 17527
rect 5825 17493 5859 17527
rect 6377 17493 6411 17527
rect 8033 17493 8067 17527
rect 8401 17493 8435 17527
rect 8953 17493 8987 17527
rect 10149 17493 10183 17527
rect 14381 17493 14415 17527
rect 15301 17493 15335 17527
rect 16681 17493 16715 17527
rect 16865 17493 16899 17527
rect 1409 17289 1443 17323
rect 2421 17289 2455 17323
rect 4169 17289 4203 17323
rect 4721 17289 4755 17323
rect 6837 17289 6871 17323
rect 7849 17289 7883 17323
rect 8677 17289 8711 17323
rect 10149 17289 10183 17323
rect 10885 17289 10919 17323
rect 14473 17289 14507 17323
rect 17417 17289 17451 17323
rect 18245 17289 18279 17323
rect 2881 17221 2915 17255
rect 4629 17221 4663 17255
rect 2053 17153 2087 17187
rect 3801 17153 3835 17187
rect 5273 17153 5307 17187
rect 6285 17153 6319 17187
rect 7389 17153 7423 17187
rect 12265 17153 12299 17187
rect 14933 17153 14967 17187
rect 3617 17085 3651 17119
rect 5733 17085 5767 17119
rect 7297 17085 7331 17119
rect 8769 17085 8803 17119
rect 9025 17085 9059 17119
rect 12541 17085 12575 17119
rect 12808 17085 12842 17119
rect 15025 17085 15059 17119
rect 16957 17085 16991 17119
rect 17693 17085 17727 17119
rect 1777 17017 1811 17051
rect 5181 17017 5215 17051
rect 15270 17017 15304 17051
rect 1869 16949 1903 16983
rect 3157 16949 3191 16983
rect 3525 16949 3559 16983
rect 5089 16949 5123 16983
rect 6561 16949 6595 16983
rect 7205 16949 7239 16983
rect 8309 16949 8343 16983
rect 11253 16949 11287 16983
rect 11713 16949 11747 16983
rect 13921 16949 13955 16983
rect 16405 16949 16439 16983
rect 17509 16949 17543 16983
rect 2881 16745 2915 16779
rect 3525 16745 3559 16779
rect 4905 16745 4939 16779
rect 5457 16745 5491 16779
rect 7573 16745 7607 16779
rect 9873 16745 9907 16779
rect 10241 16745 10275 16779
rect 10885 16745 10919 16779
rect 11161 16745 11195 16779
rect 12633 16745 12667 16779
rect 13645 16745 13679 16779
rect 15761 16745 15795 16779
rect 17233 16745 17267 16779
rect 17877 16745 17911 16779
rect 4353 16677 4387 16711
rect 6469 16677 6503 16711
rect 6929 16677 6963 16711
rect 8309 16677 8343 16711
rect 9229 16677 9263 16711
rect 13093 16677 13127 16711
rect 14105 16677 14139 16711
rect 14749 16677 14783 16711
rect 15669 16677 15703 16711
rect 1501 16609 1535 16643
rect 1768 16609 1802 16643
rect 4077 16609 4111 16643
rect 5825 16609 5859 16643
rect 7205 16609 7239 16643
rect 8217 16609 8251 16643
rect 8953 16609 8987 16643
rect 9689 16609 9723 16643
rect 11529 16609 11563 16643
rect 11621 16609 11655 16643
rect 12173 16609 12207 16643
rect 13369 16609 13403 16643
rect 13461 16609 13495 16643
rect 14013 16609 14047 16643
rect 5917 16541 5951 16575
rect 6101 16541 6135 16575
rect 8493 16541 8527 16575
rect 11805 16541 11839 16575
rect 14289 16541 14323 16575
rect 15853 16541 15887 16575
rect 17325 16541 17359 16575
rect 17509 16541 17543 16575
rect 15301 16473 15335 16507
rect 3801 16405 3835 16439
rect 5273 16405 5307 16439
rect 7849 16405 7883 16439
rect 13185 16405 13219 16439
rect 13461 16405 13495 16439
rect 15025 16405 15059 16439
rect 16497 16405 16531 16439
rect 16865 16405 16899 16439
rect 4629 16201 4663 16235
rect 7021 16201 7055 16235
rect 8033 16201 8067 16235
rect 8309 16201 8343 16235
rect 9689 16201 9723 16235
rect 10793 16201 10827 16235
rect 11805 16201 11839 16235
rect 13185 16201 13219 16235
rect 13645 16201 13679 16235
rect 17141 16201 17175 16235
rect 3617 16133 3651 16167
rect 2605 16065 2639 16099
rect 3157 16065 3191 16099
rect 4261 16065 4295 16099
rect 5825 16065 5859 16099
rect 7573 16065 7607 16099
rect 2421 15997 2455 16031
rect 4077 15997 4111 16031
rect 6101 15997 6135 16031
rect 1961 15929 1995 15963
rect 2513 15929 2547 15963
rect 5641 15929 5675 15963
rect 12725 16133 12759 16167
rect 9229 16065 9263 16099
rect 10701 16065 10735 16099
rect 11253 16065 11287 16099
rect 11345 16065 11379 16099
rect 14289 16065 14323 16099
rect 8401 15997 8435 16031
rect 9045 15997 9079 16031
rect 14013 15997 14047 16031
rect 14105 15997 14139 16031
rect 15209 15997 15243 16031
rect 6561 15929 6595 15963
rect 7481 15929 7515 15963
rect 8309 15929 8343 15963
rect 8953 15929 8987 15963
rect 13461 15929 13495 15963
rect 15476 15929 15510 15963
rect 2053 15861 2087 15895
rect 3525 15861 3559 15895
rect 3985 15861 4019 15895
rect 4997 15861 5031 15895
rect 5181 15861 5215 15895
rect 5549 15861 5583 15895
rect 6101 15861 6135 15895
rect 6285 15861 6319 15895
rect 7389 15861 7423 15895
rect 8585 15861 8619 15895
rect 9965 15861 9999 15895
rect 11161 15861 11195 15895
rect 12173 15861 12207 15895
rect 14749 15861 14783 15895
rect 15117 15861 15151 15895
rect 16589 15861 16623 15895
rect 17601 15861 17635 15895
rect 18337 15861 18371 15895
rect 1777 15657 1811 15691
rect 2145 15657 2179 15691
rect 3709 15657 3743 15691
rect 4445 15657 4479 15691
rect 5641 15657 5675 15691
rect 7205 15657 7239 15691
rect 7757 15657 7791 15691
rect 8217 15657 8251 15691
rect 9137 15657 9171 15691
rect 9689 15657 9723 15691
rect 10149 15657 10183 15691
rect 10793 15657 10827 15691
rect 11161 15657 11195 15691
rect 11437 15657 11471 15691
rect 12449 15657 12483 15691
rect 13001 15657 13035 15691
rect 13461 15657 13495 15691
rect 14105 15657 14139 15691
rect 15025 15657 15059 15691
rect 15577 15657 15611 15691
rect 15853 15657 15887 15691
rect 16405 15657 16439 15691
rect 16865 15657 16899 15691
rect 18061 15657 18095 15691
rect 18521 15657 18555 15691
rect 5181 15589 5215 15623
rect 11897 15589 11931 15623
rect 12817 15589 12851 15623
rect 16957 15589 16991 15623
rect 17509 15589 17543 15623
rect 2789 15521 2823 15555
rect 4537 15521 4571 15555
rect 6561 15521 6595 15555
rect 8125 15521 8159 15555
rect 10057 15521 10091 15555
rect 11805 15521 11839 15555
rect 13369 15521 13403 15555
rect 18429 15521 18463 15555
rect 2881 15453 2915 15487
rect 3065 15453 3099 15487
rect 4629 15453 4663 15487
rect 6009 15453 6043 15487
rect 6653 15453 6687 15487
rect 6837 15453 6871 15487
rect 8309 15453 8343 15487
rect 10333 15453 10367 15487
rect 11989 15453 12023 15487
rect 13645 15453 13679 15487
rect 17141 15453 17175 15487
rect 18613 15453 18647 15487
rect 2421 15385 2455 15419
rect 16497 15385 16531 15419
rect 4077 15317 4111 15351
rect 6193 15317 6227 15351
rect 7573 15317 7607 15351
rect 8861 15317 8895 15351
rect 14381 15317 14415 15351
rect 17877 15317 17911 15351
rect 4721 15113 4755 15147
rect 6837 15113 6871 15147
rect 8309 15113 8343 15147
rect 10793 15113 10827 15147
rect 11805 15113 11839 15147
rect 12173 15113 12207 15147
rect 12725 15113 12759 15147
rect 15025 15113 15059 15147
rect 16405 15113 16439 15147
rect 17509 15113 17543 15147
rect 13369 15045 13403 15079
rect 15945 15045 15979 15079
rect 17877 15045 17911 15079
rect 1685 14977 1719 15011
rect 5181 14977 5215 15011
rect 5365 14977 5399 15011
rect 7481 14977 7515 15011
rect 16865 14977 16899 15011
rect 16957 14977 16991 15011
rect 7205 14909 7239 14943
rect 8769 14909 8803 14943
rect 13645 14909 13679 14943
rect 13912 14909 13946 14943
rect 16313 14909 16347 14943
rect 18061 14909 18095 14943
rect 1952 14841 1986 14875
rect 4629 14841 4663 14875
rect 5089 14841 5123 14875
rect 5917 14841 5951 14875
rect 7941 14841 7975 14875
rect 8677 14841 8711 14875
rect 9014 14841 9048 14875
rect 18306 14841 18340 14875
rect 3065 14773 3099 14807
rect 3801 14773 3835 14807
rect 4169 14773 4203 14807
rect 6193 14773 6227 14807
rect 6561 14773 6595 14807
rect 7297 14773 7331 14807
rect 10149 14773 10183 14807
rect 11069 14773 11103 14807
rect 11437 14773 11471 14807
rect 13001 14773 13035 14807
rect 16773 14773 16807 14807
rect 19441 14773 19475 14807
rect 1409 14569 1443 14603
rect 2421 14569 2455 14603
rect 3801 14569 3835 14603
rect 6101 14569 6135 14603
rect 8953 14569 8987 14603
rect 10885 14569 10919 14603
rect 12633 14569 12667 14603
rect 13645 14569 13679 14603
rect 14013 14569 14047 14603
rect 18337 14569 18371 14603
rect 18889 14569 18923 14603
rect 2881 14501 2915 14535
rect 6469 14501 6503 14535
rect 9321 14501 9355 14535
rect 10057 14501 10091 14535
rect 13553 14501 13587 14535
rect 14105 14501 14139 14535
rect 15669 14501 15703 14535
rect 2789 14433 2823 14467
rect 4436 14433 4470 14467
rect 6920 14433 6954 14467
rect 9781 14433 9815 14467
rect 11437 14433 11471 14467
rect 15761 14433 15795 14467
rect 16589 14433 16623 14467
rect 17224 14433 17258 14467
rect 2329 14365 2363 14399
rect 3065 14365 3099 14399
rect 4169 14365 4203 14399
rect 6653 14365 6687 14399
rect 11529 14365 11563 14399
rect 11713 14365 11747 14399
rect 14289 14365 14323 14399
rect 15025 14365 15059 14399
rect 15945 14365 15979 14399
rect 16957 14365 16991 14399
rect 3433 14297 3467 14331
rect 8033 14297 8067 14331
rect 11069 14297 11103 14331
rect 13185 14297 13219 14331
rect 1869 14229 1903 14263
rect 5549 14229 5583 14263
rect 8677 14229 8711 14263
rect 12081 14229 12115 14263
rect 12449 14229 12483 14263
rect 15301 14229 15335 14263
rect 1409 14025 1443 14059
rect 2513 14025 2547 14059
rect 4169 14025 4203 14059
rect 6009 14025 6043 14059
rect 6377 14025 6411 14059
rect 7481 14025 7515 14059
rect 8953 14025 8987 14059
rect 9781 14025 9815 14059
rect 10793 14025 10827 14059
rect 11805 14025 11839 14059
rect 13829 14025 13863 14059
rect 14381 14025 14415 14059
rect 15945 14025 15979 14059
rect 17417 14025 17451 14059
rect 25513 14025 25547 14059
rect 2789 13957 2823 13991
rect 5733 13957 5767 13991
rect 16313 13957 16347 13991
rect 2053 13889 2087 13923
rect 4721 13889 4755 13923
rect 4905 13889 4939 13923
rect 10333 13889 10367 13923
rect 11345 13889 11379 13923
rect 12173 13889 12207 13923
rect 15393 13889 15427 13923
rect 15577 13889 15611 13923
rect 16773 13889 16807 13923
rect 24041 13889 24075 13923
rect 2973 13821 3007 13855
rect 3249 13821 3283 13855
rect 5273 13821 5307 13855
rect 7113 13821 7147 13855
rect 7573 13821 7607 13855
rect 7840 13821 7874 13855
rect 10701 13821 10735 13855
rect 11253 13821 11287 13855
rect 12449 13821 12483 13855
rect 12716 13821 12750 13855
rect 17141 13821 17175 13855
rect 18337 13821 18371 13855
rect 18705 13821 18739 13855
rect 24133 13821 24167 13855
rect 24400 13821 24434 13855
rect 4629 13753 4663 13787
rect 11161 13753 11195 13787
rect 14749 13753 14783 13787
rect 15301 13753 15335 13787
rect 1777 13685 1811 13719
rect 1869 13685 1903 13719
rect 3709 13685 3743 13719
rect 4261 13685 4295 13719
rect 14933 13685 14967 13719
rect 17785 13685 17819 13719
rect 2421 13481 2455 13515
rect 3525 13481 3559 13515
rect 5549 13481 5583 13515
rect 7113 13481 7147 13515
rect 8585 13481 8619 13515
rect 8861 13481 8895 13515
rect 9229 13481 9263 13515
rect 11621 13481 11655 13515
rect 12081 13481 12115 13515
rect 14289 13481 14323 13515
rect 15025 13481 15059 13515
rect 16681 13481 16715 13515
rect 24133 13481 24167 13515
rect 2789 13413 2823 13447
rect 5089 13413 5123 13447
rect 6285 13413 6319 13447
rect 2053 13345 2087 13379
rect 2881 13345 2915 13379
rect 3801 13345 3835 13379
rect 4445 13345 4479 13379
rect 4537 13345 4571 13379
rect 5641 13345 5675 13379
rect 7481 13345 7515 13379
rect 9689 13345 9723 13379
rect 9956 13345 9990 13379
rect 12817 13345 12851 13379
rect 15301 13345 15335 13379
rect 15568 13345 15602 13379
rect 18153 13345 18187 13379
rect 2973 13277 3007 13311
rect 4629 13277 4663 13311
rect 7573 13277 7607 13311
rect 7665 13277 7699 13311
rect 18245 13277 18279 13311
rect 18337 13277 18371 13311
rect 4077 13209 4111 13243
rect 5825 13209 5859 13243
rect 1685 13141 1719 13175
rect 6561 13141 6595 13175
rect 7021 13141 7055 13175
rect 8125 13141 8159 13175
rect 11069 13141 11103 13175
rect 12449 13141 12483 13175
rect 17233 13141 17267 13175
rect 17601 13141 17635 13175
rect 17785 13141 17819 13175
rect 18797 13141 18831 13175
rect 1409 12937 1443 12971
rect 2513 12937 2547 12971
rect 2881 12937 2915 12971
rect 5273 12937 5307 12971
rect 6193 12937 6227 12971
rect 6653 12937 6687 12971
rect 9505 12937 9539 12971
rect 10057 12937 10091 12971
rect 12265 12937 12299 12971
rect 13829 12937 13863 12971
rect 17509 12937 17543 12971
rect 18061 12937 18095 12971
rect 1869 12801 1903 12835
rect 2053 12801 2087 12835
rect 5733 12801 5767 12835
rect 7573 12801 7607 12835
rect 8125 12801 8159 12835
rect 11345 12801 11379 12835
rect 16589 12801 16623 12835
rect 18613 12801 18647 12835
rect 2973 12733 3007 12767
rect 11253 12733 11287 12767
rect 12449 12733 12483 12767
rect 12705 12733 12739 12767
rect 14197 12733 14231 12767
rect 18429 12733 18463 12767
rect 1777 12665 1811 12699
rect 3229 12665 3263 12699
rect 8033 12665 8067 12699
rect 8370 12665 8404 12699
rect 10701 12665 10735 12699
rect 11161 12665 11195 12699
rect 14464 12665 14498 12699
rect 17785 12665 17819 12699
rect 4353 12597 4387 12631
rect 4905 12597 4939 12631
rect 7021 12597 7055 12631
rect 10793 12597 10827 12631
rect 11897 12597 11931 12631
rect 15577 12597 15611 12631
rect 16129 12597 16163 12631
rect 17049 12597 17083 12631
rect 18521 12597 18555 12631
rect 19073 12597 19107 12631
rect 2881 12393 2915 12427
rect 4077 12393 4111 12427
rect 5457 12393 5491 12427
rect 6101 12393 6135 12427
rect 6469 12393 6503 12427
rect 7021 12393 7055 12427
rect 9689 12393 9723 12427
rect 11161 12393 11195 12427
rect 11345 12393 11379 12427
rect 12909 12393 12943 12427
rect 13645 12393 13679 12427
rect 14657 12393 14691 12427
rect 15025 12393 15059 12427
rect 15761 12393 15795 12427
rect 17969 12393 18003 12427
rect 18613 12393 18647 12427
rect 12817 12325 12851 12359
rect 18889 12325 18923 12359
rect 1501 12257 1535 12291
rect 1768 12257 1802 12291
rect 3893 12257 3927 12291
rect 4445 12257 4479 12291
rect 5089 12257 5123 12291
rect 7389 12257 7423 12291
rect 10057 12257 10091 12291
rect 11713 12257 11747 12291
rect 14013 12257 14047 12291
rect 16589 12257 16623 12291
rect 16856 12257 16890 12291
rect 4537 12189 4571 12223
rect 4629 12189 4663 12223
rect 5641 12189 5675 12223
rect 7481 12189 7515 12223
rect 7573 12189 7607 12223
rect 10149 12189 10183 12223
rect 10333 12189 10367 12223
rect 11805 12189 11839 12223
rect 11989 12189 12023 12223
rect 13093 12189 13127 12223
rect 13277 12189 13311 12223
rect 14105 12189 14139 12223
rect 14289 12189 14323 12223
rect 15301 12189 15335 12223
rect 9505 12121 9539 12155
rect 12449 12121 12483 12155
rect 3525 12053 3559 12087
rect 6837 12053 6871 12087
rect 8033 12053 8067 12087
rect 8401 12053 8435 12087
rect 8769 12053 8803 12087
rect 10885 12053 10919 12087
rect 13277 12053 13311 12087
rect 13553 12053 13587 12087
rect 16221 12053 16255 12087
rect 3433 11849 3467 11883
rect 4537 11849 4571 11883
rect 6285 11849 6319 11883
rect 6653 11849 6687 11883
rect 8861 11849 8895 11883
rect 9689 11849 9723 11883
rect 12081 11849 12115 11883
rect 13185 11849 13219 11883
rect 14657 11849 14691 11883
rect 15209 11849 15243 11883
rect 16129 11849 16163 11883
rect 18521 11849 18555 11883
rect 7021 11781 7055 11815
rect 4445 11713 4479 11747
rect 5089 11713 5123 11747
rect 5549 11713 5583 11747
rect 10517 11713 10551 11747
rect 13284 11713 13318 11747
rect 15669 11713 15703 11747
rect 16681 11713 16715 11747
rect 17141 11713 17175 11747
rect 2053 11645 2087 11679
rect 4077 11645 4111 11679
rect 4905 11645 4939 11679
rect 7481 11645 7515 11679
rect 10977 11645 11011 11679
rect 11437 11645 11471 11679
rect 1961 11577 1995 11611
rect 2320 11577 2354 11611
rect 4997 11577 5031 11611
rect 7748 11577 7782 11611
rect 10425 11577 10459 11611
rect 12817 11577 12851 11611
rect 13544 11577 13578 11611
rect 15945 11577 15979 11611
rect 16497 11577 16531 11611
rect 17693 11577 17727 11611
rect 9965 11509 9999 11543
rect 10333 11509 10367 11543
rect 11805 11509 11839 11543
rect 16589 11509 16623 11543
rect 18061 11509 18095 11543
rect 1961 11305 1995 11339
rect 3801 11305 3835 11339
rect 4077 11305 4111 11339
rect 5089 11305 5123 11339
rect 6101 11305 6135 11339
rect 7849 11305 7883 11339
rect 9505 11305 9539 11339
rect 11253 11305 11287 11339
rect 12725 11305 12759 11339
rect 13185 11305 13219 11339
rect 13277 11305 13311 11339
rect 15025 11305 15059 11339
rect 15485 11305 15519 11339
rect 16405 11305 16439 11339
rect 17141 11305 17175 11339
rect 1685 11237 1719 11271
rect 6714 11237 6748 11271
rect 10149 11237 10183 11271
rect 10793 11237 10827 11271
rect 14381 11237 14415 11271
rect 2789 11169 2823 11203
rect 4445 11169 4479 11203
rect 6469 11169 6503 11203
rect 8769 11169 8803 11203
rect 10057 11169 10091 11203
rect 12081 11169 12115 11203
rect 13645 11169 13679 11203
rect 17969 11169 18003 11203
rect 2881 11101 2915 11135
rect 3065 11101 3099 11135
rect 4537 11101 4571 11135
rect 4721 11101 4755 11135
rect 10333 11101 10367 11135
rect 12173 11101 12207 11135
rect 12357 11101 12391 11135
rect 13737 11101 13771 11135
rect 13829 11101 13863 11135
rect 16497 11101 16531 11135
rect 16589 11101 16623 11135
rect 18061 11101 18095 11135
rect 18153 11101 18187 11135
rect 18613 11101 18647 11135
rect 2421 11033 2455 11067
rect 3525 11033 3559 11067
rect 9689 11033 9723 11067
rect 11621 11033 11655 11067
rect 16037 11033 16071 11067
rect 17417 11033 17451 11067
rect 17601 11033 17635 11067
rect 5641 10965 5675 10999
rect 8401 10965 8435 10999
rect 11713 10965 11747 10999
rect 14657 10965 14691 10999
rect 15853 10965 15887 10999
rect 2697 10761 2731 10795
rect 5181 10761 5215 10795
rect 5549 10761 5583 10795
rect 8033 10761 8067 10795
rect 9229 10761 9263 10795
rect 11069 10761 11103 10795
rect 11713 10761 11747 10795
rect 12173 10761 12207 10795
rect 14013 10761 14047 10795
rect 16129 10761 16163 10795
rect 17693 10761 17727 10795
rect 5825 10693 5859 10727
rect 13921 10693 13955 10727
rect 2237 10625 2271 10659
rect 8585 10625 8619 10659
rect 9597 10625 9631 10659
rect 12909 10625 12943 10659
rect 13001 10625 13035 10659
rect 13553 10625 13587 10659
rect 14565 10625 14599 10659
rect 15761 10625 15795 10659
rect 16773 10625 16807 10659
rect 16957 10625 16991 10659
rect 18613 10625 18647 10659
rect 3157 10557 3191 10591
rect 5641 10557 5675 10591
rect 7573 10557 7607 10591
rect 8493 10557 8527 10591
rect 9689 10557 9723 10591
rect 9945 10557 9979 10591
rect 14381 10557 14415 10591
rect 16681 10557 16715 10591
rect 18521 10557 18555 10591
rect 3402 10489 3436 10523
rect 6837 10489 6871 10523
rect 12817 10489 12851 10523
rect 14473 10489 14507 10523
rect 18429 10489 18463 10523
rect 19073 10489 19107 10523
rect 1593 10421 1627 10455
rect 1961 10421 1995 10455
rect 2053 10421 2087 10455
rect 3065 10421 3099 10455
rect 4537 10421 4571 10455
rect 6561 10421 6595 10455
rect 7941 10421 7975 10455
rect 8401 10421 8435 10455
rect 12449 10421 12483 10455
rect 15301 10421 15335 10455
rect 16313 10421 16347 10455
rect 18061 10421 18095 10455
rect 3433 10217 3467 10251
rect 3801 10217 3835 10251
rect 5549 10217 5583 10251
rect 7757 10217 7791 10251
rect 9873 10217 9907 10251
rect 10241 10217 10275 10251
rect 13461 10217 13495 10251
rect 14105 10217 14139 10251
rect 14841 10217 14875 10251
rect 18797 10217 18831 10251
rect 2881 10149 2915 10183
rect 6000 10149 6034 10183
rect 8125 10149 8159 10183
rect 9229 10149 9263 10183
rect 10762 10149 10796 10183
rect 14381 10149 14415 10183
rect 18061 10149 18095 10183
rect 18889 10149 18923 10183
rect 2329 10081 2363 10115
rect 2789 10081 2823 10115
rect 4445 10081 4479 10115
rect 10517 10081 10551 10115
rect 13369 10081 13403 10115
rect 16201 10081 16235 10115
rect 2973 10013 3007 10047
rect 4537 10013 4571 10047
rect 4721 10013 4755 10047
rect 5733 10013 5767 10047
rect 13645 10013 13679 10047
rect 15945 10013 15979 10047
rect 18981 10013 19015 10047
rect 1685 9945 1719 9979
rect 7113 9945 7147 9979
rect 12909 9945 12943 9979
rect 18429 9945 18463 9979
rect 2421 9877 2455 9911
rect 4077 9877 4111 9911
rect 5089 9877 5123 9911
rect 8493 9877 8527 9911
rect 8861 9877 8895 9911
rect 11897 9877 11931 9911
rect 12449 9877 12483 9911
rect 13001 9877 13035 9911
rect 15761 9877 15795 9911
rect 17325 9877 17359 9911
rect 19441 9877 19475 9911
rect 19809 9877 19843 9911
rect 2513 9673 2547 9707
rect 4721 9673 4755 9707
rect 6101 9673 6135 9707
rect 6377 9605 6411 9639
rect 7113 9605 7147 9639
rect 7573 9605 7607 9639
rect 9137 9605 9171 9639
rect 15577 9605 15611 9639
rect 17509 9605 17543 9639
rect 19993 9605 20027 9639
rect 2789 9537 2823 9571
rect 5089 9537 5123 9571
rect 5549 9537 5583 9571
rect 7481 9537 7515 9571
rect 8125 9537 8159 9571
rect 9597 9537 9631 9571
rect 9781 9537 9815 9571
rect 10241 9537 10275 9571
rect 11253 9537 11287 9571
rect 16497 9537 16531 9571
rect 16589 9537 16623 9571
rect 17785 9537 17819 9571
rect 1409 9469 1443 9503
rect 1685 9469 1719 9503
rect 3056 9469 3090 9503
rect 4997 9469 5031 9503
rect 5273 9469 5307 9503
rect 8033 9469 8067 9503
rect 10609 9469 10643 9503
rect 11713 9469 11747 9503
rect 13277 9469 13311 9503
rect 16405 9469 16439 9503
rect 18061 9469 18095 9503
rect 18317 9469 18351 9503
rect 7941 9401 7975 9435
rect 8677 9401 8711 9435
rect 11161 9401 11195 9435
rect 12265 9401 12299 9435
rect 13544 9401 13578 9435
rect 4169 9333 4203 9367
rect 4997 9333 5031 9367
rect 8953 9333 8987 9367
rect 9505 9333 9539 9367
rect 10701 9333 10735 9367
rect 11069 9333 11103 9367
rect 12817 9333 12851 9367
rect 13185 9333 13219 9367
rect 14657 9333 14691 9367
rect 15853 9333 15887 9367
rect 16037 9333 16071 9367
rect 17141 9333 17175 9367
rect 19441 9333 19475 9367
rect 2789 9129 2823 9163
rect 5641 9129 5675 9163
rect 8493 9129 8527 9163
rect 9229 9129 9263 9163
rect 9873 9129 9907 9163
rect 13093 9129 13127 9163
rect 13645 9129 13679 9163
rect 16405 9129 16439 9163
rect 17969 9129 18003 9163
rect 18613 9129 18647 9163
rect 1676 9061 1710 9095
rect 4537 9061 4571 9095
rect 11406 9061 11440 9095
rect 15577 9061 15611 9095
rect 16856 9061 16890 9095
rect 1409 8993 1443 9027
rect 4445 8993 4479 9027
rect 5825 8993 5859 9027
rect 7380 8993 7414 9027
rect 14013 8993 14047 9027
rect 16589 8993 16623 9027
rect 19441 8993 19475 9027
rect 4629 8925 4663 8959
rect 7113 8925 7147 8959
rect 10057 8925 10091 8959
rect 11161 8925 11195 8959
rect 14105 8925 14139 8959
rect 14289 8925 14323 8959
rect 19533 8925 19567 8959
rect 19625 8925 19659 8959
rect 3433 8857 3467 8891
rect 5089 8857 5123 8891
rect 20085 8857 20119 8891
rect 3801 8789 3835 8823
rect 4077 8789 4111 8823
rect 5549 8789 5583 8823
rect 6193 8789 6227 8823
rect 6561 8789 6595 8823
rect 6929 8789 6963 8823
rect 10793 8789 10827 8823
rect 12541 8789 12575 8823
rect 13553 8789 13587 8823
rect 14749 8789 14783 8823
rect 15025 8789 15059 8823
rect 16037 8789 16071 8823
rect 18889 8789 18923 8823
rect 19073 8789 19107 8823
rect 20453 8789 20487 8823
rect 21189 8789 21223 8823
rect 1501 8585 1535 8619
rect 3065 8585 3099 8619
rect 9873 8585 9907 8619
rect 9965 8585 9999 8619
rect 11253 8585 11287 8619
rect 11621 8585 11655 8619
rect 13277 8585 13311 8619
rect 13553 8585 13587 8619
rect 15761 8585 15795 8619
rect 16129 8585 16163 8619
rect 17233 8585 17267 8619
rect 21189 8585 21223 8619
rect 2605 8517 2639 8551
rect 4629 8517 4663 8551
rect 6009 8517 6043 8551
rect 6469 8517 6503 8551
rect 8217 8517 8251 8551
rect 8861 8517 8895 8551
rect 13461 8517 13495 8551
rect 19073 8517 19107 8551
rect 19625 8517 19659 8551
rect 21005 8517 21039 8551
rect 1961 8449 1995 8483
rect 2145 8449 2179 8483
rect 3525 8449 3559 8483
rect 3709 8449 3743 8483
rect 5181 8449 5215 8483
rect 5641 8449 5675 8483
rect 9505 8449 9539 8483
rect 10517 8449 10551 8483
rect 12725 8449 12759 8483
rect 16865 8449 16899 8483
rect 18613 8449 18647 8483
rect 19441 8449 19475 8483
rect 20177 8449 20211 8483
rect 21741 8449 21775 8483
rect 2973 8381 3007 8415
rect 4537 8381 4571 8415
rect 6653 8381 6687 8415
rect 6837 8381 6871 8415
rect 10333 8381 10367 8415
rect 11989 8381 12023 8415
rect 12265 8381 12299 8415
rect 13461 8381 13495 8415
rect 13737 8381 13771 8415
rect 16589 8381 16623 8415
rect 19993 8381 20027 8415
rect 20085 8381 20119 8415
rect 21557 8381 21591 8415
rect 1869 8313 1903 8347
rect 4169 8313 4203 8347
rect 7082 8313 7116 8347
rect 10425 8313 10459 8347
rect 13982 8313 14016 8347
rect 16681 8313 16715 8347
rect 18429 8313 18463 8347
rect 3433 8245 3467 8279
rect 4997 8245 5031 8279
rect 5089 8245 5123 8279
rect 12081 8245 12115 8279
rect 15117 8245 15151 8279
rect 16221 8245 16255 8279
rect 17785 8245 17819 8279
rect 18061 8245 18095 8279
rect 18521 8245 18555 8279
rect 20637 8245 20671 8279
rect 21649 8245 21683 8279
rect 1685 8041 1719 8075
rect 2421 8041 2455 8075
rect 3525 8041 3559 8075
rect 3893 8041 3927 8075
rect 4629 8041 4663 8075
rect 7297 8041 7331 8075
rect 8861 8041 8895 8075
rect 10149 8041 10183 8075
rect 11069 8041 11103 8075
rect 13553 8041 13587 8075
rect 15117 8041 15151 8075
rect 19073 8041 19107 8075
rect 19165 8041 19199 8075
rect 19533 8041 19567 8075
rect 2881 7973 2915 8007
rect 2789 7905 2823 7939
rect 4077 7905 4111 7939
rect 5273 7905 5307 7939
rect 5540 7905 5574 7939
rect 8125 7905 8159 7939
rect 9689 7905 9723 7939
rect 2973 7837 3007 7871
rect 8217 7837 8251 7871
rect 8401 7837 8435 7871
rect 4905 7769 4939 7803
rect 7757 7769 7791 7803
rect 9321 7769 9355 7803
rect 14013 7973 14047 8007
rect 14933 7973 14967 8007
rect 19625 7973 19659 8007
rect 11161 7905 11195 7939
rect 11428 7905 11462 7939
rect 14105 7837 14139 7871
rect 14289 7837 14323 7871
rect 14657 7837 14691 7871
rect 15301 7905 15335 7939
rect 16681 7905 16715 7939
rect 16937 7905 16971 7939
rect 21189 7905 21223 7939
rect 19717 7837 19751 7871
rect 13185 7769 13219 7803
rect 13645 7769 13679 7803
rect 14933 7769 14967 7803
rect 15485 7769 15519 7803
rect 2329 7701 2363 7735
rect 6653 7701 6687 7735
rect 7573 7701 7607 7735
rect 10793 7701 10827 7735
rect 11069 7701 11103 7735
rect 12541 7701 12575 7735
rect 15853 7701 15887 7735
rect 16221 7701 16255 7735
rect 18061 7701 18095 7735
rect 18705 7701 18739 7735
rect 20177 7701 20211 7735
rect 20545 7701 20579 7735
rect 1685 7497 1719 7531
rect 4169 7497 4203 7531
rect 6285 7497 6319 7531
rect 6653 7497 6687 7531
rect 7849 7497 7883 7531
rect 8677 7497 8711 7531
rect 11897 7497 11931 7531
rect 13093 7497 13127 7531
rect 14197 7497 14231 7531
rect 19073 7497 19107 7531
rect 19625 7497 19659 7531
rect 21189 7497 21223 7531
rect 3617 7429 3651 7463
rect 5181 7429 5215 7463
rect 2237 7361 2271 7395
rect 5825 7361 5859 7395
rect 7389 7361 7423 7395
rect 9137 7361 9171 7395
rect 9873 7361 9907 7395
rect 10333 7361 10367 7395
rect 11345 7361 11379 7395
rect 13645 7361 13679 7395
rect 13829 7361 13863 7395
rect 17877 7361 17911 7395
rect 18613 7361 18647 7395
rect 20177 7361 20211 7395
rect 20637 7361 20671 7395
rect 21005 7361 21039 7395
rect 21741 7361 21775 7395
rect 2493 7293 2527 7327
rect 4997 7293 5031 7327
rect 5641 7293 5675 7327
rect 7205 7293 7239 7327
rect 9689 7293 9723 7327
rect 10517 7293 10551 7327
rect 11253 7293 11287 7327
rect 12725 7293 12759 7327
rect 14657 7293 14691 7327
rect 14749 7293 14783 7327
rect 17417 7293 17451 7327
rect 5549 7225 5583 7259
rect 7297 7225 7331 7259
rect 11161 7225 11195 7259
rect 14994 7225 15028 7259
rect 17141 7225 17175 7259
rect 18429 7225 18463 7259
rect 19533 7225 19567 7259
rect 19993 7225 20027 7259
rect 21649 7225 21683 7259
rect 2053 7157 2087 7191
rect 4629 7157 4663 7191
rect 6837 7157 6871 7191
rect 8217 7157 8251 7191
rect 9229 7157 9263 7191
rect 9597 7157 9631 7191
rect 10517 7157 10551 7191
rect 10609 7157 10643 7191
rect 10793 7157 10827 7191
rect 12173 7157 12207 7191
rect 13185 7157 13219 7191
rect 13553 7157 13587 7191
rect 16129 7157 16163 7191
rect 16681 7157 16715 7191
rect 17233 7157 17267 7191
rect 18061 7157 18095 7191
rect 18521 7157 18555 7191
rect 20085 7157 20119 7191
rect 21557 7157 21591 7191
rect 1777 6953 1811 6987
rect 2789 6953 2823 6987
rect 7113 6953 7147 6987
rect 8677 6953 8711 6987
rect 9321 6953 9355 6987
rect 11621 6953 11655 6987
rect 11989 6953 12023 6987
rect 12817 6953 12851 6987
rect 12909 6953 12943 6987
rect 14013 6953 14047 6987
rect 15761 6953 15795 6987
rect 19257 6953 19291 6987
rect 20177 6953 20211 6987
rect 1869 6885 1903 6919
rect 2421 6885 2455 6919
rect 7941 6885 7975 6919
rect 16681 6885 16715 6919
rect 19901 6885 19935 6919
rect 4997 6817 5031 6851
rect 5356 6817 5390 6851
rect 8033 6817 8067 6851
rect 9956 6817 9990 6851
rect 12449 6817 12483 6851
rect 13277 6817 13311 6851
rect 16129 6817 16163 6851
rect 17785 6817 17819 6851
rect 18144 6817 18178 6851
rect 1961 6749 1995 6783
rect 2973 6749 3007 6783
rect 5089 6749 5123 6783
rect 8125 6749 8159 6783
rect 9689 6749 9723 6783
rect 13369 6749 13403 6783
rect 13553 6749 13587 6783
rect 15301 6749 15335 6783
rect 16773 6749 16807 6783
rect 16865 6749 16899 6783
rect 17325 6749 17359 6783
rect 17877 6749 17911 6783
rect 21189 6749 21223 6783
rect 7573 6681 7607 6715
rect 11069 6681 11103 6715
rect 14565 6681 14599 6715
rect 16313 6681 16347 6715
rect 1409 6613 1443 6647
rect 3525 6613 3559 6647
rect 3893 6613 3927 6647
rect 4629 6613 4663 6647
rect 6469 6613 6503 6647
rect 7389 6613 7423 6647
rect 14841 6613 14875 6647
rect 20545 6613 20579 6647
rect 21557 6613 21591 6647
rect 2973 6409 3007 6443
rect 4997 6409 5031 6443
rect 7941 6409 7975 6443
rect 8309 6409 8343 6443
rect 10333 6409 10367 6443
rect 11069 6409 11103 6443
rect 11437 6409 11471 6443
rect 11805 6409 11839 6443
rect 12265 6409 12299 6443
rect 14289 6409 14323 6443
rect 16221 6409 16255 6443
rect 16405 6409 16439 6443
rect 17877 6409 17911 6443
rect 18429 6409 18463 6443
rect 20453 6409 20487 6443
rect 6561 6341 6595 6375
rect 6837 6341 6871 6375
rect 14749 6341 14783 6375
rect 20821 6341 20855 6375
rect 21005 6341 21039 6375
rect 1593 6273 1627 6307
rect 4629 6273 4663 6307
rect 5733 6273 5767 6307
rect 7297 6273 7331 6307
rect 7481 6273 7515 6307
rect 8401 6273 8435 6307
rect 10701 6273 10735 6307
rect 13737 6273 13771 6307
rect 13921 6273 13955 6307
rect 15393 6273 15427 6307
rect 15945 6273 15979 6307
rect 16957 6273 16991 6307
rect 21465 6273 21499 6307
rect 21649 6273 21683 6307
rect 6193 6205 6227 6239
rect 8668 6205 8702 6239
rect 13645 6205 13679 6239
rect 15209 6205 15243 6239
rect 18521 6205 18555 6239
rect 18777 6205 18811 6239
rect 21373 6205 21407 6239
rect 1860 6137 1894 6171
rect 3893 6137 3927 6171
rect 5549 6137 5583 6171
rect 16865 6137 16899 6171
rect 3617 6069 3651 6103
rect 4077 6069 4111 6103
rect 5089 6069 5123 6103
rect 5457 6069 5491 6103
rect 7205 6069 7239 6103
rect 9781 6069 9815 6103
rect 12909 6069 12943 6103
rect 13277 6069 13311 6103
rect 14841 6069 14875 6103
rect 15301 6069 15335 6103
rect 16773 6069 16807 6103
rect 17417 6069 17451 6103
rect 19901 6069 19935 6103
rect 22109 6069 22143 6103
rect 2881 5865 2915 5899
rect 4445 5865 4479 5899
rect 5641 5865 5675 5899
rect 6009 5865 6043 5899
rect 6929 5865 6963 5899
rect 7573 5865 7607 5899
rect 8033 5865 8067 5899
rect 10149 5865 10183 5899
rect 11345 5865 11379 5899
rect 11529 5865 11563 5899
rect 13001 5865 13035 5899
rect 13553 5865 13587 5899
rect 14105 5865 14139 5899
rect 15853 5865 15887 5899
rect 15945 5865 15979 5899
rect 16589 5865 16623 5899
rect 16865 5865 16899 5899
rect 19349 5865 19383 5899
rect 20453 5865 20487 5899
rect 1768 5797 1802 5831
rect 3801 5797 3835 5831
rect 9505 5797 9539 5831
rect 10057 5797 10091 5831
rect 10701 5797 10735 5831
rect 17294 5797 17328 5831
rect 1501 5729 1535 5763
rect 4537 5729 4571 5763
rect 6101 5729 6135 5763
rect 8401 5729 8435 5763
rect 11897 5729 11931 5763
rect 13461 5729 13495 5763
rect 14841 5729 14875 5763
rect 19533 5729 19567 5763
rect 20085 5729 20119 5763
rect 4629 5661 4663 5695
rect 6285 5661 6319 5695
rect 8493 5661 8527 5695
rect 8585 5661 8619 5695
rect 10241 5661 10275 5695
rect 11989 5661 12023 5695
rect 12081 5661 12115 5695
rect 13645 5661 13679 5695
rect 16129 5661 16163 5695
rect 17049 5661 17083 5695
rect 4077 5593 4111 5627
rect 9045 5593 9079 5627
rect 12633 5593 12667 5627
rect 3433 5525 3467 5559
rect 5273 5525 5307 5559
rect 7849 5525 7883 5559
rect 9689 5525 9723 5559
rect 13093 5525 13127 5559
rect 14565 5525 14599 5559
rect 15485 5525 15519 5559
rect 18429 5525 18463 5559
rect 18981 5525 19015 5559
rect 19717 5525 19751 5559
rect 21097 5525 21131 5559
rect 1409 5321 1443 5355
rect 2973 5321 3007 5355
rect 4169 5321 4203 5355
rect 5181 5321 5215 5355
rect 6653 5321 6687 5355
rect 11161 5321 11195 5355
rect 12173 5321 12207 5355
rect 13461 5321 13495 5355
rect 13921 5321 13955 5355
rect 14933 5321 14967 5355
rect 16313 5321 16347 5355
rect 18061 5321 18095 5355
rect 19625 5321 19659 5355
rect 20637 5321 20671 5355
rect 14197 5253 14231 5287
rect 16037 5253 16071 5287
rect 1961 5185 1995 5219
rect 2421 5185 2455 5219
rect 3617 5185 3651 5219
rect 4721 5185 4755 5219
rect 5825 5185 5859 5219
rect 7389 5185 7423 5219
rect 8585 5185 8619 5219
rect 12909 5185 12943 5219
rect 13093 5185 13127 5219
rect 15577 5185 15611 5219
rect 16773 5185 16807 5219
rect 18613 5185 18647 5219
rect 20177 5185 20211 5219
rect 1869 5117 1903 5151
rect 5089 5117 5123 5151
rect 5549 5117 5583 5151
rect 7205 5117 7239 5151
rect 11253 5117 11287 5151
rect 12817 5117 12851 5151
rect 16497 5117 16531 5151
rect 17877 5117 17911 5151
rect 18429 5117 18463 5151
rect 21189 5117 21223 5151
rect 21925 5117 21959 5151
rect 1777 5049 1811 5083
rect 8830 5049 8864 5083
rect 10517 5049 10551 5083
rect 11805 5049 11839 5083
rect 14749 5049 14783 5083
rect 15393 5049 15427 5083
rect 19993 5049 20027 5083
rect 21465 5049 21499 5083
rect 2881 4981 2915 5015
rect 3341 4981 3375 5015
rect 3433 4981 3467 5015
rect 5641 4981 5675 5015
rect 6285 4981 6319 5015
rect 6837 4981 6871 5015
rect 7297 4981 7331 5015
rect 8033 4981 8067 5015
rect 8401 4981 8435 5015
rect 9965 4981 9999 5015
rect 11437 4981 11471 5015
rect 12449 4981 12483 5015
rect 15301 4981 15335 5015
rect 17233 4981 17267 5015
rect 18521 4981 18555 5015
rect 19073 4981 19107 5015
rect 19441 4981 19475 5015
rect 20085 4981 20119 5015
rect 1685 4777 1719 4811
rect 2329 4777 2363 4811
rect 3433 4777 3467 4811
rect 3801 4777 3835 4811
rect 5641 4777 5675 4811
rect 6285 4777 6319 4811
rect 7205 4777 7239 4811
rect 8677 4777 8711 4811
rect 9505 4777 9539 4811
rect 10057 4777 10091 4811
rect 10149 4777 10183 4811
rect 13001 4777 13035 4811
rect 13645 4777 13679 4811
rect 14565 4777 14599 4811
rect 17693 4777 17727 4811
rect 18337 4777 18371 4811
rect 18613 4777 18647 4811
rect 18797 4777 18831 4811
rect 20545 4777 20579 4811
rect 3065 4709 3099 4743
rect 4506 4709 4540 4743
rect 14933 4709 14967 4743
rect 2237 4641 2271 4675
rect 4261 4641 4295 4675
rect 6929 4641 6963 4675
rect 7941 4641 7975 4675
rect 8033 4641 8067 4675
rect 11989 4641 12023 4675
rect 13553 4641 13587 4675
rect 15301 4641 15335 4675
rect 16569 4641 16603 4675
rect 19165 4641 19199 4675
rect 20913 4641 20947 4675
rect 22385 4641 22419 4675
rect 2421 4573 2455 4607
rect 8125 4573 8159 4607
rect 10241 4573 10275 4607
rect 12081 4573 12115 4607
rect 12265 4573 12299 4607
rect 13829 4573 13863 4607
rect 16313 4573 16347 4607
rect 19257 4573 19291 4607
rect 19349 4573 19383 4607
rect 19809 4573 19843 4607
rect 22661 4573 22695 4607
rect 1869 4505 1903 4539
rect 12633 4505 12667 4539
rect 7573 4437 7607 4471
rect 9045 4437 9079 4471
rect 9689 4437 9723 4471
rect 10701 4437 10735 4471
rect 11253 4437 11287 4471
rect 11621 4437 11655 4471
rect 13185 4437 13219 4471
rect 14197 4437 14231 4471
rect 15853 4437 15887 4471
rect 16221 4437 16255 4471
rect 20269 4437 20303 4471
rect 21097 4437 21131 4471
rect 6285 4233 6319 4267
rect 10701 4233 10735 4267
rect 13001 4233 13035 4267
rect 13461 4233 13495 4267
rect 16405 4233 16439 4267
rect 19165 4233 19199 4267
rect 21649 4233 21683 4267
rect 22385 4233 22419 4267
rect 2421 4097 2455 4131
rect 2881 4097 2915 4131
rect 3249 4097 3283 4131
rect 4077 4097 4111 4131
rect 5089 4097 5123 4131
rect 5641 4097 5675 4131
rect 5825 4097 5859 4131
rect 7297 4097 7331 4131
rect 7389 4097 7423 4131
rect 8769 4097 8803 4131
rect 16129 4097 16163 4131
rect 16221 4097 16255 4131
rect 16957 4097 16991 4131
rect 17417 4097 17451 4131
rect 17693 4097 17727 4131
rect 17877 4097 17911 4131
rect 18521 4097 18555 4131
rect 18705 4097 18739 4131
rect 1777 4029 1811 4063
rect 7849 4029 7883 4063
rect 11253 4029 11287 4063
rect 11805 4029 11839 4063
rect 12455 4029 12489 4063
rect 13829 4029 13863 4063
rect 15853 4029 15887 4063
rect 16865 4029 16899 4063
rect 19625 4029 19659 4063
rect 20177 4029 20211 4063
rect 20545 4029 20579 4063
rect 20729 4029 20763 4063
rect 21281 4029 21315 4063
rect 21833 4029 21867 4063
rect 23673 4029 23707 4063
rect 24225 4029 24259 4063
rect 3801 3961 3835 3995
rect 4721 3961 4755 3995
rect 5549 3961 5583 3995
rect 8677 3961 8711 3995
rect 9036 3961 9070 3995
rect 11161 3961 11195 3995
rect 12265 3961 12299 3995
rect 14074 3961 14108 3995
rect 16129 3961 16163 3995
rect 16773 3961 16807 3995
rect 17693 3961 17727 3995
rect 18429 3961 18463 3995
rect 1869 3893 1903 3927
rect 2237 3893 2271 3927
rect 2329 3893 2363 3927
rect 3433 3893 3467 3927
rect 3893 3893 3927 3927
rect 5181 3893 5215 3927
rect 6653 3893 6687 3927
rect 6837 3893 6871 3927
rect 7205 3893 7239 3927
rect 8309 3893 8343 3927
rect 10149 3893 10183 3927
rect 11437 3893 11471 3927
rect 12633 3893 12667 3927
rect 15209 3893 15243 3927
rect 18061 3893 18095 3927
rect 19533 3893 19567 3927
rect 19809 3893 19843 3927
rect 20913 3893 20947 3927
rect 22017 3893 22051 3927
rect 23857 3893 23891 3927
rect 1961 3689 1995 3723
rect 2237 3689 2271 3723
rect 2421 3689 2455 3723
rect 2789 3689 2823 3723
rect 6561 3689 6595 3723
rect 7573 3689 7607 3723
rect 8033 3689 8067 3723
rect 9689 3689 9723 3723
rect 10057 3689 10091 3723
rect 11253 3689 11287 3723
rect 11713 3689 11747 3723
rect 13737 3689 13771 3723
rect 18153 3689 18187 3723
rect 18889 3689 18923 3723
rect 19993 3689 20027 3723
rect 20361 3689 20395 3723
rect 20729 3689 20763 3723
rect 21465 3689 21499 3723
rect 2881 3621 2915 3655
rect 4322 3621 4356 3655
rect 7849 3621 7883 3655
rect 10885 3621 10919 3655
rect 15546 3621 15580 3655
rect 4077 3553 4111 3587
rect 6745 3553 6779 3587
rect 7021 3553 7055 3587
rect 8401 3553 8435 3587
rect 8493 3553 8527 3587
rect 11621 3553 11655 3587
rect 13829 3553 13863 3587
rect 15301 3553 15335 3587
rect 19165 3553 19199 3587
rect 19349 3553 19383 3587
rect 20913 3553 20947 3587
rect 22017 3553 22051 3587
rect 3065 3485 3099 3519
rect 6101 3485 6135 3519
rect 8585 3485 8619 3519
rect 9045 3485 9079 3519
rect 10149 3485 10183 3519
rect 10241 3485 10275 3519
rect 11805 3485 11839 3519
rect 12541 3485 12575 3519
rect 13921 3485 13955 3519
rect 17233 3485 17267 3519
rect 18245 3485 18279 3519
rect 18337 3485 18371 3519
rect 12817 3417 12851 3451
rect 17785 3417 17819 3451
rect 3433 3349 3467 3383
rect 3893 3349 3927 3383
rect 5457 3349 5491 3383
rect 9505 3349 9539 3383
rect 13277 3349 13311 3383
rect 13369 3349 13403 3383
rect 14565 3349 14599 3383
rect 14933 3349 14967 3383
rect 16681 3349 16715 3383
rect 17601 3349 17635 3383
rect 19533 3349 19567 3383
rect 21097 3349 21131 3383
rect 21833 3349 21867 3383
rect 22201 3349 22235 3383
rect 2513 3145 2547 3179
rect 5181 3145 5215 3179
rect 6285 3145 6319 3179
rect 9137 3145 9171 3179
rect 9321 3145 9355 3179
rect 10793 3145 10827 3179
rect 15945 3145 15979 3179
rect 16313 3145 16347 3179
rect 19073 3145 19107 3179
rect 19441 3145 19475 3179
rect 20821 3145 20855 3179
rect 21833 3145 21867 3179
rect 22569 3145 22603 3179
rect 4261 3077 4295 3111
rect 4813 3077 4847 3111
rect 5641 3077 5675 3111
rect 6561 3077 6595 3111
rect 11989 3077 12023 3111
rect 14933 3077 14967 3111
rect 22201 3077 22235 3111
rect 1685 3009 1719 3043
rect 5733 3009 5767 3043
rect 9781 3009 9815 3043
rect 9965 3009 9999 3043
rect 10333 3009 10367 3043
rect 11161 3009 11195 3043
rect 14841 3009 14875 3043
rect 15485 3009 15519 3043
rect 16773 3009 16807 3043
rect 18613 3009 18647 3043
rect 19901 3009 19935 3043
rect 1501 2941 1535 2975
rect 2881 2941 2915 2975
rect 6837 2941 6871 2975
rect 7093 2941 7127 2975
rect 9689 2941 9723 2975
rect 10885 2941 10919 2975
rect 12449 2941 12483 2975
rect 14381 2941 14415 2975
rect 15301 2941 15335 2975
rect 16497 2941 16531 2975
rect 17509 2941 17543 2975
rect 18521 2941 18555 2975
rect 19625 2941 19659 2975
rect 20361 2941 20395 2975
rect 20913 2941 20947 2975
rect 21465 2941 21499 2975
rect 22017 2941 22051 2975
rect 3126 2873 3160 2907
rect 12694 2873 12728 2907
rect 15393 2873 15427 2907
rect 17877 2873 17911 2907
rect 18429 2873 18463 2907
rect 8217 2805 8251 2839
rect 8769 2805 8803 2839
rect 11621 2805 11655 2839
rect 13829 2805 13863 2839
rect 18061 2805 18095 2839
rect 21097 2805 21131 2839
rect 2421 2601 2455 2635
rect 2881 2601 2915 2635
rect 3801 2601 3835 2635
rect 4077 2601 4111 2635
rect 4721 2601 4755 2635
rect 5641 2601 5675 2635
rect 6745 2601 6779 2635
rect 11805 2601 11839 2635
rect 13185 2601 13219 2635
rect 14197 2601 14231 2635
rect 15209 2601 15243 2635
rect 16589 2601 16623 2635
rect 18153 2601 18187 2635
rect 18797 2601 18831 2635
rect 21373 2601 21407 2635
rect 22109 2601 22143 2635
rect 1961 2533 1995 2567
rect 7472 2533 7506 2567
rect 12173 2533 12207 2567
rect 16957 2533 16991 2567
rect 19717 2533 19751 2567
rect 2329 2465 2363 2499
rect 2789 2465 2823 2499
rect 5181 2465 5215 2499
rect 5733 2465 5767 2499
rect 7205 2465 7239 2499
rect 9873 2465 9907 2499
rect 10129 2465 10163 2499
rect 13553 2465 13587 2499
rect 13645 2465 13679 2499
rect 15853 2465 15887 2499
rect 17141 2465 17175 2499
rect 18705 2465 18739 2499
rect 19901 2465 19935 2499
rect 20453 2465 20487 2499
rect 21189 2465 21223 2499
rect 21741 2465 21775 2499
rect 22293 2465 22327 2499
rect 22845 2465 22879 2499
rect 24041 2465 24075 2499
rect 24593 2465 24627 2499
rect 3065 2397 3099 2431
rect 3433 2397 3467 2431
rect 5917 2397 5951 2431
rect 6377 2397 6411 2431
rect 13737 2397 13771 2431
rect 14933 2397 14967 2431
rect 15945 2397 15979 2431
rect 16037 2397 16071 2431
rect 17693 2397 17727 2431
rect 18889 2397 18923 2431
rect 19349 2397 19383 2431
rect 5273 2329 5307 2363
rect 8585 2329 8619 2363
rect 9321 2329 9355 2363
rect 11253 2329 11287 2363
rect 13093 2329 13127 2363
rect 15485 2329 15519 2363
rect 17325 2329 17359 2363
rect 20085 2329 20119 2363
rect 22477 2329 22511 2363
rect 18337 2261 18371 2295
rect 20821 2261 20855 2295
rect 24225 2261 24259 2295
<< metal1 >>
rect 5258 27412 5264 27464
rect 5316 27452 5322 27464
rect 5350 27452 5356 27464
rect 5316 27424 5356 27452
rect 5316 27412 5322 27424
rect 5350 27412 5356 27424
rect 5408 27412 5414 27464
rect 8938 27412 8944 27464
rect 8996 27452 9002 27464
rect 9398 27452 9404 27464
rect 8996 27424 9404 27452
rect 8996 27412 9002 27424
rect 9398 27412 9404 27424
rect 9456 27412 9462 27464
rect 3510 27208 3516 27260
rect 3568 27248 3574 27260
rect 7006 27248 7012 27260
rect 3568 27220 7012 27248
rect 3568 27208 3574 27220
rect 7006 27208 7012 27220
rect 7064 27208 7070 27260
rect 4062 26528 4068 26580
rect 4120 26568 4126 26580
rect 8110 26568 8116 26580
rect 4120 26540 8116 26568
rect 4120 26528 4126 26540
rect 8110 26528 8116 26540
rect 8168 26528 8174 26580
rect 3510 26256 3516 26308
rect 3568 26296 3574 26308
rect 7190 26296 7196 26308
rect 3568 26268 7196 26296
rect 3568 26256 3574 26268
rect 7190 26256 7196 26268
rect 7248 26256 7254 26308
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1581 25483 1639 25489
rect 1581 25449 1593 25483
rect 1627 25480 1639 25483
rect 3050 25480 3056 25492
rect 1627 25452 3056 25480
rect 1627 25449 1639 25452
rect 1581 25443 1639 25449
rect 3050 25440 3056 25452
rect 3108 25440 3114 25492
rect 4062 25440 4068 25492
rect 4120 25480 4126 25492
rect 7101 25483 7159 25489
rect 7101 25480 7113 25483
rect 4120 25452 7113 25480
rect 4120 25440 4126 25452
rect 7101 25449 7113 25452
rect 7147 25449 7159 25483
rect 7101 25443 7159 25449
rect 7190 25440 7196 25492
rect 7248 25480 7254 25492
rect 8205 25483 8263 25489
rect 8205 25480 8217 25483
rect 7248 25452 8217 25480
rect 7248 25440 7254 25452
rect 8205 25449 8217 25452
rect 8251 25449 8263 25483
rect 8205 25443 8263 25449
rect 2038 25372 2044 25424
rect 2096 25412 2102 25424
rect 9490 25412 9496 25424
rect 2096 25384 9496 25412
rect 2096 25372 2102 25384
rect 9490 25372 9496 25384
rect 9548 25412 9554 25424
rect 9548 25384 9812 25412
rect 9548 25372 9554 25384
rect 1397 25347 1455 25353
rect 1397 25313 1409 25347
rect 1443 25344 1455 25347
rect 1578 25344 1584 25356
rect 1443 25316 1584 25344
rect 1443 25313 1455 25316
rect 1397 25307 1455 25313
rect 1578 25304 1584 25316
rect 1636 25304 1642 25356
rect 2501 25347 2559 25353
rect 2501 25313 2513 25347
rect 2547 25344 2559 25347
rect 2590 25344 2596 25356
rect 2547 25316 2596 25344
rect 2547 25313 2559 25316
rect 2501 25307 2559 25313
rect 2590 25304 2596 25316
rect 2648 25304 2654 25356
rect 4065 25347 4123 25353
rect 4065 25313 4077 25347
rect 4111 25344 4123 25347
rect 4430 25344 4436 25356
rect 4111 25316 4436 25344
rect 4111 25313 4123 25316
rect 4065 25307 4123 25313
rect 4430 25304 4436 25316
rect 4488 25304 4494 25356
rect 5169 25347 5227 25353
rect 5169 25313 5181 25347
rect 5215 25313 5227 25347
rect 6914 25344 6920 25356
rect 6875 25316 6920 25344
rect 5169 25307 5227 25313
rect 2866 25276 2872 25288
rect 2700 25248 2872 25276
rect 2700 25217 2728 25248
rect 2866 25236 2872 25248
rect 2924 25236 2930 25288
rect 5184 25276 5212 25307
rect 6914 25304 6920 25316
rect 6972 25304 6978 25356
rect 7742 25304 7748 25356
rect 7800 25344 7806 25356
rect 9784 25353 9812 25384
rect 8021 25347 8079 25353
rect 8021 25344 8033 25347
rect 7800 25316 8033 25344
rect 7800 25304 7806 25316
rect 8021 25313 8033 25316
rect 8067 25313 8079 25347
rect 8021 25307 8079 25313
rect 9769 25347 9827 25353
rect 9769 25313 9781 25347
rect 9815 25313 9827 25347
rect 9769 25307 9827 25313
rect 15473 25347 15531 25353
rect 15473 25313 15485 25347
rect 15519 25344 15531 25347
rect 15654 25344 15660 25356
rect 15519 25316 15660 25344
rect 15519 25313 15531 25316
rect 15473 25307 15531 25313
rect 15654 25304 15660 25316
rect 15712 25304 15718 25356
rect 5813 25279 5871 25285
rect 5813 25276 5825 25279
rect 5184 25248 5825 25276
rect 5813 25245 5825 25248
rect 5859 25276 5871 25279
rect 12618 25276 12624 25288
rect 5859 25248 12624 25276
rect 5859 25245 5871 25248
rect 5813 25239 5871 25245
rect 12618 25236 12624 25248
rect 12676 25236 12682 25288
rect 2685 25211 2743 25217
rect 2685 25177 2697 25211
rect 2731 25177 2743 25211
rect 2685 25171 2743 25177
rect 4062 25168 4068 25220
rect 4120 25208 4126 25220
rect 5353 25211 5411 25217
rect 5353 25208 5365 25211
rect 4120 25180 5365 25208
rect 4120 25168 4126 25180
rect 5353 25177 5365 25180
rect 5399 25177 5411 25211
rect 5353 25171 5411 25177
rect 7006 25168 7012 25220
rect 7064 25208 7070 25220
rect 9953 25211 10011 25217
rect 9953 25208 9965 25211
rect 7064 25180 9965 25208
rect 7064 25168 7070 25180
rect 9953 25177 9965 25180
rect 9999 25177 10011 25211
rect 9953 25171 10011 25177
rect 2041 25143 2099 25149
rect 2041 25109 2053 25143
rect 2087 25140 2099 25143
rect 2130 25140 2136 25152
rect 2087 25112 2136 25140
rect 2087 25109 2099 25112
rect 2041 25103 2099 25109
rect 2130 25100 2136 25112
rect 2188 25100 2194 25152
rect 3510 25100 3516 25152
rect 3568 25140 3574 25152
rect 4249 25143 4307 25149
rect 4249 25140 4261 25143
rect 3568 25112 4261 25140
rect 3568 25100 3574 25112
rect 4249 25109 4261 25112
rect 4295 25109 4307 25143
rect 4249 25103 4307 25109
rect 15657 25143 15715 25149
rect 15657 25109 15669 25143
rect 15703 25140 15715 25143
rect 26510 25140 26516 25152
rect 15703 25112 26516 25140
rect 15703 25109 15715 25112
rect 15657 25103 15715 25109
rect 26510 25100 26516 25112
rect 26568 25100 26574 25152
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 3326 24896 3332 24948
rect 3384 24936 3390 24948
rect 7009 24939 7067 24945
rect 7009 24936 7021 24939
rect 3384 24908 7021 24936
rect 3384 24896 3390 24908
rect 7009 24905 7021 24908
rect 7055 24905 7067 24939
rect 8110 24936 8116 24948
rect 8071 24908 8116 24936
rect 7009 24899 7067 24905
rect 8110 24896 8116 24908
rect 8168 24896 8174 24948
rect 6914 24828 6920 24880
rect 6972 24868 6978 24880
rect 7745 24871 7803 24877
rect 7745 24868 7757 24871
rect 6972 24840 7757 24868
rect 6972 24828 6978 24840
rect 7745 24837 7757 24840
rect 7791 24837 7803 24871
rect 7745 24831 7803 24837
rect 2130 24800 2136 24812
rect 1504 24772 2136 24800
rect 1504 24741 1532 24772
rect 2130 24760 2136 24772
rect 2188 24760 2194 24812
rect 5813 24803 5871 24809
rect 5813 24769 5825 24803
rect 5859 24800 5871 24803
rect 6270 24800 6276 24812
rect 5859 24772 6276 24800
rect 5859 24769 5871 24772
rect 5813 24763 5871 24769
rect 6270 24760 6276 24772
rect 6328 24760 6334 24812
rect 7469 24803 7527 24809
rect 7469 24800 7481 24803
rect 6840 24772 7481 24800
rect 1489 24735 1547 24741
rect 1489 24701 1501 24735
rect 1535 24701 1547 24735
rect 1489 24695 1547 24701
rect 1578 24692 1584 24744
rect 1636 24732 1642 24744
rect 2317 24735 2375 24741
rect 2317 24732 2329 24735
rect 1636 24704 2329 24732
rect 1636 24692 1642 24704
rect 2317 24701 2329 24704
rect 2363 24732 2375 24735
rect 2682 24732 2688 24744
rect 2363 24704 2688 24732
rect 2363 24701 2375 24704
rect 2317 24695 2375 24701
rect 2682 24692 2688 24704
rect 2740 24692 2746 24744
rect 2777 24735 2835 24741
rect 2777 24701 2789 24735
rect 2823 24732 2835 24735
rect 2958 24732 2964 24744
rect 2823 24704 2964 24732
rect 2823 24701 2835 24704
rect 2777 24695 2835 24701
rect 2958 24692 2964 24704
rect 3016 24732 3022 24744
rect 6840 24741 6868 24772
rect 7469 24769 7481 24772
rect 7515 24800 7527 24803
rect 9769 24803 9827 24809
rect 9769 24800 9781 24803
rect 7515 24772 9781 24800
rect 7515 24769 7527 24772
rect 7469 24763 7527 24769
rect 9769 24769 9781 24772
rect 9815 24769 9827 24803
rect 12618 24800 12624 24812
rect 12579 24772 12624 24800
rect 9769 24763 9827 24769
rect 12618 24760 12624 24772
rect 12676 24760 12682 24812
rect 3329 24735 3387 24741
rect 3329 24732 3341 24735
rect 3016 24704 3341 24732
rect 3016 24692 3022 24704
rect 3329 24701 3341 24704
rect 3375 24701 3387 24735
rect 3329 24695 3387 24701
rect 3881 24735 3939 24741
rect 3881 24701 3893 24735
rect 3927 24701 3939 24735
rect 3881 24695 3939 24701
rect 6825 24735 6883 24741
rect 6825 24701 6837 24735
rect 6871 24701 6883 24735
rect 6825 24695 6883 24701
rect 1762 24664 1768 24676
rect 1723 24636 1768 24664
rect 1762 24624 1768 24636
rect 1820 24624 1826 24676
rect 2498 24624 2504 24676
rect 2556 24664 2562 24676
rect 3697 24667 3755 24673
rect 3697 24664 3709 24667
rect 2556 24636 3709 24664
rect 2556 24624 2562 24636
rect 3697 24633 3709 24636
rect 3743 24664 3755 24667
rect 3896 24664 3924 24695
rect 7834 24692 7840 24744
rect 7892 24732 7898 24744
rect 7929 24735 7987 24741
rect 7929 24732 7941 24735
rect 7892 24704 7941 24732
rect 7892 24692 7898 24704
rect 7929 24701 7941 24704
rect 7975 24732 7987 24735
rect 8481 24735 8539 24741
rect 8481 24732 8493 24735
rect 7975 24704 8493 24732
rect 7975 24701 7987 24704
rect 7929 24695 7987 24701
rect 8481 24701 8493 24704
rect 8527 24701 8539 24735
rect 9490 24732 9496 24744
rect 9451 24704 9496 24732
rect 8481 24695 8539 24701
rect 9490 24692 9496 24704
rect 9548 24692 9554 24744
rect 9585 24735 9643 24741
rect 9585 24701 9597 24735
rect 9631 24732 9643 24735
rect 9950 24732 9956 24744
rect 9631 24704 9956 24732
rect 9631 24701 9643 24704
rect 9585 24695 9643 24701
rect 9950 24692 9956 24704
rect 10008 24732 10014 24744
rect 10321 24735 10379 24741
rect 10321 24732 10333 24735
rect 10008 24704 10333 24732
rect 10008 24692 10014 24704
rect 10321 24701 10333 24704
rect 10367 24701 10379 24735
rect 10321 24695 10379 24701
rect 12437 24735 12495 24741
rect 12437 24701 12449 24735
rect 12483 24732 12495 24735
rect 15105 24735 15163 24741
rect 12483 24704 13124 24732
rect 12483 24701 12495 24704
rect 12437 24695 12495 24701
rect 3743 24636 3924 24664
rect 5077 24667 5135 24673
rect 3743 24633 3755 24636
rect 3697 24627 3755 24633
rect 5077 24633 5089 24667
rect 5123 24664 5135 24667
rect 5629 24667 5687 24673
rect 5123 24636 5580 24664
rect 5123 24633 5135 24636
rect 5077 24627 5135 24633
rect 5552 24608 5580 24636
rect 5629 24633 5641 24667
rect 5675 24664 5687 24667
rect 5675 24636 6684 24664
rect 5675 24633 5687 24636
rect 5629 24627 5687 24633
rect 2590 24596 2596 24608
rect 2551 24568 2596 24596
rect 2590 24556 2596 24568
rect 2648 24556 2654 24608
rect 2961 24599 3019 24605
rect 2961 24565 2973 24599
rect 3007 24596 3019 24599
rect 3234 24596 3240 24608
rect 3007 24568 3240 24596
rect 3007 24565 3019 24568
rect 2961 24559 3019 24565
rect 3234 24556 3240 24568
rect 3292 24556 3298 24608
rect 4062 24596 4068 24608
rect 4023 24568 4068 24596
rect 4062 24556 4068 24568
rect 4120 24556 4126 24608
rect 4430 24596 4436 24608
rect 4391 24568 4436 24596
rect 4430 24556 4436 24568
rect 4488 24556 4494 24608
rect 5166 24596 5172 24608
rect 5127 24568 5172 24596
rect 5166 24556 5172 24568
rect 5224 24556 5230 24608
rect 5534 24596 5540 24608
rect 5495 24568 5540 24596
rect 5534 24556 5540 24568
rect 5592 24556 5598 24608
rect 6270 24596 6276 24608
rect 6231 24568 6276 24596
rect 6270 24556 6276 24568
rect 6328 24556 6334 24608
rect 6656 24605 6684 24636
rect 13096 24608 13124 24704
rect 15105 24701 15117 24735
rect 15151 24732 15163 24735
rect 15151 24704 15185 24732
rect 15151 24701 15163 24704
rect 15105 24695 15163 24701
rect 15013 24667 15071 24673
rect 15013 24633 15025 24667
rect 15059 24664 15071 24667
rect 15120 24664 15148 24695
rect 16114 24692 16120 24744
rect 16172 24732 16178 24744
rect 16209 24735 16267 24741
rect 16209 24732 16221 24735
rect 16172 24704 16221 24732
rect 16172 24692 16178 24704
rect 16209 24701 16221 24704
rect 16255 24732 16267 24735
rect 16761 24735 16819 24741
rect 16761 24732 16773 24735
rect 16255 24704 16773 24732
rect 16255 24701 16267 24704
rect 16209 24695 16267 24701
rect 16761 24701 16773 24704
rect 16807 24701 16819 24735
rect 16761 24695 16819 24701
rect 18049 24735 18107 24741
rect 18049 24701 18061 24735
rect 18095 24732 18107 24735
rect 18138 24732 18144 24744
rect 18095 24704 18144 24732
rect 18095 24701 18107 24704
rect 18049 24695 18107 24701
rect 18138 24692 18144 24704
rect 18196 24732 18202 24744
rect 18601 24735 18659 24741
rect 18601 24732 18613 24735
rect 18196 24704 18613 24732
rect 18196 24692 18202 24704
rect 18601 24701 18613 24704
rect 18647 24701 18659 24735
rect 18601 24695 18659 24701
rect 15378 24664 15384 24676
rect 15059 24636 15384 24664
rect 15059 24633 15071 24636
rect 15013 24627 15071 24633
rect 15378 24624 15384 24636
rect 15436 24624 15442 24676
rect 16482 24664 16488 24676
rect 15488 24636 16488 24664
rect 6641 24599 6699 24605
rect 6641 24565 6653 24599
rect 6687 24596 6699 24599
rect 6822 24596 6828 24608
rect 6687 24568 6828 24596
rect 6687 24565 6699 24568
rect 6641 24559 6699 24565
rect 6822 24556 6828 24568
rect 6880 24556 6886 24608
rect 8846 24596 8852 24608
rect 8807 24568 8852 24596
rect 8846 24556 8852 24568
rect 8904 24556 8910 24608
rect 13078 24556 13084 24608
rect 13136 24596 13142 24608
rect 13173 24599 13231 24605
rect 13173 24596 13185 24599
rect 13136 24568 13185 24596
rect 13136 24556 13142 24568
rect 13173 24565 13185 24568
rect 13219 24565 13231 24599
rect 13630 24596 13636 24608
rect 13591 24568 13636 24596
rect 13173 24559 13231 24565
rect 13630 24556 13636 24568
rect 13688 24556 13694 24608
rect 15289 24599 15347 24605
rect 15289 24565 15301 24599
rect 15335 24596 15347 24599
rect 15488 24596 15516 24636
rect 16482 24624 16488 24636
rect 16540 24624 16546 24676
rect 15654 24596 15660 24608
rect 15335 24568 15516 24596
rect 15615 24568 15660 24596
rect 15335 24565 15347 24568
rect 15289 24559 15347 24565
rect 15654 24556 15660 24568
rect 15712 24556 15718 24608
rect 16390 24596 16396 24608
rect 16351 24568 16396 24596
rect 16390 24556 16396 24568
rect 16448 24556 16454 24608
rect 18230 24596 18236 24608
rect 18191 24568 18236 24596
rect 18230 24556 18236 24568
rect 18288 24556 18294 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 2866 24352 2872 24404
rect 2924 24392 2930 24404
rect 3142 24392 3148 24404
rect 2924 24364 3148 24392
rect 2924 24352 2930 24364
rect 3142 24352 3148 24364
rect 3200 24352 3206 24404
rect 4890 24352 4896 24404
rect 4948 24392 4954 24404
rect 8389 24395 8447 24401
rect 8389 24392 8401 24395
rect 4948 24364 8401 24392
rect 4948 24352 4954 24364
rect 8389 24361 8401 24364
rect 8435 24392 8447 24395
rect 9306 24392 9312 24404
rect 8435 24364 9312 24392
rect 8435 24361 8447 24364
rect 8389 24355 8447 24361
rect 9306 24352 9312 24364
rect 9364 24352 9370 24404
rect 9493 24395 9551 24401
rect 9493 24361 9505 24395
rect 9539 24392 9551 24395
rect 10413 24395 10471 24401
rect 10413 24392 10425 24395
rect 9539 24364 10425 24392
rect 9539 24361 9551 24364
rect 9493 24355 9551 24361
rect 10413 24361 10425 24364
rect 10459 24392 10471 24395
rect 11517 24395 11575 24401
rect 11517 24392 11529 24395
rect 10459 24364 11529 24392
rect 10459 24361 10471 24364
rect 10413 24355 10471 24361
rect 11517 24361 11529 24364
rect 11563 24361 11575 24395
rect 11517 24355 11575 24361
rect 11977 24395 12035 24401
rect 11977 24361 11989 24395
rect 12023 24392 12035 24395
rect 12066 24392 12072 24404
rect 12023 24364 12072 24392
rect 12023 24361 12035 24364
rect 11977 24355 12035 24361
rect 12066 24352 12072 24364
rect 12124 24352 12130 24404
rect 13078 24392 13084 24404
rect 13039 24364 13084 24392
rect 13078 24352 13084 24364
rect 13136 24352 13142 24404
rect 15473 24395 15531 24401
rect 15473 24361 15485 24395
rect 15519 24392 15531 24395
rect 16206 24392 16212 24404
rect 15519 24364 16212 24392
rect 15519 24361 15531 24364
rect 15473 24355 15531 24361
rect 16206 24352 16212 24364
rect 16264 24352 16270 24404
rect 17681 24395 17739 24401
rect 17681 24361 17693 24395
rect 17727 24392 17739 24395
rect 18506 24392 18512 24404
rect 17727 24364 18512 24392
rect 17727 24361 17739 24364
rect 17681 24355 17739 24361
rect 18506 24352 18512 24364
rect 18564 24352 18570 24404
rect 18782 24392 18788 24404
rect 18743 24364 18788 24392
rect 18782 24352 18788 24364
rect 18840 24352 18846 24404
rect 22189 24395 22247 24401
rect 22189 24361 22201 24395
rect 22235 24392 22247 24395
rect 23106 24392 23112 24404
rect 22235 24364 23112 24392
rect 22235 24361 22247 24364
rect 22189 24355 22247 24361
rect 23106 24352 23112 24364
rect 23164 24352 23170 24404
rect 23290 24392 23296 24404
rect 23251 24364 23296 24392
rect 23290 24352 23296 24364
rect 23348 24352 23354 24404
rect 1946 24324 1952 24336
rect 1907 24296 1952 24324
rect 1946 24284 1952 24296
rect 2004 24284 2010 24336
rect 1670 24256 1676 24268
rect 1631 24228 1676 24256
rect 1670 24216 1676 24228
rect 1728 24216 1734 24268
rect 2222 24216 2228 24268
rect 2280 24256 2286 24268
rect 4065 24259 4123 24265
rect 4065 24256 4077 24259
rect 2280 24228 4077 24256
rect 2280 24216 2286 24228
rect 4065 24225 4077 24228
rect 4111 24256 4123 24259
rect 4617 24259 4675 24265
rect 4617 24256 4629 24259
rect 4111 24228 4629 24256
rect 4111 24225 4123 24228
rect 4065 24219 4123 24225
rect 4617 24225 4629 24228
rect 4663 24225 4675 24259
rect 4617 24219 4675 24225
rect 5528 24259 5586 24265
rect 5528 24225 5540 24259
rect 5574 24256 5586 24259
rect 6270 24256 6276 24268
rect 5574 24228 6276 24256
rect 5574 24225 5586 24228
rect 5528 24219 5586 24225
rect 6270 24216 6276 24228
rect 6328 24216 6334 24268
rect 8481 24259 8539 24265
rect 8481 24225 8493 24259
rect 8527 24256 8539 24259
rect 9030 24256 9036 24268
rect 8527 24228 9036 24256
rect 8527 24225 8539 24228
rect 8481 24219 8539 24225
rect 9030 24216 9036 24228
rect 9088 24216 9094 24268
rect 10318 24256 10324 24268
rect 10279 24228 10324 24256
rect 10318 24216 10324 24228
rect 10376 24216 10382 24268
rect 11885 24259 11943 24265
rect 11885 24225 11897 24259
rect 11931 24256 11943 24259
rect 12250 24256 12256 24268
rect 11931 24228 12256 24256
rect 11931 24225 11943 24228
rect 11885 24219 11943 24225
rect 12250 24216 12256 24228
rect 12308 24216 12314 24268
rect 13354 24216 13360 24268
rect 13412 24256 13418 24268
rect 13449 24259 13507 24265
rect 13449 24256 13461 24259
rect 13412 24228 13461 24256
rect 13412 24216 13418 24228
rect 13449 24225 13461 24228
rect 13495 24225 13507 24259
rect 15286 24256 15292 24268
rect 15247 24228 15292 24256
rect 13449 24219 13507 24225
rect 15286 24216 15292 24228
rect 15344 24216 15350 24268
rect 16390 24256 16396 24268
rect 16351 24228 16396 24256
rect 16390 24216 16396 24228
rect 16448 24216 16454 24268
rect 17494 24256 17500 24268
rect 17455 24228 17500 24256
rect 17494 24216 17500 24228
rect 17552 24216 17558 24268
rect 18506 24216 18512 24268
rect 18564 24256 18570 24268
rect 18601 24259 18659 24265
rect 18601 24256 18613 24259
rect 18564 24228 18613 24256
rect 18564 24216 18570 24228
rect 18601 24225 18613 24228
rect 18647 24225 18659 24259
rect 18601 24219 18659 24225
rect 20806 24216 20812 24268
rect 20864 24256 20870 24268
rect 20901 24259 20959 24265
rect 20901 24256 20913 24259
rect 20864 24228 20913 24256
rect 20864 24216 20870 24228
rect 20901 24225 20913 24228
rect 20947 24225 20959 24259
rect 22002 24256 22008 24268
rect 21963 24228 22008 24256
rect 20901 24219 20959 24225
rect 22002 24216 22008 24228
rect 22060 24216 22066 24268
rect 23109 24259 23167 24265
rect 23109 24225 23121 24259
rect 23155 24256 23167 24259
rect 23290 24256 23296 24268
rect 23155 24228 23296 24256
rect 23155 24225 23167 24228
rect 23109 24219 23167 24225
rect 23290 24216 23296 24228
rect 23348 24216 23354 24268
rect 3237 24191 3295 24197
rect 3237 24157 3249 24191
rect 3283 24188 3295 24191
rect 3326 24188 3332 24200
rect 3283 24160 3332 24188
rect 3283 24157 3295 24160
rect 3237 24151 3295 24157
rect 3326 24148 3332 24160
rect 3384 24188 3390 24200
rect 5261 24191 5319 24197
rect 5261 24188 5273 24191
rect 3384 24160 5273 24188
rect 3384 24148 3390 24160
rect 5261 24157 5273 24160
rect 5307 24157 5319 24191
rect 5261 24151 5319 24157
rect 7929 24191 7987 24197
rect 7929 24157 7941 24191
rect 7975 24188 7987 24191
rect 8662 24188 8668 24200
rect 7975 24160 8668 24188
rect 7975 24157 7987 24160
rect 7929 24151 7987 24157
rect 8662 24148 8668 24160
rect 8720 24148 8726 24200
rect 10134 24148 10140 24200
rect 10192 24188 10198 24200
rect 10505 24191 10563 24197
rect 10505 24188 10517 24191
rect 10192 24160 10517 24188
rect 10192 24148 10198 24160
rect 10505 24157 10517 24160
rect 10551 24157 10563 24191
rect 10505 24151 10563 24157
rect 12161 24191 12219 24197
rect 12161 24157 12173 24191
rect 12207 24188 12219 24191
rect 12342 24188 12348 24200
rect 12207 24160 12348 24188
rect 12207 24157 12219 24160
rect 12161 24151 12219 24157
rect 12342 24148 12348 24160
rect 12400 24148 12406 24200
rect 13538 24188 13544 24200
rect 13499 24160 13544 24188
rect 13538 24148 13544 24160
rect 13596 24148 13602 24200
rect 13722 24188 13728 24200
rect 13683 24160 13728 24188
rect 13722 24148 13728 24160
rect 13780 24148 13786 24200
rect 9950 24120 9956 24132
rect 9911 24092 9956 24120
rect 9950 24080 9956 24092
rect 10008 24080 10014 24132
rect 12986 24120 12992 24132
rect 12899 24092 12992 24120
rect 12986 24080 12992 24092
rect 13044 24120 13050 24132
rect 13740 24120 13768 24148
rect 13044 24092 13768 24120
rect 16577 24123 16635 24129
rect 13044 24080 13050 24092
rect 16577 24089 16589 24123
rect 16623 24120 16635 24123
rect 17862 24120 17868 24132
rect 16623 24092 17868 24120
rect 16623 24089 16635 24092
rect 16577 24083 16635 24089
rect 17862 24080 17868 24092
rect 17920 24080 17926 24132
rect 21085 24123 21143 24129
rect 21085 24089 21097 24123
rect 21131 24120 21143 24123
rect 22462 24120 22468 24132
rect 21131 24092 22468 24120
rect 21131 24089 21143 24092
rect 21085 24083 21143 24089
rect 22462 24080 22468 24092
rect 22520 24080 22526 24132
rect 3970 24012 3976 24064
rect 4028 24052 4034 24064
rect 4249 24055 4307 24061
rect 4249 24052 4261 24055
rect 4028 24024 4261 24052
rect 4028 24012 4034 24024
rect 4249 24021 4261 24024
rect 4295 24021 4307 24055
rect 6638 24052 6644 24064
rect 6599 24024 6644 24052
rect 4249 24015 4307 24021
rect 6638 24012 6644 24024
rect 6696 24012 6702 24064
rect 7006 24012 7012 24064
rect 7064 24052 7070 24064
rect 7193 24055 7251 24061
rect 7193 24052 7205 24055
rect 7064 24024 7205 24052
rect 7064 24012 7070 24024
rect 7193 24021 7205 24024
rect 7239 24021 7251 24055
rect 7193 24015 7251 24021
rect 8021 24055 8079 24061
rect 8021 24021 8033 24055
rect 8067 24052 8079 24055
rect 8110 24052 8116 24064
rect 8067 24024 8116 24052
rect 8067 24021 8079 24024
rect 8021 24015 8079 24021
rect 8110 24012 8116 24024
rect 8168 24012 8174 24064
rect 13814 24012 13820 24064
rect 13872 24052 13878 24064
rect 14093 24055 14151 24061
rect 14093 24052 14105 24055
rect 13872 24024 14105 24052
rect 13872 24012 13878 24024
rect 14093 24021 14105 24024
rect 14139 24021 14151 24055
rect 14093 24015 14151 24021
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 2317 23851 2375 23857
rect 2317 23817 2329 23851
rect 2363 23848 2375 23851
rect 2406 23848 2412 23860
rect 2363 23820 2412 23848
rect 2363 23817 2375 23820
rect 2317 23811 2375 23817
rect 1762 23712 1768 23724
rect 1723 23684 1768 23712
rect 1762 23672 1768 23684
rect 1820 23672 1826 23724
rect 1489 23647 1547 23653
rect 1489 23613 1501 23647
rect 1535 23644 1547 23647
rect 2332 23644 2360 23811
rect 2406 23808 2412 23820
rect 2464 23808 2470 23860
rect 3326 23848 3332 23860
rect 3160 23820 3332 23848
rect 3160 23721 3188 23820
rect 3326 23808 3332 23820
rect 3384 23808 3390 23860
rect 5353 23851 5411 23857
rect 5353 23817 5365 23851
rect 5399 23848 5411 23851
rect 6270 23848 6276 23860
rect 5399 23820 6276 23848
rect 5399 23817 5411 23820
rect 5353 23811 5411 23817
rect 6270 23808 6276 23820
rect 6328 23848 6334 23860
rect 8389 23851 8447 23857
rect 8389 23848 8401 23851
rect 6328 23820 8401 23848
rect 6328 23808 6334 23820
rect 8389 23817 8401 23820
rect 8435 23817 8447 23851
rect 9030 23848 9036 23860
rect 8991 23820 9036 23848
rect 8389 23811 8447 23817
rect 9030 23808 9036 23820
rect 9088 23808 9094 23860
rect 9306 23848 9312 23860
rect 9267 23820 9312 23848
rect 9306 23808 9312 23820
rect 9364 23808 9370 23860
rect 11238 23848 11244 23860
rect 11199 23820 11244 23848
rect 11238 23808 11244 23820
rect 11296 23808 11302 23860
rect 11885 23851 11943 23857
rect 11885 23817 11897 23851
rect 11931 23848 11943 23851
rect 12066 23848 12072 23860
rect 11931 23820 12072 23848
rect 11931 23817 11943 23820
rect 11885 23811 11943 23817
rect 12066 23808 12072 23820
rect 12124 23808 12130 23860
rect 13722 23808 13728 23860
rect 13780 23848 13786 23860
rect 14921 23851 14979 23857
rect 14921 23848 14933 23851
rect 13780 23820 14933 23848
rect 13780 23808 13786 23820
rect 14921 23817 14933 23820
rect 14967 23817 14979 23851
rect 14921 23811 14979 23817
rect 16390 23808 16396 23860
rect 16448 23848 16454 23860
rect 16761 23851 16819 23857
rect 16761 23848 16773 23851
rect 16448 23820 16773 23848
rect 16448 23808 16454 23820
rect 16761 23817 16773 23820
rect 16807 23817 16819 23851
rect 16761 23811 16819 23817
rect 18233 23851 18291 23857
rect 18233 23817 18245 23851
rect 18279 23848 18291 23851
rect 19058 23848 19064 23860
rect 18279 23820 19064 23848
rect 18279 23817 18291 23820
rect 18233 23811 18291 23817
rect 19058 23808 19064 23820
rect 19116 23808 19122 23860
rect 19337 23851 19395 23857
rect 19337 23817 19349 23851
rect 19383 23848 19395 23851
rect 19518 23848 19524 23860
rect 19383 23820 19524 23848
rect 19383 23817 19395 23820
rect 19337 23811 19395 23817
rect 19518 23808 19524 23820
rect 19576 23808 19582 23860
rect 20441 23851 20499 23857
rect 20441 23817 20453 23851
rect 20487 23848 20499 23851
rect 21358 23848 21364 23860
rect 20487 23820 21364 23848
rect 20487 23817 20499 23820
rect 20441 23811 20499 23817
rect 21358 23808 21364 23820
rect 21416 23808 21422 23860
rect 21545 23851 21603 23857
rect 21545 23817 21557 23851
rect 21591 23848 21603 23851
rect 21910 23848 21916 23860
rect 21591 23820 21916 23848
rect 21591 23817 21603 23820
rect 21545 23811 21603 23817
rect 21910 23808 21916 23820
rect 21968 23808 21974 23860
rect 22649 23851 22707 23857
rect 22649 23817 22661 23851
rect 22695 23848 22707 23851
rect 23658 23848 23664 23860
rect 22695 23820 23664 23848
rect 22695 23817 22707 23820
rect 22649 23811 22707 23817
rect 23658 23808 23664 23820
rect 23716 23808 23722 23860
rect 23845 23851 23903 23857
rect 23845 23817 23857 23851
rect 23891 23848 23903 23851
rect 25314 23848 25320 23860
rect 23891 23820 25320 23848
rect 23891 23817 23903 23820
rect 23845 23811 23903 23817
rect 25314 23808 25320 23820
rect 25372 23808 25378 23860
rect 12618 23780 12624 23792
rect 12579 23752 12624 23780
rect 12618 23740 12624 23752
rect 12676 23740 12682 23792
rect 3145 23715 3203 23721
rect 3145 23681 3157 23715
rect 3191 23681 3203 23715
rect 7006 23712 7012 23724
rect 6967 23684 7012 23712
rect 3145 23675 3203 23681
rect 7006 23672 7012 23684
rect 7064 23672 7070 23724
rect 15378 23672 15384 23724
rect 15436 23712 15442 23724
rect 16209 23715 16267 23721
rect 16209 23712 16221 23715
rect 15436 23684 16221 23712
rect 15436 23672 15442 23684
rect 16209 23681 16221 23684
rect 16255 23681 16267 23715
rect 18601 23715 18659 23721
rect 18601 23712 18613 23715
rect 16209 23675 16267 23681
rect 18064 23684 18613 23712
rect 18064 23656 18092 23684
rect 18601 23681 18613 23684
rect 18647 23681 18659 23715
rect 18601 23675 18659 23681
rect 1535 23616 2360 23644
rect 5629 23647 5687 23653
rect 1535 23613 1547 23616
rect 1489 23607 1547 23613
rect 5629 23613 5641 23647
rect 5675 23644 5687 23647
rect 9861 23647 9919 23653
rect 5675 23616 6132 23644
rect 5675 23613 5687 23616
rect 5629 23607 5687 23613
rect 3053 23579 3111 23585
rect 3053 23545 3065 23579
rect 3099 23576 3111 23579
rect 3412 23579 3470 23585
rect 3412 23576 3424 23579
rect 3099 23548 3424 23576
rect 3099 23545 3111 23548
rect 3053 23539 3111 23545
rect 3412 23545 3424 23548
rect 3458 23576 3470 23579
rect 3458 23548 4108 23576
rect 3458 23545 3470 23548
rect 3412 23539 3470 23545
rect 4080 23520 4108 23548
rect 6104 23520 6132 23616
rect 9861 23613 9873 23647
rect 9907 23644 9919 23647
rect 9950 23644 9956 23656
rect 9907 23616 9956 23644
rect 9907 23613 9919 23616
rect 9861 23607 9919 23613
rect 9950 23604 9956 23616
rect 10008 23604 10014 23656
rect 12066 23604 12072 23656
rect 12124 23644 12130 23656
rect 12437 23647 12495 23653
rect 12437 23644 12449 23647
rect 12124 23616 12449 23644
rect 12124 23604 12130 23616
rect 12437 23613 12449 23616
rect 12483 23644 12495 23647
rect 12989 23647 13047 23653
rect 12989 23644 13001 23647
rect 12483 23616 13001 23644
rect 12483 23613 12495 23616
rect 12437 23607 12495 23613
rect 12989 23613 13001 23616
rect 13035 23613 13047 23647
rect 12989 23607 13047 23613
rect 13541 23647 13599 23653
rect 13541 23613 13553 23647
rect 13587 23644 13599 23647
rect 13630 23644 13636 23656
rect 13587 23616 13636 23644
rect 13587 23613 13599 23616
rect 13541 23607 13599 23613
rect 13630 23604 13636 23616
rect 13688 23604 13694 23656
rect 16025 23647 16083 23653
rect 16025 23613 16037 23647
rect 16071 23613 16083 23647
rect 18046 23644 18052 23656
rect 18007 23616 18052 23644
rect 16025 23607 16083 23613
rect 6641 23579 6699 23585
rect 6641 23545 6653 23579
rect 6687 23576 6699 23579
rect 7254 23579 7312 23585
rect 7254 23576 7266 23579
rect 6687 23548 7266 23576
rect 6687 23545 6699 23548
rect 6641 23539 6699 23545
rect 7254 23545 7266 23548
rect 7300 23576 7312 23579
rect 7558 23576 7564 23588
rect 7300 23548 7564 23576
rect 7300 23545 7312 23548
rect 7254 23539 7312 23545
rect 7558 23536 7564 23548
rect 7616 23536 7622 23588
rect 10134 23585 10140 23588
rect 10128 23576 10140 23585
rect 10095 23548 10140 23576
rect 10128 23539 10140 23548
rect 10134 23536 10140 23539
rect 10192 23536 10198 23588
rect 10318 23536 10324 23588
rect 10376 23536 10382 23588
rect 13808 23579 13866 23585
rect 13808 23545 13820 23579
rect 13854 23576 13866 23579
rect 13906 23576 13912 23588
rect 13854 23548 13912 23576
rect 13854 23545 13866 23548
rect 13808 23539 13866 23545
rect 13906 23536 13912 23548
rect 13964 23536 13970 23588
rect 15841 23579 15899 23585
rect 15841 23576 15853 23579
rect 14660 23548 15853 23576
rect 2682 23508 2688 23520
rect 2643 23480 2688 23508
rect 2682 23468 2688 23480
rect 2740 23468 2746 23520
rect 4062 23468 4068 23520
rect 4120 23468 4126 23520
rect 4338 23468 4344 23520
rect 4396 23508 4402 23520
rect 4525 23511 4583 23517
rect 4525 23508 4537 23511
rect 4396 23480 4537 23508
rect 4396 23468 4402 23480
rect 4525 23477 4537 23480
rect 4571 23477 4583 23511
rect 5810 23508 5816 23520
rect 5771 23480 5816 23508
rect 4525 23471 4583 23477
rect 5810 23468 5816 23480
rect 5868 23468 5874 23520
rect 6086 23468 6092 23520
rect 6144 23508 6150 23520
rect 6181 23511 6239 23517
rect 6181 23508 6193 23511
rect 6144 23480 6193 23508
rect 6144 23468 6150 23480
rect 6181 23477 6193 23480
rect 6227 23477 6239 23511
rect 6181 23471 6239 23477
rect 9769 23511 9827 23517
rect 9769 23477 9781 23511
rect 9815 23508 9827 23511
rect 10336 23508 10364 23536
rect 10962 23508 10968 23520
rect 9815 23480 10968 23508
rect 9815 23477 9827 23480
rect 9769 23471 9827 23477
rect 10962 23468 10968 23480
rect 11020 23468 11026 23520
rect 12250 23508 12256 23520
rect 12211 23480 12256 23508
rect 12250 23468 12256 23480
rect 12308 23468 12314 23520
rect 13354 23508 13360 23520
rect 13315 23480 13360 23508
rect 13354 23468 13360 23480
rect 13412 23468 13418 23520
rect 13446 23468 13452 23520
rect 13504 23508 13510 23520
rect 14660 23508 14688 23548
rect 15841 23545 15853 23548
rect 15887 23576 15899 23579
rect 16040 23576 16068 23607
rect 18046 23604 18052 23616
rect 18104 23604 18110 23656
rect 18414 23604 18420 23656
rect 18472 23644 18478 23656
rect 19153 23647 19211 23653
rect 19153 23644 19165 23647
rect 18472 23616 19165 23644
rect 18472 23604 18478 23616
rect 19153 23613 19165 23616
rect 19199 23644 19211 23647
rect 19705 23647 19763 23653
rect 19705 23644 19717 23647
rect 19199 23616 19717 23644
rect 19199 23613 19211 23616
rect 19153 23607 19211 23613
rect 19705 23613 19717 23616
rect 19751 23613 19763 23647
rect 20257 23647 20315 23653
rect 20257 23644 20269 23647
rect 19705 23607 19763 23613
rect 20088 23616 20269 23644
rect 15887 23548 16068 23576
rect 15887 23545 15899 23548
rect 15841 23539 15899 23545
rect 18506 23536 18512 23588
rect 18564 23576 18570 23588
rect 18969 23579 19027 23585
rect 18969 23576 18981 23579
rect 18564 23548 18981 23576
rect 18564 23536 18570 23548
rect 18969 23545 18981 23548
rect 19015 23545 19027 23579
rect 18969 23539 19027 23545
rect 20088 23520 20116 23616
rect 20257 23613 20269 23616
rect 20303 23613 20315 23647
rect 21358 23644 21364 23656
rect 21319 23616 21364 23644
rect 20257 23607 20315 23613
rect 21358 23604 21364 23616
rect 21416 23644 21422 23656
rect 21913 23647 21971 23653
rect 21913 23644 21925 23647
rect 21416 23616 21925 23644
rect 21416 23604 21422 23616
rect 21913 23613 21925 23616
rect 21959 23613 21971 23647
rect 21913 23607 21971 23613
rect 22370 23604 22376 23656
rect 22428 23644 22434 23656
rect 22465 23647 22523 23653
rect 22465 23644 22477 23647
rect 22428 23616 22477 23644
rect 22428 23604 22434 23616
rect 22465 23613 22477 23616
rect 22511 23644 22523 23647
rect 23017 23647 23075 23653
rect 23017 23644 23029 23647
rect 22511 23616 23029 23644
rect 22511 23613 22523 23616
rect 22465 23607 22523 23613
rect 23017 23613 23029 23616
rect 23063 23613 23075 23647
rect 23017 23607 23075 23613
rect 23474 23604 23480 23656
rect 23532 23644 23538 23656
rect 23661 23647 23719 23653
rect 23661 23644 23673 23647
rect 23532 23616 23673 23644
rect 23532 23604 23538 23616
rect 23661 23613 23673 23616
rect 23707 23644 23719 23647
rect 24213 23647 24271 23653
rect 24213 23644 24225 23647
rect 23707 23616 24225 23644
rect 23707 23613 23719 23616
rect 23661 23607 23719 23613
rect 24213 23613 24225 23616
rect 24259 23613 24271 23647
rect 24213 23607 24271 23613
rect 13504 23480 14688 23508
rect 13504 23468 13510 23480
rect 15194 23468 15200 23520
rect 15252 23508 15258 23520
rect 15473 23511 15531 23517
rect 15473 23508 15485 23511
rect 15252 23480 15485 23508
rect 15252 23468 15258 23480
rect 15473 23477 15485 23480
rect 15519 23477 15531 23511
rect 15473 23471 15531 23477
rect 17126 23468 17132 23520
rect 17184 23508 17190 23520
rect 17494 23508 17500 23520
rect 17184 23480 17500 23508
rect 17184 23468 17190 23480
rect 17494 23468 17500 23480
rect 17552 23468 17558 23520
rect 20070 23508 20076 23520
rect 20031 23480 20076 23508
rect 20070 23468 20076 23480
rect 20128 23468 20134 23520
rect 20806 23468 20812 23520
rect 20864 23508 20870 23520
rect 20901 23511 20959 23517
rect 20901 23508 20913 23511
rect 20864 23480 20913 23508
rect 20864 23468 20870 23480
rect 20901 23477 20913 23480
rect 20947 23477 20959 23511
rect 20901 23471 20959 23477
rect 21174 23468 21180 23520
rect 21232 23508 21238 23520
rect 22002 23508 22008 23520
rect 21232 23480 22008 23508
rect 21232 23468 21238 23480
rect 22002 23468 22008 23480
rect 22060 23508 22066 23520
rect 22281 23511 22339 23517
rect 22281 23508 22293 23511
rect 22060 23480 22293 23508
rect 22060 23468 22066 23480
rect 22281 23477 22293 23480
rect 22327 23477 22339 23511
rect 22281 23471 22339 23477
rect 23290 23468 23296 23520
rect 23348 23508 23354 23520
rect 23385 23511 23443 23517
rect 23385 23508 23397 23511
rect 23348 23480 23397 23508
rect 23348 23468 23354 23480
rect 23385 23477 23397 23480
rect 23431 23477 23443 23511
rect 23385 23471 23443 23477
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 1670 23264 1676 23316
rect 1728 23304 1734 23316
rect 1857 23307 1915 23313
rect 1857 23304 1869 23307
rect 1728 23276 1869 23304
rect 1728 23264 1734 23276
rect 1857 23273 1869 23276
rect 1903 23304 1915 23307
rect 2409 23307 2467 23313
rect 2409 23304 2421 23307
rect 1903 23276 2421 23304
rect 1903 23273 1915 23276
rect 1857 23267 1915 23273
rect 2409 23273 2421 23276
rect 2455 23273 2467 23307
rect 7006 23304 7012 23316
rect 6967 23276 7012 23304
rect 2409 23267 2467 23273
rect 7006 23264 7012 23276
rect 7064 23264 7070 23316
rect 7558 23264 7564 23316
rect 7616 23304 7622 23316
rect 8481 23307 8539 23313
rect 8481 23304 8493 23307
rect 7616 23276 8493 23304
rect 7616 23264 7622 23276
rect 8481 23273 8493 23276
rect 8527 23273 8539 23307
rect 8481 23267 8539 23273
rect 9493 23307 9551 23313
rect 9493 23273 9505 23307
rect 9539 23304 9551 23307
rect 10045 23307 10103 23313
rect 10045 23304 10057 23307
rect 9539 23276 10057 23304
rect 9539 23273 9551 23276
rect 9493 23267 9551 23273
rect 10045 23273 10057 23276
rect 10091 23304 10103 23307
rect 10134 23304 10140 23316
rect 10091 23276 10140 23304
rect 10091 23273 10103 23276
rect 10045 23267 10103 23273
rect 10134 23264 10140 23276
rect 10192 23304 10198 23316
rect 11609 23307 11667 23313
rect 11609 23304 11621 23307
rect 10192 23276 11621 23304
rect 10192 23264 10198 23276
rect 11609 23273 11621 23276
rect 11655 23273 11667 23307
rect 12342 23304 12348 23316
rect 12255 23276 12348 23304
rect 11609 23267 11667 23273
rect 1397 23171 1455 23177
rect 1397 23137 1409 23171
rect 1443 23168 1455 23171
rect 2406 23168 2412 23180
rect 1443 23140 2412 23168
rect 1443 23137 1455 23140
rect 1397 23131 1455 23137
rect 2406 23128 2412 23140
rect 2464 23168 2470 23180
rect 4338 23177 4344 23180
rect 2777 23171 2835 23177
rect 2777 23168 2789 23171
rect 2464 23140 2789 23168
rect 2464 23128 2470 23140
rect 2777 23137 2789 23140
rect 2823 23137 2835 23171
rect 4321 23171 4344 23177
rect 4321 23168 4333 23171
rect 2777 23131 2835 23137
rect 2976 23140 4333 23168
rect 2317 23103 2375 23109
rect 2317 23069 2329 23103
rect 2363 23100 2375 23103
rect 2866 23100 2872 23112
rect 2363 23072 2872 23100
rect 2363 23069 2375 23072
rect 2317 23063 2375 23069
rect 2866 23060 2872 23072
rect 2924 23060 2930 23112
rect 2976 23109 3004 23140
rect 4321 23137 4333 23140
rect 4396 23168 4402 23180
rect 6089 23171 6147 23177
rect 4396 23140 4469 23168
rect 4321 23131 4344 23137
rect 4338 23128 4344 23131
rect 4396 23128 4402 23140
rect 6089 23137 6101 23171
rect 6135 23168 6147 23171
rect 6546 23168 6552 23180
rect 6135 23140 6552 23168
rect 6135 23137 6147 23140
rect 6089 23131 6147 23137
rect 6546 23128 6552 23140
rect 6604 23168 6610 23180
rect 7024 23168 7052 23264
rect 10502 23245 10508 23248
rect 10496 23236 10508 23245
rect 10463 23208 10508 23236
rect 10496 23199 10508 23208
rect 10560 23236 10566 23248
rect 12268 23245 12296 23276
rect 12342 23264 12348 23276
rect 12400 23304 12406 23316
rect 14093 23307 14151 23313
rect 14093 23304 14105 23307
rect 12400 23276 14105 23304
rect 12400 23264 12406 23276
rect 14093 23273 14105 23276
rect 14139 23273 14151 23307
rect 14093 23267 14151 23273
rect 14734 23264 14740 23316
rect 14792 23304 14798 23316
rect 15749 23307 15807 23313
rect 15749 23304 15761 23307
rect 14792 23276 15761 23304
rect 14792 23264 14798 23276
rect 15749 23273 15761 23276
rect 15795 23273 15807 23307
rect 15749 23267 15807 23273
rect 19613 23307 19671 23313
rect 19613 23273 19625 23307
rect 19659 23304 19671 23307
rect 20622 23304 20628 23316
rect 19659 23276 20628 23304
rect 19659 23273 19671 23276
rect 19613 23267 19671 23273
rect 20622 23264 20628 23276
rect 20680 23264 20686 23316
rect 12253 23239 12311 23245
rect 12253 23236 12265 23239
rect 10560 23208 12265 23236
rect 10502 23196 10508 23199
rect 10560 23196 10566 23208
rect 12253 23205 12265 23208
rect 12299 23205 12311 23239
rect 12253 23199 12311 23205
rect 12621 23239 12679 23245
rect 12621 23205 12633 23239
rect 12667 23236 12679 23239
rect 13538 23236 13544 23248
rect 12667 23208 13544 23236
rect 12667 23205 12679 23208
rect 12621 23199 12679 23205
rect 13538 23196 13544 23208
rect 13596 23196 13602 23248
rect 17126 23236 17132 23248
rect 17087 23208 17132 23236
rect 17126 23196 17132 23208
rect 17184 23196 17190 23248
rect 21174 23236 21180 23248
rect 21135 23208 21180 23236
rect 21174 23196 21180 23208
rect 21232 23196 21238 23248
rect 22741 23239 22799 23245
rect 22741 23205 22753 23239
rect 22787 23236 22799 23239
rect 23382 23236 23388 23248
rect 22787 23208 23388 23236
rect 22787 23205 22799 23208
rect 22741 23199 22799 23205
rect 23382 23196 23388 23208
rect 23440 23196 23446 23248
rect 7101 23171 7159 23177
rect 7101 23168 7113 23171
rect 6604 23140 7113 23168
rect 6604 23128 6610 23140
rect 7101 23137 7113 23140
rect 7147 23137 7159 23171
rect 7101 23131 7159 23137
rect 7368 23171 7426 23177
rect 7368 23137 7380 23171
rect 7414 23168 7426 23171
rect 7650 23168 7656 23180
rect 7414 23140 7656 23168
rect 7414 23137 7426 23140
rect 7368 23131 7426 23137
rect 7650 23128 7656 23140
rect 7708 23128 7714 23180
rect 12986 23177 12992 23180
rect 12980 23168 12992 23177
rect 12947 23140 12992 23168
rect 12980 23131 12992 23140
rect 12986 23128 12992 23131
rect 13044 23128 13050 23180
rect 15562 23128 15568 23180
rect 15620 23168 15626 23180
rect 15657 23171 15715 23177
rect 15657 23168 15669 23171
rect 15620 23140 15669 23168
rect 15620 23128 15626 23140
rect 15657 23137 15669 23140
rect 15703 23168 15715 23171
rect 16114 23168 16120 23180
rect 15703 23140 16120 23168
rect 15703 23137 15715 23140
rect 15657 23131 15715 23137
rect 16114 23128 16120 23140
rect 16172 23128 16178 23180
rect 16758 23128 16764 23180
rect 16816 23168 16822 23180
rect 16853 23171 16911 23177
rect 16853 23168 16865 23171
rect 16816 23140 16865 23168
rect 16816 23128 16822 23140
rect 16853 23137 16865 23140
rect 16899 23137 16911 23171
rect 16853 23131 16911 23137
rect 18141 23171 18199 23177
rect 18141 23137 18153 23171
rect 18187 23168 18199 23171
rect 18230 23168 18236 23180
rect 18187 23140 18236 23168
rect 18187 23137 18199 23140
rect 18141 23131 18199 23137
rect 18230 23128 18236 23140
rect 18288 23128 18294 23180
rect 18417 23171 18475 23177
rect 18417 23137 18429 23171
rect 18463 23168 18475 23171
rect 19426 23168 19432 23180
rect 18463 23140 19432 23168
rect 18463 23137 18475 23140
rect 18417 23131 18475 23137
rect 19426 23128 19432 23140
rect 19484 23128 19490 23180
rect 20898 23168 20904 23180
rect 20859 23140 20904 23168
rect 20898 23128 20904 23140
rect 20956 23128 20962 23180
rect 22462 23168 22468 23180
rect 22423 23140 22468 23168
rect 22462 23128 22468 23140
rect 22520 23128 22526 23180
rect 2961 23103 3019 23109
rect 2961 23069 2973 23103
rect 3007 23069 3019 23103
rect 2961 23063 3019 23069
rect 2774 22992 2780 23044
rect 2832 23032 2838 23044
rect 2976 23032 3004 23063
rect 3326 23060 3332 23112
rect 3384 23100 3390 23112
rect 3878 23100 3884 23112
rect 3384 23072 3884 23100
rect 3384 23060 3390 23072
rect 3878 23060 3884 23072
rect 3936 23100 3942 23112
rect 4065 23103 4123 23109
rect 4065 23100 4077 23103
rect 3936 23072 4077 23100
rect 3936 23060 3942 23072
rect 4065 23069 4077 23072
rect 4111 23069 4123 23103
rect 4065 23063 4123 23069
rect 9030 23060 9036 23112
rect 9088 23100 9094 23112
rect 9125 23103 9183 23109
rect 9125 23100 9137 23103
rect 9088 23072 9137 23100
rect 9088 23060 9094 23072
rect 9125 23069 9137 23072
rect 9171 23100 9183 23103
rect 9950 23100 9956 23112
rect 9171 23072 9956 23100
rect 9171 23069 9183 23072
rect 9125 23063 9183 23069
rect 9950 23060 9956 23072
rect 10008 23100 10014 23112
rect 10226 23100 10232 23112
rect 10008 23072 10232 23100
rect 10008 23060 10014 23072
rect 10226 23060 10232 23072
rect 10284 23060 10290 23112
rect 12526 23060 12532 23112
rect 12584 23100 12590 23112
rect 12713 23103 12771 23109
rect 12713 23100 12725 23103
rect 12584 23072 12725 23100
rect 12584 23060 12590 23072
rect 12713 23069 12725 23072
rect 12759 23069 12771 23103
rect 15930 23100 15936 23112
rect 15891 23072 15936 23100
rect 12713 23063 12771 23069
rect 15930 23060 15936 23072
rect 15988 23060 15994 23112
rect 2832 23004 3004 23032
rect 2832 22992 2838 23004
rect 3510 22964 3516 22976
rect 3471 22936 3516 22964
rect 3510 22924 3516 22936
rect 3568 22924 3574 22976
rect 5442 22964 5448 22976
rect 5403 22936 5448 22964
rect 5442 22924 5448 22936
rect 5500 22924 5506 22976
rect 15286 22964 15292 22976
rect 15247 22936 15292 22964
rect 15286 22924 15292 22936
rect 15344 22924 15350 22976
rect 15470 22924 15476 22976
rect 15528 22964 15534 22976
rect 16301 22967 16359 22973
rect 16301 22964 16313 22967
rect 15528 22936 16313 22964
rect 15528 22924 15534 22936
rect 16301 22933 16313 22936
rect 16347 22933 16359 22967
rect 16301 22927 16359 22933
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 2406 22760 2412 22772
rect 2367 22732 2412 22760
rect 2406 22720 2412 22732
rect 2464 22720 2470 22772
rect 2682 22720 2688 22772
rect 2740 22760 2746 22772
rect 2961 22763 3019 22769
rect 2961 22760 2973 22763
rect 2740 22732 2973 22760
rect 2740 22720 2746 22732
rect 2961 22729 2973 22732
rect 3007 22729 3019 22763
rect 2961 22723 3019 22729
rect 5629 22763 5687 22769
rect 5629 22729 5641 22763
rect 5675 22760 5687 22763
rect 6638 22760 6644 22772
rect 5675 22732 6644 22760
rect 5675 22729 5687 22732
rect 5629 22723 5687 22729
rect 2777 22695 2835 22701
rect 2777 22661 2789 22695
rect 2823 22661 2835 22695
rect 2777 22655 2835 22661
rect 1949 22627 2007 22633
rect 1949 22593 1961 22627
rect 1995 22624 2007 22627
rect 2038 22624 2044 22636
rect 1995 22596 2044 22624
rect 1995 22593 2007 22596
rect 1949 22587 2007 22593
rect 2038 22584 2044 22596
rect 2096 22584 2102 22636
rect 2792 22624 2820 22655
rect 2866 22652 2872 22704
rect 2924 22692 2930 22704
rect 4525 22695 4583 22701
rect 4525 22692 4537 22695
rect 2924 22664 4537 22692
rect 2924 22652 2930 22664
rect 4525 22661 4537 22664
rect 4571 22661 4583 22695
rect 4525 22655 4583 22661
rect 3602 22624 3608 22636
rect 2792 22596 3608 22624
rect 3602 22584 3608 22596
rect 3660 22584 3666 22636
rect 4154 22584 4160 22636
rect 4212 22624 4218 22636
rect 5169 22627 5227 22633
rect 5169 22624 5181 22627
rect 4212 22596 5181 22624
rect 4212 22584 4218 22596
rect 5169 22593 5181 22596
rect 5215 22624 5227 22627
rect 5644 22624 5672 22723
rect 6638 22720 6644 22732
rect 6696 22720 6702 22772
rect 6822 22720 6828 22772
rect 6880 22760 6886 22772
rect 7009 22763 7067 22769
rect 7009 22760 7021 22763
rect 6880 22732 7021 22760
rect 6880 22720 6886 22732
rect 7009 22729 7021 22732
rect 7055 22729 7067 22763
rect 7009 22723 7067 22729
rect 8481 22763 8539 22769
rect 8481 22729 8493 22763
rect 8527 22760 8539 22763
rect 8570 22760 8576 22772
rect 8527 22732 8576 22760
rect 8527 22729 8539 22732
rect 8481 22723 8539 22729
rect 8570 22720 8576 22732
rect 8628 22720 8634 22772
rect 10502 22760 10508 22772
rect 10463 22732 10508 22760
rect 10502 22720 10508 22732
rect 10560 22720 10566 22772
rect 12805 22763 12863 22769
rect 12805 22729 12817 22763
rect 12851 22760 12863 22763
rect 12986 22760 12992 22772
rect 12851 22732 12992 22760
rect 12851 22729 12863 22732
rect 12805 22723 12863 22729
rect 12986 22720 12992 22732
rect 13044 22720 13050 22772
rect 13265 22763 13323 22769
rect 13265 22729 13277 22763
rect 13311 22760 13323 22763
rect 13538 22760 13544 22772
rect 13311 22732 13544 22760
rect 13311 22729 13323 22732
rect 13265 22723 13323 22729
rect 13538 22720 13544 22732
rect 13596 22720 13602 22772
rect 14458 22720 14464 22772
rect 14516 22760 14522 22772
rect 14734 22760 14740 22772
rect 14516 22732 14740 22760
rect 14516 22720 14522 22732
rect 14734 22720 14740 22732
rect 14792 22760 14798 22772
rect 14921 22763 14979 22769
rect 14921 22760 14933 22763
rect 14792 22732 14933 22760
rect 14792 22720 14798 22732
rect 14921 22729 14933 22732
rect 14967 22729 14979 22763
rect 19426 22760 19432 22772
rect 19387 22732 19432 22760
rect 14921 22723 14979 22729
rect 19426 22720 19432 22732
rect 19484 22720 19490 22772
rect 20898 22760 20904 22772
rect 20859 22732 20904 22760
rect 20898 22720 20904 22732
rect 20956 22720 20962 22772
rect 16850 22692 16856 22704
rect 16811 22664 16856 22692
rect 16850 22652 16856 22664
rect 16908 22652 16914 22704
rect 7558 22624 7564 22636
rect 5215 22596 5672 22624
rect 7519 22596 7564 22624
rect 5215 22593 5227 22596
rect 5169 22587 5227 22593
rect 7558 22584 7564 22596
rect 7616 22624 7622 22636
rect 8021 22627 8079 22633
rect 8021 22624 8033 22627
rect 7616 22596 8033 22624
rect 7616 22584 7622 22596
rect 8021 22593 8033 22596
rect 8067 22593 8079 22627
rect 8021 22587 8079 22593
rect 13173 22627 13231 22633
rect 13173 22593 13185 22627
rect 13219 22624 13231 22627
rect 13722 22624 13728 22636
rect 13219 22596 13728 22624
rect 13219 22593 13231 22596
rect 13173 22587 13231 22593
rect 13722 22584 13728 22596
rect 13780 22584 13786 22636
rect 13906 22624 13912 22636
rect 13867 22596 13912 22624
rect 13906 22584 13912 22596
rect 13964 22584 13970 22636
rect 15470 22624 15476 22636
rect 15431 22596 15476 22624
rect 15470 22584 15476 22596
rect 15528 22584 15534 22636
rect 1673 22559 1731 22565
rect 1673 22525 1685 22559
rect 1719 22556 1731 22559
rect 2682 22556 2688 22568
rect 1719 22528 2688 22556
rect 1719 22525 1731 22528
rect 1673 22519 1731 22525
rect 2682 22516 2688 22528
rect 2740 22516 2746 22568
rect 2774 22516 2780 22568
rect 2832 22556 2838 22568
rect 3973 22559 4031 22565
rect 3973 22556 3985 22559
rect 2832 22528 3985 22556
rect 2832 22516 2838 22528
rect 3973 22525 3985 22528
rect 4019 22525 4031 22559
rect 4982 22556 4988 22568
rect 4943 22528 4988 22556
rect 3973 22519 4031 22525
rect 4982 22516 4988 22528
rect 5040 22516 5046 22568
rect 6273 22559 6331 22565
rect 6273 22525 6285 22559
rect 6319 22556 6331 22559
rect 7650 22556 7656 22568
rect 6319 22528 7656 22556
rect 6319 22525 6331 22528
rect 6273 22519 6331 22525
rect 7650 22516 7656 22528
rect 7708 22516 7714 22568
rect 8573 22559 8631 22565
rect 8573 22525 8585 22559
rect 8619 22525 8631 22559
rect 8573 22519 8631 22525
rect 2866 22448 2872 22500
rect 2924 22488 2930 22500
rect 3050 22488 3056 22500
rect 2924 22460 3056 22488
rect 2924 22448 2930 22460
rect 3050 22448 3056 22460
rect 3108 22448 3114 22500
rect 4433 22491 4491 22497
rect 4433 22457 4445 22491
rect 4479 22488 4491 22491
rect 5000 22488 5028 22516
rect 4479 22460 5028 22488
rect 6641 22491 6699 22497
rect 4479 22457 4491 22460
rect 4433 22451 4491 22457
rect 6641 22457 6653 22491
rect 6687 22488 6699 22491
rect 8588 22488 8616 22519
rect 8662 22516 8668 22568
rect 8720 22556 8726 22568
rect 8829 22559 8887 22565
rect 8829 22556 8841 22559
rect 8720 22528 8841 22556
rect 8720 22516 8726 22528
rect 8829 22525 8841 22528
rect 8875 22525 8887 22559
rect 8829 22519 8887 22525
rect 13262 22516 13268 22568
rect 13320 22556 13326 22568
rect 13633 22559 13691 22565
rect 13633 22556 13645 22559
rect 13320 22528 13645 22556
rect 13320 22516 13326 22528
rect 13633 22525 13645 22528
rect 13679 22525 13691 22559
rect 22462 22556 22468 22568
rect 22423 22528 22468 22556
rect 13633 22519 13691 22525
rect 22462 22516 22468 22528
rect 22520 22516 22526 22568
rect 9030 22488 9036 22500
rect 6687 22460 7512 22488
rect 8588 22460 9036 22488
rect 6687 22457 6699 22460
rect 6641 22451 6699 22457
rect 3326 22420 3332 22432
rect 3287 22392 3332 22420
rect 3326 22380 3332 22392
rect 3384 22380 3390 22432
rect 3421 22423 3479 22429
rect 3421 22389 3433 22423
rect 3467 22420 3479 22423
rect 3510 22420 3516 22432
rect 3467 22392 3516 22420
rect 3467 22389 3479 22392
rect 3421 22383 3479 22389
rect 3510 22380 3516 22392
rect 3568 22420 3574 22432
rect 4062 22420 4068 22432
rect 3568 22392 4068 22420
rect 3568 22380 3574 22392
rect 4062 22380 4068 22392
rect 4120 22380 4126 22432
rect 4522 22380 4528 22432
rect 4580 22420 4586 22432
rect 4893 22423 4951 22429
rect 4893 22420 4905 22423
rect 4580 22392 4905 22420
rect 4580 22380 4586 22392
rect 4893 22389 4905 22392
rect 4939 22389 4951 22423
rect 4893 22383 4951 22389
rect 7098 22380 7104 22432
rect 7156 22420 7162 22432
rect 7484 22429 7512 22460
rect 9030 22448 9036 22460
rect 9088 22448 9094 22500
rect 10226 22448 10232 22500
rect 10284 22488 10290 22500
rect 15746 22497 15752 22500
rect 10965 22491 11023 22497
rect 10965 22488 10977 22491
rect 10284 22460 10977 22488
rect 10284 22448 10290 22460
rect 10965 22457 10977 22460
rect 11011 22488 11023 22491
rect 14645 22491 14703 22497
rect 11011 22460 12296 22488
rect 11011 22457 11023 22460
rect 10965 22451 11023 22457
rect 7377 22423 7435 22429
rect 7377 22420 7389 22423
rect 7156 22392 7389 22420
rect 7156 22380 7162 22392
rect 7377 22389 7389 22392
rect 7423 22389 7435 22423
rect 7377 22383 7435 22389
rect 7469 22423 7527 22429
rect 7469 22389 7481 22423
rect 7515 22420 7527 22423
rect 8754 22420 8760 22432
rect 7515 22392 8760 22420
rect 7515 22389 7527 22392
rect 7469 22383 7527 22389
rect 8754 22380 8760 22392
rect 8812 22380 8818 22432
rect 9582 22380 9588 22432
rect 9640 22420 9646 22432
rect 9953 22423 10011 22429
rect 9953 22420 9965 22423
rect 9640 22392 9965 22420
rect 9640 22380 9646 22392
rect 9953 22389 9965 22392
rect 9999 22389 10011 22423
rect 11054 22420 11060 22432
rect 11015 22392 11060 22420
rect 9953 22383 10011 22389
rect 11054 22380 11060 22392
rect 11112 22380 11118 22432
rect 12268 22429 12296 22460
rect 14645 22457 14657 22491
rect 14691 22488 14703 22491
rect 15718 22491 15752 22497
rect 15718 22488 15730 22491
rect 14691 22460 15730 22488
rect 14691 22457 14703 22460
rect 14645 22451 14703 22457
rect 15718 22457 15730 22460
rect 15804 22488 15810 22500
rect 15804 22460 15866 22488
rect 15718 22451 15752 22457
rect 15746 22448 15752 22451
rect 15804 22448 15810 22460
rect 16114 22448 16120 22500
rect 16172 22488 16178 22500
rect 16758 22488 16764 22500
rect 16172 22460 16764 22488
rect 16172 22448 16178 22460
rect 16758 22448 16764 22460
rect 16816 22488 16822 22500
rect 17405 22491 17463 22497
rect 17405 22488 17417 22491
rect 16816 22460 17417 22488
rect 16816 22448 16822 22460
rect 17405 22457 17417 22460
rect 17451 22457 17463 22491
rect 17405 22451 17463 22457
rect 12253 22423 12311 22429
rect 12253 22389 12265 22423
rect 12299 22420 12311 22423
rect 12526 22420 12532 22432
rect 12299 22392 12532 22420
rect 12299 22389 12311 22392
rect 12253 22383 12311 22389
rect 12526 22380 12532 22392
rect 12584 22380 12590 22432
rect 14182 22380 14188 22432
rect 14240 22420 14246 22432
rect 15289 22423 15347 22429
rect 15289 22420 15301 22423
rect 14240 22392 15301 22420
rect 14240 22380 14246 22392
rect 15289 22389 15301 22392
rect 15335 22420 15347 22423
rect 15562 22420 15568 22432
rect 15335 22392 15568 22420
rect 15335 22389 15347 22392
rect 15289 22383 15347 22389
rect 15562 22380 15568 22392
rect 15620 22380 15626 22432
rect 18230 22420 18236 22432
rect 18191 22392 18236 22420
rect 18230 22380 18236 22392
rect 18288 22380 18294 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 10962 22176 10968 22228
rect 11020 22216 11026 22228
rect 11333 22219 11391 22225
rect 11333 22216 11345 22219
rect 11020 22188 11345 22216
rect 11020 22176 11026 22188
rect 11333 22185 11345 22188
rect 11379 22185 11391 22219
rect 11333 22179 11391 22185
rect 12621 22219 12679 22225
rect 12621 22185 12633 22219
rect 12667 22216 12679 22219
rect 13354 22216 13360 22228
rect 12667 22188 13360 22216
rect 12667 22185 12679 22188
rect 12621 22179 12679 22185
rect 13354 22176 13360 22188
rect 13412 22176 13418 22228
rect 13722 22216 13728 22228
rect 13683 22188 13728 22216
rect 13722 22176 13728 22188
rect 13780 22176 13786 22228
rect 15289 22219 15347 22225
rect 15289 22185 15301 22219
rect 15335 22216 15347 22219
rect 15470 22216 15476 22228
rect 15335 22188 15476 22216
rect 15335 22185 15347 22188
rect 15289 22179 15347 22185
rect 15470 22176 15476 22188
rect 15528 22176 15534 22228
rect 3326 22108 3332 22160
rect 3384 22148 3390 22160
rect 3421 22151 3479 22157
rect 3421 22148 3433 22151
rect 3384 22120 3433 22148
rect 3384 22108 3390 22120
rect 3421 22117 3433 22120
rect 3467 22117 3479 22151
rect 3421 22111 3479 22117
rect 5160 22151 5218 22157
rect 5160 22117 5172 22151
rect 5206 22148 5218 22151
rect 5442 22148 5448 22160
rect 5206 22120 5448 22148
rect 5206 22117 5218 22120
rect 5160 22111 5218 22117
rect 5442 22108 5448 22120
rect 5500 22108 5506 22160
rect 7374 22108 7380 22160
rect 7432 22148 7438 22160
rect 8018 22148 8024 22160
rect 7432 22120 8024 22148
rect 7432 22108 7438 22120
rect 8018 22108 8024 22120
rect 8076 22108 8082 22160
rect 1578 22080 1584 22092
rect 1539 22052 1584 22080
rect 1578 22040 1584 22052
rect 1636 22040 1642 22092
rect 1857 22083 1915 22089
rect 1857 22049 1869 22083
rect 1903 22080 1915 22083
rect 2406 22080 2412 22092
rect 1903 22052 2412 22080
rect 1903 22049 1915 22052
rect 1857 22043 1915 22049
rect 2406 22040 2412 22052
rect 2464 22040 2470 22092
rect 2501 22083 2559 22089
rect 2501 22049 2513 22083
rect 2547 22080 2559 22083
rect 2682 22080 2688 22092
rect 2547 22052 2688 22080
rect 2547 22049 2559 22052
rect 2501 22043 2559 22049
rect 2682 22040 2688 22052
rect 2740 22040 2746 22092
rect 2774 22040 2780 22092
rect 2832 22080 2838 22092
rect 2869 22083 2927 22089
rect 2869 22080 2881 22083
rect 2832 22052 2881 22080
rect 2832 22040 2838 22052
rect 2869 22049 2881 22052
rect 2915 22049 2927 22083
rect 2869 22043 2927 22049
rect 7650 22040 7656 22092
rect 7708 22080 7714 22092
rect 8386 22080 8392 22092
rect 7708 22052 8392 22080
rect 7708 22040 7714 22052
rect 4893 22015 4951 22021
rect 4893 22012 4905 22015
rect 3896 21984 4905 22012
rect 3896 21888 3924 21984
rect 4893 21981 4905 21984
rect 4939 21981 4951 22015
rect 4893 21975 4951 21981
rect 6638 21972 6644 22024
rect 6696 22012 6702 22024
rect 8110 22012 8116 22024
rect 6696 21984 8116 22012
rect 6696 21972 6702 21984
rect 8110 21972 8116 21984
rect 8168 21972 8174 22024
rect 8312 22021 8340 22052
rect 8386 22040 8392 22052
rect 8444 22080 8450 22092
rect 9582 22080 9588 22092
rect 8444 22052 9588 22080
rect 8444 22040 8450 22052
rect 9582 22040 9588 22052
rect 9640 22040 9646 22092
rect 10042 22040 10048 22092
rect 10100 22080 10106 22092
rect 10137 22083 10195 22089
rect 10137 22080 10149 22083
rect 10100 22052 10149 22080
rect 10100 22040 10106 22052
rect 10137 22049 10149 22052
rect 10183 22049 10195 22083
rect 10137 22043 10195 22049
rect 13446 22040 13452 22092
rect 13504 22080 13510 22092
rect 13817 22083 13875 22089
rect 13817 22080 13829 22083
rect 13504 22052 13829 22080
rect 13504 22040 13510 22052
rect 13817 22049 13829 22052
rect 13863 22049 13875 22083
rect 13817 22043 13875 22049
rect 14093 22083 14151 22089
rect 14093 22049 14105 22083
rect 14139 22080 14151 22083
rect 14826 22080 14832 22092
rect 14139 22052 14832 22080
rect 14139 22049 14151 22052
rect 14093 22043 14151 22049
rect 14826 22040 14832 22052
rect 14884 22040 14890 22092
rect 15289 22083 15347 22089
rect 15289 22049 15301 22083
rect 15335 22080 15347 22083
rect 15381 22083 15439 22089
rect 15381 22080 15393 22083
rect 15335 22052 15393 22080
rect 15335 22049 15347 22052
rect 15289 22043 15347 22049
rect 15381 22049 15393 22052
rect 15427 22049 15439 22083
rect 15648 22083 15706 22089
rect 15648 22080 15660 22083
rect 15381 22043 15439 22049
rect 15488 22052 15660 22080
rect 8297 22015 8355 22021
rect 8297 21981 8309 22015
rect 8343 22012 8355 22015
rect 8343 21984 8377 22012
rect 8343 21981 8355 21984
rect 8297 21975 8355 21981
rect 9122 21972 9128 22024
rect 9180 22012 9186 22024
rect 10226 22012 10232 22024
rect 9180 21984 10232 22012
rect 9180 21972 9186 21984
rect 10226 21972 10232 21984
rect 10284 21972 10290 22024
rect 10410 22012 10416 22024
rect 10371 21984 10416 22012
rect 10410 21972 10416 21984
rect 10468 21972 10474 22024
rect 15105 22015 15163 22021
rect 15105 21981 15117 22015
rect 15151 22012 15163 22015
rect 15488 22012 15516 22052
rect 15648 22049 15660 22052
rect 15694 22080 15706 22083
rect 15930 22080 15936 22092
rect 15694 22052 15936 22080
rect 15694 22049 15706 22052
rect 15648 22043 15706 22049
rect 15930 22040 15936 22052
rect 15988 22040 15994 22092
rect 15151 21984 15516 22012
rect 15151 21981 15163 21984
rect 15105 21975 15163 21981
rect 6270 21944 6276 21956
rect 6231 21916 6276 21944
rect 6270 21904 6276 21916
rect 6328 21904 6334 21956
rect 7561 21947 7619 21953
rect 7561 21913 7573 21947
rect 7607 21944 7619 21947
rect 8018 21944 8024 21956
rect 7607 21916 8024 21944
rect 7607 21913 7619 21916
rect 7561 21907 7619 21913
rect 8018 21904 8024 21916
rect 8076 21904 8082 21956
rect 9769 21947 9827 21953
rect 9769 21913 9781 21947
rect 9815 21944 9827 21947
rect 10962 21944 10968 21956
rect 9815 21916 10968 21944
rect 9815 21913 9827 21916
rect 9769 21907 9827 21913
rect 10962 21904 10968 21916
rect 11020 21904 11026 21956
rect 3050 21876 3056 21888
rect 3011 21848 3056 21876
rect 3050 21836 3056 21848
rect 3108 21836 3114 21888
rect 3878 21876 3884 21888
rect 3839 21848 3884 21876
rect 3878 21836 3884 21848
rect 3936 21836 3942 21888
rect 4522 21876 4528 21888
rect 4483 21848 4528 21876
rect 4522 21836 4528 21848
rect 4580 21836 4586 21888
rect 7098 21876 7104 21888
rect 7059 21848 7104 21876
rect 7098 21836 7104 21848
rect 7156 21836 7162 21888
rect 7650 21876 7656 21888
rect 7611 21848 7656 21876
rect 7650 21836 7656 21848
rect 7708 21836 7714 21888
rect 8757 21879 8815 21885
rect 8757 21845 8769 21879
rect 8803 21876 8815 21879
rect 9030 21876 9036 21888
rect 8803 21848 9036 21876
rect 8803 21845 8815 21848
rect 8757 21839 8815 21845
rect 9030 21836 9036 21848
rect 9088 21836 9094 21888
rect 10686 21836 10692 21888
rect 10744 21876 10750 21888
rect 10781 21879 10839 21885
rect 10781 21876 10793 21879
rect 10744 21848 10793 21876
rect 10744 21836 10750 21848
rect 10781 21845 10793 21848
rect 10827 21845 10839 21879
rect 10781 21839 10839 21845
rect 12529 21879 12587 21885
rect 12529 21845 12541 21879
rect 12575 21876 12587 21879
rect 12802 21876 12808 21888
rect 12575 21848 12808 21876
rect 12575 21845 12587 21848
rect 12529 21839 12587 21845
rect 12802 21836 12808 21848
rect 12860 21836 12866 21888
rect 13262 21876 13268 21888
rect 13223 21848 13268 21876
rect 13262 21836 13268 21848
rect 13320 21836 13326 21888
rect 15746 21836 15752 21888
rect 15804 21876 15810 21888
rect 16761 21879 16819 21885
rect 16761 21876 16773 21879
rect 15804 21848 16773 21876
rect 15804 21836 15810 21848
rect 16761 21845 16773 21848
rect 16807 21845 16819 21879
rect 16761 21839 16819 21845
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 2774 21632 2780 21684
rect 2832 21672 2838 21684
rect 2869 21675 2927 21681
rect 2869 21672 2881 21675
rect 2832 21644 2881 21672
rect 2832 21632 2838 21644
rect 2869 21641 2881 21644
rect 2915 21641 2927 21675
rect 4154 21672 4160 21684
rect 4115 21644 4160 21672
rect 2869 21635 2927 21641
rect 4154 21632 4160 21644
rect 4212 21632 4218 21684
rect 5261 21675 5319 21681
rect 5261 21641 5273 21675
rect 5307 21672 5319 21675
rect 5442 21672 5448 21684
rect 5307 21644 5448 21672
rect 5307 21641 5319 21644
rect 5261 21635 5319 21641
rect 2133 21539 2191 21545
rect 2133 21505 2145 21539
rect 2179 21536 2191 21539
rect 2222 21536 2228 21548
rect 2179 21508 2228 21536
rect 2179 21505 2191 21508
rect 2133 21499 2191 21505
rect 2222 21496 2228 21508
rect 2280 21496 2286 21548
rect 3145 21539 3203 21545
rect 3145 21505 3157 21539
rect 3191 21536 3203 21539
rect 3326 21536 3332 21548
rect 3191 21508 3332 21536
rect 3191 21505 3203 21508
rect 3145 21499 3203 21505
rect 3326 21496 3332 21508
rect 3384 21496 3390 21548
rect 4338 21496 4344 21548
rect 4396 21536 4402 21548
rect 4801 21539 4859 21545
rect 4801 21536 4813 21539
rect 4396 21508 4813 21536
rect 4396 21496 4402 21508
rect 4801 21505 4813 21508
rect 4847 21536 4859 21539
rect 5276 21536 5304 21635
rect 5442 21632 5448 21644
rect 5500 21632 5506 21684
rect 6638 21672 6644 21684
rect 6599 21644 6644 21672
rect 6638 21632 6644 21644
rect 6696 21632 6702 21684
rect 7374 21672 7380 21684
rect 7335 21644 7380 21672
rect 7374 21632 7380 21644
rect 7432 21632 7438 21684
rect 10134 21632 10140 21684
rect 10192 21672 10198 21684
rect 10410 21672 10416 21684
rect 10192 21644 10416 21672
rect 10192 21632 10198 21644
rect 10410 21632 10416 21644
rect 10468 21672 10474 21684
rect 11333 21675 11391 21681
rect 11333 21672 11345 21675
rect 10468 21644 11345 21672
rect 10468 21632 10474 21644
rect 11333 21641 11345 21644
rect 11379 21641 11391 21675
rect 11333 21635 11391 21641
rect 12158 21604 12164 21616
rect 12119 21576 12164 21604
rect 12158 21564 12164 21576
rect 12216 21564 12222 21616
rect 4847 21508 5304 21536
rect 4847 21505 4859 21508
rect 4801 21499 4859 21505
rect 5534 21496 5540 21548
rect 5592 21536 5598 21548
rect 5721 21539 5779 21545
rect 5721 21536 5733 21539
rect 5592 21508 5733 21536
rect 5592 21496 5598 21508
rect 5721 21505 5733 21508
rect 5767 21505 5779 21539
rect 5721 21499 5779 21505
rect 10597 21539 10655 21545
rect 10597 21505 10609 21539
rect 10643 21536 10655 21539
rect 10686 21536 10692 21548
rect 10643 21508 10692 21536
rect 10643 21505 10655 21508
rect 10597 21499 10655 21505
rect 10686 21496 10692 21508
rect 10744 21496 10750 21548
rect 11882 21496 11888 21548
rect 11940 21536 11946 21548
rect 12989 21539 13047 21545
rect 12989 21536 13001 21539
rect 11940 21508 13001 21536
rect 11940 21496 11946 21508
rect 12989 21505 13001 21508
rect 13035 21505 13047 21539
rect 12989 21499 13047 21505
rect 13630 21496 13636 21548
rect 13688 21536 13694 21548
rect 13906 21536 13912 21548
rect 13688 21508 13912 21536
rect 13688 21496 13694 21508
rect 13906 21496 13912 21508
rect 13964 21536 13970 21548
rect 14001 21539 14059 21545
rect 14001 21536 14013 21539
rect 13964 21508 14013 21536
rect 13964 21496 13970 21508
rect 14001 21505 14013 21508
rect 14047 21505 14059 21539
rect 14001 21499 14059 21505
rect 1857 21471 1915 21477
rect 1857 21468 1869 21471
rect 1780 21440 1869 21468
rect 1780 21344 1808 21440
rect 1857 21437 1869 21440
rect 1903 21437 1915 21471
rect 1857 21431 1915 21437
rect 4065 21471 4123 21477
rect 4065 21437 4077 21471
rect 4111 21468 4123 21471
rect 4617 21471 4675 21477
rect 4617 21468 4629 21471
rect 4111 21440 4629 21468
rect 4111 21437 4123 21440
rect 4065 21431 4123 21437
rect 4617 21437 4629 21440
rect 4663 21468 4675 21471
rect 5166 21468 5172 21480
rect 4663 21440 5172 21468
rect 4663 21437 4675 21440
rect 4617 21431 4675 21437
rect 5166 21428 5172 21440
rect 5224 21428 5230 21480
rect 7469 21471 7527 21477
rect 7469 21437 7481 21471
rect 7515 21468 7527 21471
rect 9030 21468 9036 21480
rect 7515 21440 9036 21468
rect 7515 21437 7527 21440
rect 7469 21431 7527 21437
rect 9030 21428 9036 21440
rect 9088 21428 9094 21480
rect 9766 21428 9772 21480
rect 9824 21468 9830 21480
rect 10413 21471 10471 21477
rect 10413 21468 10425 21471
rect 9824 21440 10425 21468
rect 9824 21428 9830 21440
rect 10413 21437 10425 21440
rect 10459 21437 10471 21471
rect 10413 21431 10471 21437
rect 6270 21400 6276 21412
rect 4540 21372 6276 21400
rect 1762 21332 1768 21344
rect 1723 21304 1768 21332
rect 1762 21292 1768 21304
rect 1820 21292 1826 21344
rect 3418 21292 3424 21344
rect 3476 21332 3482 21344
rect 4540 21341 4568 21372
rect 6270 21360 6276 21372
rect 6328 21360 6334 21412
rect 7736 21403 7794 21409
rect 7736 21369 7748 21403
rect 7782 21400 7794 21403
rect 8018 21400 8024 21412
rect 7782 21372 8024 21400
rect 7782 21369 7794 21372
rect 7736 21363 7794 21369
rect 8018 21360 8024 21372
rect 8076 21360 8082 21412
rect 9122 21360 9128 21412
rect 9180 21400 9186 21412
rect 9401 21403 9459 21409
rect 9401 21400 9413 21403
rect 9180 21372 9413 21400
rect 9180 21360 9186 21372
rect 9401 21369 9413 21372
rect 9447 21369 9459 21403
rect 9401 21363 9459 21369
rect 9674 21360 9680 21412
rect 9732 21400 9738 21412
rect 10321 21403 10379 21409
rect 10321 21400 10333 21403
rect 9732 21372 10333 21400
rect 9732 21360 9738 21372
rect 10321 21369 10333 21372
rect 10367 21400 10379 21403
rect 10965 21403 11023 21409
rect 10965 21400 10977 21403
rect 10367 21372 10977 21400
rect 10367 21369 10379 21372
rect 10321 21363 10379 21369
rect 10965 21369 10977 21372
rect 11011 21369 11023 21403
rect 10965 21363 11023 21369
rect 12158 21360 12164 21412
rect 12216 21400 12222 21412
rect 12897 21403 12955 21409
rect 12897 21400 12909 21403
rect 12216 21372 12909 21400
rect 12216 21360 12222 21372
rect 12897 21369 12909 21372
rect 12943 21369 12955 21403
rect 14246 21403 14304 21409
rect 14246 21400 14258 21403
rect 12897 21363 12955 21369
rect 13832 21372 14258 21400
rect 13832 21344 13860 21372
rect 14246 21369 14258 21372
rect 14292 21369 14304 21403
rect 14246 21363 14304 21369
rect 15470 21360 15476 21412
rect 15528 21400 15534 21412
rect 15528 21372 16436 21400
rect 15528 21360 15534 21372
rect 16408 21344 16436 21372
rect 3605 21335 3663 21341
rect 3605 21332 3617 21335
rect 3476 21304 3617 21332
rect 3476 21292 3482 21304
rect 3605 21301 3617 21304
rect 3651 21332 3663 21335
rect 4525 21335 4583 21341
rect 4525 21332 4537 21335
rect 3651 21304 4537 21332
rect 3651 21301 3663 21304
rect 3605 21295 3663 21301
rect 4525 21301 4537 21304
rect 4571 21301 4583 21335
rect 5626 21332 5632 21344
rect 5587 21304 5632 21332
rect 4525 21295 4583 21301
rect 5626 21292 5632 21304
rect 5684 21332 5690 21344
rect 6181 21335 6239 21341
rect 6181 21332 6193 21335
rect 5684 21304 6193 21332
rect 5684 21292 5690 21304
rect 6181 21301 6193 21304
rect 6227 21332 6239 21335
rect 6546 21332 6552 21344
rect 6227 21304 6552 21332
rect 6227 21301 6239 21304
rect 6181 21295 6239 21301
rect 6546 21292 6552 21304
rect 6604 21292 6610 21344
rect 8849 21335 8907 21341
rect 8849 21301 8861 21335
rect 8895 21332 8907 21335
rect 9306 21332 9312 21344
rect 8895 21304 9312 21332
rect 8895 21301 8907 21304
rect 8849 21295 8907 21301
rect 9306 21292 9312 21304
rect 9364 21292 9370 21344
rect 9766 21332 9772 21344
rect 9727 21304 9772 21332
rect 9766 21292 9772 21304
rect 9824 21292 9830 21344
rect 9950 21332 9956 21344
rect 9911 21304 9956 21332
rect 9950 21292 9956 21304
rect 10008 21292 10014 21344
rect 11882 21332 11888 21344
rect 11843 21304 11888 21332
rect 11882 21292 11888 21304
rect 11940 21292 11946 21344
rect 12434 21292 12440 21344
rect 12492 21332 12498 21344
rect 12802 21332 12808 21344
rect 12492 21304 12537 21332
rect 12763 21304 12808 21332
rect 12492 21292 12498 21304
rect 12802 21292 12808 21304
rect 12860 21292 12866 21344
rect 13446 21332 13452 21344
rect 13407 21304 13452 21332
rect 13446 21292 13452 21304
rect 13504 21292 13510 21344
rect 13814 21332 13820 21344
rect 13775 21304 13820 21332
rect 13814 21292 13820 21304
rect 13872 21292 13878 21344
rect 15381 21335 15439 21341
rect 15381 21301 15393 21335
rect 15427 21332 15439 21335
rect 15930 21332 15936 21344
rect 15427 21304 15936 21332
rect 15427 21301 15439 21304
rect 15381 21295 15439 21301
rect 15930 21292 15936 21304
rect 15988 21292 15994 21344
rect 16390 21332 16396 21344
rect 16351 21304 16396 21332
rect 16390 21292 16396 21304
rect 16448 21292 16454 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 1578 21128 1584 21140
rect 1539 21100 1584 21128
rect 1578 21088 1584 21100
rect 1636 21088 1642 21140
rect 4338 21128 4344 21140
rect 4299 21100 4344 21128
rect 4338 21088 4344 21100
rect 4396 21088 4402 21140
rect 8386 21128 8392 21140
rect 8347 21100 8392 21128
rect 8386 21088 8392 21100
rect 8444 21088 8450 21140
rect 12069 21131 12127 21137
rect 12069 21097 12081 21131
rect 12115 21128 12127 21131
rect 12434 21128 12440 21140
rect 12115 21100 12440 21128
rect 12115 21097 12127 21100
rect 12069 21091 12127 21097
rect 12434 21088 12440 21100
rect 12492 21128 12498 21140
rect 12897 21131 12955 21137
rect 12897 21128 12909 21131
rect 12492 21100 12909 21128
rect 12492 21088 12498 21100
rect 12897 21097 12909 21100
rect 12943 21097 12955 21131
rect 12897 21091 12955 21097
rect 13906 21088 13912 21140
rect 13964 21128 13970 21140
rect 14001 21131 14059 21137
rect 14001 21128 14013 21131
rect 13964 21100 14013 21128
rect 13964 21088 13970 21100
rect 14001 21097 14013 21100
rect 14047 21097 14059 21131
rect 14001 21091 14059 21097
rect 15286 21088 15292 21140
rect 15344 21128 15350 21140
rect 15749 21131 15807 21137
rect 15749 21128 15761 21131
rect 15344 21100 15761 21128
rect 15344 21088 15350 21100
rect 15749 21097 15761 21100
rect 15795 21128 15807 21131
rect 16022 21128 16028 21140
rect 15795 21100 16028 21128
rect 15795 21097 15807 21100
rect 15749 21091 15807 21097
rect 16022 21088 16028 21100
rect 16080 21088 16086 21140
rect 2225 21063 2283 21069
rect 2225 21029 2237 21063
rect 2271 21060 2283 21063
rect 2590 21060 2596 21072
rect 2271 21032 2596 21060
rect 2271 21029 2283 21032
rect 2225 21023 2283 21029
rect 2590 21020 2596 21032
rect 2648 21020 2654 21072
rect 5074 21020 5080 21072
rect 5132 21069 5138 21072
rect 5132 21063 5196 21069
rect 5132 21029 5150 21063
rect 5184 21029 5196 21063
rect 5132 21023 5196 21029
rect 9953 21063 10011 21069
rect 9953 21029 9965 21063
rect 9999 21060 10011 21063
rect 10042 21060 10048 21072
rect 9999 21032 10048 21060
rect 9999 21029 10011 21032
rect 9953 21023 10011 21029
rect 5132 21020 5138 21023
rect 10042 21020 10048 21032
rect 10100 21060 10106 21072
rect 10870 21060 10876 21072
rect 10100 21032 10876 21060
rect 10100 21020 10106 21032
rect 10870 21020 10876 21032
rect 10928 21020 10934 21072
rect 1946 20992 1952 21004
rect 1907 20964 1952 20992
rect 1946 20952 1952 20964
rect 2004 20952 2010 21004
rect 2777 20995 2835 21001
rect 2777 20961 2789 20995
rect 2823 20992 2835 20995
rect 3145 20995 3203 21001
rect 3145 20992 3157 20995
rect 2823 20964 3157 20992
rect 2823 20961 2835 20964
rect 2777 20955 2835 20961
rect 3145 20961 3157 20964
rect 3191 20992 3203 20995
rect 3878 20992 3884 21004
rect 3191 20964 3884 20992
rect 3191 20961 3203 20964
rect 3145 20955 3203 20961
rect 3878 20952 3884 20964
rect 3936 20992 3942 21004
rect 4801 20995 4859 21001
rect 4801 20992 4813 20995
rect 3936 20964 4813 20992
rect 3936 20952 3942 20964
rect 4801 20961 4813 20964
rect 4847 20992 4859 20995
rect 4893 20995 4951 21001
rect 4893 20992 4905 20995
rect 4847 20964 4905 20992
rect 4847 20961 4859 20964
rect 4801 20955 4859 20961
rect 4893 20961 4905 20964
rect 4939 20992 4951 20995
rect 5626 20992 5632 21004
rect 4939 20964 5632 20992
rect 4939 20961 4951 20964
rect 4893 20955 4951 20961
rect 5626 20952 5632 20964
rect 5684 20992 5690 21004
rect 6270 20992 6276 21004
rect 5684 20964 6276 20992
rect 5684 20952 5690 20964
rect 6270 20952 6276 20964
rect 6328 20952 6334 21004
rect 7745 20995 7803 21001
rect 7745 20961 7757 20995
rect 7791 20992 7803 20995
rect 8202 20992 8208 21004
rect 7791 20964 8208 20992
rect 7791 20961 7803 20964
rect 7745 20955 7803 20961
rect 8202 20952 8208 20964
rect 8260 20952 8266 21004
rect 10312 20995 10370 21001
rect 10312 20961 10324 20995
rect 10358 20992 10370 20995
rect 10686 20992 10692 21004
rect 10358 20964 10692 20992
rect 10358 20961 10370 20964
rect 10312 20955 10370 20961
rect 10686 20952 10692 20964
rect 10744 20952 10750 21004
rect 12526 20952 12532 21004
rect 12584 20992 12590 21004
rect 13814 20992 13820 21004
rect 12584 20964 13820 20992
rect 12584 20952 12590 20964
rect 7098 20884 7104 20936
rect 7156 20924 7162 20936
rect 7834 20924 7840 20936
rect 7156 20896 7840 20924
rect 7156 20884 7162 20896
rect 7834 20884 7840 20896
rect 7892 20884 7898 20936
rect 8018 20924 8024 20936
rect 7979 20896 8024 20924
rect 8018 20884 8024 20896
rect 8076 20884 8082 20936
rect 10045 20927 10103 20933
rect 10045 20924 10057 20927
rect 9048 20896 10057 20924
rect 7285 20859 7343 20865
rect 7285 20825 7297 20859
rect 7331 20856 7343 20859
rect 8036 20856 8064 20884
rect 7331 20828 8064 20856
rect 7331 20825 7343 20828
rect 7285 20819 7343 20825
rect 9048 20800 9076 20896
rect 10045 20893 10057 20896
rect 10091 20893 10103 20927
rect 10045 20887 10103 20893
rect 12437 20927 12495 20933
rect 12437 20893 12449 20927
rect 12483 20924 12495 20927
rect 12986 20924 12992 20936
rect 12483 20896 12992 20924
rect 12483 20893 12495 20896
rect 12437 20887 12495 20893
rect 12986 20884 12992 20896
rect 13044 20884 13050 20936
rect 13096 20933 13124 20964
rect 13814 20952 13820 20964
rect 13872 20952 13878 21004
rect 15286 20952 15292 21004
rect 15344 20992 15350 21004
rect 15657 20995 15715 21001
rect 15657 20992 15669 20995
rect 15344 20964 15669 20992
rect 15344 20952 15350 20964
rect 15657 20961 15669 20964
rect 15703 20961 15715 20995
rect 15657 20955 15715 20961
rect 13081 20927 13139 20933
rect 13081 20893 13093 20927
rect 13127 20893 13139 20927
rect 13081 20887 13139 20893
rect 14185 20927 14243 20933
rect 14185 20893 14197 20927
rect 14231 20924 14243 20927
rect 14550 20924 14556 20936
rect 14231 20896 14556 20924
rect 14231 20893 14243 20896
rect 14185 20887 14243 20893
rect 14550 20884 14556 20896
rect 14608 20884 14614 20936
rect 15838 20924 15844 20936
rect 15799 20896 15844 20924
rect 15838 20884 15844 20896
rect 15896 20884 15902 20936
rect 12526 20856 12532 20868
rect 12487 20828 12532 20856
rect 12526 20816 12532 20828
rect 12584 20816 12590 20868
rect 15289 20859 15347 20865
rect 15289 20825 15301 20859
rect 15335 20856 15347 20859
rect 15378 20856 15384 20868
rect 15335 20828 15384 20856
rect 15335 20825 15347 20828
rect 15289 20819 15347 20825
rect 15378 20816 15384 20828
rect 15436 20816 15442 20868
rect 5534 20748 5540 20800
rect 5592 20788 5598 20800
rect 6273 20791 6331 20797
rect 6273 20788 6285 20791
rect 5592 20760 6285 20788
rect 5592 20748 5598 20760
rect 6273 20757 6285 20760
rect 6319 20788 6331 20791
rect 6825 20791 6883 20797
rect 6825 20788 6837 20791
rect 6319 20760 6837 20788
rect 6319 20757 6331 20760
rect 6273 20751 6331 20757
rect 6825 20757 6837 20760
rect 6871 20788 6883 20791
rect 6914 20788 6920 20800
rect 6871 20760 6920 20788
rect 6871 20757 6883 20760
rect 6825 20751 6883 20757
rect 6914 20748 6920 20760
rect 6972 20748 6978 20800
rect 7374 20788 7380 20800
rect 7335 20760 7380 20788
rect 7374 20748 7380 20760
rect 7432 20748 7438 20800
rect 9030 20788 9036 20800
rect 8991 20760 9036 20788
rect 9030 20748 9036 20760
rect 9088 20748 9094 20800
rect 9398 20788 9404 20800
rect 9359 20760 9404 20788
rect 9398 20748 9404 20760
rect 9456 20748 9462 20800
rect 11425 20791 11483 20797
rect 11425 20757 11437 20791
rect 11471 20788 11483 20791
rect 11606 20788 11612 20800
rect 11471 20760 11612 20788
rect 11471 20757 11483 20760
rect 11425 20751 11483 20757
rect 11606 20748 11612 20760
rect 11664 20748 11670 20800
rect 13354 20748 13360 20800
rect 13412 20788 13418 20800
rect 13541 20791 13599 20797
rect 13541 20788 13553 20791
rect 13412 20760 13553 20788
rect 13412 20748 13418 20760
rect 13541 20757 13553 20760
rect 13587 20757 13599 20791
rect 13541 20751 13599 20757
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 1670 20584 1676 20596
rect 1631 20556 1676 20584
rect 1670 20544 1676 20556
rect 1728 20544 1734 20596
rect 1946 20544 1952 20596
rect 2004 20584 2010 20596
rect 2498 20584 2504 20596
rect 2004 20556 2504 20584
rect 2004 20544 2010 20556
rect 2498 20544 2504 20556
rect 2556 20544 2562 20596
rect 8202 20544 8208 20596
rect 8260 20584 8266 20596
rect 8941 20587 8999 20593
rect 8941 20584 8953 20587
rect 8260 20556 8953 20584
rect 8260 20544 8266 20556
rect 8941 20553 8953 20556
rect 8987 20553 8999 20587
rect 11882 20584 11888 20596
rect 11843 20556 11888 20584
rect 8941 20547 8999 20553
rect 11882 20544 11888 20556
rect 11940 20544 11946 20596
rect 12253 20587 12311 20593
rect 12253 20553 12265 20587
rect 12299 20584 12311 20587
rect 12342 20584 12348 20596
rect 12299 20556 12348 20584
rect 12299 20553 12311 20556
rect 12253 20547 12311 20553
rect 12342 20544 12348 20556
rect 12400 20544 12406 20596
rect 13814 20544 13820 20596
rect 13872 20584 13878 20596
rect 14001 20587 14059 20593
rect 14001 20584 14013 20587
rect 13872 20556 14013 20584
rect 13872 20544 13878 20556
rect 14001 20553 14013 20556
rect 14047 20553 14059 20587
rect 14550 20584 14556 20596
rect 14511 20556 14556 20584
rect 14001 20547 14059 20553
rect 14550 20544 14556 20556
rect 14608 20544 14614 20596
rect 15838 20544 15844 20596
rect 15896 20584 15902 20596
rect 16117 20587 16175 20593
rect 16117 20584 16129 20587
rect 15896 20556 16129 20584
rect 15896 20544 15902 20556
rect 16117 20553 16129 20556
rect 16163 20553 16175 20587
rect 16117 20547 16175 20553
rect 4341 20519 4399 20525
rect 4341 20485 4353 20519
rect 4387 20516 4399 20519
rect 5074 20516 5080 20528
rect 4387 20488 5080 20516
rect 4387 20485 4399 20488
rect 4341 20479 4399 20485
rect 5074 20476 5080 20488
rect 5132 20476 5138 20528
rect 7834 20476 7840 20528
rect 7892 20516 7898 20528
rect 8757 20519 8815 20525
rect 8757 20516 8769 20519
rect 7892 20488 8769 20516
rect 7892 20476 7898 20488
rect 8757 20485 8769 20488
rect 8803 20485 8815 20519
rect 8757 20479 8815 20485
rect 2038 20448 2044 20460
rect 1999 20420 2044 20448
rect 2038 20408 2044 20420
rect 2096 20408 2102 20460
rect 4709 20451 4767 20457
rect 4709 20417 4721 20451
rect 4755 20448 4767 20451
rect 5353 20451 5411 20457
rect 5353 20448 5365 20451
rect 4755 20420 5365 20448
rect 4755 20417 4767 20420
rect 4709 20411 4767 20417
rect 5353 20417 5365 20420
rect 5399 20448 5411 20451
rect 5442 20448 5448 20460
rect 5399 20420 5448 20448
rect 5399 20417 5411 20420
rect 5353 20411 5411 20417
rect 5442 20408 5448 20420
rect 5500 20408 5506 20460
rect 11900 20448 11928 20544
rect 15105 20519 15163 20525
rect 15105 20485 15117 20519
rect 15151 20516 15163 20519
rect 15286 20516 15292 20528
rect 15151 20488 15292 20516
rect 15151 20485 15163 20488
rect 15105 20479 15163 20485
rect 15286 20476 15292 20488
rect 15344 20476 15350 20528
rect 12437 20451 12495 20457
rect 12437 20448 12449 20451
rect 11900 20420 12449 20448
rect 12437 20417 12449 20420
rect 12483 20417 12495 20451
rect 12437 20411 12495 20417
rect 15749 20451 15807 20457
rect 15749 20417 15761 20451
rect 15795 20448 15807 20451
rect 15930 20448 15936 20460
rect 15795 20420 15936 20448
rect 15795 20417 15807 20420
rect 15749 20411 15807 20417
rect 15930 20408 15936 20420
rect 15988 20448 15994 20460
rect 16485 20451 16543 20457
rect 16485 20448 16497 20451
rect 15988 20420 16497 20448
rect 15988 20408 15994 20420
rect 16485 20417 16497 20420
rect 16531 20417 16543 20451
rect 16666 20448 16672 20460
rect 16627 20420 16672 20448
rect 16485 20411 16543 20417
rect 16666 20408 16672 20420
rect 16724 20408 16730 20460
rect 1670 20340 1676 20392
rect 1728 20380 1734 20392
rect 1765 20383 1823 20389
rect 1765 20380 1777 20383
rect 1728 20352 1777 20380
rect 1728 20340 1734 20352
rect 1765 20349 1777 20352
rect 1811 20349 1823 20383
rect 3053 20383 3111 20389
rect 3053 20380 3065 20383
rect 1765 20343 1823 20349
rect 2884 20352 3065 20380
rect 2884 20256 2912 20352
rect 3053 20349 3065 20352
rect 3099 20349 3111 20383
rect 3053 20343 3111 20349
rect 3973 20383 4031 20389
rect 3973 20349 3985 20383
rect 4019 20380 4031 20383
rect 5261 20383 5319 20389
rect 5261 20380 5273 20383
rect 4019 20352 5273 20380
rect 4019 20349 4031 20352
rect 3973 20343 4031 20349
rect 5261 20349 5273 20352
rect 5307 20380 5319 20383
rect 5902 20380 5908 20392
rect 5307 20352 5908 20380
rect 5307 20349 5319 20352
rect 5261 20343 5319 20349
rect 5902 20340 5908 20352
rect 5960 20340 5966 20392
rect 6273 20383 6331 20389
rect 6273 20349 6285 20383
rect 6319 20380 6331 20383
rect 6546 20380 6552 20392
rect 6319 20352 6552 20380
rect 6319 20349 6331 20352
rect 6273 20343 6331 20349
rect 6546 20340 6552 20352
rect 6604 20340 6610 20392
rect 6825 20383 6883 20389
rect 6825 20349 6837 20383
rect 6871 20349 6883 20383
rect 6825 20343 6883 20349
rect 4338 20272 4344 20324
rect 4396 20312 4402 20324
rect 5169 20315 5227 20321
rect 5169 20312 5181 20315
rect 4396 20284 5181 20312
rect 4396 20272 4402 20284
rect 5169 20281 5181 20284
rect 5215 20312 5227 20315
rect 5813 20315 5871 20321
rect 5813 20312 5825 20315
rect 5215 20284 5825 20312
rect 5215 20281 5227 20284
rect 5169 20275 5227 20281
rect 5813 20281 5825 20284
rect 5859 20281 5871 20315
rect 6840 20312 6868 20343
rect 6914 20340 6920 20392
rect 6972 20380 6978 20392
rect 7081 20383 7139 20389
rect 7081 20380 7093 20383
rect 6972 20352 7093 20380
rect 6972 20340 6978 20352
rect 7081 20349 7093 20352
rect 7127 20349 7139 20383
rect 7081 20343 7139 20349
rect 9030 20340 9036 20392
rect 9088 20380 9094 20392
rect 9309 20383 9367 20389
rect 9309 20380 9321 20383
rect 9088 20352 9321 20380
rect 9088 20340 9094 20352
rect 9309 20349 9321 20352
rect 9355 20349 9367 20383
rect 9309 20343 9367 20349
rect 11330 20340 11336 20392
rect 11388 20380 11394 20392
rect 12621 20383 12679 20389
rect 12621 20380 12633 20383
rect 11388 20352 12633 20380
rect 11388 20340 11394 20352
rect 12621 20349 12633 20352
rect 12667 20380 12679 20383
rect 13354 20380 13360 20392
rect 12667 20352 13360 20380
rect 12667 20349 12679 20352
rect 12621 20343 12679 20349
rect 13354 20340 13360 20352
rect 13412 20340 13418 20392
rect 14550 20340 14556 20392
rect 14608 20380 14614 20392
rect 15473 20383 15531 20389
rect 15473 20380 15485 20383
rect 14608 20352 15485 20380
rect 14608 20340 14614 20352
rect 15473 20349 15485 20352
rect 15519 20349 15531 20383
rect 15473 20343 15531 20349
rect 5813 20275 5871 20281
rect 6380 20284 6868 20312
rect 2866 20244 2872 20256
rect 2827 20216 2872 20244
rect 2866 20204 2872 20216
rect 2924 20204 2930 20256
rect 3234 20244 3240 20256
rect 3195 20216 3240 20244
rect 3234 20204 3240 20216
rect 3292 20204 3298 20256
rect 4798 20244 4804 20256
rect 4759 20216 4804 20244
rect 4798 20204 4804 20216
rect 4856 20204 4862 20256
rect 6270 20204 6276 20256
rect 6328 20244 6334 20256
rect 6380 20253 6408 20284
rect 7742 20272 7748 20324
rect 7800 20312 7806 20324
rect 9398 20312 9404 20324
rect 7800 20284 9404 20312
rect 7800 20272 7806 20284
rect 9398 20272 9404 20284
rect 9456 20312 9462 20324
rect 9554 20315 9612 20321
rect 9554 20312 9566 20315
rect 9456 20284 9566 20312
rect 9456 20272 9462 20284
rect 9554 20281 9566 20284
rect 9600 20281 9612 20315
rect 9554 20275 9612 20281
rect 12437 20315 12495 20321
rect 12437 20281 12449 20315
rect 12483 20312 12495 20315
rect 12710 20312 12716 20324
rect 12483 20284 12716 20312
rect 12483 20281 12495 20284
rect 12437 20275 12495 20281
rect 12710 20272 12716 20284
rect 12768 20312 12774 20324
rect 12866 20315 12924 20321
rect 12866 20312 12878 20315
rect 12768 20284 12878 20312
rect 12768 20272 12774 20284
rect 12866 20281 12878 20284
rect 12912 20281 12924 20315
rect 12866 20275 12924 20281
rect 6365 20247 6423 20253
rect 6365 20244 6377 20247
rect 6328 20216 6377 20244
rect 6328 20204 6334 20216
rect 6365 20213 6377 20216
rect 6411 20213 6423 20247
rect 6365 20207 6423 20213
rect 8018 20204 8024 20256
rect 8076 20244 8082 20256
rect 8205 20247 8263 20253
rect 8205 20244 8217 20247
rect 8076 20216 8217 20244
rect 8076 20204 8082 20216
rect 8205 20213 8217 20216
rect 8251 20244 8263 20247
rect 8570 20244 8576 20256
rect 8251 20216 8576 20244
rect 8251 20213 8263 20216
rect 8205 20207 8263 20213
rect 8570 20204 8576 20216
rect 8628 20204 8634 20256
rect 8941 20247 8999 20253
rect 8941 20213 8953 20247
rect 8987 20244 8999 20247
rect 9217 20247 9275 20253
rect 9217 20244 9229 20247
rect 8987 20216 9229 20244
rect 8987 20213 8999 20216
rect 8941 20207 8999 20213
rect 9217 20213 9229 20216
rect 9263 20244 9275 20247
rect 9766 20244 9772 20256
rect 9263 20216 9772 20244
rect 9263 20213 9275 20216
rect 9217 20207 9275 20213
rect 9766 20204 9772 20216
rect 9824 20204 9830 20256
rect 10686 20244 10692 20256
rect 10647 20216 10692 20244
rect 10686 20204 10692 20216
rect 10744 20244 10750 20256
rect 11241 20247 11299 20253
rect 11241 20244 11253 20247
rect 10744 20216 11253 20244
rect 10744 20204 10750 20216
rect 11241 20213 11253 20216
rect 11287 20213 11299 20247
rect 11241 20207 11299 20213
rect 15013 20247 15071 20253
rect 15013 20213 15025 20247
rect 15059 20244 15071 20247
rect 15378 20244 15384 20256
rect 15059 20216 15384 20244
rect 15059 20213 15071 20216
rect 15013 20207 15071 20213
rect 15378 20204 15384 20216
rect 15436 20244 15442 20256
rect 15565 20247 15623 20253
rect 15565 20244 15577 20247
rect 15436 20216 15577 20244
rect 15436 20204 15442 20216
rect 15565 20213 15577 20216
rect 15611 20213 15623 20247
rect 15565 20207 15623 20213
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 3878 20040 3884 20052
rect 3839 20012 3884 20040
rect 3878 20000 3884 20012
rect 3936 20000 3942 20052
rect 4338 20040 4344 20052
rect 4299 20012 4344 20040
rect 4338 20000 4344 20012
rect 4396 20000 4402 20052
rect 5902 20040 5908 20052
rect 5863 20012 5908 20040
rect 5902 20000 5908 20012
rect 5960 20000 5966 20052
rect 6273 20043 6331 20049
rect 6273 20009 6285 20043
rect 6319 20040 6331 20043
rect 6822 20040 6828 20052
rect 6319 20012 6828 20040
rect 6319 20009 6331 20012
rect 6273 20003 6331 20009
rect 6822 20000 6828 20012
rect 6880 20000 6886 20052
rect 7374 20000 7380 20052
rect 7432 20040 7438 20052
rect 7837 20043 7895 20049
rect 7837 20040 7849 20043
rect 7432 20012 7849 20040
rect 7432 20000 7438 20012
rect 7837 20009 7849 20012
rect 7883 20040 7895 20043
rect 8849 20043 8907 20049
rect 8849 20040 8861 20043
rect 7883 20012 8861 20040
rect 7883 20009 7895 20012
rect 7837 20003 7895 20009
rect 8849 20009 8861 20012
rect 8895 20009 8907 20043
rect 8849 20003 8907 20009
rect 9950 20000 9956 20052
rect 10008 20040 10014 20052
rect 10137 20043 10195 20049
rect 10137 20040 10149 20043
rect 10008 20012 10149 20040
rect 10008 20000 10014 20012
rect 10137 20009 10149 20012
rect 10183 20009 10195 20043
rect 12710 20040 12716 20052
rect 12671 20012 12716 20040
rect 10137 20003 10195 20009
rect 12710 20000 12716 20012
rect 12768 20040 12774 20052
rect 13265 20043 13323 20049
rect 13265 20040 13277 20043
rect 12768 20012 13277 20040
rect 12768 20000 12774 20012
rect 13265 20009 13277 20012
rect 13311 20040 13323 20043
rect 13538 20040 13544 20052
rect 13311 20012 13544 20040
rect 13311 20009 13323 20012
rect 13265 20003 13323 20009
rect 13538 20000 13544 20012
rect 13596 20000 13602 20052
rect 15105 20043 15163 20049
rect 15105 20009 15117 20043
rect 15151 20040 15163 20043
rect 15286 20040 15292 20052
rect 15151 20012 15292 20040
rect 15151 20009 15163 20012
rect 15105 20003 15163 20009
rect 15286 20000 15292 20012
rect 15344 20000 15350 20052
rect 16022 20040 16028 20052
rect 15983 20012 16028 20040
rect 16022 20000 16028 20012
rect 16080 20000 16086 20052
rect 16761 20043 16819 20049
rect 16761 20009 16773 20043
rect 16807 20040 16819 20043
rect 17402 20040 17408 20052
rect 16807 20012 17408 20040
rect 16807 20009 16819 20012
rect 16761 20003 16819 20009
rect 17402 20000 17408 20012
rect 17460 20000 17466 20052
rect 1673 19975 1731 19981
rect 1673 19941 1685 19975
rect 1719 19972 1731 19975
rect 2590 19972 2596 19984
rect 1719 19944 2596 19972
rect 1719 19941 1731 19944
rect 1673 19935 1731 19941
rect 2590 19932 2596 19944
rect 2648 19932 2654 19984
rect 2958 19972 2964 19984
rect 2919 19944 2964 19972
rect 2958 19932 2964 19944
rect 3016 19932 3022 19984
rect 3694 19932 3700 19984
rect 3752 19972 3758 19984
rect 6917 19975 6975 19981
rect 6917 19972 6929 19975
rect 3752 19944 6929 19972
rect 3752 19932 3758 19944
rect 6917 19941 6929 19944
rect 6963 19972 6975 19975
rect 7282 19972 7288 19984
rect 6963 19944 7288 19972
rect 6963 19941 6975 19944
rect 6917 19935 6975 19941
rect 7282 19932 7288 19944
rect 7340 19932 7346 19984
rect 10594 19932 10600 19984
rect 10652 19972 10658 19984
rect 10870 19972 10876 19984
rect 10652 19944 10876 19972
rect 10652 19932 10658 19944
rect 10870 19932 10876 19944
rect 10928 19932 10934 19984
rect 14090 19972 14096 19984
rect 14051 19944 14096 19972
rect 14090 19932 14096 19944
rect 14148 19932 14154 19984
rect 1397 19907 1455 19913
rect 1397 19873 1409 19907
rect 1443 19904 1455 19907
rect 2682 19904 2688 19916
rect 1443 19876 2268 19904
rect 2595 19876 2688 19904
rect 1443 19873 1455 19876
rect 1397 19867 1455 19873
rect 2240 19848 2268 19876
rect 2682 19864 2688 19876
rect 2740 19904 2746 19916
rect 2774 19904 2780 19916
rect 2740 19876 2780 19904
rect 2740 19864 2746 19876
rect 2774 19864 2780 19876
rect 2832 19864 2838 19916
rect 4706 19904 4712 19916
rect 4667 19876 4712 19904
rect 4706 19864 4712 19876
rect 4764 19864 4770 19916
rect 4801 19907 4859 19913
rect 4801 19873 4813 19907
rect 4847 19873 4859 19907
rect 4801 19867 4859 19873
rect 6365 19907 6423 19913
rect 6365 19873 6377 19907
rect 6411 19904 6423 19907
rect 6638 19904 6644 19916
rect 6411 19876 6644 19904
rect 6411 19873 6423 19876
rect 6365 19867 6423 19873
rect 2222 19836 2228 19848
rect 2183 19808 2228 19836
rect 2222 19796 2228 19808
rect 2280 19796 2286 19848
rect 4338 19796 4344 19848
rect 4396 19836 4402 19848
rect 4522 19836 4528 19848
rect 4396 19808 4528 19836
rect 4396 19796 4402 19808
rect 4522 19796 4528 19808
rect 4580 19796 4586 19848
rect 4816 19780 4844 19867
rect 6638 19864 6644 19876
rect 6696 19864 6702 19916
rect 7929 19907 7987 19913
rect 7929 19873 7941 19907
rect 7975 19904 7987 19907
rect 8294 19904 8300 19916
rect 7975 19876 8300 19904
rect 7975 19873 7987 19876
rect 7929 19867 7987 19873
rect 8294 19864 8300 19876
rect 8352 19864 8358 19916
rect 9122 19864 9128 19916
rect 9180 19904 9186 19916
rect 11606 19913 11612 19916
rect 9217 19907 9275 19913
rect 9217 19904 9229 19907
rect 9180 19876 9229 19904
rect 9180 19864 9186 19876
rect 9217 19873 9229 19876
rect 9263 19873 9275 19907
rect 11589 19907 11612 19913
rect 11589 19904 11601 19907
rect 9217 19867 9275 19873
rect 10336 19876 11601 19904
rect 10336 19848 10364 19876
rect 11589 19873 11601 19876
rect 11664 19904 11670 19916
rect 13814 19904 13820 19916
rect 11664 19876 11737 19904
rect 13775 19876 13820 19904
rect 11589 19867 11612 19873
rect 11606 19864 11612 19867
rect 11664 19864 11670 19876
rect 13814 19864 13820 19876
rect 13872 19864 13878 19916
rect 15286 19904 15292 19916
rect 15247 19876 15292 19904
rect 15286 19864 15292 19876
rect 15344 19864 15350 19916
rect 15565 19907 15623 19913
rect 15565 19873 15577 19907
rect 15611 19904 15623 19907
rect 16574 19904 16580 19916
rect 15611 19876 16580 19904
rect 15611 19873 15623 19876
rect 15565 19867 15623 19873
rect 16574 19864 16580 19876
rect 16632 19864 16638 19916
rect 4985 19839 5043 19845
rect 4985 19805 4997 19839
rect 5031 19805 5043 19839
rect 6546 19836 6552 19848
rect 6507 19808 6552 19836
rect 4985 19799 5043 19805
rect 4798 19728 4804 19780
rect 4856 19728 4862 19780
rect 5000 19768 5028 19799
rect 6546 19796 6552 19808
rect 6604 19796 6610 19848
rect 7742 19796 7748 19848
rect 7800 19836 7806 19848
rect 8021 19839 8079 19845
rect 8021 19836 8033 19839
rect 7800 19808 8033 19836
rect 7800 19796 7806 19808
rect 8021 19805 8033 19808
rect 8067 19805 8079 19839
rect 10226 19836 10232 19848
rect 10187 19808 10232 19836
rect 8021 19799 8079 19805
rect 10226 19796 10232 19808
rect 10284 19796 10290 19848
rect 10318 19796 10324 19848
rect 10376 19836 10382 19848
rect 11333 19839 11391 19845
rect 10376 19808 10421 19836
rect 10376 19796 10382 19808
rect 11333 19805 11345 19839
rect 11379 19805 11391 19839
rect 11333 19799 11391 19805
rect 5074 19768 5080 19780
rect 4987 19740 5080 19768
rect 5074 19728 5080 19740
rect 5132 19768 5138 19780
rect 5813 19771 5871 19777
rect 5813 19768 5825 19771
rect 5132 19740 5825 19768
rect 5132 19728 5138 19740
rect 5813 19737 5825 19740
rect 5859 19768 5871 19771
rect 6564 19768 6592 19796
rect 5859 19740 6592 19768
rect 5859 19737 5871 19740
rect 5813 19731 5871 19737
rect 7006 19728 7012 19780
rect 7064 19768 7070 19780
rect 7469 19771 7527 19777
rect 7469 19768 7481 19771
rect 7064 19740 7481 19768
rect 7064 19728 7070 19740
rect 7469 19737 7481 19740
rect 7515 19737 7527 19771
rect 7469 19731 7527 19737
rect 9769 19771 9827 19777
rect 9769 19737 9781 19771
rect 9815 19768 9827 19771
rect 10042 19768 10048 19780
rect 9815 19740 10048 19768
rect 9815 19737 9827 19740
rect 9769 19731 9827 19737
rect 10042 19728 10048 19740
rect 10100 19728 10106 19780
rect 11348 19712 11376 19799
rect 1946 19660 1952 19712
rect 2004 19700 2010 19712
rect 2501 19703 2559 19709
rect 2501 19700 2513 19703
rect 2004 19672 2513 19700
rect 2004 19660 2010 19672
rect 2501 19669 2513 19672
rect 2547 19669 2559 19703
rect 2501 19663 2559 19669
rect 2590 19660 2596 19712
rect 2648 19700 2654 19712
rect 3421 19703 3479 19709
rect 3421 19700 3433 19703
rect 2648 19672 3433 19700
rect 2648 19660 2654 19672
rect 3421 19669 3433 19672
rect 3467 19669 3479 19703
rect 3421 19663 3479 19669
rect 5258 19660 5264 19712
rect 5316 19700 5322 19712
rect 5353 19703 5411 19709
rect 5353 19700 5365 19703
rect 5316 19672 5365 19700
rect 5316 19660 5322 19672
rect 5353 19669 5365 19672
rect 5399 19669 5411 19703
rect 7374 19700 7380 19712
rect 7335 19672 7380 19700
rect 5353 19663 5411 19669
rect 7374 19660 7380 19672
rect 7432 19660 7438 19712
rect 8570 19700 8576 19712
rect 8531 19672 8576 19700
rect 8570 19660 8576 19672
rect 8628 19660 8634 19712
rect 9030 19700 9036 19712
rect 8991 19672 9036 19700
rect 9030 19660 9036 19672
rect 9088 19660 9094 19712
rect 10870 19700 10876 19712
rect 10831 19672 10876 19700
rect 10870 19660 10876 19672
rect 10928 19660 10934 19712
rect 11241 19703 11299 19709
rect 11241 19669 11253 19703
rect 11287 19700 11299 19703
rect 11330 19700 11336 19712
rect 11287 19672 11336 19700
rect 11287 19669 11299 19672
rect 11241 19663 11299 19669
rect 11330 19660 11336 19672
rect 11388 19660 11394 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 6549 19499 6607 19505
rect 6549 19465 6561 19499
rect 6595 19496 6607 19499
rect 6638 19496 6644 19508
rect 6595 19468 6644 19496
rect 6595 19465 6607 19468
rect 6549 19459 6607 19465
rect 6638 19456 6644 19468
rect 6696 19456 6702 19508
rect 9861 19499 9919 19505
rect 9861 19465 9873 19499
rect 9907 19496 9919 19499
rect 10318 19496 10324 19508
rect 9907 19468 10324 19496
rect 9907 19465 9919 19468
rect 9861 19459 9919 19465
rect 10318 19456 10324 19468
rect 10376 19456 10382 19508
rect 11606 19456 11612 19508
rect 11664 19496 11670 19508
rect 11793 19499 11851 19505
rect 11793 19496 11805 19499
rect 11664 19468 11805 19496
rect 11664 19456 11670 19468
rect 11793 19465 11805 19468
rect 11839 19465 11851 19499
rect 12986 19496 12992 19508
rect 12947 19468 12992 19496
rect 11793 19459 11851 19465
rect 12986 19456 12992 19468
rect 13044 19456 13050 19508
rect 16574 19456 16580 19508
rect 16632 19496 16638 19508
rect 17313 19499 17371 19505
rect 17313 19496 17325 19499
rect 16632 19468 17325 19496
rect 16632 19456 16638 19468
rect 17313 19465 17325 19468
rect 17359 19465 17371 19499
rect 17313 19459 17371 19465
rect 10226 19388 10232 19440
rect 10284 19428 10290 19440
rect 10781 19431 10839 19437
rect 10781 19428 10793 19431
rect 10284 19400 10793 19428
rect 10284 19388 10290 19400
rect 10781 19397 10793 19400
rect 10827 19397 10839 19431
rect 10781 19391 10839 19397
rect 2133 19363 2191 19369
rect 2133 19329 2145 19363
rect 2179 19360 2191 19363
rect 7282 19360 7288 19372
rect 2179 19332 2636 19360
rect 7243 19332 7288 19360
rect 2179 19329 2191 19332
rect 2133 19323 2191 19329
rect 1394 19252 1400 19304
rect 1452 19292 1458 19304
rect 1857 19295 1915 19301
rect 1857 19292 1869 19295
rect 1452 19264 1869 19292
rect 1452 19252 1458 19264
rect 1857 19261 1869 19264
rect 1903 19292 1915 19295
rect 2498 19292 2504 19304
rect 1903 19264 2504 19292
rect 1903 19261 1915 19264
rect 1857 19255 1915 19261
rect 2498 19252 2504 19264
rect 2556 19252 2562 19304
rect 1486 19156 1492 19168
rect 1447 19128 1492 19156
rect 1486 19116 1492 19128
rect 1544 19116 1550 19168
rect 1946 19156 1952 19168
rect 1907 19128 1952 19156
rect 1946 19116 1952 19128
rect 2004 19116 2010 19168
rect 2608 19165 2636 19332
rect 7282 19320 7288 19332
rect 7340 19320 7346 19372
rect 7469 19363 7527 19369
rect 7469 19329 7481 19363
rect 7515 19360 7527 19363
rect 8202 19360 8208 19372
rect 7515 19332 8208 19360
rect 7515 19329 7527 19332
rect 7469 19323 7527 19329
rect 8202 19320 8208 19332
rect 8260 19320 8266 19372
rect 8570 19320 8576 19372
rect 8628 19360 8634 19372
rect 8941 19363 8999 19369
rect 8941 19360 8953 19363
rect 8628 19332 8953 19360
rect 8628 19320 8634 19332
rect 8941 19329 8953 19332
rect 8987 19329 8999 19363
rect 8941 19323 8999 19329
rect 10321 19363 10379 19369
rect 10321 19329 10333 19363
rect 10367 19360 10379 19363
rect 10686 19360 10692 19372
rect 10367 19332 10692 19360
rect 10367 19329 10379 19332
rect 10321 19323 10379 19329
rect 10686 19320 10692 19332
rect 10744 19360 10750 19372
rect 11333 19363 11391 19369
rect 11333 19360 11345 19363
rect 10744 19332 11345 19360
rect 10744 19320 10750 19332
rect 11333 19329 11345 19332
rect 11379 19329 11391 19363
rect 13538 19360 13544 19372
rect 13499 19332 13544 19360
rect 11333 19323 11391 19329
rect 13538 19320 13544 19332
rect 13596 19320 13602 19372
rect 15286 19360 15292 19372
rect 15120 19332 15292 19360
rect 3053 19295 3111 19301
rect 3053 19261 3065 19295
rect 3099 19292 3111 19295
rect 3142 19292 3148 19304
rect 3099 19264 3148 19292
rect 3099 19261 3111 19264
rect 3053 19255 3111 19261
rect 3142 19252 3148 19264
rect 3200 19292 3206 19304
rect 3878 19292 3884 19304
rect 3200 19264 3884 19292
rect 3200 19252 3206 19264
rect 3878 19252 3884 19264
rect 3936 19252 3942 19304
rect 5534 19292 5540 19304
rect 5495 19264 5540 19292
rect 5534 19252 5540 19264
rect 5592 19252 5598 19304
rect 6181 19295 6239 19301
rect 6181 19261 6193 19295
rect 6227 19292 6239 19295
rect 6822 19292 6828 19304
rect 6227 19264 6828 19292
rect 6227 19261 6239 19264
rect 6181 19255 6239 19261
rect 6822 19252 6828 19264
rect 6880 19252 6886 19304
rect 8297 19295 8355 19301
rect 8297 19261 8309 19295
rect 8343 19292 8355 19295
rect 8754 19292 8760 19304
rect 8343 19264 8760 19292
rect 8343 19261 8355 19264
rect 8297 19255 8355 19261
rect 8754 19252 8760 19264
rect 8812 19252 8818 19304
rect 9493 19295 9551 19301
rect 9493 19261 9505 19295
rect 9539 19292 9551 19295
rect 10226 19292 10232 19304
rect 9539 19264 10232 19292
rect 9539 19261 9551 19264
rect 9493 19255 9551 19261
rect 10226 19252 10232 19264
rect 10284 19252 10290 19304
rect 11238 19292 11244 19304
rect 11199 19264 11244 19292
rect 11238 19252 11244 19264
rect 11296 19252 11302 19304
rect 12434 19252 12440 19304
rect 12492 19292 12498 19304
rect 13630 19292 13636 19304
rect 12492 19264 13636 19292
rect 12492 19252 12498 19264
rect 13630 19252 13636 19264
rect 13688 19252 13694 19304
rect 13722 19252 13728 19304
rect 13780 19292 13786 19304
rect 14829 19295 14887 19301
rect 14829 19292 14841 19295
rect 13780 19264 14841 19292
rect 13780 19252 13786 19264
rect 14829 19261 14841 19264
rect 14875 19292 14887 19295
rect 15120 19292 15148 19332
rect 15286 19320 15292 19332
rect 15344 19320 15350 19372
rect 14875 19264 15148 19292
rect 15381 19295 15439 19301
rect 14875 19261 14887 19264
rect 14829 19255 14887 19261
rect 15381 19261 15393 19295
rect 15427 19292 15439 19295
rect 15470 19292 15476 19304
rect 15427 19264 15476 19292
rect 15427 19261 15439 19264
rect 15381 19255 15439 19261
rect 15470 19252 15476 19264
rect 15528 19252 15534 19304
rect 3298 19227 3356 19233
rect 3298 19224 3310 19227
rect 3068 19196 3310 19224
rect 3068 19168 3096 19196
rect 3298 19193 3310 19196
rect 3344 19193 3356 19227
rect 3298 19187 3356 19193
rect 7929 19227 7987 19233
rect 7929 19193 7941 19227
rect 7975 19224 7987 19227
rect 10689 19227 10747 19233
rect 7975 19196 8892 19224
rect 7975 19193 7987 19196
rect 7929 19187 7987 19193
rect 8864 19168 8892 19196
rect 10689 19193 10701 19227
rect 10735 19224 10747 19227
rect 11146 19224 11152 19236
rect 10735 19196 11152 19224
rect 10735 19193 10747 19196
rect 10689 19187 10747 19193
rect 11146 19184 11152 19196
rect 11204 19184 11210 19236
rect 11330 19184 11336 19236
rect 11388 19224 11394 19236
rect 12161 19227 12219 19233
rect 12161 19224 12173 19227
rect 11388 19196 12173 19224
rect 11388 19184 11394 19196
rect 12161 19193 12173 19196
rect 12207 19193 12219 19227
rect 12161 19187 12219 19193
rect 12897 19227 12955 19233
rect 12897 19193 12909 19227
rect 12943 19224 12955 19227
rect 13357 19227 13415 19233
rect 13357 19224 13369 19227
rect 12943 19196 13369 19224
rect 12943 19193 12955 19196
rect 12897 19187 12955 19193
rect 13357 19193 13369 19196
rect 13403 19224 13415 19227
rect 13906 19224 13912 19236
rect 13403 19196 13912 19224
rect 13403 19193 13415 19196
rect 13357 19187 13415 19193
rect 13906 19184 13912 19196
rect 13964 19184 13970 19236
rect 14274 19184 14280 19236
rect 14332 19224 14338 19236
rect 15289 19227 15347 19233
rect 15289 19224 15301 19227
rect 14332 19196 15301 19224
rect 14332 19184 14338 19196
rect 15289 19193 15301 19196
rect 15335 19224 15347 19227
rect 15648 19227 15706 19233
rect 15648 19224 15660 19227
rect 15335 19196 15660 19224
rect 15335 19193 15347 19196
rect 15289 19187 15347 19193
rect 15648 19193 15660 19196
rect 15694 19224 15706 19227
rect 16666 19224 16672 19236
rect 15694 19196 16672 19224
rect 15694 19193 15706 19196
rect 15648 19187 15706 19193
rect 16666 19184 16672 19196
rect 16724 19184 16730 19236
rect 2593 19159 2651 19165
rect 2593 19125 2605 19159
rect 2639 19156 2651 19159
rect 2682 19156 2688 19168
rect 2639 19128 2688 19156
rect 2639 19125 2651 19128
rect 2593 19119 2651 19125
rect 2682 19116 2688 19128
rect 2740 19116 2746 19168
rect 2961 19159 3019 19165
rect 2961 19125 2973 19159
rect 3007 19156 3019 19159
rect 3050 19156 3056 19168
rect 3007 19128 3056 19156
rect 3007 19125 3019 19128
rect 2961 19119 3019 19125
rect 3050 19116 3056 19128
rect 3108 19116 3114 19168
rect 4433 19159 4491 19165
rect 4433 19125 4445 19159
rect 4479 19156 4491 19159
rect 4522 19156 4528 19168
rect 4479 19128 4528 19156
rect 4479 19125 4491 19128
rect 4433 19119 4491 19125
rect 4522 19116 4528 19128
rect 4580 19116 4586 19168
rect 4798 19116 4804 19168
rect 4856 19156 4862 19168
rect 4985 19159 5043 19165
rect 4985 19156 4997 19159
rect 4856 19128 4997 19156
rect 4856 19116 4862 19128
rect 4985 19125 4997 19128
rect 5031 19125 5043 19159
rect 5350 19156 5356 19168
rect 5311 19128 5356 19156
rect 4985 19119 5043 19125
rect 5350 19116 5356 19128
rect 5408 19116 5414 19168
rect 5534 19116 5540 19168
rect 5592 19156 5598 19168
rect 5721 19159 5779 19165
rect 5721 19156 5733 19159
rect 5592 19128 5733 19156
rect 5592 19116 5598 19128
rect 5721 19125 5733 19128
rect 5767 19125 5779 19159
rect 6822 19156 6828 19168
rect 6783 19128 6828 19156
rect 5721 19119 5779 19125
rect 6822 19116 6828 19128
rect 6880 19116 6886 19168
rect 7006 19116 7012 19168
rect 7064 19156 7070 19168
rect 7193 19159 7251 19165
rect 7193 19156 7205 19159
rect 7064 19128 7205 19156
rect 7064 19116 7070 19128
rect 7193 19125 7205 19128
rect 7239 19156 7251 19159
rect 7374 19156 7380 19168
rect 7239 19128 7380 19156
rect 7239 19125 7251 19128
rect 7193 19119 7251 19125
rect 7374 19116 7380 19128
rect 7432 19156 7438 19168
rect 7558 19156 7564 19168
rect 7432 19128 7564 19156
rect 7432 19116 7438 19128
rect 7558 19116 7564 19128
rect 7616 19116 7622 19168
rect 8294 19116 8300 19168
rect 8352 19156 8358 19168
rect 8389 19159 8447 19165
rect 8389 19156 8401 19159
rect 8352 19128 8401 19156
rect 8352 19116 8358 19128
rect 8389 19125 8401 19128
rect 8435 19125 8447 19159
rect 8846 19156 8852 19168
rect 8807 19128 8852 19156
rect 8389 19119 8447 19125
rect 8846 19116 8852 19128
rect 8904 19116 8910 19168
rect 13449 19159 13507 19165
rect 13449 19125 13461 19159
rect 13495 19156 13507 19159
rect 13538 19156 13544 19168
rect 13495 19128 13544 19156
rect 13495 19125 13507 19128
rect 13449 19119 13507 19125
rect 13538 19116 13544 19128
rect 13596 19116 13602 19168
rect 13630 19116 13636 19168
rect 13688 19156 13694 19168
rect 13814 19156 13820 19168
rect 13688 19128 13820 19156
rect 13688 19116 13694 19128
rect 13814 19116 13820 19128
rect 13872 19156 13878 19168
rect 14001 19159 14059 19165
rect 14001 19156 14013 19159
rect 13872 19128 14013 19156
rect 13872 19116 13878 19128
rect 14001 19125 14013 19128
rect 14047 19125 14059 19159
rect 14001 19119 14059 19125
rect 14553 19159 14611 19165
rect 14553 19125 14565 19159
rect 14599 19156 14611 19159
rect 15470 19156 15476 19168
rect 14599 19128 15476 19156
rect 14599 19125 14611 19128
rect 14553 19119 14611 19125
rect 15470 19116 15476 19128
rect 15528 19116 15534 19168
rect 16758 19156 16764 19168
rect 16719 19128 16764 19156
rect 16758 19116 16764 19128
rect 16816 19116 16822 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 1394 18952 1400 18964
rect 1355 18924 1400 18952
rect 1394 18912 1400 18924
rect 1452 18912 1458 18964
rect 2774 18912 2780 18964
rect 2832 18952 2838 18964
rect 2961 18955 3019 18961
rect 2832 18924 2877 18952
rect 2832 18912 2838 18924
rect 2961 18921 2973 18955
rect 3007 18952 3019 18955
rect 4706 18952 4712 18964
rect 3007 18924 4712 18952
rect 3007 18921 3019 18924
rect 2961 18915 3019 18921
rect 4706 18912 4712 18924
rect 4764 18952 4770 18964
rect 5350 18952 5356 18964
rect 4764 18924 5356 18952
rect 4764 18912 4770 18924
rect 5350 18912 5356 18924
rect 5408 18912 5414 18964
rect 6454 18952 6460 18964
rect 5460 18924 6460 18952
rect 3421 18887 3479 18893
rect 3421 18884 3433 18887
rect 1596 18856 3433 18884
rect 1394 18708 1400 18760
rect 1452 18748 1458 18760
rect 1596 18748 1624 18856
rect 3421 18853 3433 18856
rect 3467 18853 3479 18887
rect 3421 18847 3479 18853
rect 4246 18844 4252 18896
rect 4304 18884 4310 18896
rect 4617 18887 4675 18893
rect 4617 18884 4629 18887
rect 4304 18856 4629 18884
rect 4304 18844 4310 18856
rect 4617 18853 4629 18856
rect 4663 18853 4675 18887
rect 4617 18847 4675 18853
rect 5074 18844 5080 18896
rect 5132 18884 5138 18896
rect 5169 18887 5227 18893
rect 5169 18884 5181 18887
rect 5132 18856 5181 18884
rect 5132 18844 5138 18856
rect 5169 18853 5181 18856
rect 5215 18853 5227 18887
rect 5169 18847 5227 18853
rect 1762 18816 1768 18828
rect 1723 18788 1768 18816
rect 1762 18776 1768 18788
rect 1820 18816 1826 18828
rect 3789 18819 3847 18825
rect 3789 18816 3801 18819
rect 1820 18788 3801 18816
rect 1820 18776 1826 18788
rect 3789 18785 3801 18788
rect 3835 18785 3847 18819
rect 3789 18779 3847 18785
rect 4154 18776 4160 18828
rect 4212 18816 4218 18828
rect 4525 18819 4583 18825
rect 4525 18816 4537 18819
rect 4212 18788 4537 18816
rect 4212 18776 4218 18788
rect 4525 18785 4537 18788
rect 4571 18816 4583 18819
rect 5460 18816 5488 18924
rect 6454 18912 6460 18924
rect 6512 18912 6518 18964
rect 7742 18952 7748 18964
rect 7703 18924 7748 18952
rect 7742 18912 7748 18924
rect 7800 18912 7806 18964
rect 8113 18955 8171 18961
rect 8113 18921 8125 18955
rect 8159 18952 8171 18955
rect 8202 18952 8208 18964
rect 8159 18924 8208 18952
rect 8159 18921 8171 18924
rect 8113 18915 8171 18921
rect 8202 18912 8208 18924
rect 8260 18912 8266 18964
rect 8294 18912 8300 18964
rect 8352 18952 8358 18964
rect 8757 18955 8815 18961
rect 8757 18952 8769 18955
rect 8352 18924 8769 18952
rect 8352 18912 8358 18924
rect 8757 18921 8769 18924
rect 8803 18921 8815 18955
rect 9214 18952 9220 18964
rect 9175 18924 9220 18952
rect 8757 18915 8815 18921
rect 9214 18912 9220 18924
rect 9272 18912 9278 18964
rect 9950 18952 9956 18964
rect 9911 18924 9956 18952
rect 9950 18912 9956 18924
rect 10008 18912 10014 18964
rect 10042 18912 10048 18964
rect 10100 18952 10106 18964
rect 10505 18955 10563 18961
rect 10505 18952 10517 18955
rect 10100 18924 10517 18952
rect 10100 18912 10106 18924
rect 10505 18921 10517 18924
rect 10551 18952 10563 18955
rect 11609 18955 11667 18961
rect 11609 18952 11621 18955
rect 10551 18924 11621 18952
rect 10551 18921 10563 18924
rect 10505 18915 10563 18921
rect 11609 18921 11621 18924
rect 11655 18921 11667 18955
rect 13630 18952 13636 18964
rect 13591 18924 13636 18952
rect 11609 18915 11667 18921
rect 13630 18912 13636 18924
rect 13688 18912 13694 18964
rect 14366 18912 14372 18964
rect 14424 18952 14430 18964
rect 14642 18952 14648 18964
rect 14424 18924 14648 18952
rect 14424 18912 14430 18924
rect 14642 18912 14648 18924
rect 14700 18912 14706 18964
rect 16666 18952 16672 18964
rect 16627 18924 16672 18952
rect 16666 18912 16672 18924
rect 16724 18912 16730 18964
rect 5988 18887 6046 18893
rect 5988 18853 6000 18887
rect 6034 18884 6046 18887
rect 6178 18884 6184 18896
rect 6034 18856 6184 18884
rect 6034 18853 6046 18856
rect 5988 18847 6046 18853
rect 6178 18844 6184 18856
rect 6236 18844 6242 18896
rect 10962 18844 10968 18896
rect 11020 18884 11026 18896
rect 11425 18887 11483 18893
rect 11425 18884 11437 18887
rect 11020 18856 11437 18884
rect 11020 18844 11026 18856
rect 11425 18853 11437 18856
rect 11471 18884 11483 18887
rect 12069 18887 12127 18893
rect 12069 18884 12081 18887
rect 11471 18856 12081 18884
rect 11471 18853 11483 18856
rect 11425 18847 11483 18853
rect 12069 18853 12081 18856
rect 12115 18853 12127 18887
rect 12069 18847 12127 18853
rect 12618 18844 12624 18896
rect 12676 18884 12682 18896
rect 18046 18884 18052 18896
rect 12676 18856 18052 18884
rect 12676 18844 12682 18856
rect 18046 18844 18052 18856
rect 18104 18844 18110 18896
rect 4571 18788 5488 18816
rect 5721 18819 5779 18825
rect 4571 18785 4583 18788
rect 4525 18779 4583 18785
rect 5721 18785 5733 18819
rect 5767 18816 5779 18819
rect 6270 18816 6276 18828
rect 5767 18788 6276 18816
rect 5767 18785 5779 18788
rect 5721 18779 5779 18785
rect 6270 18776 6276 18788
rect 6328 18776 6334 18828
rect 8205 18819 8263 18825
rect 8205 18785 8217 18819
rect 8251 18816 8263 18819
rect 8570 18816 8576 18828
rect 8251 18788 8576 18816
rect 8251 18785 8263 18788
rect 8205 18779 8263 18785
rect 8570 18776 8576 18788
rect 8628 18776 8634 18828
rect 10134 18776 10140 18828
rect 10192 18816 10198 18828
rect 10413 18819 10471 18825
rect 10413 18816 10425 18819
rect 10192 18788 10425 18816
rect 10192 18776 10198 18788
rect 10413 18785 10425 18788
rect 10459 18785 10471 18819
rect 10413 18779 10471 18785
rect 11698 18776 11704 18828
rect 11756 18816 11762 18828
rect 11977 18819 12035 18825
rect 11977 18816 11989 18819
rect 11756 18788 11989 18816
rect 11756 18776 11762 18788
rect 11977 18785 11989 18788
rect 12023 18785 12035 18819
rect 11977 18779 12035 18785
rect 13541 18819 13599 18825
rect 13541 18785 13553 18819
rect 13587 18816 13599 18819
rect 13998 18816 14004 18828
rect 13587 18788 14004 18816
rect 13587 18785 13599 18788
rect 13541 18779 13599 18785
rect 13998 18776 14004 18788
rect 14056 18776 14062 18828
rect 14093 18819 14151 18825
rect 14093 18785 14105 18819
rect 14139 18816 14151 18819
rect 14366 18816 14372 18828
rect 14139 18788 14372 18816
rect 14139 18785 14151 18788
rect 14093 18779 14151 18785
rect 14366 18776 14372 18788
rect 14424 18776 14430 18828
rect 15013 18819 15071 18825
rect 15013 18785 15025 18819
rect 15059 18816 15071 18819
rect 15556 18819 15614 18825
rect 15556 18816 15568 18819
rect 15059 18788 15568 18816
rect 15059 18785 15071 18788
rect 15013 18779 15071 18785
rect 15556 18785 15568 18788
rect 15602 18816 15614 18819
rect 15930 18816 15936 18828
rect 15602 18788 15936 18816
rect 15602 18785 15614 18788
rect 15556 18779 15614 18785
rect 15930 18776 15936 18788
rect 15988 18776 15994 18828
rect 1857 18751 1915 18757
rect 1857 18748 1869 18751
rect 1452 18720 1869 18748
rect 1452 18708 1458 18720
rect 1857 18717 1869 18720
rect 1903 18717 1915 18751
rect 1857 18711 1915 18717
rect 2041 18751 2099 18757
rect 2041 18717 2053 18751
rect 2087 18748 2099 18751
rect 4706 18748 4712 18760
rect 2087 18720 2544 18748
rect 4667 18720 4712 18748
rect 2087 18717 2099 18720
rect 2041 18711 2099 18717
rect 2516 18624 2544 18720
rect 4706 18708 4712 18720
rect 4764 18708 4770 18760
rect 10594 18748 10600 18760
rect 10555 18720 10600 18748
rect 10594 18708 10600 18720
rect 10652 18708 10658 18760
rect 12158 18748 12164 18760
rect 12119 18720 12164 18748
rect 12158 18708 12164 18720
rect 12216 18708 12222 18760
rect 14274 18748 14280 18760
rect 14235 18720 14280 18748
rect 14274 18708 14280 18720
rect 14332 18708 14338 18760
rect 15289 18751 15347 18757
rect 15289 18717 15301 18751
rect 15335 18717 15347 18751
rect 15289 18711 15347 18717
rect 4522 18640 4528 18692
rect 4580 18680 4586 18692
rect 4724 18680 4752 18708
rect 8386 18680 8392 18692
rect 4580 18652 4752 18680
rect 8347 18652 8392 18680
rect 4580 18640 4586 18652
rect 8386 18640 8392 18652
rect 8444 18640 8450 18692
rect 2498 18612 2504 18624
rect 2459 18584 2504 18612
rect 2498 18572 2504 18584
rect 2556 18572 2562 18624
rect 4157 18615 4215 18621
rect 4157 18581 4169 18615
rect 4203 18612 4215 18615
rect 5074 18612 5080 18624
rect 4203 18584 5080 18612
rect 4203 18581 4215 18584
rect 4157 18575 4215 18581
rect 5074 18572 5080 18584
rect 5132 18572 5138 18624
rect 5350 18572 5356 18624
rect 5408 18612 5414 18624
rect 5537 18615 5595 18621
rect 5537 18612 5549 18615
rect 5408 18584 5549 18612
rect 5408 18572 5414 18584
rect 5537 18581 5549 18584
rect 5583 18581 5595 18615
rect 5537 18575 5595 18581
rect 7006 18572 7012 18624
rect 7064 18612 7070 18624
rect 7101 18615 7159 18621
rect 7101 18612 7113 18615
rect 7064 18584 7113 18612
rect 7064 18572 7070 18584
rect 7101 18581 7113 18584
rect 7147 18581 7159 18615
rect 7101 18575 7159 18581
rect 10045 18615 10103 18621
rect 10045 18581 10057 18615
rect 10091 18612 10103 18615
rect 10870 18612 10876 18624
rect 10091 18584 10876 18612
rect 10091 18581 10103 18584
rect 10045 18575 10103 18581
rect 10870 18572 10876 18584
rect 10928 18572 10934 18624
rect 11146 18612 11152 18624
rect 11107 18584 11152 18612
rect 11146 18572 11152 18584
rect 11204 18572 11210 18624
rect 12434 18572 12440 18624
rect 12492 18612 12498 18624
rect 12621 18615 12679 18621
rect 12621 18612 12633 18615
rect 12492 18584 12633 18612
rect 12492 18572 12498 18584
rect 12621 18581 12633 18584
rect 12667 18581 12679 18615
rect 12621 18575 12679 18581
rect 13081 18615 13139 18621
rect 13081 18581 13093 18615
rect 13127 18612 13139 18615
rect 13538 18612 13544 18624
rect 13127 18584 13544 18612
rect 13127 18581 13139 18584
rect 13081 18575 13139 18581
rect 13538 18572 13544 18584
rect 13596 18612 13602 18624
rect 13906 18612 13912 18624
rect 13596 18584 13912 18612
rect 13596 18572 13602 18584
rect 13906 18572 13912 18584
rect 13964 18572 13970 18624
rect 15304 18612 15332 18711
rect 15470 18612 15476 18624
rect 15304 18584 15476 18612
rect 15470 18572 15476 18584
rect 15528 18612 15534 18624
rect 16390 18612 16396 18624
rect 15528 18584 16396 18612
rect 15528 18572 15534 18584
rect 16390 18572 16396 18584
rect 16448 18572 16454 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 4154 18408 4160 18420
rect 4115 18380 4160 18408
rect 4154 18368 4160 18380
rect 4212 18368 4218 18420
rect 4246 18368 4252 18420
rect 4304 18408 4310 18420
rect 4525 18411 4583 18417
rect 4525 18408 4537 18411
rect 4304 18380 4537 18408
rect 4304 18368 4310 18380
rect 4525 18377 4537 18380
rect 4571 18377 4583 18411
rect 5166 18408 5172 18420
rect 5127 18380 5172 18408
rect 4525 18371 4583 18377
rect 5166 18368 5172 18380
rect 5224 18368 5230 18420
rect 8202 18368 8208 18420
rect 8260 18408 8266 18420
rect 8481 18411 8539 18417
rect 8481 18408 8493 18411
rect 8260 18380 8493 18408
rect 8260 18368 8266 18380
rect 8481 18377 8493 18380
rect 8527 18408 8539 18411
rect 8662 18408 8668 18420
rect 8527 18380 8668 18408
rect 8527 18377 8539 18380
rect 8481 18371 8539 18377
rect 8662 18368 8668 18380
rect 8720 18368 8726 18420
rect 9585 18411 9643 18417
rect 9585 18377 9597 18411
rect 9631 18408 9643 18411
rect 10042 18408 10048 18420
rect 9631 18380 10048 18408
rect 9631 18377 9643 18380
rect 9585 18371 9643 18377
rect 10042 18368 10048 18380
rect 10100 18368 10106 18420
rect 11882 18408 11888 18420
rect 11795 18380 11888 18408
rect 11882 18368 11888 18380
rect 11940 18408 11946 18420
rect 12158 18408 12164 18420
rect 11940 18380 12164 18408
rect 11940 18368 11946 18380
rect 12158 18368 12164 18380
rect 12216 18368 12222 18420
rect 13998 18368 14004 18420
rect 14056 18408 14062 18420
rect 14921 18411 14979 18417
rect 14921 18408 14933 18411
rect 14056 18380 14933 18408
rect 14056 18368 14062 18380
rect 14921 18377 14933 18380
rect 14967 18377 14979 18411
rect 14921 18371 14979 18377
rect 5442 18300 5448 18352
rect 5500 18340 5506 18352
rect 6270 18340 6276 18352
rect 5500 18312 6276 18340
rect 5500 18300 5506 18312
rect 6270 18300 6276 18312
rect 6328 18300 6334 18352
rect 10686 18300 10692 18352
rect 10744 18340 10750 18352
rect 11238 18340 11244 18352
rect 10744 18312 11244 18340
rect 10744 18300 10750 18312
rect 11238 18300 11244 18312
rect 11296 18300 11302 18352
rect 14274 18300 14280 18352
rect 14332 18340 14338 18352
rect 14369 18343 14427 18349
rect 14369 18340 14381 18343
rect 14332 18312 14381 18340
rect 14332 18300 14338 18312
rect 14369 18309 14381 18312
rect 14415 18309 14427 18343
rect 14734 18340 14740 18352
rect 14695 18312 14740 18340
rect 14369 18303 14427 18309
rect 14734 18300 14740 18312
rect 14792 18340 14798 18352
rect 14792 18312 15424 18340
rect 14792 18300 14798 18312
rect 5077 18275 5135 18281
rect 5077 18241 5089 18275
rect 5123 18272 5135 18275
rect 5721 18275 5779 18281
rect 5721 18272 5733 18275
rect 5123 18244 5733 18272
rect 5123 18241 5135 18244
rect 5077 18235 5135 18241
rect 5721 18241 5733 18244
rect 5767 18272 5779 18275
rect 6549 18275 6607 18281
rect 6549 18272 6561 18275
rect 5767 18244 6561 18272
rect 5767 18241 5779 18244
rect 5721 18235 5779 18241
rect 6549 18241 6561 18244
rect 6595 18272 6607 18275
rect 7006 18272 7012 18284
rect 6595 18244 7012 18272
rect 6595 18241 6607 18244
rect 6549 18235 6607 18241
rect 7006 18232 7012 18244
rect 7064 18272 7070 18284
rect 9674 18272 9680 18284
rect 7064 18244 7236 18272
rect 9635 18244 9680 18272
rect 7064 18232 7070 18244
rect 1486 18164 1492 18216
rect 1544 18204 1550 18216
rect 2041 18207 2099 18213
rect 2041 18204 2053 18207
rect 1544 18176 2053 18204
rect 1544 18164 1550 18176
rect 2041 18173 2053 18176
rect 2087 18204 2099 18207
rect 3142 18204 3148 18216
rect 2087 18176 3148 18204
rect 2087 18173 2099 18176
rect 2041 18167 2099 18173
rect 3142 18164 3148 18176
rect 3200 18164 3206 18216
rect 5534 18164 5540 18216
rect 5592 18204 5598 18216
rect 5629 18207 5687 18213
rect 5629 18204 5641 18207
rect 5592 18176 5641 18204
rect 5592 18164 5598 18176
rect 5629 18173 5641 18176
rect 5675 18173 5687 18207
rect 5629 18167 5687 18173
rect 6270 18164 6276 18216
rect 6328 18204 6334 18216
rect 7101 18207 7159 18213
rect 7101 18204 7113 18207
rect 6328 18176 7113 18204
rect 6328 18164 6334 18176
rect 7101 18173 7113 18176
rect 7147 18173 7159 18207
rect 7208 18204 7236 18244
rect 9674 18232 9680 18244
rect 9732 18232 9738 18284
rect 10594 18232 10600 18284
rect 10652 18272 10658 18284
rect 11333 18275 11391 18281
rect 11333 18272 11345 18275
rect 10652 18244 11345 18272
rect 10652 18232 10658 18244
rect 11333 18241 11345 18244
rect 11379 18272 11391 18275
rect 12158 18272 12164 18284
rect 11379 18244 12164 18272
rect 11379 18241 11391 18244
rect 11333 18235 11391 18241
rect 12158 18232 12164 18244
rect 12216 18272 12222 18284
rect 15396 18281 15424 18312
rect 15381 18275 15439 18281
rect 12216 18244 12572 18272
rect 12216 18232 12222 18244
rect 7357 18207 7415 18213
rect 7357 18204 7369 18207
rect 7208 18176 7369 18204
rect 7101 18167 7159 18173
rect 7357 18173 7369 18176
rect 7403 18173 7415 18207
rect 11146 18204 11152 18216
rect 11107 18176 11152 18204
rect 7357 18167 7415 18173
rect 1949 18139 2007 18145
rect 1949 18105 1961 18139
rect 1995 18136 2007 18139
rect 2308 18139 2366 18145
rect 2308 18136 2320 18139
rect 1995 18108 2320 18136
rect 1995 18105 2007 18108
rect 1949 18099 2007 18105
rect 2308 18105 2320 18108
rect 2354 18136 2366 18139
rect 2682 18136 2688 18148
rect 2354 18108 2688 18136
rect 2354 18105 2366 18108
rect 2308 18099 2366 18105
rect 2682 18096 2688 18108
rect 2740 18096 2746 18148
rect 6914 18136 6920 18148
rect 5552 18108 6920 18136
rect 1854 18028 1860 18080
rect 1912 18068 1918 18080
rect 2958 18068 2964 18080
rect 1912 18040 2964 18068
rect 1912 18028 1918 18040
rect 2958 18028 2964 18040
rect 3016 18028 3022 18080
rect 3050 18028 3056 18080
rect 3108 18068 3114 18080
rect 3421 18071 3479 18077
rect 3421 18068 3433 18071
rect 3108 18040 3433 18068
rect 3108 18028 3114 18040
rect 3421 18037 3433 18040
rect 3467 18037 3479 18071
rect 3421 18031 3479 18037
rect 5258 18028 5264 18080
rect 5316 18068 5322 18080
rect 5552 18077 5580 18108
rect 6914 18096 6920 18108
rect 6972 18096 6978 18148
rect 7116 18136 7144 18167
rect 11146 18164 11152 18176
rect 11204 18164 11210 18216
rect 12434 18204 12440 18216
rect 12395 18176 12440 18204
rect 12434 18164 12440 18176
rect 12492 18164 12498 18216
rect 12544 18204 12572 18244
rect 15381 18241 15393 18275
rect 15427 18241 15439 18275
rect 15381 18235 15439 18241
rect 15565 18275 15623 18281
rect 15565 18241 15577 18275
rect 15611 18272 15623 18275
rect 15930 18272 15936 18284
rect 15611 18244 15936 18272
rect 15611 18241 15623 18244
rect 15565 18235 15623 18241
rect 15930 18232 15936 18244
rect 15988 18232 15994 18284
rect 12693 18207 12751 18213
rect 12693 18204 12705 18207
rect 12544 18176 12705 18204
rect 12693 18173 12705 18176
rect 12739 18173 12751 18207
rect 12693 18167 12751 18173
rect 7834 18136 7840 18148
rect 7116 18108 7840 18136
rect 7834 18096 7840 18108
rect 7892 18096 7898 18148
rect 10229 18139 10287 18145
rect 10229 18105 10241 18139
rect 10275 18136 10287 18139
rect 10594 18136 10600 18148
rect 10275 18108 10600 18136
rect 10275 18105 10287 18108
rect 10229 18099 10287 18105
rect 10594 18096 10600 18108
rect 10652 18096 10658 18148
rect 15102 18096 15108 18148
rect 15160 18136 15166 18148
rect 15289 18139 15347 18145
rect 15289 18136 15301 18139
rect 15160 18108 15301 18136
rect 15160 18096 15166 18108
rect 15289 18105 15301 18108
rect 15335 18136 15347 18139
rect 16485 18139 16543 18145
rect 16485 18136 16497 18139
rect 15335 18108 16497 18136
rect 15335 18105 15347 18108
rect 15289 18099 15347 18105
rect 16485 18105 16497 18108
rect 16531 18105 16543 18139
rect 16485 18099 16543 18105
rect 5537 18071 5595 18077
rect 5537 18068 5549 18071
rect 5316 18040 5549 18068
rect 5316 18028 5322 18040
rect 5537 18037 5549 18040
rect 5583 18037 5595 18071
rect 6178 18068 6184 18080
rect 6139 18040 6184 18068
rect 5537 18031 5595 18037
rect 6178 18028 6184 18040
rect 6236 18028 6242 18080
rect 7006 18028 7012 18080
rect 7064 18068 7070 18080
rect 7282 18068 7288 18080
rect 7064 18040 7288 18068
rect 7064 18028 7070 18040
rect 7282 18028 7288 18040
rect 7340 18028 7346 18080
rect 8570 18028 8576 18080
rect 8628 18068 8634 18080
rect 9125 18071 9183 18077
rect 9125 18068 9137 18071
rect 8628 18040 9137 18068
rect 8628 18028 8634 18040
rect 9125 18037 9137 18040
rect 9171 18068 9183 18071
rect 9950 18068 9956 18080
rect 9171 18040 9956 18068
rect 9171 18037 9183 18040
rect 9125 18031 9183 18037
rect 9950 18028 9956 18040
rect 10008 18028 10014 18080
rect 10778 18068 10784 18080
rect 10739 18040 10784 18068
rect 10778 18028 10784 18040
rect 10836 18028 10842 18080
rect 11054 18028 11060 18080
rect 11112 18068 11118 18080
rect 11241 18071 11299 18077
rect 11241 18068 11253 18071
rect 11112 18040 11253 18068
rect 11112 18028 11118 18040
rect 11241 18037 11253 18040
rect 11287 18037 11299 18071
rect 13814 18068 13820 18080
rect 13775 18040 13820 18068
rect 11241 18031 11299 18037
rect 13814 18028 13820 18040
rect 13872 18028 13878 18080
rect 15930 18068 15936 18080
rect 15891 18040 15936 18068
rect 15930 18028 15936 18040
rect 15988 18028 15994 18080
rect 16390 18068 16396 18080
rect 16351 18040 16396 18068
rect 16390 18028 16396 18040
rect 16448 18028 16454 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 2777 17867 2835 17873
rect 2777 17833 2789 17867
rect 2823 17864 2835 17867
rect 2958 17864 2964 17876
rect 2823 17836 2964 17864
rect 2823 17833 2835 17836
rect 2777 17827 2835 17833
rect 2958 17824 2964 17836
rect 3016 17864 3022 17876
rect 3142 17864 3148 17876
rect 3016 17836 3148 17864
rect 3016 17824 3022 17836
rect 3142 17824 3148 17836
rect 3200 17824 3206 17876
rect 6914 17864 6920 17876
rect 6875 17836 6920 17864
rect 6914 17824 6920 17836
rect 6972 17824 6978 17876
rect 9677 17867 9735 17873
rect 9677 17833 9689 17867
rect 9723 17864 9735 17867
rect 9766 17864 9772 17876
rect 9723 17836 9772 17864
rect 9723 17833 9735 17836
rect 9677 17827 9735 17833
rect 9766 17824 9772 17836
rect 9824 17824 9830 17876
rect 10689 17867 10747 17873
rect 10689 17833 10701 17867
rect 10735 17864 10747 17867
rect 10962 17864 10968 17876
rect 10735 17836 10968 17864
rect 10735 17833 10747 17836
rect 10689 17827 10747 17833
rect 10962 17824 10968 17836
rect 11020 17824 11026 17876
rect 12158 17864 12164 17876
rect 12119 17836 12164 17864
rect 12158 17824 12164 17836
rect 12216 17824 12222 17876
rect 12710 17864 12716 17876
rect 12671 17836 12716 17864
rect 12710 17824 12716 17836
rect 12768 17864 12774 17876
rect 13725 17867 13783 17873
rect 13725 17864 13737 17867
rect 12768 17836 13737 17864
rect 12768 17824 12774 17836
rect 13725 17833 13737 17836
rect 13771 17833 13783 17867
rect 13725 17827 13783 17833
rect 15013 17867 15071 17873
rect 15013 17833 15025 17867
rect 15059 17864 15071 17867
rect 15102 17864 15108 17876
rect 15059 17836 15108 17864
rect 15059 17833 15071 17836
rect 15013 17827 15071 17833
rect 15102 17824 15108 17836
rect 15160 17824 15166 17876
rect 4614 17756 4620 17808
rect 4672 17805 4678 17808
rect 4672 17799 4736 17805
rect 4672 17765 4690 17799
rect 4724 17765 4736 17799
rect 4672 17759 4736 17765
rect 4672 17756 4678 17759
rect 10870 17756 10876 17808
rect 10928 17796 10934 17808
rect 11048 17799 11106 17805
rect 11048 17796 11060 17799
rect 10928 17768 11060 17796
rect 10928 17756 10934 17768
rect 11048 17765 11060 17768
rect 11094 17796 11106 17799
rect 11882 17796 11888 17808
rect 11094 17768 11888 17796
rect 11094 17765 11106 17768
rect 11048 17759 11106 17765
rect 11882 17756 11888 17768
rect 11940 17756 11946 17808
rect 12434 17756 12440 17808
rect 12492 17796 12498 17808
rect 15654 17796 15660 17808
rect 12492 17768 15240 17796
rect 15615 17768 15660 17796
rect 12492 17756 12498 17768
rect 842 17688 848 17740
rect 900 17728 906 17740
rect 2406 17728 2412 17740
rect 900 17700 2412 17728
rect 900 17688 906 17700
rect 2406 17688 2412 17700
rect 2464 17728 2470 17740
rect 2869 17731 2927 17737
rect 2869 17728 2881 17731
rect 2464 17700 2881 17728
rect 2464 17688 2470 17700
rect 2869 17697 2881 17700
rect 2915 17728 2927 17731
rect 2958 17728 2964 17740
rect 2915 17700 2964 17728
rect 2915 17697 2927 17700
rect 2869 17691 2927 17697
rect 2958 17688 2964 17700
rect 3016 17688 3022 17740
rect 4433 17731 4491 17737
rect 4433 17697 4445 17731
rect 4479 17728 4491 17731
rect 5442 17728 5448 17740
rect 4479 17700 5448 17728
rect 4479 17697 4491 17700
rect 4433 17691 4491 17697
rect 5442 17688 5448 17700
rect 5500 17688 5506 17740
rect 7282 17728 7288 17740
rect 7243 17700 7288 17728
rect 7282 17688 7288 17700
rect 7340 17688 7346 17740
rect 11330 17728 11336 17740
rect 10888 17700 11336 17728
rect 1673 17663 1731 17669
rect 1673 17629 1685 17663
rect 1719 17660 1731 17663
rect 1854 17660 1860 17672
rect 1719 17632 1860 17660
rect 1719 17629 1731 17632
rect 1673 17623 1731 17629
rect 1854 17620 1860 17632
rect 1912 17620 1918 17672
rect 3050 17660 3056 17672
rect 3011 17632 3056 17660
rect 3050 17620 3056 17632
rect 3108 17620 3114 17672
rect 7374 17660 7380 17672
rect 7335 17632 7380 17660
rect 7374 17620 7380 17632
rect 7432 17620 7438 17672
rect 7469 17663 7527 17669
rect 7469 17629 7481 17663
rect 7515 17629 7527 17663
rect 8478 17660 8484 17672
rect 8439 17632 8484 17660
rect 7469 17623 7527 17629
rect 2038 17552 2044 17604
rect 2096 17592 2102 17604
rect 3421 17595 3479 17601
rect 3421 17592 3433 17595
rect 2096 17564 3433 17592
rect 2096 17552 2102 17564
rect 3421 17561 3433 17564
rect 3467 17561 3479 17595
rect 3421 17555 3479 17561
rect 5534 17552 5540 17604
rect 5592 17592 5598 17604
rect 6733 17595 6791 17601
rect 6733 17592 6745 17595
rect 5592 17564 6745 17592
rect 5592 17552 5598 17564
rect 6733 17561 6745 17564
rect 6779 17561 6791 17595
rect 7484 17592 7512 17623
rect 8478 17620 8484 17632
rect 8536 17620 8542 17672
rect 10781 17663 10839 17669
rect 10781 17629 10793 17663
rect 10827 17660 10839 17663
rect 10888 17660 10916 17700
rect 11330 17688 11336 17700
rect 11388 17688 11394 17740
rect 12618 17688 12624 17740
rect 12676 17728 12682 17740
rect 13633 17731 13691 17737
rect 13633 17728 13645 17731
rect 12676 17700 13645 17728
rect 12676 17688 12682 17700
rect 13633 17697 13645 17700
rect 13679 17697 13691 17731
rect 13633 17691 13691 17697
rect 13998 17688 14004 17740
rect 14056 17728 14062 17740
rect 14826 17728 14832 17740
rect 14056 17700 14832 17728
rect 14056 17688 14062 17700
rect 14826 17688 14832 17700
rect 14884 17688 14890 17740
rect 15212 17728 15240 17768
rect 15654 17756 15660 17768
rect 15712 17756 15718 17808
rect 16301 17731 16359 17737
rect 16301 17728 16313 17731
rect 15212 17700 16313 17728
rect 16301 17697 16313 17700
rect 16347 17697 16359 17731
rect 16301 17691 16359 17697
rect 17221 17731 17279 17737
rect 17221 17697 17233 17731
rect 17267 17728 17279 17731
rect 17402 17728 17408 17740
rect 17267 17700 17408 17728
rect 17267 17697 17279 17700
rect 17221 17691 17279 17697
rect 17402 17688 17408 17700
rect 17460 17688 17466 17740
rect 13170 17660 13176 17672
rect 10827 17632 10916 17660
rect 13083 17632 13176 17660
rect 10827 17629 10839 17632
rect 10781 17623 10839 17629
rect 6733 17555 6791 17561
rect 7392 17564 7512 17592
rect 1670 17484 1676 17536
rect 1728 17524 1734 17536
rect 1949 17527 2007 17533
rect 1949 17524 1961 17527
rect 1728 17496 1961 17524
rect 1728 17484 1734 17496
rect 1949 17493 1961 17496
rect 1995 17493 2007 17527
rect 1949 17487 2007 17493
rect 2409 17527 2467 17533
rect 2409 17493 2421 17527
rect 2455 17524 2467 17527
rect 3602 17524 3608 17536
rect 2455 17496 3608 17524
rect 2455 17493 2467 17496
rect 2409 17487 2467 17493
rect 3602 17484 3608 17496
rect 3660 17484 3666 17536
rect 3881 17527 3939 17533
rect 3881 17493 3893 17527
rect 3927 17524 3939 17527
rect 4341 17527 4399 17533
rect 4341 17524 4353 17527
rect 3927 17496 4353 17524
rect 3927 17493 3939 17496
rect 3881 17487 3939 17493
rect 4341 17493 4353 17496
rect 4387 17524 4399 17527
rect 4614 17524 4620 17536
rect 4387 17496 4620 17524
rect 4387 17493 4399 17496
rect 4341 17487 4399 17493
rect 4614 17484 4620 17496
rect 4672 17484 4678 17536
rect 5442 17484 5448 17536
rect 5500 17524 5506 17536
rect 5813 17527 5871 17533
rect 5813 17524 5825 17527
rect 5500 17496 5825 17524
rect 5500 17484 5506 17496
rect 5813 17493 5825 17496
rect 5859 17524 5871 17527
rect 6178 17524 6184 17536
rect 5859 17496 6184 17524
rect 5859 17493 5871 17496
rect 5813 17487 5871 17493
rect 6178 17484 6184 17496
rect 6236 17484 6242 17536
rect 6362 17524 6368 17536
rect 6323 17496 6368 17524
rect 6362 17484 6368 17496
rect 6420 17484 6426 17536
rect 6638 17484 6644 17536
rect 6696 17524 6702 17536
rect 7392 17524 7420 17564
rect 8754 17552 8760 17604
rect 8812 17592 8818 17604
rect 9030 17592 9036 17604
rect 8812 17564 9036 17592
rect 8812 17552 8818 17564
rect 9030 17552 9036 17564
rect 9088 17592 9094 17604
rect 9309 17595 9367 17601
rect 9309 17592 9321 17595
rect 9088 17564 9321 17592
rect 9088 17552 9094 17564
rect 9309 17561 9321 17564
rect 9355 17592 9367 17595
rect 10796 17592 10824 17623
rect 13170 17620 13176 17632
rect 13228 17660 13234 17672
rect 13814 17660 13820 17672
rect 13228 17632 13820 17660
rect 13228 17620 13234 17632
rect 13814 17620 13820 17632
rect 13872 17620 13878 17672
rect 15746 17660 15752 17672
rect 15707 17632 15752 17660
rect 15746 17620 15752 17632
rect 15804 17620 15810 17672
rect 15933 17663 15991 17669
rect 15933 17629 15945 17663
rect 15979 17629 15991 17663
rect 15933 17623 15991 17629
rect 9355 17564 10824 17592
rect 13265 17595 13323 17601
rect 9355 17561 9367 17564
rect 9309 17555 9367 17561
rect 13265 17561 13277 17595
rect 13311 17592 13323 17595
rect 13722 17592 13728 17604
rect 13311 17564 13728 17592
rect 13311 17561 13323 17564
rect 13265 17555 13323 17561
rect 13722 17552 13728 17564
rect 13780 17552 13786 17604
rect 14826 17552 14832 17604
rect 14884 17592 14890 17604
rect 15948 17592 15976 17623
rect 16758 17620 16764 17672
rect 16816 17660 16822 17672
rect 17313 17663 17371 17669
rect 17313 17660 17325 17663
rect 16816 17632 17325 17660
rect 16816 17620 16822 17632
rect 17313 17629 17325 17632
rect 17359 17629 17371 17663
rect 17494 17660 17500 17672
rect 17455 17632 17500 17660
rect 17313 17623 17371 17629
rect 17494 17620 17500 17632
rect 17552 17620 17558 17672
rect 17512 17592 17540 17620
rect 14884 17564 17540 17592
rect 14884 17552 14890 17564
rect 6696 17496 7420 17524
rect 6696 17484 6702 17496
rect 7834 17484 7840 17536
rect 7892 17524 7898 17536
rect 8021 17527 8079 17533
rect 8021 17524 8033 17527
rect 7892 17496 8033 17524
rect 7892 17484 7898 17496
rect 8021 17493 8033 17496
rect 8067 17524 8079 17527
rect 8386 17524 8392 17536
rect 8067 17496 8392 17524
rect 8067 17493 8079 17496
rect 8021 17487 8079 17493
rect 8386 17484 8392 17496
rect 8444 17524 8450 17536
rect 8941 17527 8999 17533
rect 8941 17524 8953 17527
rect 8444 17496 8953 17524
rect 8444 17484 8450 17496
rect 8941 17493 8953 17496
rect 8987 17493 8999 17527
rect 8941 17487 8999 17493
rect 9674 17484 9680 17536
rect 9732 17524 9738 17536
rect 10134 17524 10140 17536
rect 9732 17496 10140 17524
rect 9732 17484 9738 17496
rect 10134 17484 10140 17496
rect 10192 17484 10198 17536
rect 14366 17524 14372 17536
rect 14327 17496 14372 17524
rect 14366 17484 14372 17496
rect 14424 17484 14430 17536
rect 15286 17524 15292 17536
rect 15247 17496 15292 17524
rect 15286 17484 15292 17496
rect 15344 17484 15350 17536
rect 16390 17484 16396 17536
rect 16448 17524 16454 17536
rect 16666 17524 16672 17536
rect 16448 17496 16672 17524
rect 16448 17484 16454 17496
rect 16666 17484 16672 17496
rect 16724 17484 16730 17536
rect 16850 17524 16856 17536
rect 16811 17496 16856 17524
rect 16850 17484 16856 17496
rect 16908 17484 16914 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 1397 17323 1455 17329
rect 1397 17289 1409 17323
rect 1443 17320 1455 17323
rect 1762 17320 1768 17332
rect 1443 17292 1768 17320
rect 1443 17289 1455 17292
rect 1397 17283 1455 17289
rect 1762 17280 1768 17292
rect 1820 17280 1826 17332
rect 2406 17320 2412 17332
rect 2367 17292 2412 17320
rect 2406 17280 2412 17292
rect 2464 17280 2470 17332
rect 3050 17280 3056 17332
rect 3108 17320 3114 17332
rect 4157 17323 4215 17329
rect 4157 17320 4169 17323
rect 3108 17292 4169 17320
rect 3108 17280 3114 17292
rect 4157 17289 4169 17292
rect 4203 17289 4215 17323
rect 4157 17283 4215 17289
rect 4709 17323 4767 17329
rect 4709 17289 4721 17323
rect 4755 17320 4767 17323
rect 5534 17320 5540 17332
rect 4755 17292 5540 17320
rect 4755 17289 4767 17292
rect 4709 17283 4767 17289
rect 5534 17280 5540 17292
rect 5592 17280 5598 17332
rect 6825 17323 6883 17329
rect 6825 17289 6837 17323
rect 6871 17320 6883 17323
rect 7374 17320 7380 17332
rect 6871 17292 7380 17320
rect 6871 17289 6883 17292
rect 6825 17283 6883 17289
rect 7374 17280 7380 17292
rect 7432 17320 7438 17332
rect 7837 17323 7895 17329
rect 7837 17320 7849 17323
rect 7432 17292 7849 17320
rect 7432 17280 7438 17292
rect 7837 17289 7849 17292
rect 7883 17289 7895 17323
rect 8662 17320 8668 17332
rect 8623 17292 8668 17320
rect 7837 17283 7895 17289
rect 8662 17280 8668 17292
rect 8720 17280 8726 17332
rect 10137 17323 10195 17329
rect 10137 17289 10149 17323
rect 10183 17320 10195 17323
rect 10870 17320 10876 17332
rect 10183 17292 10876 17320
rect 10183 17289 10195 17292
rect 10137 17283 10195 17289
rect 10870 17280 10876 17292
rect 10928 17280 10934 17332
rect 12526 17280 12532 17332
rect 12584 17320 12590 17332
rect 14461 17323 14519 17329
rect 14461 17320 14473 17323
rect 12584 17292 14473 17320
rect 12584 17280 12590 17292
rect 14461 17289 14473 17292
rect 14507 17320 14519 17323
rect 15746 17320 15752 17332
rect 14507 17292 15752 17320
rect 14507 17289 14519 17292
rect 14461 17283 14519 17289
rect 15746 17280 15752 17292
rect 15804 17280 15810 17332
rect 17402 17320 17408 17332
rect 17363 17292 17408 17320
rect 17402 17280 17408 17292
rect 17460 17280 17466 17332
rect 17494 17280 17500 17332
rect 17552 17320 17558 17332
rect 18233 17323 18291 17329
rect 18233 17320 18245 17323
rect 17552 17292 18245 17320
rect 17552 17280 17558 17292
rect 18233 17289 18245 17292
rect 18279 17289 18291 17323
rect 18233 17283 18291 17289
rect 2869 17255 2927 17261
rect 2869 17221 2881 17255
rect 2915 17252 2927 17255
rect 3142 17252 3148 17264
rect 2915 17224 3148 17252
rect 2915 17221 2927 17224
rect 2869 17215 2927 17221
rect 3142 17212 3148 17224
rect 3200 17212 3206 17264
rect 4614 17252 4620 17264
rect 3804 17224 4620 17252
rect 2038 17184 2044 17196
rect 1999 17156 2044 17184
rect 2038 17144 2044 17156
rect 2096 17144 2102 17196
rect 3804 17193 3832 17224
rect 4614 17212 4620 17224
rect 4672 17252 4678 17264
rect 4672 17224 6132 17252
rect 4672 17212 4678 17224
rect 6104 17196 6132 17224
rect 6178 17212 6184 17264
rect 6236 17252 6242 17264
rect 6638 17252 6644 17264
rect 6236 17224 6644 17252
rect 6236 17212 6242 17224
rect 6638 17212 6644 17224
rect 6696 17212 6702 17264
rect 3789 17187 3847 17193
rect 3789 17153 3801 17187
rect 3835 17153 3847 17187
rect 3789 17147 3847 17153
rect 4890 17144 4896 17196
rect 4948 17184 4954 17196
rect 5261 17187 5319 17193
rect 5261 17184 5273 17187
rect 4948 17156 5273 17184
rect 4948 17144 4954 17156
rect 5261 17153 5273 17156
rect 5307 17184 5319 17187
rect 5442 17184 5448 17196
rect 5307 17156 5448 17184
rect 5307 17153 5319 17156
rect 5261 17147 5319 17153
rect 5442 17144 5448 17156
rect 5500 17144 5506 17196
rect 6086 17144 6092 17196
rect 6144 17184 6150 17196
rect 6273 17187 6331 17193
rect 6273 17184 6285 17187
rect 6144 17156 6285 17184
rect 6144 17144 6150 17156
rect 6273 17153 6285 17156
rect 6319 17184 6331 17187
rect 7377 17187 7435 17193
rect 7377 17184 7389 17187
rect 6319 17156 7389 17184
rect 6319 17153 6331 17156
rect 6273 17147 6331 17153
rect 7377 17153 7389 17156
rect 7423 17153 7435 17187
rect 8680 17184 8708 17280
rect 12253 17187 12311 17193
rect 8680 17156 8892 17184
rect 7377 17147 7435 17153
rect 3602 17116 3608 17128
rect 3515 17088 3608 17116
rect 3602 17076 3608 17088
rect 3660 17116 3666 17128
rect 5721 17119 5779 17125
rect 5721 17116 5733 17119
rect 3660 17088 5733 17116
rect 3660 17076 3666 17088
rect 5721 17085 5733 17088
rect 5767 17085 5779 17119
rect 5721 17079 5779 17085
rect 5994 17076 6000 17128
rect 6052 17116 6058 17128
rect 6546 17116 6552 17128
rect 6052 17088 6552 17116
rect 6052 17076 6058 17088
rect 6546 17076 6552 17088
rect 6604 17076 6610 17128
rect 6914 17076 6920 17128
rect 6972 17116 6978 17128
rect 7285 17119 7343 17125
rect 7285 17116 7297 17119
rect 6972 17088 7297 17116
rect 6972 17076 6978 17088
rect 7285 17085 7297 17088
rect 7331 17116 7343 17119
rect 7834 17116 7840 17128
rect 7331 17088 7840 17116
rect 7331 17085 7343 17088
rect 7285 17079 7343 17085
rect 7834 17076 7840 17088
rect 7892 17076 7898 17128
rect 8754 17116 8760 17128
rect 8715 17088 8760 17116
rect 8754 17076 8760 17088
rect 8812 17076 8818 17128
rect 8864 17116 8892 17156
rect 12253 17153 12265 17187
rect 12299 17184 12311 17187
rect 14921 17187 14979 17193
rect 12299 17156 12664 17184
rect 12299 17153 12311 17156
rect 12253 17147 12311 17153
rect 9013 17119 9071 17125
rect 9013 17116 9025 17119
rect 8864 17088 9025 17116
rect 9013 17085 9025 17088
rect 9059 17116 9071 17119
rect 9582 17116 9588 17128
rect 9059 17088 9588 17116
rect 9059 17085 9071 17088
rect 9013 17079 9071 17085
rect 9582 17076 9588 17088
rect 9640 17076 9646 17128
rect 12434 17076 12440 17128
rect 12492 17116 12498 17128
rect 12529 17119 12587 17125
rect 12529 17116 12541 17119
rect 12492 17088 12541 17116
rect 12492 17076 12498 17088
rect 12529 17085 12541 17088
rect 12575 17085 12587 17119
rect 12636 17116 12664 17156
rect 14921 17153 14933 17187
rect 14967 17184 14979 17187
rect 14967 17156 15148 17184
rect 14967 17153 14979 17156
rect 14921 17147 14979 17153
rect 12796 17119 12854 17125
rect 12796 17116 12808 17119
rect 12636 17088 12808 17116
rect 12529 17079 12587 17085
rect 12796 17085 12808 17088
rect 12842 17116 12854 17119
rect 13170 17116 13176 17128
rect 12842 17088 13176 17116
rect 12842 17085 12854 17088
rect 12796 17079 12854 17085
rect 1670 17008 1676 17060
rect 1728 17048 1734 17060
rect 1765 17051 1823 17057
rect 1765 17048 1777 17051
rect 1728 17020 1777 17048
rect 1728 17008 1734 17020
rect 1765 17017 1777 17020
rect 1811 17017 1823 17051
rect 5169 17051 5227 17057
rect 5169 17048 5181 17051
rect 1765 17011 1823 17017
rect 3160 17020 5181 17048
rect 1854 16980 1860 16992
rect 1815 16952 1860 16980
rect 1854 16940 1860 16952
rect 1912 16940 1918 16992
rect 3160 16989 3188 17020
rect 5169 17017 5181 17020
rect 5215 17048 5227 17051
rect 6362 17048 6368 17060
rect 5215 17020 6368 17048
rect 5215 17017 5227 17020
rect 5169 17011 5227 17017
rect 6362 17008 6368 17020
rect 6420 17008 6426 17060
rect 12544 17048 12572 17079
rect 13170 17076 13176 17088
rect 13228 17076 13234 17128
rect 15010 17116 15016 17128
rect 14971 17088 15016 17116
rect 15010 17076 15016 17088
rect 15068 17076 15074 17128
rect 15120 17116 15148 17156
rect 15562 17116 15568 17128
rect 15120 17088 15568 17116
rect 15562 17076 15568 17088
rect 15620 17076 15626 17128
rect 16758 17076 16764 17128
rect 16816 17116 16822 17128
rect 16945 17119 17003 17125
rect 16945 17116 16957 17119
rect 16816 17088 16957 17116
rect 16816 17076 16822 17088
rect 16945 17085 16957 17088
rect 16991 17085 17003 17119
rect 16945 17079 17003 17085
rect 17678 17076 17684 17128
rect 17736 17116 17742 17128
rect 17736 17088 17781 17116
rect 17736 17076 17742 17088
rect 13078 17048 13084 17060
rect 12544 17020 13084 17048
rect 13078 17008 13084 17020
rect 13136 17008 13142 17060
rect 14734 17008 14740 17060
rect 14792 17048 14798 17060
rect 15258 17051 15316 17057
rect 15258 17048 15270 17051
rect 14792 17020 15270 17048
rect 14792 17008 14798 17020
rect 15258 17017 15270 17020
rect 15304 17017 15316 17051
rect 17696 17048 17724 17076
rect 15258 17011 15316 17017
rect 15396 17020 17724 17048
rect 3145 16983 3203 16989
rect 3145 16949 3157 16983
rect 3191 16949 3203 16983
rect 3510 16980 3516 16992
rect 3471 16952 3516 16980
rect 3145 16943 3203 16949
rect 3510 16940 3516 16952
rect 3568 16940 3574 16992
rect 5074 16980 5080 16992
rect 5035 16952 5080 16980
rect 5074 16940 5080 16952
rect 5132 16940 5138 16992
rect 6454 16940 6460 16992
rect 6512 16980 6518 16992
rect 6549 16983 6607 16989
rect 6549 16980 6561 16983
rect 6512 16952 6561 16980
rect 6512 16940 6518 16952
rect 6549 16949 6561 16952
rect 6595 16980 6607 16983
rect 7193 16983 7251 16989
rect 7193 16980 7205 16983
rect 6595 16952 7205 16980
rect 6595 16949 6607 16952
rect 6549 16943 6607 16949
rect 7193 16949 7205 16952
rect 7239 16949 7251 16983
rect 8294 16980 8300 16992
rect 8255 16952 8300 16980
rect 7193 16943 7251 16949
rect 8294 16940 8300 16952
rect 8352 16940 8358 16992
rect 11241 16983 11299 16989
rect 11241 16949 11253 16983
rect 11287 16980 11299 16983
rect 11514 16980 11520 16992
rect 11287 16952 11520 16980
rect 11287 16949 11299 16952
rect 11241 16943 11299 16949
rect 11514 16940 11520 16952
rect 11572 16940 11578 16992
rect 11698 16980 11704 16992
rect 11659 16952 11704 16980
rect 11698 16940 11704 16952
rect 11756 16940 11762 16992
rect 13538 16940 13544 16992
rect 13596 16980 13602 16992
rect 13906 16980 13912 16992
rect 13596 16952 13912 16980
rect 13596 16940 13602 16952
rect 13906 16940 13912 16952
rect 13964 16940 13970 16992
rect 14274 16940 14280 16992
rect 14332 16980 14338 16992
rect 15396 16980 15424 17020
rect 14332 16952 15424 16980
rect 14332 16940 14338 16952
rect 15562 16940 15568 16992
rect 15620 16980 15626 16992
rect 15930 16980 15936 16992
rect 15620 16952 15936 16980
rect 15620 16940 15626 16952
rect 15930 16940 15936 16952
rect 15988 16980 15994 16992
rect 16393 16983 16451 16989
rect 16393 16980 16405 16983
rect 15988 16952 16405 16980
rect 15988 16940 15994 16952
rect 16393 16949 16405 16952
rect 16439 16949 16451 16983
rect 16393 16943 16451 16949
rect 16666 16940 16672 16992
rect 16724 16980 16730 16992
rect 17497 16983 17555 16989
rect 17497 16980 17509 16983
rect 16724 16952 17509 16980
rect 16724 16940 16730 16952
rect 17497 16949 17509 16952
rect 17543 16980 17555 16983
rect 17862 16980 17868 16992
rect 17543 16952 17868 16980
rect 17543 16949 17555 16952
rect 17497 16943 17555 16949
rect 17862 16940 17868 16952
rect 17920 16940 17926 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 2774 16736 2780 16788
rect 2832 16776 2838 16788
rect 2869 16779 2927 16785
rect 2869 16776 2881 16779
rect 2832 16748 2881 16776
rect 2832 16736 2838 16748
rect 2869 16745 2881 16748
rect 2915 16745 2927 16779
rect 3510 16776 3516 16788
rect 3471 16748 3516 16776
rect 2869 16739 2927 16745
rect 3510 16736 3516 16748
rect 3568 16736 3574 16788
rect 4890 16776 4896 16788
rect 4851 16748 4896 16776
rect 4890 16736 4896 16748
rect 4948 16736 4954 16788
rect 5445 16779 5503 16785
rect 5445 16745 5457 16779
rect 5491 16776 5503 16779
rect 7282 16776 7288 16788
rect 5491 16748 7288 16776
rect 5491 16745 5503 16748
rect 5445 16739 5503 16745
rect 7282 16736 7288 16748
rect 7340 16776 7346 16788
rect 7561 16779 7619 16785
rect 7561 16776 7573 16779
rect 7340 16748 7573 16776
rect 7340 16736 7346 16748
rect 7561 16745 7573 16748
rect 7607 16745 7619 16779
rect 7561 16739 7619 16745
rect 9766 16736 9772 16788
rect 9824 16776 9830 16788
rect 9861 16779 9919 16785
rect 9861 16776 9873 16779
rect 9824 16748 9873 16776
rect 9824 16736 9830 16748
rect 9861 16745 9873 16748
rect 9907 16745 9919 16779
rect 9861 16739 9919 16745
rect 10042 16736 10048 16788
rect 10100 16776 10106 16788
rect 10229 16779 10287 16785
rect 10229 16776 10241 16779
rect 10100 16748 10241 16776
rect 10100 16736 10106 16748
rect 10229 16745 10241 16748
rect 10275 16745 10287 16779
rect 10870 16776 10876 16788
rect 10831 16748 10876 16776
rect 10229 16739 10287 16745
rect 10870 16736 10876 16748
rect 10928 16736 10934 16788
rect 11146 16776 11152 16788
rect 11107 16748 11152 16776
rect 11146 16736 11152 16748
rect 11204 16736 11210 16788
rect 12618 16776 12624 16788
rect 12579 16748 12624 16776
rect 12618 16736 12624 16748
rect 12676 16736 12682 16788
rect 13538 16736 13544 16788
rect 13596 16736 13602 16788
rect 13633 16779 13691 16785
rect 13633 16745 13645 16779
rect 13679 16776 13691 16779
rect 14826 16776 14832 16788
rect 13679 16748 14832 16776
rect 13679 16745 13691 16748
rect 13633 16739 13691 16745
rect 14826 16736 14832 16748
rect 14884 16776 14890 16788
rect 15749 16779 15807 16785
rect 15749 16776 15761 16779
rect 14884 16748 15761 16776
rect 14884 16736 14890 16748
rect 15749 16745 15761 16748
rect 15795 16745 15807 16779
rect 15749 16739 15807 16745
rect 15838 16736 15844 16788
rect 15896 16776 15902 16788
rect 17126 16776 17132 16788
rect 15896 16748 17132 16776
rect 15896 16736 15902 16748
rect 17126 16736 17132 16748
rect 17184 16776 17190 16788
rect 17221 16779 17279 16785
rect 17221 16776 17233 16779
rect 17184 16748 17233 16776
rect 17184 16736 17190 16748
rect 17221 16745 17233 16748
rect 17267 16745 17279 16779
rect 17221 16739 17279 16745
rect 17678 16736 17684 16788
rect 17736 16776 17742 16788
rect 17865 16779 17923 16785
rect 17865 16776 17877 16779
rect 17736 16748 17877 16776
rect 17736 16736 17742 16748
rect 17865 16745 17877 16748
rect 17911 16745 17923 16779
rect 17865 16739 17923 16745
rect 4341 16711 4399 16717
rect 4341 16677 4353 16711
rect 4387 16708 4399 16711
rect 5350 16708 5356 16720
rect 4387 16680 5356 16708
rect 4387 16677 4399 16680
rect 4341 16671 4399 16677
rect 5350 16668 5356 16680
rect 5408 16668 5414 16720
rect 6457 16711 6515 16717
rect 6457 16708 6469 16711
rect 5460 16680 6469 16708
rect 1486 16640 1492 16652
rect 1447 16612 1492 16640
rect 1486 16600 1492 16612
rect 1544 16600 1550 16652
rect 1756 16643 1814 16649
rect 1756 16609 1768 16643
rect 1802 16640 1814 16643
rect 2498 16640 2504 16652
rect 1802 16612 2504 16640
rect 1802 16609 1814 16612
rect 1756 16603 1814 16609
rect 2498 16600 2504 16612
rect 2556 16640 2562 16652
rect 3050 16640 3056 16652
rect 2556 16612 3056 16640
rect 2556 16600 2562 16612
rect 3050 16600 3056 16612
rect 3108 16600 3114 16652
rect 3786 16600 3792 16652
rect 3844 16640 3850 16652
rect 4065 16643 4123 16649
rect 4065 16640 4077 16643
rect 3844 16612 4077 16640
rect 3844 16600 3850 16612
rect 4065 16609 4077 16612
rect 4111 16609 4123 16643
rect 4065 16603 4123 16609
rect 5074 16600 5080 16652
rect 5132 16640 5138 16652
rect 5460 16640 5488 16680
rect 6457 16677 6469 16680
rect 6503 16677 6515 16711
rect 6457 16671 6515 16677
rect 6822 16668 6828 16720
rect 6880 16708 6886 16720
rect 6917 16711 6975 16717
rect 6917 16708 6929 16711
rect 6880 16680 6929 16708
rect 6880 16668 6886 16680
rect 6917 16677 6929 16680
rect 6963 16677 6975 16711
rect 6917 16671 6975 16677
rect 7006 16668 7012 16720
rect 7064 16708 7070 16720
rect 8294 16708 8300 16720
rect 7064 16680 8300 16708
rect 7064 16668 7070 16680
rect 8294 16668 8300 16680
rect 8352 16668 8358 16720
rect 8754 16668 8760 16720
rect 8812 16708 8818 16720
rect 9217 16711 9275 16717
rect 9217 16708 9229 16711
rect 8812 16680 9229 16708
rect 8812 16668 8818 16680
rect 9217 16677 9229 16680
rect 9263 16708 9275 16711
rect 12434 16708 12440 16720
rect 9263 16680 12440 16708
rect 9263 16677 9275 16680
rect 9217 16671 9275 16677
rect 12434 16668 12440 16680
rect 12492 16668 12498 16720
rect 13081 16711 13139 16717
rect 13081 16677 13093 16711
rect 13127 16708 13139 16711
rect 13556 16708 13584 16736
rect 13127 16680 13584 16708
rect 14093 16711 14151 16717
rect 13127 16677 13139 16680
rect 13081 16671 13139 16677
rect 14093 16677 14105 16711
rect 14139 16708 14151 16711
rect 14642 16708 14648 16720
rect 14139 16680 14648 16708
rect 14139 16677 14151 16680
rect 14093 16671 14151 16677
rect 5810 16640 5816 16652
rect 5132 16612 5488 16640
rect 5771 16612 5816 16640
rect 5132 16600 5138 16612
rect 5810 16600 5816 16612
rect 5868 16600 5874 16652
rect 6638 16600 6644 16652
rect 6696 16640 6702 16652
rect 7193 16643 7251 16649
rect 7193 16640 7205 16643
rect 6696 16612 7205 16640
rect 6696 16600 6702 16612
rect 7193 16609 7205 16612
rect 7239 16609 7251 16643
rect 7193 16603 7251 16609
rect 8205 16643 8263 16649
rect 8205 16609 8217 16643
rect 8251 16640 8263 16643
rect 8938 16640 8944 16652
rect 8251 16612 8944 16640
rect 8251 16609 8263 16612
rect 8205 16603 8263 16609
rect 8938 16600 8944 16612
rect 8996 16600 9002 16652
rect 9677 16643 9735 16649
rect 9677 16609 9689 16643
rect 9723 16640 9735 16643
rect 10042 16640 10048 16652
rect 9723 16612 10048 16640
rect 9723 16609 9735 16612
rect 9677 16603 9735 16609
rect 10042 16600 10048 16612
rect 10100 16600 10106 16652
rect 11514 16640 11520 16652
rect 11475 16612 11520 16640
rect 11514 16600 11520 16612
rect 11572 16600 11578 16652
rect 11606 16600 11612 16652
rect 11664 16640 11670 16652
rect 12161 16643 12219 16649
rect 12161 16640 12173 16643
rect 11664 16612 12173 16640
rect 11664 16600 11670 16612
rect 12161 16609 12173 16612
rect 12207 16609 12219 16643
rect 12161 16603 12219 16609
rect 12802 16600 12808 16652
rect 12860 16640 12866 16652
rect 13357 16643 13415 16649
rect 13357 16640 13369 16643
rect 12860 16612 13369 16640
rect 12860 16600 12866 16612
rect 13357 16609 13369 16612
rect 13403 16640 13415 16643
rect 13449 16643 13507 16649
rect 13449 16640 13461 16643
rect 13403 16612 13461 16640
rect 13403 16609 13415 16612
rect 13357 16603 13415 16609
rect 13449 16609 13461 16612
rect 13495 16609 13507 16643
rect 13449 16603 13507 16609
rect 13538 16600 13544 16652
rect 13596 16640 13602 16652
rect 13998 16640 14004 16652
rect 13596 16612 14004 16640
rect 13596 16600 13602 16612
rect 13998 16600 14004 16612
rect 14056 16600 14062 16652
rect 5905 16575 5963 16581
rect 5905 16541 5917 16575
rect 5951 16541 5963 16575
rect 6086 16572 6092 16584
rect 6047 16544 6092 16572
rect 5905 16535 5963 16541
rect 5920 16504 5948 16535
rect 6086 16532 6092 16544
rect 6144 16532 6150 16584
rect 8478 16572 8484 16584
rect 8391 16544 8484 16572
rect 8478 16532 8484 16544
rect 8536 16572 8542 16584
rect 9766 16572 9772 16584
rect 8536 16544 9772 16572
rect 8536 16532 8542 16544
rect 9766 16532 9772 16544
rect 9824 16532 9830 16584
rect 11793 16575 11851 16581
rect 11793 16541 11805 16575
rect 11839 16572 11851 16575
rect 11882 16572 11888 16584
rect 11839 16544 11888 16572
rect 11839 16541 11851 16544
rect 11793 16535 11851 16541
rect 11882 16532 11888 16544
rect 11940 16532 11946 16584
rect 13170 16532 13176 16584
rect 13228 16572 13234 16584
rect 14108 16572 14136 16671
rect 14642 16668 14648 16680
rect 14700 16668 14706 16720
rect 14737 16711 14795 16717
rect 14737 16677 14749 16711
rect 14783 16708 14795 16711
rect 14918 16708 14924 16720
rect 14783 16680 14924 16708
rect 14783 16677 14795 16680
rect 14737 16671 14795 16677
rect 14918 16668 14924 16680
rect 14976 16668 14982 16720
rect 15286 16668 15292 16720
rect 15344 16708 15350 16720
rect 15657 16711 15715 16717
rect 15657 16708 15669 16711
rect 15344 16680 15669 16708
rect 15344 16668 15350 16680
rect 15657 16677 15669 16680
rect 15703 16677 15715 16711
rect 15657 16671 15715 16677
rect 14366 16600 14372 16652
rect 14424 16640 14430 16652
rect 14424 16612 15332 16640
rect 14424 16600 14430 16612
rect 13228 16544 14136 16572
rect 14277 16575 14335 16581
rect 13228 16532 13234 16544
rect 14277 16541 14289 16575
rect 14323 16572 14335 16575
rect 14323 16544 14780 16572
rect 14323 16541 14335 16544
rect 14277 16535 14335 16541
rect 6270 16504 6276 16516
rect 5920 16476 6276 16504
rect 6270 16464 6276 16476
rect 6328 16464 6334 16516
rect 14752 16448 14780 16544
rect 15304 16513 15332 16612
rect 15562 16532 15568 16584
rect 15620 16572 15626 16584
rect 15841 16575 15899 16581
rect 15841 16572 15853 16575
rect 15620 16544 15853 16572
rect 15620 16532 15626 16544
rect 15841 16541 15853 16544
rect 15887 16541 15899 16575
rect 17310 16572 17316 16584
rect 17271 16544 17316 16572
rect 15841 16535 15899 16541
rect 17310 16532 17316 16544
rect 17368 16532 17374 16584
rect 17494 16572 17500 16584
rect 17455 16544 17500 16572
rect 17494 16532 17500 16544
rect 17552 16532 17558 16584
rect 15289 16507 15347 16513
rect 15289 16473 15301 16507
rect 15335 16473 15347 16507
rect 15289 16467 15347 16473
rect 3050 16396 3056 16448
rect 3108 16436 3114 16448
rect 3789 16439 3847 16445
rect 3789 16436 3801 16439
rect 3108 16408 3801 16436
rect 3108 16396 3114 16408
rect 3789 16405 3801 16408
rect 3835 16405 3847 16439
rect 3789 16399 3847 16405
rect 5261 16439 5319 16445
rect 5261 16405 5273 16439
rect 5307 16436 5319 16439
rect 6454 16436 6460 16448
rect 5307 16408 6460 16436
rect 5307 16405 5319 16408
rect 5261 16399 5319 16405
rect 6454 16396 6460 16408
rect 6512 16396 6518 16448
rect 7834 16436 7840 16448
rect 7795 16408 7840 16436
rect 7834 16396 7840 16408
rect 7892 16396 7898 16448
rect 13078 16396 13084 16448
rect 13136 16436 13142 16448
rect 13173 16439 13231 16445
rect 13173 16436 13185 16439
rect 13136 16408 13185 16436
rect 13136 16396 13142 16408
rect 13173 16405 13185 16408
rect 13219 16405 13231 16439
rect 13173 16399 13231 16405
rect 13449 16439 13507 16445
rect 13449 16405 13461 16439
rect 13495 16436 13507 16439
rect 14274 16436 14280 16448
rect 13495 16408 14280 16436
rect 13495 16405 13507 16408
rect 13449 16399 13507 16405
rect 14274 16396 14280 16408
rect 14332 16396 14338 16448
rect 14734 16396 14740 16448
rect 14792 16436 14798 16448
rect 15013 16439 15071 16445
rect 15013 16436 15025 16439
rect 14792 16408 15025 16436
rect 14792 16396 14798 16408
rect 15013 16405 15025 16408
rect 15059 16405 15071 16439
rect 16482 16436 16488 16448
rect 16443 16408 16488 16436
rect 15013 16399 15071 16405
rect 16482 16396 16488 16408
rect 16540 16396 16546 16448
rect 16853 16439 16911 16445
rect 16853 16405 16865 16439
rect 16899 16436 16911 16439
rect 16942 16436 16948 16448
rect 16899 16408 16948 16436
rect 16899 16405 16911 16408
rect 16853 16399 16911 16405
rect 16942 16396 16948 16408
rect 17000 16396 17006 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 4614 16232 4620 16244
rect 4575 16204 4620 16232
rect 4614 16192 4620 16204
rect 4672 16192 4678 16244
rect 7006 16232 7012 16244
rect 6967 16204 7012 16232
rect 7006 16192 7012 16204
rect 7064 16192 7070 16244
rect 7558 16192 7564 16244
rect 7616 16232 7622 16244
rect 8021 16235 8079 16241
rect 8021 16232 8033 16235
rect 7616 16204 8033 16232
rect 7616 16192 7622 16204
rect 8021 16201 8033 16204
rect 8067 16232 8079 16235
rect 8297 16235 8355 16241
rect 8297 16232 8309 16235
rect 8067 16204 8309 16232
rect 8067 16201 8079 16204
rect 8021 16195 8079 16201
rect 8297 16201 8309 16204
rect 8343 16201 8355 16235
rect 8297 16195 8355 16201
rect 9677 16235 9735 16241
rect 9677 16201 9689 16235
rect 9723 16232 9735 16235
rect 9766 16232 9772 16244
rect 9723 16204 9772 16232
rect 9723 16201 9735 16204
rect 9677 16195 9735 16201
rect 9766 16192 9772 16204
rect 9824 16192 9830 16244
rect 10781 16235 10839 16241
rect 10781 16201 10793 16235
rect 10827 16232 10839 16235
rect 10962 16232 10968 16244
rect 10827 16204 10968 16232
rect 10827 16201 10839 16204
rect 10781 16195 10839 16201
rect 10962 16192 10968 16204
rect 11020 16192 11026 16244
rect 11514 16192 11520 16244
rect 11572 16232 11578 16244
rect 11793 16235 11851 16241
rect 11793 16232 11805 16235
rect 11572 16204 11805 16232
rect 11572 16192 11578 16204
rect 11793 16201 11805 16204
rect 11839 16201 11851 16235
rect 13170 16232 13176 16244
rect 13131 16204 13176 16232
rect 11793 16195 11851 16201
rect 13170 16192 13176 16204
rect 13228 16192 13234 16244
rect 13630 16232 13636 16244
rect 13591 16204 13636 16232
rect 13630 16192 13636 16204
rect 13688 16192 13694 16244
rect 16758 16232 16764 16244
rect 13832 16204 16764 16232
rect 3605 16167 3663 16173
rect 3605 16133 3617 16167
rect 3651 16164 3663 16167
rect 4062 16164 4068 16176
rect 3651 16136 4068 16164
rect 3651 16133 3663 16136
rect 3605 16127 3663 16133
rect 4062 16124 4068 16136
rect 4120 16124 4126 16176
rect 11146 16164 11152 16176
rect 10796 16136 11152 16164
rect 10796 16108 10824 16136
rect 11146 16124 11152 16136
rect 11204 16164 11210 16176
rect 11204 16136 11376 16164
rect 11204 16124 11210 16136
rect 1762 16056 1768 16108
rect 1820 16096 1826 16108
rect 2593 16099 2651 16105
rect 2593 16096 2605 16099
rect 1820 16068 2605 16096
rect 1820 16056 1826 16068
rect 2593 16065 2605 16068
rect 2639 16096 2651 16099
rect 3145 16099 3203 16105
rect 3145 16096 3157 16099
rect 2639 16068 3157 16096
rect 2639 16065 2651 16068
rect 2593 16059 2651 16065
rect 3145 16065 3157 16068
rect 3191 16096 3203 16099
rect 4246 16096 4252 16108
rect 3191 16068 4252 16096
rect 3191 16065 3203 16068
rect 3145 16059 3203 16065
rect 4246 16056 4252 16068
rect 4304 16056 4310 16108
rect 5813 16099 5871 16105
rect 5813 16065 5825 16099
rect 5859 16096 5871 16099
rect 6454 16096 6460 16108
rect 5859 16068 6460 16096
rect 5859 16065 5871 16068
rect 5813 16059 5871 16065
rect 6454 16056 6460 16068
rect 6512 16056 6518 16108
rect 7558 16096 7564 16108
rect 7519 16068 7564 16096
rect 7558 16056 7564 16068
rect 7616 16056 7622 16108
rect 9214 16096 9220 16108
rect 9175 16068 9220 16096
rect 9214 16056 9220 16068
rect 9272 16056 9278 16108
rect 10689 16099 10747 16105
rect 10689 16065 10701 16099
rect 10735 16096 10747 16099
rect 10778 16096 10784 16108
rect 10735 16068 10784 16096
rect 10735 16065 10747 16068
rect 10689 16059 10747 16065
rect 10778 16056 10784 16068
rect 10836 16056 10842 16108
rect 11238 16096 11244 16108
rect 11199 16068 11244 16096
rect 11238 16056 11244 16068
rect 11296 16056 11302 16108
rect 11348 16105 11376 16136
rect 12618 16124 12624 16176
rect 12676 16164 12682 16176
rect 12713 16167 12771 16173
rect 12713 16164 12725 16167
rect 12676 16136 12725 16164
rect 12676 16124 12682 16136
rect 12713 16133 12725 16136
rect 12759 16133 12771 16167
rect 12713 16127 12771 16133
rect 11333 16099 11391 16105
rect 11333 16065 11345 16099
rect 11379 16065 11391 16099
rect 11333 16059 11391 16065
rect 2406 16028 2412 16040
rect 2367 16000 2412 16028
rect 2406 15988 2412 16000
rect 2464 16028 2470 16040
rect 3602 16028 3608 16040
rect 2464 16000 3608 16028
rect 2464 15988 2470 16000
rect 3602 15988 3608 16000
rect 3660 15988 3666 16040
rect 4065 16031 4123 16037
rect 4065 15997 4077 16031
rect 4111 16028 4123 16031
rect 4154 16028 4160 16040
rect 4111 16000 4160 16028
rect 4111 15997 4123 16000
rect 4065 15991 4123 15997
rect 4154 15988 4160 16000
rect 4212 15988 4218 16040
rect 6089 16031 6147 16037
rect 6089 15997 6101 16031
rect 6135 16028 6147 16031
rect 8389 16031 8447 16037
rect 8389 16028 8401 16031
rect 6135 16000 8401 16028
rect 6135 15997 6147 16000
rect 6089 15991 6147 15997
rect 8389 15997 8401 16000
rect 8435 16028 8447 16031
rect 9033 16031 9091 16037
rect 9033 16028 9045 16031
rect 8435 16000 9045 16028
rect 8435 15997 8447 16000
rect 8389 15991 8447 15997
rect 9033 15997 9045 16000
rect 9079 15997 9091 16031
rect 12728 16028 12756 16127
rect 13832 16028 13860 16204
rect 16758 16192 16764 16204
rect 16816 16192 16822 16244
rect 17126 16232 17132 16244
rect 17087 16204 17132 16232
rect 17126 16192 17132 16204
rect 17184 16192 17190 16244
rect 13906 16056 13912 16108
rect 13964 16096 13970 16108
rect 14277 16099 14335 16105
rect 14277 16096 14289 16099
rect 13964 16068 14289 16096
rect 13964 16056 13970 16068
rect 14277 16065 14289 16068
rect 14323 16096 14335 16099
rect 14323 16068 14504 16096
rect 14323 16065 14335 16068
rect 14277 16059 14335 16065
rect 14001 16031 14059 16037
rect 14001 16028 14013 16031
rect 12728 16000 14013 16028
rect 9033 15991 9091 15997
rect 14001 15997 14013 16000
rect 14047 15997 14059 16031
rect 14001 15991 14059 15997
rect 14090 15988 14096 16040
rect 14148 16028 14154 16040
rect 14148 16000 14193 16028
rect 14148 15988 14154 16000
rect 1949 15963 2007 15969
rect 1949 15929 1961 15963
rect 1995 15960 2007 15963
rect 2314 15960 2320 15972
rect 1995 15932 2320 15960
rect 1995 15929 2007 15932
rect 1949 15923 2007 15929
rect 2314 15920 2320 15932
rect 2372 15960 2378 15972
rect 2498 15960 2504 15972
rect 2372 15932 2504 15960
rect 2372 15920 2378 15932
rect 2498 15920 2504 15932
rect 2556 15920 2562 15972
rect 4430 15920 4436 15972
rect 4488 15960 4494 15972
rect 4890 15960 4896 15972
rect 4488 15932 4896 15960
rect 4488 15920 4494 15932
rect 4890 15920 4896 15932
rect 4948 15920 4954 15972
rect 5629 15963 5687 15969
rect 5629 15960 5641 15963
rect 5000 15932 5641 15960
rect 2038 15892 2044 15904
rect 1999 15864 2044 15892
rect 2038 15852 2044 15864
rect 2096 15852 2102 15904
rect 3513 15895 3571 15901
rect 3513 15861 3525 15895
rect 3559 15892 3571 15895
rect 3878 15892 3884 15904
rect 3559 15864 3884 15892
rect 3559 15861 3571 15864
rect 3513 15855 3571 15861
rect 3878 15852 3884 15864
rect 3936 15892 3942 15904
rect 3973 15895 4031 15901
rect 3973 15892 3985 15895
rect 3936 15864 3985 15892
rect 3936 15852 3942 15864
rect 3973 15861 3985 15864
rect 4019 15861 4031 15895
rect 3973 15855 4031 15861
rect 4706 15852 4712 15904
rect 4764 15892 4770 15904
rect 5000 15901 5028 15932
rect 5629 15929 5641 15932
rect 5675 15960 5687 15963
rect 6549 15963 6607 15969
rect 6549 15960 6561 15963
rect 5675 15932 6561 15960
rect 5675 15929 5687 15932
rect 5629 15923 5687 15929
rect 6549 15929 6561 15932
rect 6595 15960 6607 15963
rect 7469 15963 7527 15969
rect 7469 15960 7481 15963
rect 6595 15932 7481 15960
rect 6595 15929 6607 15932
rect 6549 15923 6607 15929
rect 7469 15929 7481 15932
rect 7515 15929 7527 15963
rect 7469 15923 7527 15929
rect 8297 15963 8355 15969
rect 8297 15929 8309 15963
rect 8343 15960 8355 15963
rect 8941 15963 8999 15969
rect 8941 15960 8953 15963
rect 8343 15932 8953 15960
rect 8343 15929 8355 15932
rect 8297 15923 8355 15929
rect 8941 15929 8953 15932
rect 8987 15929 8999 15963
rect 8941 15923 8999 15929
rect 11514 15920 11520 15972
rect 11572 15960 11578 15972
rect 13449 15963 13507 15969
rect 13449 15960 13461 15963
rect 11572 15932 13461 15960
rect 11572 15920 11578 15932
rect 13449 15929 13461 15932
rect 13495 15960 13507 15963
rect 13538 15960 13544 15972
rect 13495 15932 13544 15960
rect 13495 15929 13507 15932
rect 13449 15923 13507 15929
rect 13538 15920 13544 15932
rect 13596 15920 13602 15972
rect 14476 15960 14504 16068
rect 15197 16031 15255 16037
rect 15197 15997 15209 16031
rect 15243 16028 15255 16031
rect 16390 16028 16396 16040
rect 15243 16000 16396 16028
rect 15243 15997 15255 16000
rect 15197 15991 15255 15997
rect 16390 15988 16396 16000
rect 16448 15988 16454 16040
rect 15464 15963 15522 15969
rect 15464 15960 15476 15963
rect 14476 15932 15476 15960
rect 15464 15929 15476 15932
rect 15510 15960 15522 15963
rect 15838 15960 15844 15972
rect 15510 15932 15844 15960
rect 15510 15929 15522 15932
rect 15464 15923 15522 15929
rect 15838 15920 15844 15932
rect 15896 15920 15902 15972
rect 17494 15960 17500 15972
rect 16592 15932 17500 15960
rect 4985 15895 5043 15901
rect 4985 15892 4997 15895
rect 4764 15864 4997 15892
rect 4764 15852 4770 15864
rect 4985 15861 4997 15864
rect 5031 15861 5043 15895
rect 5166 15892 5172 15904
rect 5127 15864 5172 15892
rect 4985 15855 5043 15861
rect 5166 15852 5172 15864
rect 5224 15852 5230 15904
rect 5350 15852 5356 15904
rect 5408 15892 5414 15904
rect 5537 15895 5595 15901
rect 5537 15892 5549 15895
rect 5408 15864 5549 15892
rect 5408 15852 5414 15864
rect 5537 15861 5549 15864
rect 5583 15892 5595 15895
rect 6089 15895 6147 15901
rect 6089 15892 6101 15895
rect 5583 15864 6101 15892
rect 5583 15861 5595 15864
rect 5537 15855 5595 15861
rect 6089 15861 6101 15864
rect 6135 15861 6147 15895
rect 6270 15892 6276 15904
rect 6183 15864 6276 15892
rect 6089 15855 6147 15861
rect 6270 15852 6276 15864
rect 6328 15892 6334 15904
rect 6730 15892 6736 15904
rect 6328 15864 6736 15892
rect 6328 15852 6334 15864
rect 6730 15852 6736 15864
rect 6788 15852 6794 15904
rect 6914 15852 6920 15904
rect 6972 15892 6978 15904
rect 7377 15895 7435 15901
rect 7377 15892 7389 15895
rect 6972 15864 7389 15892
rect 6972 15852 6978 15864
rect 7377 15861 7389 15864
rect 7423 15861 7435 15895
rect 7377 15855 7435 15861
rect 8573 15895 8631 15901
rect 8573 15861 8585 15895
rect 8619 15892 8631 15895
rect 9122 15892 9128 15904
rect 8619 15864 9128 15892
rect 8619 15861 8631 15864
rect 8573 15855 8631 15861
rect 9122 15852 9128 15864
rect 9180 15852 9186 15904
rect 9766 15852 9772 15904
rect 9824 15892 9830 15904
rect 9953 15895 10011 15901
rect 9953 15892 9965 15895
rect 9824 15864 9965 15892
rect 9824 15852 9830 15864
rect 9953 15861 9965 15864
rect 9999 15892 10011 15895
rect 10042 15892 10048 15904
rect 9999 15864 10048 15892
rect 9999 15861 10011 15864
rect 9953 15855 10011 15861
rect 10042 15852 10048 15864
rect 10100 15852 10106 15904
rect 11149 15895 11207 15901
rect 11149 15861 11161 15895
rect 11195 15892 11207 15895
rect 12161 15895 12219 15901
rect 12161 15892 12173 15895
rect 11195 15864 12173 15892
rect 11195 15861 11207 15864
rect 11149 15855 11207 15861
rect 12161 15861 12173 15864
rect 12207 15892 12219 15895
rect 12618 15892 12624 15904
rect 12207 15864 12624 15892
rect 12207 15861 12219 15864
rect 12161 15855 12219 15861
rect 12618 15852 12624 15864
rect 12676 15852 12682 15904
rect 14734 15892 14740 15904
rect 14695 15864 14740 15892
rect 14734 15852 14740 15864
rect 14792 15852 14798 15904
rect 15105 15895 15163 15901
rect 15105 15861 15117 15895
rect 15151 15892 15163 15895
rect 15286 15892 15292 15904
rect 15151 15864 15292 15892
rect 15151 15861 15163 15864
rect 15105 15855 15163 15861
rect 15286 15852 15292 15864
rect 15344 15852 15350 15904
rect 16592 15901 16620 15932
rect 17494 15920 17500 15932
rect 17552 15960 17558 15972
rect 17552 15932 17632 15960
rect 17552 15920 17558 15932
rect 17604 15901 17632 15932
rect 16577 15895 16635 15901
rect 16577 15861 16589 15895
rect 16623 15861 16635 15895
rect 16577 15855 16635 15861
rect 17589 15895 17647 15901
rect 17589 15861 17601 15895
rect 17635 15892 17647 15895
rect 17862 15892 17868 15904
rect 17635 15864 17868 15892
rect 17635 15861 17647 15864
rect 17589 15855 17647 15861
rect 17862 15852 17868 15864
rect 17920 15852 17926 15904
rect 17954 15852 17960 15904
rect 18012 15892 18018 15904
rect 18325 15895 18383 15901
rect 18325 15892 18337 15895
rect 18012 15864 18337 15892
rect 18012 15852 18018 15864
rect 18325 15861 18337 15864
rect 18371 15892 18383 15895
rect 18690 15892 18696 15904
rect 18371 15864 18696 15892
rect 18371 15861 18383 15864
rect 18325 15855 18383 15861
rect 18690 15852 18696 15864
rect 18748 15852 18754 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1762 15688 1768 15700
rect 1723 15660 1768 15688
rect 1762 15648 1768 15660
rect 1820 15648 1826 15700
rect 2133 15691 2191 15697
rect 2133 15657 2145 15691
rect 2179 15688 2191 15691
rect 2406 15688 2412 15700
rect 2179 15660 2412 15688
rect 2179 15657 2191 15660
rect 2133 15651 2191 15657
rect 2406 15648 2412 15660
rect 2464 15648 2470 15700
rect 3697 15691 3755 15697
rect 3697 15657 3709 15691
rect 3743 15688 3755 15691
rect 4154 15688 4160 15700
rect 3743 15660 4160 15688
rect 3743 15657 3755 15660
rect 3697 15651 3755 15657
rect 4154 15648 4160 15660
rect 4212 15648 4218 15700
rect 4430 15688 4436 15700
rect 4343 15660 4436 15688
rect 4430 15648 4436 15660
rect 4488 15688 4494 15700
rect 5442 15688 5448 15700
rect 4488 15660 5448 15688
rect 4488 15648 4494 15660
rect 5442 15648 5448 15660
rect 5500 15648 5506 15700
rect 5629 15691 5687 15697
rect 5629 15657 5641 15691
rect 5675 15688 5687 15691
rect 5994 15688 6000 15700
rect 5675 15660 6000 15688
rect 5675 15657 5687 15660
rect 5629 15651 5687 15657
rect 5994 15648 6000 15660
rect 6052 15648 6058 15700
rect 6914 15648 6920 15700
rect 6972 15688 6978 15700
rect 7193 15691 7251 15697
rect 7193 15688 7205 15691
rect 6972 15660 7205 15688
rect 6972 15648 6978 15660
rect 7193 15657 7205 15660
rect 7239 15657 7251 15691
rect 7742 15688 7748 15700
rect 7703 15660 7748 15688
rect 7193 15651 7251 15657
rect 7742 15648 7748 15660
rect 7800 15648 7806 15700
rect 7834 15648 7840 15700
rect 7892 15688 7898 15700
rect 8205 15691 8263 15697
rect 8205 15688 8217 15691
rect 7892 15660 8217 15688
rect 7892 15648 7898 15660
rect 8205 15657 8217 15660
rect 8251 15688 8263 15691
rect 9125 15691 9183 15697
rect 9125 15688 9137 15691
rect 8251 15660 9137 15688
rect 8251 15657 8263 15660
rect 8205 15651 8263 15657
rect 9125 15657 9137 15660
rect 9171 15657 9183 15691
rect 9674 15688 9680 15700
rect 9635 15660 9680 15688
rect 9125 15651 9183 15657
rect 9674 15648 9680 15660
rect 9732 15648 9738 15700
rect 10137 15691 10195 15697
rect 10137 15657 10149 15691
rect 10183 15688 10195 15691
rect 10778 15688 10784 15700
rect 10183 15660 10784 15688
rect 10183 15657 10195 15660
rect 10137 15651 10195 15657
rect 10778 15648 10784 15660
rect 10836 15648 10842 15700
rect 11146 15688 11152 15700
rect 11107 15660 11152 15688
rect 11146 15648 11152 15660
rect 11204 15648 11210 15700
rect 11425 15691 11483 15697
rect 11425 15657 11437 15691
rect 11471 15688 11483 15691
rect 11606 15688 11612 15700
rect 11471 15660 11612 15688
rect 11471 15657 11483 15660
rect 11425 15651 11483 15657
rect 11606 15648 11612 15660
rect 11664 15648 11670 15700
rect 12434 15688 12440 15700
rect 12395 15660 12440 15688
rect 12434 15648 12440 15660
rect 12492 15648 12498 15700
rect 12618 15648 12624 15700
rect 12676 15688 12682 15700
rect 12989 15691 13047 15697
rect 12989 15688 13001 15691
rect 12676 15660 13001 15688
rect 12676 15648 12682 15660
rect 12989 15657 13001 15660
rect 13035 15657 13047 15691
rect 12989 15651 13047 15657
rect 13170 15648 13176 15700
rect 13228 15688 13234 15700
rect 13446 15688 13452 15700
rect 13228 15660 13452 15688
rect 13228 15648 13234 15660
rect 13446 15648 13452 15660
rect 13504 15648 13510 15700
rect 14090 15688 14096 15700
rect 14051 15660 14096 15688
rect 14090 15648 14096 15660
rect 14148 15648 14154 15700
rect 14826 15648 14832 15700
rect 14884 15688 14890 15700
rect 15013 15691 15071 15697
rect 15013 15688 15025 15691
rect 14884 15660 15025 15688
rect 14884 15648 14890 15660
rect 15013 15657 15025 15660
rect 15059 15657 15071 15691
rect 15562 15688 15568 15700
rect 15523 15660 15568 15688
rect 15013 15651 15071 15657
rect 15562 15648 15568 15660
rect 15620 15648 15626 15700
rect 15838 15688 15844 15700
rect 15799 15660 15844 15688
rect 15838 15648 15844 15660
rect 15896 15648 15902 15700
rect 16393 15691 16451 15697
rect 16393 15657 16405 15691
rect 16439 15688 16451 15691
rect 16853 15691 16911 15697
rect 16853 15688 16865 15691
rect 16439 15660 16865 15688
rect 16439 15657 16451 15660
rect 16393 15651 16451 15657
rect 16853 15657 16865 15660
rect 16899 15688 16911 15691
rect 18049 15691 18107 15697
rect 18049 15688 18061 15691
rect 16899 15660 18061 15688
rect 16899 15657 16911 15660
rect 16853 15651 16911 15657
rect 18049 15657 18061 15660
rect 18095 15657 18107 15691
rect 18506 15688 18512 15700
rect 18467 15660 18512 15688
rect 18049 15651 18107 15657
rect 18506 15648 18512 15660
rect 18564 15648 18570 15700
rect 3142 15580 3148 15632
rect 3200 15620 3206 15632
rect 5169 15623 5227 15629
rect 5169 15620 5181 15623
rect 3200 15592 5181 15620
rect 3200 15580 3206 15592
rect 5169 15589 5181 15592
rect 5215 15620 5227 15623
rect 5350 15620 5356 15632
rect 5215 15592 5356 15620
rect 5215 15589 5227 15592
rect 5169 15583 5227 15589
rect 5350 15580 5356 15592
rect 5408 15580 5414 15632
rect 11885 15623 11943 15629
rect 11885 15620 11897 15623
rect 11440 15592 11897 15620
rect 11440 15564 11468 15592
rect 11885 15589 11897 15592
rect 11931 15589 11943 15623
rect 12802 15620 12808 15632
rect 12763 15592 12808 15620
rect 11885 15583 11943 15589
rect 12802 15580 12808 15592
rect 12860 15580 12866 15632
rect 16298 15580 16304 15632
rect 16356 15620 16362 15632
rect 16942 15620 16948 15632
rect 16356 15592 16948 15620
rect 16356 15580 16362 15592
rect 16942 15580 16948 15592
rect 17000 15580 17006 15632
rect 17310 15580 17316 15632
rect 17368 15620 17374 15632
rect 17497 15623 17555 15629
rect 17497 15620 17509 15623
rect 17368 15592 17509 15620
rect 17368 15580 17374 15592
rect 17497 15589 17509 15592
rect 17543 15589 17555 15623
rect 17497 15583 17555 15589
rect 17954 15580 17960 15632
rect 18012 15620 18018 15632
rect 18524 15620 18552 15648
rect 18012 15592 18552 15620
rect 18012 15580 18018 15592
rect 2777 15555 2835 15561
rect 2777 15521 2789 15555
rect 2823 15552 2835 15555
rect 3234 15552 3240 15564
rect 2823 15524 3240 15552
rect 2823 15521 2835 15524
rect 2777 15515 2835 15521
rect 3234 15512 3240 15524
rect 3292 15512 3298 15564
rect 4522 15512 4528 15564
rect 4580 15552 4586 15564
rect 5442 15552 5448 15564
rect 4580 15524 5448 15552
rect 4580 15512 4586 15524
rect 5442 15512 5448 15524
rect 5500 15512 5506 15564
rect 6454 15512 6460 15564
rect 6512 15552 6518 15564
rect 6549 15555 6607 15561
rect 6549 15552 6561 15555
rect 6512 15524 6561 15552
rect 6512 15512 6518 15524
rect 6549 15521 6561 15524
rect 6595 15521 6607 15555
rect 6549 15515 6607 15521
rect 6914 15512 6920 15564
rect 6972 15552 6978 15564
rect 8113 15555 8171 15561
rect 8113 15552 8125 15555
rect 6972 15524 8125 15552
rect 6972 15512 6978 15524
rect 8113 15521 8125 15524
rect 8159 15552 8171 15555
rect 8202 15552 8208 15564
rect 8159 15524 8208 15552
rect 8159 15521 8171 15524
rect 8113 15515 8171 15521
rect 8202 15512 8208 15524
rect 8260 15512 8266 15564
rect 10045 15555 10103 15561
rect 10045 15521 10057 15555
rect 10091 15552 10103 15555
rect 10134 15552 10140 15564
rect 10091 15524 10140 15552
rect 10091 15521 10103 15524
rect 10045 15515 10103 15521
rect 10134 15512 10140 15524
rect 10192 15512 10198 15564
rect 11422 15512 11428 15564
rect 11480 15512 11486 15564
rect 11698 15512 11704 15564
rect 11756 15552 11762 15564
rect 11793 15555 11851 15561
rect 11793 15552 11805 15555
rect 11756 15524 11805 15552
rect 11756 15512 11762 15524
rect 11793 15521 11805 15524
rect 11839 15521 11851 15555
rect 11793 15515 11851 15521
rect 12710 15512 12716 15564
rect 12768 15552 12774 15564
rect 13357 15555 13415 15561
rect 13357 15552 13369 15555
rect 12768 15524 13369 15552
rect 12768 15512 12774 15524
rect 13357 15521 13369 15524
rect 13403 15521 13415 15555
rect 13357 15515 13415 15521
rect 18046 15512 18052 15564
rect 18104 15552 18110 15564
rect 18230 15552 18236 15564
rect 18104 15524 18236 15552
rect 18104 15512 18110 15524
rect 18230 15512 18236 15524
rect 18288 15552 18294 15564
rect 18417 15555 18475 15561
rect 18417 15552 18429 15555
rect 18288 15524 18429 15552
rect 18288 15512 18294 15524
rect 18417 15521 18429 15524
rect 18463 15521 18475 15555
rect 18417 15515 18475 15521
rect 2869 15487 2927 15493
rect 2869 15453 2881 15487
rect 2915 15453 2927 15487
rect 3050 15484 3056 15496
rect 3011 15456 3056 15484
rect 2869 15447 2927 15453
rect 1946 15376 1952 15428
rect 2004 15416 2010 15428
rect 2409 15419 2467 15425
rect 2409 15416 2421 15419
rect 2004 15388 2421 15416
rect 2004 15376 2010 15388
rect 2409 15385 2421 15388
rect 2455 15385 2467 15419
rect 2884 15416 2912 15447
rect 3050 15444 3056 15456
rect 3108 15444 3114 15496
rect 4430 15444 4436 15496
rect 4488 15484 4494 15496
rect 4617 15487 4675 15493
rect 4617 15484 4629 15487
rect 4488 15456 4629 15484
rect 4488 15444 4494 15456
rect 4617 15453 4629 15456
rect 4663 15453 4675 15487
rect 5994 15484 6000 15496
rect 5955 15456 6000 15484
rect 4617 15447 4675 15453
rect 5994 15444 6000 15456
rect 6052 15444 6058 15496
rect 6178 15444 6184 15496
rect 6236 15484 6242 15496
rect 6641 15487 6699 15493
rect 6641 15484 6653 15487
rect 6236 15456 6653 15484
rect 6236 15444 6242 15456
rect 6641 15453 6653 15456
rect 6687 15453 6699 15487
rect 6641 15447 6699 15453
rect 6825 15487 6883 15493
rect 6825 15453 6837 15487
rect 6871 15484 6883 15487
rect 8297 15487 8355 15493
rect 6871 15456 7604 15484
rect 6871 15453 6883 15456
rect 6825 15447 6883 15453
rect 2884 15388 4016 15416
rect 2409 15379 2467 15385
rect 3988 15360 4016 15388
rect 7576 15360 7604 15456
rect 8297 15453 8309 15487
rect 8343 15453 8355 15487
rect 8297 15447 8355 15453
rect 10321 15487 10379 15493
rect 10321 15453 10333 15487
rect 10367 15484 10379 15487
rect 10778 15484 10784 15496
rect 10367 15456 10784 15484
rect 10367 15453 10379 15456
rect 10321 15447 10379 15453
rect 8110 15376 8116 15428
rect 8168 15416 8174 15428
rect 8312 15416 8340 15447
rect 10778 15444 10784 15456
rect 10836 15484 10842 15496
rect 11146 15484 11152 15496
rect 10836 15456 11152 15484
rect 10836 15444 10842 15456
rect 11146 15444 11152 15456
rect 11204 15444 11210 15496
rect 11974 15484 11980 15496
rect 11935 15456 11980 15484
rect 11974 15444 11980 15456
rect 12032 15444 12038 15496
rect 13633 15487 13691 15493
rect 13633 15453 13645 15487
rect 13679 15484 13691 15487
rect 13722 15484 13728 15496
rect 13679 15456 13728 15484
rect 13679 15453 13691 15456
rect 13633 15447 13691 15453
rect 13722 15444 13728 15456
rect 13780 15444 13786 15496
rect 17129 15487 17187 15493
rect 17129 15453 17141 15487
rect 17175 15484 17187 15487
rect 17218 15484 17224 15496
rect 17175 15456 17224 15484
rect 17175 15453 17187 15456
rect 17129 15447 17187 15453
rect 17218 15444 17224 15456
rect 17276 15444 17282 15496
rect 18601 15487 18659 15493
rect 18601 15453 18613 15487
rect 18647 15453 18659 15487
rect 18601 15447 18659 15453
rect 16482 15416 16488 15428
rect 8168 15388 8340 15416
rect 16443 15388 16488 15416
rect 8168 15376 8174 15388
rect 16482 15376 16488 15388
rect 16540 15376 16546 15428
rect 18616 15416 18644 15447
rect 17880 15388 18644 15416
rect 17880 15360 17908 15388
rect 3970 15308 3976 15360
rect 4028 15348 4034 15360
rect 4065 15351 4123 15357
rect 4065 15348 4077 15351
rect 4028 15320 4077 15348
rect 4028 15308 4034 15320
rect 4065 15317 4077 15320
rect 4111 15317 4123 15351
rect 4065 15311 4123 15317
rect 6181 15351 6239 15357
rect 6181 15317 6193 15351
rect 6227 15348 6239 15351
rect 6822 15348 6828 15360
rect 6227 15320 6828 15348
rect 6227 15317 6239 15320
rect 6181 15311 6239 15317
rect 6822 15308 6828 15320
rect 6880 15308 6886 15360
rect 7558 15348 7564 15360
rect 7519 15320 7564 15348
rect 7558 15308 7564 15320
rect 7616 15308 7622 15360
rect 8849 15351 8907 15357
rect 8849 15317 8861 15351
rect 8895 15348 8907 15351
rect 9214 15348 9220 15360
rect 8895 15320 9220 15348
rect 8895 15317 8907 15320
rect 8849 15311 8907 15317
rect 9214 15308 9220 15320
rect 9272 15348 9278 15360
rect 9582 15348 9588 15360
rect 9272 15320 9588 15348
rect 9272 15308 9278 15320
rect 9582 15308 9588 15320
rect 9640 15308 9646 15360
rect 14366 15348 14372 15360
rect 14327 15320 14372 15348
rect 14366 15308 14372 15320
rect 14424 15308 14430 15360
rect 17862 15348 17868 15360
rect 17823 15320 17868 15348
rect 17862 15308 17868 15320
rect 17920 15308 17926 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 3234 15104 3240 15156
rect 3292 15144 3298 15156
rect 4709 15147 4767 15153
rect 4709 15144 4721 15147
rect 3292 15116 4721 15144
rect 3292 15104 3298 15116
rect 4709 15113 4721 15116
rect 4755 15144 4767 15147
rect 5350 15144 5356 15156
rect 4755 15116 5356 15144
rect 4755 15113 4767 15116
rect 4709 15107 4767 15113
rect 5350 15104 5356 15116
rect 5408 15104 5414 15156
rect 6825 15147 6883 15153
rect 6825 15113 6837 15147
rect 6871 15144 6883 15147
rect 6914 15144 6920 15156
rect 6871 15116 6920 15144
rect 6871 15113 6883 15116
rect 6825 15107 6883 15113
rect 6914 15104 6920 15116
rect 6972 15104 6978 15156
rect 8297 15147 8355 15153
rect 8297 15113 8309 15147
rect 8343 15144 8355 15147
rect 8478 15144 8484 15156
rect 8343 15116 8484 15144
rect 8343 15113 8355 15116
rect 8297 15107 8355 15113
rect 1486 14968 1492 15020
rect 1544 15008 1550 15020
rect 1673 15011 1731 15017
rect 1673 15008 1685 15011
rect 1544 14980 1685 15008
rect 1544 14968 1550 14980
rect 1673 14977 1685 14980
rect 1719 14977 1731 15011
rect 1673 14971 1731 14977
rect 4154 14968 4160 15020
rect 4212 15008 4218 15020
rect 5166 15008 5172 15020
rect 4212 14980 5172 15008
rect 4212 14968 4218 14980
rect 5166 14968 5172 14980
rect 5224 14968 5230 15020
rect 5353 15011 5411 15017
rect 5353 14977 5365 15011
rect 5399 14977 5411 15011
rect 5353 14971 5411 14977
rect 7469 15011 7527 15017
rect 7469 14977 7481 15011
rect 7515 15008 7527 15011
rect 8312 15008 8340 15107
rect 8478 15104 8484 15116
rect 8536 15104 8542 15156
rect 10778 15144 10784 15156
rect 10739 15116 10784 15144
rect 10778 15104 10784 15116
rect 10836 15104 10842 15156
rect 11698 15104 11704 15156
rect 11756 15144 11762 15156
rect 11793 15147 11851 15153
rect 11793 15144 11805 15147
rect 11756 15116 11805 15144
rect 11756 15104 11762 15116
rect 11793 15113 11805 15116
rect 11839 15144 11851 15147
rect 11882 15144 11888 15156
rect 11839 15116 11888 15144
rect 11839 15113 11851 15116
rect 11793 15107 11851 15113
rect 11882 15104 11888 15116
rect 11940 15104 11946 15156
rect 11974 15104 11980 15156
rect 12032 15144 12038 15156
rect 12161 15147 12219 15153
rect 12161 15144 12173 15147
rect 12032 15116 12173 15144
rect 12032 15104 12038 15116
rect 12161 15113 12173 15116
rect 12207 15144 12219 15147
rect 12713 15147 12771 15153
rect 12713 15144 12725 15147
rect 12207 15116 12725 15144
rect 12207 15113 12219 15116
rect 12161 15107 12219 15113
rect 12713 15113 12725 15116
rect 12759 15144 12771 15147
rect 13630 15144 13636 15156
rect 12759 15116 13636 15144
rect 12759 15113 12771 15116
rect 12713 15107 12771 15113
rect 13630 15104 13636 15116
rect 13688 15104 13694 15156
rect 14734 15104 14740 15156
rect 14792 15144 14798 15156
rect 15013 15147 15071 15153
rect 15013 15144 15025 15147
rect 14792 15116 15025 15144
rect 14792 15104 14798 15116
rect 15013 15113 15025 15116
rect 15059 15113 15071 15147
rect 15013 15107 15071 15113
rect 16114 15104 16120 15156
rect 16172 15144 16178 15156
rect 16393 15147 16451 15153
rect 16393 15144 16405 15147
rect 16172 15116 16405 15144
rect 16172 15104 16178 15116
rect 16393 15113 16405 15116
rect 16439 15113 16451 15147
rect 17494 15144 17500 15156
rect 17407 15116 17500 15144
rect 16393 15107 16451 15113
rect 17494 15104 17500 15116
rect 17552 15144 17558 15156
rect 17954 15144 17960 15156
rect 17552 15116 17960 15144
rect 17552 15104 17558 15116
rect 17954 15104 17960 15116
rect 18012 15104 18018 15156
rect 12618 15036 12624 15088
rect 12676 15076 12682 15088
rect 13170 15076 13176 15088
rect 12676 15048 13176 15076
rect 12676 15036 12682 15048
rect 13170 15036 13176 15048
rect 13228 15076 13234 15088
rect 13357 15079 13415 15085
rect 13357 15076 13369 15079
rect 13228 15048 13369 15076
rect 13228 15036 13234 15048
rect 13357 15045 13369 15048
rect 13403 15045 13415 15079
rect 13357 15039 13415 15045
rect 15933 15079 15991 15085
rect 15933 15045 15945 15079
rect 15979 15076 15991 15079
rect 16298 15076 16304 15088
rect 15979 15048 16304 15076
rect 15979 15045 15991 15048
rect 15933 15039 15991 15045
rect 16298 15036 16304 15048
rect 16356 15036 16362 15088
rect 17586 15036 17592 15088
rect 17644 15076 17650 15088
rect 17865 15079 17923 15085
rect 17865 15076 17877 15079
rect 17644 15048 17877 15076
rect 17644 15036 17650 15048
rect 17865 15045 17877 15048
rect 17911 15076 17923 15079
rect 18046 15076 18052 15088
rect 17911 15048 18052 15076
rect 17911 15045 17923 15048
rect 17865 15039 17923 15045
rect 18046 15036 18052 15048
rect 18104 15036 18110 15088
rect 7515 14980 8340 15008
rect 7515 14977 7527 14980
rect 7469 14971 7527 14977
rect 1940 14875 1998 14881
rect 1940 14841 1952 14875
rect 1986 14872 1998 14875
rect 2130 14872 2136 14884
rect 1986 14844 2136 14872
rect 1986 14841 1998 14844
rect 1940 14835 1998 14841
rect 2130 14832 2136 14844
rect 2188 14832 2194 14884
rect 4617 14875 4675 14881
rect 4617 14841 4629 14875
rect 4663 14872 4675 14875
rect 5074 14872 5080 14884
rect 4663 14844 5080 14872
rect 4663 14841 4675 14844
rect 4617 14835 4675 14841
rect 5074 14832 5080 14844
rect 5132 14832 5138 14884
rect 3050 14804 3056 14816
rect 3011 14776 3056 14804
rect 3050 14764 3056 14776
rect 3108 14764 3114 14816
rect 3786 14804 3792 14816
rect 3747 14776 3792 14804
rect 3786 14764 3792 14776
rect 3844 14804 3850 14816
rect 4157 14807 4215 14813
rect 4157 14804 4169 14807
rect 3844 14776 4169 14804
rect 3844 14764 3850 14776
rect 4157 14773 4169 14776
rect 4203 14804 4215 14807
rect 4430 14804 4436 14816
rect 4203 14776 4436 14804
rect 4203 14773 4215 14776
rect 4157 14767 4215 14773
rect 4430 14764 4436 14776
rect 4488 14804 4494 14816
rect 5368 14804 5396 14971
rect 16574 14968 16580 15020
rect 16632 15008 16638 15020
rect 16853 15011 16911 15017
rect 16853 15008 16865 15011
rect 16632 14980 16865 15008
rect 16632 14968 16638 14980
rect 16853 14977 16865 14980
rect 16899 14977 16911 15011
rect 16853 14971 16911 14977
rect 16945 15011 17003 15017
rect 16945 14977 16957 15011
rect 16991 14977 17003 15011
rect 16945 14971 17003 14977
rect 6914 14900 6920 14952
rect 6972 14940 6978 14952
rect 7193 14943 7251 14949
rect 7193 14940 7205 14943
rect 6972 14912 7205 14940
rect 6972 14900 6978 14912
rect 7193 14909 7205 14912
rect 7239 14909 7251 14943
rect 8754 14940 8760 14952
rect 8715 14912 8760 14940
rect 7193 14903 7251 14909
rect 8754 14900 8760 14912
rect 8812 14900 8818 14952
rect 12434 14900 12440 14952
rect 12492 14940 12498 14952
rect 13078 14940 13084 14952
rect 12492 14912 13084 14940
rect 12492 14900 12498 14912
rect 13078 14900 13084 14912
rect 13136 14940 13142 14952
rect 13906 14949 13912 14952
rect 13633 14943 13691 14949
rect 13633 14940 13645 14943
rect 13136 14912 13645 14940
rect 13136 14900 13142 14912
rect 13633 14909 13645 14912
rect 13679 14909 13691 14943
rect 13900 14940 13912 14949
rect 13819 14912 13912 14940
rect 13633 14903 13691 14909
rect 13900 14903 13912 14912
rect 13964 14940 13970 14952
rect 14366 14940 14372 14952
rect 13964 14912 14372 14940
rect 13906 14900 13912 14903
rect 13964 14900 13970 14912
rect 14366 14900 14372 14912
rect 14424 14900 14430 14952
rect 16301 14943 16359 14949
rect 16301 14909 16313 14943
rect 16347 14940 16359 14943
rect 16960 14940 16988 14971
rect 16347 14912 16988 14940
rect 16347 14909 16359 14912
rect 16301 14903 16359 14909
rect 5905 14875 5963 14881
rect 5905 14841 5917 14875
rect 5951 14872 5963 14875
rect 7098 14872 7104 14884
rect 5951 14844 7104 14872
rect 5951 14841 5963 14844
rect 5905 14835 5963 14841
rect 7098 14832 7104 14844
rect 7156 14832 7162 14884
rect 7929 14875 7987 14881
rect 7929 14841 7941 14875
rect 7975 14872 7987 14875
rect 8110 14872 8116 14884
rect 7975 14844 8116 14872
rect 7975 14841 7987 14844
rect 7929 14835 7987 14841
rect 8110 14832 8116 14844
rect 8168 14872 8174 14884
rect 8665 14875 8723 14881
rect 8665 14872 8677 14875
rect 8168 14844 8677 14872
rect 8168 14832 8174 14844
rect 8665 14841 8677 14844
rect 8711 14872 8723 14875
rect 8938 14872 8944 14884
rect 8711 14844 8944 14872
rect 8711 14841 8723 14844
rect 8665 14835 8723 14841
rect 8938 14832 8944 14844
rect 8996 14881 9002 14884
rect 8996 14875 9060 14881
rect 8996 14841 9014 14875
rect 9048 14841 9060 14875
rect 16960 14872 16988 14912
rect 18049 14943 18107 14949
rect 18049 14909 18061 14943
rect 18095 14940 18107 14943
rect 18690 14940 18696 14952
rect 18095 14912 18696 14940
rect 18095 14909 18107 14912
rect 18049 14903 18107 14909
rect 18690 14900 18696 14912
rect 18748 14900 18754 14952
rect 18322 14881 18328 14884
rect 18294 14875 18328 14881
rect 18294 14872 18306 14875
rect 16960 14844 18306 14872
rect 8996 14835 9060 14841
rect 18294 14841 18306 14844
rect 18380 14872 18386 14884
rect 18380 14844 18442 14872
rect 18294 14835 18328 14841
rect 8996 14832 9002 14835
rect 18322 14832 18328 14835
rect 18380 14832 18386 14844
rect 6178 14804 6184 14816
rect 4488 14776 5396 14804
rect 6139 14776 6184 14804
rect 4488 14764 4494 14776
rect 6178 14764 6184 14776
rect 6236 14764 6242 14816
rect 6454 14764 6460 14816
rect 6512 14804 6518 14816
rect 6549 14807 6607 14813
rect 6549 14804 6561 14807
rect 6512 14776 6561 14804
rect 6512 14764 6518 14776
rect 6549 14773 6561 14776
rect 6595 14773 6607 14807
rect 6549 14767 6607 14773
rect 7285 14807 7343 14813
rect 7285 14773 7297 14807
rect 7331 14804 7343 14807
rect 8294 14804 8300 14816
rect 7331 14776 8300 14804
rect 7331 14773 7343 14776
rect 7285 14767 7343 14773
rect 8294 14764 8300 14776
rect 8352 14764 8358 14816
rect 9582 14764 9588 14816
rect 9640 14804 9646 14816
rect 10042 14804 10048 14816
rect 9640 14776 10048 14804
rect 9640 14764 9646 14776
rect 10042 14764 10048 14776
rect 10100 14804 10106 14816
rect 10137 14807 10195 14813
rect 10137 14804 10149 14807
rect 10100 14776 10149 14804
rect 10100 14764 10106 14776
rect 10137 14773 10149 14776
rect 10183 14773 10195 14807
rect 11054 14804 11060 14816
rect 11015 14776 11060 14804
rect 10137 14767 10195 14773
rect 11054 14764 11060 14776
rect 11112 14764 11118 14816
rect 11422 14804 11428 14816
rect 11383 14776 11428 14804
rect 11422 14764 11428 14776
rect 11480 14764 11486 14816
rect 12710 14764 12716 14816
rect 12768 14804 12774 14816
rect 12989 14807 13047 14813
rect 12989 14804 13001 14807
rect 12768 14776 13001 14804
rect 12768 14764 12774 14776
rect 12989 14773 13001 14776
rect 13035 14773 13047 14807
rect 12989 14767 13047 14773
rect 13354 14764 13360 14816
rect 13412 14804 13418 14816
rect 15378 14804 15384 14816
rect 13412 14776 15384 14804
rect 13412 14764 13418 14776
rect 15378 14764 15384 14776
rect 15436 14764 15442 14816
rect 16758 14804 16764 14816
rect 16719 14776 16764 14804
rect 16758 14764 16764 14776
rect 16816 14764 16822 14816
rect 19426 14804 19432 14816
rect 19387 14776 19432 14804
rect 19426 14764 19432 14776
rect 19484 14764 19490 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1397 14603 1455 14609
rect 1397 14569 1409 14603
rect 1443 14600 1455 14603
rect 1670 14600 1676 14612
rect 1443 14572 1676 14600
rect 1443 14569 1455 14572
rect 1397 14563 1455 14569
rect 1670 14560 1676 14572
rect 1728 14560 1734 14612
rect 2406 14600 2412 14612
rect 2367 14572 2412 14600
rect 2406 14560 2412 14572
rect 2464 14560 2470 14612
rect 3050 14560 3056 14612
rect 3108 14600 3114 14612
rect 3789 14603 3847 14609
rect 3789 14600 3801 14603
rect 3108 14572 3801 14600
rect 3108 14560 3114 14572
rect 3789 14569 3801 14572
rect 3835 14569 3847 14603
rect 3789 14563 3847 14569
rect 5442 14560 5448 14612
rect 5500 14600 5506 14612
rect 6089 14603 6147 14609
rect 6089 14600 6101 14603
rect 5500 14572 6101 14600
rect 5500 14560 5506 14572
rect 6089 14569 6101 14572
rect 6135 14569 6147 14603
rect 6089 14563 6147 14569
rect 6914 14560 6920 14612
rect 6972 14600 6978 14612
rect 8941 14603 8999 14609
rect 8941 14600 8953 14603
rect 6972 14572 8953 14600
rect 6972 14560 6978 14572
rect 8941 14569 8953 14572
rect 8987 14569 8999 14603
rect 8941 14563 8999 14569
rect 10873 14603 10931 14609
rect 10873 14569 10885 14603
rect 10919 14600 10931 14603
rect 11146 14600 11152 14612
rect 10919 14572 11152 14600
rect 10919 14569 10931 14572
rect 10873 14563 10931 14569
rect 11146 14560 11152 14572
rect 11204 14600 11210 14612
rect 12621 14603 12679 14609
rect 12621 14600 12633 14603
rect 11204 14572 12633 14600
rect 11204 14560 11210 14572
rect 12621 14569 12633 14572
rect 12667 14569 12679 14603
rect 12621 14563 12679 14569
rect 12986 14560 12992 14612
rect 13044 14600 13050 14612
rect 13633 14603 13691 14609
rect 13633 14600 13645 14603
rect 13044 14572 13645 14600
rect 13044 14560 13050 14572
rect 13633 14569 13645 14572
rect 13679 14569 13691 14603
rect 13633 14563 13691 14569
rect 14001 14603 14059 14609
rect 14001 14569 14013 14603
rect 14047 14600 14059 14603
rect 14182 14600 14188 14612
rect 14047 14572 14188 14600
rect 14047 14569 14059 14572
rect 14001 14563 14059 14569
rect 14182 14560 14188 14572
rect 14240 14560 14246 14612
rect 18322 14600 18328 14612
rect 18283 14572 18328 14600
rect 18322 14560 18328 14572
rect 18380 14600 18386 14612
rect 18877 14603 18935 14609
rect 18877 14600 18889 14603
rect 18380 14572 18889 14600
rect 18380 14560 18386 14572
rect 18877 14569 18889 14572
rect 18923 14569 18935 14603
rect 18877 14563 18935 14569
rect 2869 14535 2927 14541
rect 2869 14501 2881 14535
rect 2915 14532 2927 14535
rect 3142 14532 3148 14544
rect 2915 14504 3148 14532
rect 2915 14501 2927 14504
rect 2869 14495 2927 14501
rect 3142 14492 3148 14504
rect 3200 14532 3206 14544
rect 3326 14532 3332 14544
rect 3200 14504 3332 14532
rect 3200 14492 3206 14504
rect 3326 14492 3332 14504
rect 3384 14492 3390 14544
rect 5534 14492 5540 14544
rect 5592 14532 5598 14544
rect 6457 14535 6515 14541
rect 6457 14532 6469 14535
rect 5592 14504 6469 14532
rect 5592 14492 5598 14504
rect 6457 14501 6469 14504
rect 6503 14501 6515 14535
rect 6457 14495 6515 14501
rect 7098 14492 7104 14544
rect 7156 14532 7162 14544
rect 7558 14532 7564 14544
rect 7156 14504 7564 14532
rect 7156 14492 7162 14504
rect 7558 14492 7564 14504
rect 7616 14492 7622 14544
rect 8202 14492 8208 14544
rect 8260 14532 8266 14544
rect 9309 14535 9367 14541
rect 9309 14532 9321 14535
rect 8260 14504 9321 14532
rect 8260 14492 8266 14504
rect 9309 14501 9321 14504
rect 9355 14501 9367 14535
rect 9309 14495 9367 14501
rect 9950 14492 9956 14544
rect 10008 14532 10014 14544
rect 10045 14535 10103 14541
rect 10045 14532 10057 14535
rect 10008 14504 10057 14532
rect 10008 14492 10014 14504
rect 10045 14501 10057 14504
rect 10091 14501 10103 14535
rect 10045 14495 10103 14501
rect 12526 14492 12532 14544
rect 12584 14532 12590 14544
rect 13541 14535 13599 14541
rect 13541 14532 13553 14535
rect 12584 14504 13553 14532
rect 12584 14492 12590 14504
rect 13541 14501 13553 14504
rect 13587 14532 13599 14535
rect 14093 14535 14151 14541
rect 14093 14532 14105 14535
rect 13587 14504 14105 14532
rect 13587 14501 13599 14504
rect 13541 14495 13599 14501
rect 14093 14501 14105 14504
rect 14139 14532 14151 14535
rect 14550 14532 14556 14544
rect 14139 14504 14556 14532
rect 14139 14501 14151 14504
rect 14093 14495 14151 14501
rect 14550 14492 14556 14504
rect 14608 14492 14614 14544
rect 15654 14532 15660 14544
rect 15615 14504 15660 14532
rect 15654 14492 15660 14504
rect 15712 14492 15718 14544
rect 2774 14424 2780 14476
rect 2832 14464 2838 14476
rect 4246 14464 4252 14476
rect 2832 14436 2877 14464
rect 3068 14436 4252 14464
rect 2832 14424 2838 14436
rect 3068 14405 3096 14436
rect 4246 14424 4252 14436
rect 4304 14464 4310 14476
rect 4424 14467 4482 14473
rect 4424 14464 4436 14467
rect 4304 14436 4436 14464
rect 4304 14424 4310 14436
rect 4424 14433 4436 14436
rect 4470 14464 4482 14467
rect 6546 14464 6552 14476
rect 4470 14436 6552 14464
rect 4470 14433 4482 14436
rect 4424 14427 4482 14433
rect 6546 14424 6552 14436
rect 6604 14424 6610 14476
rect 6908 14467 6966 14473
rect 6908 14433 6920 14467
rect 6954 14464 6966 14467
rect 7116 14464 7144 14492
rect 6954 14436 7144 14464
rect 9769 14467 9827 14473
rect 6954 14433 6966 14436
rect 6908 14427 6966 14433
rect 9769 14433 9781 14467
rect 9815 14433 9827 14467
rect 9769 14427 9827 14433
rect 2317 14399 2375 14405
rect 2317 14365 2329 14399
rect 2363 14396 2375 14399
rect 3053 14399 3111 14405
rect 3053 14396 3065 14399
rect 2363 14368 3065 14396
rect 2363 14365 2375 14368
rect 2317 14359 2375 14365
rect 3053 14365 3065 14368
rect 3099 14365 3111 14399
rect 4154 14396 4160 14408
rect 4115 14368 4160 14396
rect 3053 14359 3111 14365
rect 4154 14356 4160 14368
rect 4212 14356 4218 14408
rect 6641 14399 6699 14405
rect 6641 14365 6653 14399
rect 6687 14365 6699 14399
rect 6641 14359 6699 14365
rect 2130 14288 2136 14340
rect 2188 14328 2194 14340
rect 3421 14331 3479 14337
rect 3421 14328 3433 14331
rect 2188 14300 3433 14328
rect 2188 14288 2194 14300
rect 3421 14297 3433 14300
rect 3467 14328 3479 14331
rect 3786 14328 3792 14340
rect 3467 14300 3792 14328
rect 3467 14297 3479 14300
rect 3421 14291 3479 14297
rect 3786 14288 3792 14300
rect 3844 14288 3850 14340
rect 1762 14220 1768 14272
rect 1820 14260 1826 14272
rect 1857 14263 1915 14269
rect 1857 14260 1869 14263
rect 1820 14232 1869 14260
rect 1820 14220 1826 14232
rect 1857 14229 1869 14232
rect 1903 14229 1915 14263
rect 3804 14260 3832 14288
rect 5537 14263 5595 14269
rect 5537 14260 5549 14263
rect 3804 14232 5549 14260
rect 1857 14223 1915 14229
rect 5537 14229 5549 14232
rect 5583 14229 5595 14263
rect 6656 14260 6684 14359
rect 9784 14340 9812 14427
rect 11054 14424 11060 14476
rect 11112 14464 11118 14476
rect 11425 14467 11483 14473
rect 11425 14464 11437 14467
rect 11112 14436 11437 14464
rect 11112 14424 11118 14436
rect 11425 14433 11437 14436
rect 11471 14433 11483 14467
rect 11425 14427 11483 14433
rect 12342 14424 12348 14476
rect 12400 14464 12406 14476
rect 15746 14464 15752 14476
rect 12400 14436 15752 14464
rect 12400 14424 12406 14436
rect 15746 14424 15752 14436
rect 15804 14424 15810 14476
rect 17218 14473 17224 14476
rect 16577 14467 16635 14473
rect 16577 14433 16589 14467
rect 16623 14464 16635 14467
rect 17212 14464 17224 14473
rect 16623 14436 17224 14464
rect 16623 14433 16635 14436
rect 16577 14427 16635 14433
rect 17212 14427 17224 14436
rect 17218 14424 17224 14427
rect 17276 14424 17282 14476
rect 11514 14396 11520 14408
rect 11475 14368 11520 14396
rect 11514 14356 11520 14368
rect 11572 14356 11578 14408
rect 11698 14396 11704 14408
rect 11659 14368 11704 14396
rect 11698 14356 11704 14368
rect 11756 14356 11762 14408
rect 14274 14396 14280 14408
rect 14235 14368 14280 14396
rect 14274 14356 14280 14368
rect 14332 14356 14338 14408
rect 14550 14356 14556 14408
rect 14608 14396 14614 14408
rect 15013 14399 15071 14405
rect 15013 14396 15025 14399
rect 14608 14368 15025 14396
rect 14608 14356 14614 14368
rect 15013 14365 15025 14368
rect 15059 14396 15071 14399
rect 15930 14396 15936 14408
rect 15059 14368 15936 14396
rect 15059 14365 15071 14368
rect 15013 14359 15071 14365
rect 15930 14356 15936 14368
rect 15988 14356 15994 14408
rect 16945 14399 17003 14405
rect 16945 14365 16957 14399
rect 16991 14365 17003 14399
rect 16945 14359 17003 14365
rect 7742 14288 7748 14340
rect 7800 14328 7806 14340
rect 8021 14331 8079 14337
rect 8021 14328 8033 14331
rect 7800 14300 8033 14328
rect 7800 14288 7806 14300
rect 8021 14297 8033 14300
rect 8067 14328 8079 14331
rect 8478 14328 8484 14340
rect 8067 14300 8484 14328
rect 8067 14297 8079 14300
rect 8021 14291 8079 14297
rect 8478 14288 8484 14300
rect 8536 14288 8542 14340
rect 9766 14328 9772 14340
rect 9679 14300 9772 14328
rect 9766 14288 9772 14300
rect 9824 14328 9830 14340
rect 11057 14331 11115 14337
rect 11057 14328 11069 14331
rect 9824 14300 11069 14328
rect 9824 14288 9830 14300
rect 11057 14297 11069 14300
rect 11103 14297 11115 14331
rect 13170 14328 13176 14340
rect 13083 14300 13176 14328
rect 11057 14291 11115 14297
rect 13170 14288 13176 14300
rect 13228 14328 13234 14340
rect 14292 14328 14320 14356
rect 13228 14300 14320 14328
rect 13228 14288 13234 14300
rect 8202 14260 8208 14272
rect 6656 14232 8208 14260
rect 5537 14223 5595 14229
rect 8202 14220 8208 14232
rect 8260 14220 8266 14272
rect 8294 14220 8300 14272
rect 8352 14260 8358 14272
rect 8665 14263 8723 14269
rect 8665 14260 8677 14263
rect 8352 14232 8677 14260
rect 8352 14220 8358 14232
rect 8665 14229 8677 14232
rect 8711 14260 8723 14263
rect 9398 14260 9404 14272
rect 8711 14232 9404 14260
rect 8711 14229 8723 14232
rect 8665 14223 8723 14229
rect 9398 14220 9404 14232
rect 9456 14220 9462 14272
rect 12066 14260 12072 14272
rect 12027 14232 12072 14260
rect 12066 14220 12072 14232
rect 12124 14220 12130 14272
rect 12434 14260 12440 14272
rect 12395 14232 12440 14260
rect 12434 14220 12440 14232
rect 12492 14220 12498 14272
rect 15289 14263 15347 14269
rect 15289 14229 15301 14263
rect 15335 14260 15347 14263
rect 15378 14260 15384 14272
rect 15335 14232 15384 14260
rect 15335 14229 15347 14232
rect 15289 14223 15347 14229
rect 15378 14220 15384 14232
rect 15436 14220 15442 14272
rect 16482 14220 16488 14272
rect 16540 14260 16546 14272
rect 16960 14260 16988 14359
rect 18690 14260 18696 14272
rect 16540 14232 18696 14260
rect 16540 14220 16546 14232
rect 18690 14220 18696 14232
rect 18748 14220 18754 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 1394 14056 1400 14068
rect 1355 14028 1400 14056
rect 1394 14016 1400 14028
rect 1452 14016 1458 14068
rect 2501 14059 2559 14065
rect 2501 14025 2513 14059
rect 2547 14056 2559 14059
rect 3142 14056 3148 14068
rect 2547 14028 3148 14056
rect 2547 14025 2559 14028
rect 2501 14019 2559 14025
rect 3142 14016 3148 14028
rect 3200 14016 3206 14068
rect 4157 14059 4215 14065
rect 4157 14025 4169 14059
rect 4203 14056 4215 14059
rect 4338 14056 4344 14068
rect 4203 14028 4344 14056
rect 4203 14025 4215 14028
rect 4157 14019 4215 14025
rect 4338 14016 4344 14028
rect 4396 14056 4402 14068
rect 4396 14028 4752 14056
rect 4396 14016 4402 14028
rect 2774 13948 2780 14000
rect 2832 13988 2838 14000
rect 4724 13988 4752 14028
rect 5166 14016 5172 14068
rect 5224 14056 5230 14068
rect 5997 14059 6055 14065
rect 5997 14056 6009 14059
rect 5224 14028 6009 14056
rect 5224 14016 5230 14028
rect 5997 14025 6009 14028
rect 6043 14025 6055 14059
rect 5997 14019 6055 14025
rect 6086 14016 6092 14068
rect 6144 14056 6150 14068
rect 6365 14059 6423 14065
rect 6365 14056 6377 14059
rect 6144 14028 6377 14056
rect 6144 14016 6150 14028
rect 6365 14025 6377 14028
rect 6411 14025 6423 14059
rect 6365 14019 6423 14025
rect 7469 14059 7527 14065
rect 7469 14025 7481 14059
rect 7515 14056 7527 14059
rect 7742 14056 7748 14068
rect 7515 14028 7748 14056
rect 7515 14025 7527 14028
rect 7469 14019 7527 14025
rect 7742 14016 7748 14028
rect 7800 14016 7806 14068
rect 8938 14056 8944 14068
rect 8899 14028 8944 14056
rect 8938 14016 8944 14028
rect 8996 14016 9002 14068
rect 9766 14056 9772 14068
rect 9727 14028 9772 14056
rect 9766 14016 9772 14028
rect 9824 14016 9830 14068
rect 10781 14059 10839 14065
rect 10781 14025 10793 14059
rect 10827 14056 10839 14059
rect 11054 14056 11060 14068
rect 10827 14028 11060 14056
rect 10827 14025 10839 14028
rect 10781 14019 10839 14025
rect 11054 14016 11060 14028
rect 11112 14016 11118 14068
rect 11698 14016 11704 14068
rect 11756 14056 11762 14068
rect 11793 14059 11851 14065
rect 11793 14056 11805 14059
rect 11756 14028 11805 14056
rect 11756 14016 11762 14028
rect 11793 14025 11805 14028
rect 11839 14056 11851 14059
rect 13817 14059 13875 14065
rect 13817 14056 13829 14059
rect 11839 14028 13829 14056
rect 11839 14025 11851 14028
rect 11793 14019 11851 14025
rect 13817 14025 13829 14028
rect 13863 14056 13875 14059
rect 13906 14056 13912 14068
rect 13863 14028 13912 14056
rect 13863 14025 13875 14028
rect 13817 14019 13875 14025
rect 13906 14016 13912 14028
rect 13964 14016 13970 14068
rect 14182 14016 14188 14068
rect 14240 14056 14246 14068
rect 14366 14056 14372 14068
rect 14240 14028 14372 14056
rect 14240 14016 14246 14028
rect 14366 14016 14372 14028
rect 14424 14016 14430 14068
rect 15746 14016 15752 14068
rect 15804 14056 15810 14068
rect 15933 14059 15991 14065
rect 15933 14056 15945 14059
rect 15804 14028 15945 14056
rect 15804 14016 15810 14028
rect 15933 14025 15945 14028
rect 15979 14025 15991 14059
rect 15933 14019 15991 14025
rect 16758 14016 16764 14068
rect 16816 14056 16822 14068
rect 17405 14059 17463 14065
rect 17405 14056 17417 14059
rect 16816 14028 17417 14056
rect 16816 14016 16822 14028
rect 17405 14025 17417 14028
rect 17451 14056 17463 14059
rect 17954 14056 17960 14068
rect 17451 14028 17960 14056
rect 17451 14025 17463 14028
rect 17405 14019 17463 14025
rect 17954 14016 17960 14028
rect 18012 14016 18018 14068
rect 25498 14056 25504 14068
rect 25459 14028 25504 14056
rect 25498 14016 25504 14028
rect 25556 14016 25562 14068
rect 5721 13991 5779 13997
rect 2832 13960 2877 13988
rect 4724 13960 5396 13988
rect 2832 13948 2838 13960
rect 2041 13923 2099 13929
rect 2041 13889 2053 13923
rect 2087 13920 2099 13923
rect 2130 13920 2136 13932
rect 2087 13892 2136 13920
rect 2087 13889 2099 13892
rect 2041 13883 2099 13889
rect 2130 13880 2136 13892
rect 2188 13880 2194 13932
rect 4724 13929 4752 13960
rect 4709 13923 4767 13929
rect 4709 13889 4721 13923
rect 4755 13889 4767 13923
rect 4709 13883 4767 13889
rect 4893 13923 4951 13929
rect 4893 13889 4905 13923
rect 4939 13889 4951 13923
rect 5368 13920 5396 13960
rect 5721 13957 5733 13991
rect 5767 13988 5779 13991
rect 6546 13988 6552 14000
rect 5767 13960 6552 13988
rect 5767 13957 5779 13960
rect 5721 13951 5779 13957
rect 6546 13948 6552 13960
rect 6604 13948 6610 14000
rect 15654 13948 15660 14000
rect 15712 13988 15718 14000
rect 16301 13991 16359 13997
rect 16301 13988 16313 13991
rect 15712 13960 16313 13988
rect 15712 13948 15718 13960
rect 16301 13957 16313 13960
rect 16347 13957 16359 13991
rect 16301 13951 16359 13957
rect 6086 13920 6092 13932
rect 5368 13892 6092 13920
rect 4893 13883 4951 13889
rect 2958 13852 2964 13864
rect 2919 13824 2964 13852
rect 2958 13812 2964 13824
rect 3016 13812 3022 13864
rect 3234 13852 3240 13864
rect 3195 13824 3240 13852
rect 3234 13812 3240 13824
rect 3292 13812 3298 13864
rect 4908 13852 4936 13883
rect 6086 13880 6092 13892
rect 6144 13880 6150 13932
rect 10321 13923 10379 13929
rect 10321 13889 10333 13923
rect 10367 13920 10379 13923
rect 11333 13923 11391 13929
rect 11333 13920 11345 13923
rect 10367 13892 11345 13920
rect 10367 13889 10379 13892
rect 10321 13883 10379 13889
rect 11333 13889 11345 13892
rect 11379 13920 11391 13923
rect 11974 13920 11980 13932
rect 11379 13892 11980 13920
rect 11379 13889 11391 13892
rect 11333 13883 11391 13889
rect 11974 13880 11980 13892
rect 12032 13920 12038 13932
rect 12161 13923 12219 13929
rect 12161 13920 12173 13923
rect 12032 13892 12173 13920
rect 12032 13880 12038 13892
rect 12161 13889 12173 13892
rect 12207 13920 12219 13923
rect 15381 13923 15439 13929
rect 12207 13892 12572 13920
rect 12207 13889 12219 13892
rect 12161 13883 12219 13889
rect 5074 13852 5080 13864
rect 4908 13824 5080 13852
rect 5074 13812 5080 13824
rect 5132 13852 5138 13864
rect 5261 13855 5319 13861
rect 5261 13852 5273 13855
rect 5132 13824 5273 13852
rect 5132 13812 5138 13824
rect 5261 13821 5273 13824
rect 5307 13821 5319 13855
rect 7098 13852 7104 13864
rect 7059 13824 7104 13852
rect 5261 13815 5319 13821
rect 7098 13812 7104 13824
rect 7156 13812 7162 13864
rect 7834 13861 7840 13864
rect 7561 13855 7619 13861
rect 7561 13821 7573 13855
rect 7607 13852 7619 13855
rect 7828 13852 7840 13861
rect 7607 13824 7696 13852
rect 7795 13824 7840 13852
rect 7607 13821 7619 13824
rect 7561 13815 7619 13821
rect 4617 13787 4675 13793
rect 4617 13784 4629 13787
rect 3712 13756 4629 13784
rect 1762 13716 1768 13728
rect 1723 13688 1768 13716
rect 1762 13676 1768 13688
rect 1820 13676 1826 13728
rect 1857 13719 1915 13725
rect 1857 13685 1869 13719
rect 1903 13716 1915 13719
rect 2314 13716 2320 13728
rect 1903 13688 2320 13716
rect 1903 13685 1915 13688
rect 1857 13679 1915 13685
rect 2314 13676 2320 13688
rect 2372 13676 2378 13728
rect 3510 13676 3516 13728
rect 3568 13716 3574 13728
rect 3712 13725 3740 13756
rect 4617 13753 4629 13756
rect 4663 13784 4675 13787
rect 7374 13784 7380 13796
rect 4663 13756 7380 13784
rect 4663 13753 4675 13756
rect 4617 13747 4675 13753
rect 7374 13744 7380 13756
rect 7432 13744 7438 13796
rect 7668 13784 7696 13824
rect 7828 13815 7840 13824
rect 7834 13812 7840 13815
rect 7892 13812 7898 13864
rect 8754 13852 8760 13864
rect 7944 13824 8760 13852
rect 7944 13784 7972 13824
rect 8754 13812 8760 13824
rect 8812 13852 8818 13864
rect 9214 13852 9220 13864
rect 8812 13824 9220 13852
rect 8812 13812 8818 13824
rect 9214 13812 9220 13824
rect 9272 13812 9278 13864
rect 10686 13852 10692 13864
rect 10599 13824 10692 13852
rect 10686 13812 10692 13824
rect 10744 13852 10750 13864
rect 11238 13852 11244 13864
rect 10744 13824 11244 13852
rect 10744 13812 10750 13824
rect 11238 13812 11244 13824
rect 11296 13812 11302 13864
rect 12434 13852 12440 13864
rect 12395 13824 12440 13852
rect 12434 13812 12440 13824
rect 12492 13812 12498 13864
rect 12544 13852 12572 13892
rect 15381 13889 15393 13923
rect 15427 13920 15439 13923
rect 15470 13920 15476 13932
rect 15427 13892 15476 13920
rect 15427 13889 15439 13892
rect 15381 13883 15439 13889
rect 15470 13880 15476 13892
rect 15528 13880 15534 13932
rect 15565 13923 15623 13929
rect 15565 13889 15577 13923
rect 15611 13920 15623 13923
rect 15930 13920 15936 13932
rect 15611 13892 15936 13920
rect 15611 13889 15623 13892
rect 15565 13883 15623 13889
rect 15930 13880 15936 13892
rect 15988 13920 15994 13932
rect 16758 13920 16764 13932
rect 15988 13892 16764 13920
rect 15988 13880 15994 13892
rect 16758 13880 16764 13892
rect 16816 13880 16822 13932
rect 24029 13923 24087 13929
rect 24029 13889 24041 13923
rect 24075 13920 24087 13923
rect 24075 13892 24256 13920
rect 24075 13889 24087 13892
rect 24029 13883 24087 13889
rect 12704 13855 12762 13861
rect 12704 13852 12716 13855
rect 12544 13824 12716 13852
rect 12704 13821 12716 13824
rect 12750 13852 12762 13855
rect 13722 13852 13728 13864
rect 12750 13824 13728 13852
rect 12750 13821 12762 13824
rect 12704 13815 12762 13821
rect 13722 13812 13728 13824
rect 13780 13812 13786 13864
rect 17129 13855 17187 13861
rect 17129 13821 17141 13855
rect 17175 13852 17187 13855
rect 17218 13852 17224 13864
rect 17175 13824 17224 13852
rect 17175 13821 17187 13824
rect 17129 13815 17187 13821
rect 17218 13812 17224 13824
rect 17276 13852 17282 13864
rect 18325 13855 18383 13861
rect 17276 13824 17908 13852
rect 17276 13812 17282 13824
rect 11146 13784 11152 13796
rect 7668 13756 7972 13784
rect 11107 13756 11152 13784
rect 11146 13744 11152 13756
rect 11204 13744 11210 13796
rect 14182 13744 14188 13796
rect 14240 13784 14246 13796
rect 14737 13787 14795 13793
rect 14737 13784 14749 13787
rect 14240 13756 14749 13784
rect 14240 13744 14246 13756
rect 14737 13753 14749 13756
rect 14783 13784 14795 13787
rect 15289 13787 15347 13793
rect 15289 13784 15301 13787
rect 14783 13756 15301 13784
rect 14783 13753 14795 13756
rect 14737 13747 14795 13753
rect 15289 13753 15301 13756
rect 15335 13784 15347 13787
rect 16022 13784 16028 13796
rect 15335 13756 16028 13784
rect 15335 13753 15347 13756
rect 15289 13747 15347 13753
rect 16022 13744 16028 13756
rect 16080 13744 16086 13796
rect 17880 13784 17908 13824
rect 18325 13821 18337 13855
rect 18371 13852 18383 13855
rect 18690 13852 18696 13864
rect 18371 13824 18696 13852
rect 18371 13821 18383 13824
rect 18325 13815 18383 13821
rect 18690 13812 18696 13824
rect 18748 13812 18754 13864
rect 24118 13852 24124 13864
rect 24079 13824 24124 13852
rect 24118 13812 24124 13824
rect 24176 13812 24182 13864
rect 24228 13852 24256 13892
rect 24394 13861 24400 13864
rect 24388 13852 24400 13861
rect 24228 13824 24400 13852
rect 24388 13815 24400 13824
rect 24394 13812 24400 13815
rect 24452 13812 24458 13864
rect 18506 13784 18512 13796
rect 17880 13756 18512 13784
rect 18506 13744 18512 13756
rect 18564 13744 18570 13796
rect 3697 13719 3755 13725
rect 3697 13716 3709 13719
rect 3568 13688 3709 13716
rect 3568 13676 3574 13688
rect 3697 13685 3709 13688
rect 3743 13685 3755 13719
rect 4246 13716 4252 13728
rect 4207 13688 4252 13716
rect 3697 13679 3755 13685
rect 4246 13676 4252 13688
rect 4304 13676 4310 13728
rect 10962 13676 10968 13728
rect 11020 13716 11026 13728
rect 11790 13716 11796 13728
rect 11020 13688 11796 13716
rect 11020 13676 11026 13688
rect 11790 13676 11796 13688
rect 11848 13676 11854 13728
rect 13998 13676 14004 13728
rect 14056 13716 14062 13728
rect 14921 13719 14979 13725
rect 14921 13716 14933 13719
rect 14056 13688 14933 13716
rect 14056 13676 14062 13688
rect 14921 13685 14933 13688
rect 14967 13685 14979 13719
rect 14921 13679 14979 13685
rect 17218 13676 17224 13728
rect 17276 13716 17282 13728
rect 17773 13719 17831 13725
rect 17773 13716 17785 13719
rect 17276 13688 17785 13716
rect 17276 13676 17282 13688
rect 17773 13685 17785 13688
rect 17819 13685 17831 13719
rect 17773 13679 17831 13685
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 2406 13512 2412 13524
rect 2367 13484 2412 13512
rect 2406 13472 2412 13484
rect 2464 13472 2470 13524
rect 3513 13515 3571 13521
rect 3513 13481 3525 13515
rect 3559 13512 3571 13515
rect 3786 13512 3792 13524
rect 3559 13484 3792 13512
rect 3559 13481 3571 13484
rect 3513 13475 3571 13481
rect 3786 13472 3792 13484
rect 3844 13472 3850 13524
rect 5534 13512 5540 13524
rect 5495 13484 5540 13512
rect 5534 13472 5540 13484
rect 5592 13472 5598 13524
rect 7101 13515 7159 13521
rect 7101 13481 7113 13515
rect 7147 13512 7159 13515
rect 8018 13512 8024 13524
rect 7147 13484 8024 13512
rect 7147 13481 7159 13484
rect 7101 13475 7159 13481
rect 8018 13472 8024 13484
rect 8076 13472 8082 13524
rect 8294 13472 8300 13524
rect 8352 13512 8358 13524
rect 8573 13515 8631 13521
rect 8573 13512 8585 13515
rect 8352 13484 8585 13512
rect 8352 13472 8358 13484
rect 8573 13481 8585 13484
rect 8619 13512 8631 13515
rect 8849 13515 8907 13521
rect 8849 13512 8861 13515
rect 8619 13484 8861 13512
rect 8619 13481 8631 13484
rect 8573 13475 8631 13481
rect 8849 13481 8861 13484
rect 8895 13481 8907 13515
rect 9214 13512 9220 13524
rect 9175 13484 9220 13512
rect 8849 13475 8907 13481
rect 9214 13472 9220 13484
rect 9272 13472 9278 13524
rect 11514 13472 11520 13524
rect 11572 13512 11578 13524
rect 11609 13515 11667 13521
rect 11609 13512 11621 13515
rect 11572 13484 11621 13512
rect 11572 13472 11578 13484
rect 11609 13481 11621 13484
rect 11655 13481 11667 13515
rect 12066 13512 12072 13524
rect 12027 13484 12072 13512
rect 11609 13475 11667 13481
rect 12066 13472 12072 13484
rect 12124 13512 12130 13524
rect 13262 13512 13268 13524
rect 12124 13484 13268 13512
rect 12124 13472 12130 13484
rect 13262 13472 13268 13484
rect 13320 13472 13326 13524
rect 14274 13512 14280 13524
rect 14235 13484 14280 13512
rect 14274 13472 14280 13484
rect 14332 13472 14338 13524
rect 15013 13515 15071 13521
rect 15013 13481 15025 13515
rect 15059 13512 15071 13515
rect 15470 13512 15476 13524
rect 15059 13484 15476 13512
rect 15059 13481 15071 13484
rect 15013 13475 15071 13481
rect 15470 13472 15476 13484
rect 15528 13472 15534 13524
rect 16666 13512 16672 13524
rect 16627 13484 16672 13512
rect 16666 13472 16672 13484
rect 16724 13472 16730 13524
rect 24118 13512 24124 13524
rect 24079 13484 24124 13512
rect 24118 13472 24124 13484
rect 24176 13472 24182 13524
rect 2777 13447 2835 13453
rect 2777 13413 2789 13447
rect 2823 13444 2835 13447
rect 3970 13444 3976 13456
rect 2823 13416 3976 13444
rect 2823 13413 2835 13416
rect 2777 13407 2835 13413
rect 3970 13404 3976 13416
rect 4028 13444 4034 13456
rect 5077 13447 5135 13453
rect 5077 13444 5089 13447
rect 4028 13416 5089 13444
rect 4028 13404 4034 13416
rect 5077 13413 5089 13416
rect 5123 13413 5135 13447
rect 5077 13407 5135 13413
rect 5350 13404 5356 13456
rect 5408 13444 5414 13456
rect 6273 13447 6331 13453
rect 6273 13444 6285 13447
rect 5408 13416 6285 13444
rect 5408 13404 5414 13416
rect 6273 13413 6285 13416
rect 6319 13413 6331 13447
rect 12158 13444 12164 13456
rect 6273 13407 6331 13413
rect 9692 13416 12164 13444
rect 2038 13376 2044 13388
rect 1999 13348 2044 13376
rect 2038 13336 2044 13348
rect 2096 13336 2102 13388
rect 2869 13379 2927 13385
rect 2869 13345 2881 13379
rect 2915 13376 2927 13379
rect 3789 13379 3847 13385
rect 3789 13376 3801 13379
rect 2915 13348 3801 13376
rect 2915 13345 2927 13348
rect 2869 13339 2927 13345
rect 3789 13345 3801 13348
rect 3835 13345 3847 13379
rect 3789 13339 3847 13345
rect 2958 13308 2964 13320
rect 2919 13280 2964 13308
rect 2958 13268 2964 13280
rect 3016 13268 3022 13320
rect 3804 13240 3832 13339
rect 4246 13336 4252 13388
rect 4304 13376 4310 13388
rect 4433 13379 4491 13385
rect 4433 13376 4445 13379
rect 4304 13348 4445 13376
rect 4304 13336 4310 13348
rect 4433 13345 4445 13348
rect 4479 13345 4491 13379
rect 4433 13339 4491 13345
rect 4522 13336 4528 13388
rect 4580 13376 4586 13388
rect 5626 13376 5632 13388
rect 4580 13348 4625 13376
rect 5587 13348 5632 13376
rect 4580 13336 4586 13348
rect 5626 13336 5632 13348
rect 5684 13376 5690 13388
rect 6178 13376 6184 13388
rect 5684 13348 6184 13376
rect 5684 13336 5690 13348
rect 6178 13336 6184 13348
rect 6236 13336 6242 13388
rect 7098 13336 7104 13388
rect 7156 13376 7162 13388
rect 9692 13385 9720 13416
rect 12158 13404 12164 13416
rect 12216 13444 12222 13456
rect 12434 13444 12440 13456
rect 12216 13416 12440 13444
rect 12216 13404 12222 13416
rect 12434 13404 12440 13416
rect 12492 13404 12498 13456
rect 16482 13444 16488 13456
rect 15304 13416 16488 13444
rect 9950 13385 9956 13388
rect 7469 13379 7527 13385
rect 7469 13376 7481 13379
rect 7156 13348 7481 13376
rect 7156 13336 7162 13348
rect 7469 13345 7481 13348
rect 7515 13345 7527 13379
rect 7469 13339 7527 13345
rect 9677 13379 9735 13385
rect 9677 13345 9689 13379
rect 9723 13345 9735 13379
rect 9944 13376 9956 13385
rect 9911 13348 9956 13376
rect 9677 13339 9735 13345
rect 9944 13339 9956 13348
rect 9950 13336 9956 13339
rect 10008 13336 10014 13388
rect 12802 13376 12808 13388
rect 12763 13348 12808 13376
rect 12802 13336 12808 13348
rect 12860 13336 12866 13388
rect 15304 13385 15332 13416
rect 16482 13404 16488 13416
rect 16540 13404 16546 13456
rect 15562 13385 15568 13388
rect 15289 13379 15347 13385
rect 15289 13345 15301 13379
rect 15335 13345 15347 13379
rect 15556 13376 15568 13385
rect 15523 13348 15568 13376
rect 15289 13339 15347 13345
rect 15556 13339 15568 13348
rect 15562 13336 15568 13339
rect 15620 13336 15626 13388
rect 17494 13336 17500 13388
rect 17552 13376 17558 13388
rect 18141 13379 18199 13385
rect 18141 13376 18153 13379
rect 17552 13348 18153 13376
rect 17552 13336 17558 13348
rect 18141 13345 18153 13348
rect 18187 13345 18199 13379
rect 18141 13339 18199 13345
rect 4614 13308 4620 13320
rect 4575 13280 4620 13308
rect 4614 13268 4620 13280
rect 4672 13268 4678 13320
rect 7558 13308 7564 13320
rect 7519 13280 7564 13308
rect 7558 13268 7564 13280
rect 7616 13268 7622 13320
rect 7650 13268 7656 13320
rect 7708 13308 7714 13320
rect 18230 13308 18236 13320
rect 7708 13280 7753 13308
rect 18191 13280 18236 13308
rect 7708 13268 7714 13280
rect 18230 13268 18236 13280
rect 18288 13268 18294 13320
rect 18322 13268 18328 13320
rect 18380 13308 18386 13320
rect 18380 13280 18425 13308
rect 18380 13268 18386 13280
rect 4065 13243 4123 13249
rect 4065 13240 4077 13243
rect 3804 13212 4077 13240
rect 4065 13209 4077 13212
rect 4111 13209 4123 13243
rect 5810 13240 5816 13252
rect 5771 13212 5816 13240
rect 4065 13203 4123 13209
rect 5810 13200 5816 13212
rect 5868 13200 5874 13252
rect 1673 13175 1731 13181
rect 1673 13141 1685 13175
rect 1719 13172 1731 13175
rect 2314 13172 2320 13184
rect 1719 13144 2320 13172
rect 1719 13141 1731 13144
rect 1673 13135 1731 13141
rect 2314 13132 2320 13144
rect 2372 13132 2378 13184
rect 6546 13172 6552 13184
rect 6507 13144 6552 13172
rect 6546 13132 6552 13144
rect 6604 13132 6610 13184
rect 7009 13175 7067 13181
rect 7009 13141 7021 13175
rect 7055 13172 7067 13175
rect 7098 13172 7104 13184
rect 7055 13144 7104 13172
rect 7055 13141 7067 13144
rect 7009 13135 7067 13141
rect 7098 13132 7104 13144
rect 7156 13132 7162 13184
rect 8110 13172 8116 13184
rect 8071 13144 8116 13172
rect 8110 13132 8116 13144
rect 8168 13132 8174 13184
rect 11054 13172 11060 13184
rect 11015 13144 11060 13172
rect 11054 13132 11060 13144
rect 11112 13132 11118 13184
rect 12434 13132 12440 13184
rect 12492 13172 12498 13184
rect 12492 13144 12537 13172
rect 12492 13132 12498 13144
rect 15286 13132 15292 13184
rect 15344 13172 15350 13184
rect 15654 13172 15660 13184
rect 15344 13144 15660 13172
rect 15344 13132 15350 13144
rect 15654 13132 15660 13144
rect 15712 13132 15718 13184
rect 17218 13172 17224 13184
rect 17179 13144 17224 13172
rect 17218 13132 17224 13144
rect 17276 13172 17282 13184
rect 17589 13175 17647 13181
rect 17589 13172 17601 13175
rect 17276 13144 17601 13172
rect 17276 13132 17282 13144
rect 17589 13141 17601 13144
rect 17635 13141 17647 13175
rect 17589 13135 17647 13141
rect 17773 13175 17831 13181
rect 17773 13141 17785 13175
rect 17819 13172 17831 13175
rect 18782 13172 18788 13184
rect 17819 13144 18788 13172
rect 17819 13141 17831 13144
rect 17773 13135 17831 13141
rect 18782 13132 18788 13144
rect 18840 13132 18846 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1394 12968 1400 12980
rect 1355 12940 1400 12968
rect 1394 12928 1400 12940
rect 1452 12928 1458 12980
rect 2501 12971 2559 12977
rect 2501 12937 2513 12971
rect 2547 12968 2559 12971
rect 2590 12968 2596 12980
rect 2547 12940 2596 12968
rect 2547 12937 2559 12940
rect 2501 12931 2559 12937
rect 2516 12900 2544 12931
rect 2590 12928 2596 12940
rect 2648 12928 2654 12980
rect 2869 12971 2927 12977
rect 2869 12937 2881 12971
rect 2915 12968 2927 12971
rect 2958 12968 2964 12980
rect 2915 12940 2964 12968
rect 2915 12937 2927 12940
rect 2869 12931 2927 12937
rect 2958 12928 2964 12940
rect 3016 12928 3022 12980
rect 4522 12928 4528 12980
rect 4580 12968 4586 12980
rect 5261 12971 5319 12977
rect 5261 12968 5273 12971
rect 4580 12940 5273 12968
rect 4580 12928 4586 12940
rect 5261 12937 5273 12940
rect 5307 12937 5319 12971
rect 6178 12968 6184 12980
rect 6139 12940 6184 12968
rect 5261 12931 5319 12937
rect 6178 12928 6184 12940
rect 6236 12928 6242 12980
rect 6641 12971 6699 12977
rect 6641 12937 6653 12971
rect 6687 12968 6699 12971
rect 7558 12968 7564 12980
rect 6687 12940 7564 12968
rect 6687 12937 6699 12940
rect 6641 12931 6699 12937
rect 7558 12928 7564 12940
rect 7616 12928 7622 12980
rect 7650 12928 7656 12980
rect 7708 12968 7714 12980
rect 9493 12971 9551 12977
rect 9493 12968 9505 12971
rect 7708 12940 9505 12968
rect 7708 12928 7714 12940
rect 9493 12937 9505 12940
rect 9539 12968 9551 12971
rect 9950 12968 9956 12980
rect 9539 12940 9956 12968
rect 9539 12937 9551 12940
rect 9493 12931 9551 12937
rect 9950 12928 9956 12940
rect 10008 12968 10014 12980
rect 10045 12971 10103 12977
rect 10045 12968 10057 12971
rect 10008 12940 10057 12968
rect 10008 12928 10014 12940
rect 10045 12937 10057 12940
rect 10091 12937 10103 12971
rect 10045 12931 10103 12937
rect 12253 12971 12311 12977
rect 12253 12937 12265 12971
rect 12299 12968 12311 12971
rect 12802 12968 12808 12980
rect 12299 12940 12808 12968
rect 12299 12937 12311 12940
rect 12253 12931 12311 12937
rect 12802 12928 12808 12940
rect 12860 12968 12866 12980
rect 13630 12968 13636 12980
rect 12860 12940 13636 12968
rect 12860 12928 12866 12940
rect 13630 12928 13636 12940
rect 13688 12928 13694 12980
rect 13814 12968 13820 12980
rect 13775 12940 13820 12968
rect 13814 12928 13820 12940
rect 13872 12928 13878 12980
rect 17494 12968 17500 12980
rect 17455 12940 17500 12968
rect 17494 12928 17500 12940
rect 17552 12928 17558 12980
rect 17954 12928 17960 12980
rect 18012 12968 18018 12980
rect 18049 12971 18107 12977
rect 18049 12968 18061 12971
rect 18012 12940 18061 12968
rect 18012 12928 18018 12940
rect 18049 12937 18061 12940
rect 18095 12937 18107 12971
rect 18049 12931 18107 12937
rect 1872 12872 2544 12900
rect 1872 12841 1900 12872
rect 12434 12860 12440 12912
rect 12492 12860 12498 12912
rect 1857 12835 1915 12841
rect 1857 12801 1869 12835
rect 1903 12801 1915 12835
rect 1857 12795 1915 12801
rect 2041 12835 2099 12841
rect 2041 12801 2053 12835
rect 2087 12832 2099 12835
rect 5721 12835 5779 12841
rect 2087 12804 2912 12832
rect 2087 12801 2099 12804
rect 2041 12795 2099 12801
rect 1765 12699 1823 12705
rect 1765 12665 1777 12699
rect 1811 12696 1823 12699
rect 2038 12696 2044 12708
rect 1811 12668 2044 12696
rect 1811 12665 1823 12668
rect 1765 12659 1823 12665
rect 2038 12656 2044 12668
rect 2096 12656 2102 12708
rect 2884 12628 2912 12804
rect 5721 12801 5733 12835
rect 5767 12832 5779 12835
rect 6454 12832 6460 12844
rect 5767 12804 6460 12832
rect 5767 12801 5779 12804
rect 5721 12795 5779 12801
rect 6454 12792 6460 12804
rect 6512 12792 6518 12844
rect 7561 12835 7619 12841
rect 7561 12801 7573 12835
rect 7607 12832 7619 12835
rect 7650 12832 7656 12844
rect 7607 12804 7656 12832
rect 7607 12801 7619 12804
rect 7561 12795 7619 12801
rect 7650 12792 7656 12804
rect 7708 12792 7714 12844
rect 8110 12832 8116 12844
rect 8071 12804 8116 12832
rect 8110 12792 8116 12804
rect 8168 12792 8174 12844
rect 11054 12792 11060 12844
rect 11112 12832 11118 12844
rect 11333 12835 11391 12841
rect 11333 12832 11345 12835
rect 11112 12804 11345 12832
rect 11112 12792 11118 12804
rect 11333 12801 11345 12804
rect 11379 12832 11391 12835
rect 12452 12832 12480 12860
rect 16577 12835 16635 12841
rect 11379 12804 12572 12832
rect 11379 12801 11391 12804
rect 11333 12795 11391 12801
rect 2961 12767 3019 12773
rect 2961 12733 2973 12767
rect 3007 12764 3019 12767
rect 3050 12764 3056 12776
rect 3007 12736 3056 12764
rect 3007 12733 3019 12736
rect 2961 12727 3019 12733
rect 3050 12724 3056 12736
rect 3108 12764 3114 12776
rect 4154 12764 4160 12776
rect 3108 12736 4160 12764
rect 3108 12724 3114 12736
rect 4154 12724 4160 12736
rect 4212 12764 4218 12776
rect 5442 12764 5448 12776
rect 4212 12736 5448 12764
rect 4212 12724 4218 12736
rect 5442 12724 5448 12736
rect 5500 12724 5506 12776
rect 10870 12724 10876 12776
rect 10928 12764 10934 12776
rect 11241 12767 11299 12773
rect 11241 12764 11253 12767
rect 10928 12736 11253 12764
rect 10928 12724 10934 12736
rect 11241 12733 11253 12736
rect 11287 12733 11299 12767
rect 11241 12727 11299 12733
rect 12158 12724 12164 12776
rect 12216 12764 12222 12776
rect 12437 12767 12495 12773
rect 12437 12764 12449 12767
rect 12216 12736 12449 12764
rect 12216 12724 12222 12736
rect 12437 12733 12449 12736
rect 12483 12733 12495 12767
rect 12544 12764 12572 12804
rect 16577 12801 16589 12835
rect 16623 12832 16635 12835
rect 17512 12832 17540 12928
rect 18598 12832 18604 12844
rect 16623 12804 17540 12832
rect 18559 12804 18604 12832
rect 16623 12801 16635 12804
rect 16577 12795 16635 12801
rect 18598 12792 18604 12804
rect 18656 12792 18662 12844
rect 12693 12767 12751 12773
rect 12693 12764 12705 12767
rect 12544 12736 12705 12764
rect 12437 12727 12495 12733
rect 12693 12733 12705 12736
rect 12739 12733 12751 12767
rect 12693 12727 12751 12733
rect 14185 12767 14243 12773
rect 14185 12733 14197 12767
rect 14231 12764 14243 12767
rect 15746 12764 15752 12776
rect 14231 12736 15752 12764
rect 14231 12733 14243 12736
rect 14185 12727 14243 12733
rect 3217 12699 3275 12705
rect 3217 12665 3229 12699
rect 3263 12696 3275 12699
rect 8018 12696 8024 12708
rect 3263 12665 3280 12696
rect 7931 12668 8024 12696
rect 3217 12659 3280 12665
rect 3252 12628 3280 12659
rect 8018 12656 8024 12668
rect 8076 12696 8082 12708
rect 8358 12699 8416 12705
rect 8358 12696 8370 12699
rect 8076 12668 8370 12696
rect 8076 12656 8082 12668
rect 8358 12665 8370 12668
rect 8404 12665 8416 12699
rect 8358 12659 8416 12665
rect 10689 12699 10747 12705
rect 10689 12665 10701 12699
rect 10735 12696 10747 12699
rect 10962 12696 10968 12708
rect 10735 12668 10968 12696
rect 10735 12665 10747 12668
rect 10689 12659 10747 12665
rect 10962 12656 10968 12668
rect 11020 12696 11026 12708
rect 11149 12699 11207 12705
rect 11149 12696 11161 12699
rect 11020 12668 11161 12696
rect 11020 12656 11026 12668
rect 11149 12665 11161 12668
rect 11195 12665 11207 12699
rect 12452 12696 12480 12727
rect 14200 12696 14228 12727
rect 15746 12724 15752 12736
rect 15804 12764 15810 12776
rect 17218 12764 17224 12776
rect 15804 12736 17224 12764
rect 15804 12724 15810 12736
rect 17218 12724 17224 12736
rect 17276 12724 17282 12776
rect 18417 12767 18475 12773
rect 18417 12733 18429 12767
rect 18463 12764 18475 12767
rect 18782 12764 18788 12776
rect 18463 12736 18788 12764
rect 18463 12733 18475 12736
rect 18417 12727 18475 12733
rect 18782 12724 18788 12736
rect 18840 12724 18846 12776
rect 12452 12668 14228 12696
rect 14452 12699 14510 12705
rect 11149 12659 11207 12665
rect 14452 12665 14464 12699
rect 14498 12696 14510 12699
rect 14642 12696 14648 12708
rect 14498 12668 14648 12696
rect 14498 12665 14510 12668
rect 14452 12659 14510 12665
rect 14642 12656 14648 12668
rect 14700 12656 14706 12708
rect 16758 12656 16764 12708
rect 16816 12696 16822 12708
rect 17773 12699 17831 12705
rect 17773 12696 17785 12699
rect 16816 12668 17785 12696
rect 16816 12656 16822 12668
rect 17773 12665 17785 12668
rect 17819 12696 17831 12699
rect 18230 12696 18236 12708
rect 17819 12668 18236 12696
rect 17819 12665 17831 12668
rect 17773 12659 17831 12665
rect 18230 12656 18236 12668
rect 18288 12656 18294 12708
rect 3510 12628 3516 12640
rect 2884 12600 3516 12628
rect 3510 12588 3516 12600
rect 3568 12588 3574 12640
rect 4338 12628 4344 12640
rect 4299 12600 4344 12628
rect 4338 12588 4344 12600
rect 4396 12628 4402 12640
rect 4614 12628 4620 12640
rect 4396 12600 4620 12628
rect 4396 12588 4402 12600
rect 4614 12588 4620 12600
rect 4672 12628 4678 12640
rect 4893 12631 4951 12637
rect 4893 12628 4905 12631
rect 4672 12600 4905 12628
rect 4672 12588 4678 12600
rect 4893 12597 4905 12600
rect 4939 12597 4951 12631
rect 7006 12628 7012 12640
rect 6967 12600 7012 12628
rect 4893 12591 4951 12597
rect 7006 12588 7012 12600
rect 7064 12588 7070 12640
rect 10781 12631 10839 12637
rect 10781 12597 10793 12631
rect 10827 12628 10839 12631
rect 11054 12628 11060 12640
rect 10827 12600 11060 12628
rect 10827 12597 10839 12600
rect 10781 12591 10839 12597
rect 11054 12588 11060 12600
rect 11112 12588 11118 12640
rect 11882 12628 11888 12640
rect 11843 12600 11888 12628
rect 11882 12588 11888 12600
rect 11940 12588 11946 12640
rect 13262 12588 13268 12640
rect 13320 12628 13326 12640
rect 15010 12628 15016 12640
rect 13320 12600 15016 12628
rect 13320 12588 13326 12600
rect 15010 12588 15016 12600
rect 15068 12588 15074 12640
rect 15194 12588 15200 12640
rect 15252 12628 15258 12640
rect 15562 12628 15568 12640
rect 15252 12600 15568 12628
rect 15252 12588 15258 12600
rect 15562 12588 15568 12600
rect 15620 12628 15626 12640
rect 16117 12631 16175 12637
rect 16117 12628 16129 12631
rect 15620 12600 16129 12628
rect 15620 12588 15626 12600
rect 16117 12597 16129 12600
rect 16163 12597 16175 12631
rect 16117 12591 16175 12597
rect 16850 12588 16856 12640
rect 16908 12628 16914 12640
rect 17037 12631 17095 12637
rect 17037 12628 17049 12631
rect 16908 12600 17049 12628
rect 16908 12588 16914 12600
rect 17037 12597 17049 12600
rect 17083 12628 17095 12631
rect 17862 12628 17868 12640
rect 17083 12600 17868 12628
rect 17083 12597 17095 12600
rect 17037 12591 17095 12597
rect 17862 12588 17868 12600
rect 17920 12628 17926 12640
rect 18322 12628 18328 12640
rect 17920 12600 18328 12628
rect 17920 12588 17926 12600
rect 18322 12588 18328 12600
rect 18380 12588 18386 12640
rect 18414 12588 18420 12640
rect 18472 12628 18478 12640
rect 18509 12631 18567 12637
rect 18509 12628 18521 12631
rect 18472 12600 18521 12628
rect 18472 12588 18478 12600
rect 18509 12597 18521 12600
rect 18555 12628 18567 12631
rect 19061 12631 19119 12637
rect 19061 12628 19073 12631
rect 18555 12600 19073 12628
rect 18555 12597 18567 12600
rect 18509 12591 18567 12597
rect 19061 12597 19073 12600
rect 19107 12597 19119 12631
rect 19061 12591 19119 12597
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 2866 12424 2872 12436
rect 2827 12396 2872 12424
rect 2866 12384 2872 12396
rect 2924 12384 2930 12436
rect 3970 12384 3976 12436
rect 4028 12424 4034 12436
rect 4065 12427 4123 12433
rect 4065 12424 4077 12427
rect 4028 12396 4077 12424
rect 4028 12384 4034 12396
rect 4065 12393 4077 12396
rect 4111 12393 4123 12427
rect 5442 12424 5448 12436
rect 5403 12396 5448 12424
rect 4065 12387 4123 12393
rect 5442 12384 5448 12396
rect 5500 12424 5506 12436
rect 6086 12424 6092 12436
rect 5500 12396 6092 12424
rect 5500 12384 5506 12396
rect 6086 12384 6092 12396
rect 6144 12424 6150 12436
rect 6457 12427 6515 12433
rect 6457 12424 6469 12427
rect 6144 12396 6469 12424
rect 6144 12384 6150 12396
rect 6457 12393 6469 12396
rect 6503 12424 6515 12427
rect 6546 12424 6552 12436
rect 6503 12396 6552 12424
rect 6503 12393 6515 12396
rect 6457 12387 6515 12393
rect 6546 12384 6552 12396
rect 6604 12384 6610 12436
rect 7009 12427 7067 12433
rect 7009 12393 7021 12427
rect 7055 12424 7067 12427
rect 7098 12424 7104 12436
rect 7055 12396 7104 12424
rect 7055 12393 7067 12396
rect 7009 12387 7067 12393
rect 7098 12384 7104 12396
rect 7156 12384 7162 12436
rect 9674 12424 9680 12436
rect 9635 12396 9680 12424
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 11146 12424 11152 12436
rect 11107 12396 11152 12424
rect 11146 12384 11152 12396
rect 11204 12384 11210 12436
rect 11333 12427 11391 12433
rect 11333 12393 11345 12427
rect 11379 12424 11391 12427
rect 11514 12424 11520 12436
rect 11379 12396 11520 12424
rect 11379 12393 11391 12396
rect 11333 12387 11391 12393
rect 11514 12384 11520 12396
rect 11572 12384 11578 12436
rect 12894 12424 12900 12436
rect 12855 12396 12900 12424
rect 12894 12384 12900 12396
rect 12952 12384 12958 12436
rect 13538 12384 13544 12436
rect 13596 12424 13602 12436
rect 13633 12427 13691 12433
rect 13633 12424 13645 12427
rect 13596 12396 13645 12424
rect 13596 12384 13602 12396
rect 13633 12393 13645 12396
rect 13679 12393 13691 12427
rect 13633 12387 13691 12393
rect 13998 12384 14004 12436
rect 14056 12424 14062 12436
rect 14642 12424 14648 12436
rect 14056 12396 14412 12424
rect 14603 12396 14648 12424
rect 14056 12384 14062 12396
rect 2038 12356 2044 12368
rect 1504 12328 2044 12356
rect 1504 12297 1532 12328
rect 2038 12316 2044 12328
rect 2096 12356 2102 12368
rect 3050 12356 3056 12368
rect 2096 12328 3056 12356
rect 2096 12316 2102 12328
rect 3050 12316 3056 12328
rect 3108 12316 3114 12368
rect 3326 12316 3332 12368
rect 3384 12356 3390 12368
rect 8846 12356 8852 12368
rect 3384 12328 8852 12356
rect 3384 12316 3390 12328
rect 8846 12316 8852 12328
rect 8904 12316 8910 12368
rect 12805 12359 12863 12365
rect 12805 12325 12817 12359
rect 12851 12356 12863 12359
rect 14016 12356 14044 12384
rect 12851 12328 14044 12356
rect 12851 12325 12863 12328
rect 12805 12319 12863 12325
rect 1762 12297 1768 12300
rect 1489 12291 1547 12297
rect 1489 12257 1501 12291
rect 1535 12257 1547 12291
rect 1489 12251 1547 12257
rect 1756 12251 1768 12297
rect 1820 12288 1826 12300
rect 3881 12291 3939 12297
rect 1820 12260 1856 12288
rect 1762 12248 1768 12251
rect 1820 12248 1826 12260
rect 3881 12257 3893 12291
rect 3927 12288 3939 12291
rect 4246 12288 4252 12300
rect 3927 12260 4252 12288
rect 3927 12257 3939 12260
rect 3881 12251 3939 12257
rect 4246 12248 4252 12260
rect 4304 12248 4310 12300
rect 4430 12288 4436 12300
rect 4343 12260 4436 12288
rect 4430 12248 4436 12260
rect 4488 12288 4494 12300
rect 5077 12291 5135 12297
rect 5077 12288 5089 12291
rect 4488 12260 5089 12288
rect 4488 12248 4494 12260
rect 5077 12257 5089 12260
rect 5123 12257 5135 12291
rect 5077 12251 5135 12257
rect 7006 12248 7012 12300
rect 7064 12288 7070 12300
rect 7374 12288 7380 12300
rect 7064 12260 7380 12288
rect 7064 12248 7070 12260
rect 7374 12248 7380 12260
rect 7432 12248 7438 12300
rect 10042 12288 10048 12300
rect 10003 12260 10048 12288
rect 10042 12248 10048 12260
rect 10100 12248 10106 12300
rect 11701 12291 11759 12297
rect 11701 12257 11713 12291
rect 11747 12288 11759 12291
rect 12066 12288 12072 12300
rect 11747 12260 12072 12288
rect 11747 12257 11759 12260
rect 11701 12251 11759 12257
rect 12066 12248 12072 12260
rect 12124 12248 12130 12300
rect 13998 12288 14004 12300
rect 13959 12260 14004 12288
rect 13998 12248 14004 12260
rect 14056 12248 14062 12300
rect 14384 12232 14412 12396
rect 14642 12384 14648 12396
rect 14700 12384 14706 12436
rect 15010 12424 15016 12436
rect 14971 12396 15016 12424
rect 15010 12384 15016 12396
rect 15068 12384 15074 12436
rect 15746 12424 15752 12436
rect 15707 12396 15752 12424
rect 15746 12384 15752 12396
rect 15804 12384 15810 12436
rect 17957 12427 18015 12433
rect 17957 12393 17969 12427
rect 18003 12424 18015 12427
rect 18598 12424 18604 12436
rect 18003 12396 18604 12424
rect 18003 12393 18015 12396
rect 17957 12387 18015 12393
rect 18598 12384 18604 12396
rect 18656 12384 18662 12436
rect 15028 12288 15056 12384
rect 18506 12356 18512 12368
rect 16592 12328 18512 12356
rect 16592 12300 16620 12328
rect 18506 12316 18512 12328
rect 18564 12356 18570 12368
rect 18877 12359 18935 12365
rect 18877 12356 18889 12359
rect 18564 12328 18889 12356
rect 18564 12316 18570 12328
rect 18877 12325 18889 12328
rect 18923 12325 18935 12359
rect 18877 12319 18935 12325
rect 15746 12288 15752 12300
rect 15028 12260 15752 12288
rect 15746 12248 15752 12260
rect 15804 12248 15810 12300
rect 16574 12288 16580 12300
rect 16535 12260 16580 12288
rect 16574 12248 16580 12260
rect 16632 12248 16638 12300
rect 16850 12297 16856 12300
rect 16844 12288 16856 12297
rect 16811 12260 16856 12288
rect 16844 12251 16856 12260
rect 16850 12248 16856 12251
rect 16908 12248 16914 12300
rect 4522 12220 4528 12232
rect 4483 12192 4528 12220
rect 4522 12180 4528 12192
rect 4580 12180 4586 12232
rect 4617 12223 4675 12229
rect 4617 12189 4629 12223
rect 4663 12189 4675 12223
rect 4617 12183 4675 12189
rect 3786 12112 3792 12164
rect 3844 12152 3850 12164
rect 4338 12152 4344 12164
rect 3844 12124 4344 12152
rect 3844 12112 3850 12124
rect 4338 12112 4344 12124
rect 4396 12152 4402 12164
rect 4632 12152 4660 12183
rect 4890 12180 4896 12232
rect 4948 12220 4954 12232
rect 5629 12223 5687 12229
rect 5629 12220 5641 12223
rect 4948 12192 5641 12220
rect 4948 12180 4954 12192
rect 5629 12189 5641 12192
rect 5675 12189 5687 12223
rect 5629 12183 5687 12189
rect 7190 12180 7196 12232
rect 7248 12220 7254 12232
rect 7469 12223 7527 12229
rect 7469 12220 7481 12223
rect 7248 12192 7481 12220
rect 7248 12180 7254 12192
rect 7469 12189 7481 12192
rect 7515 12189 7527 12223
rect 7469 12183 7527 12189
rect 7561 12223 7619 12229
rect 7561 12189 7573 12223
rect 7607 12220 7619 12223
rect 8018 12220 8024 12232
rect 7607 12192 8024 12220
rect 7607 12189 7619 12192
rect 7561 12183 7619 12189
rect 4396 12124 4660 12152
rect 4396 12112 4402 12124
rect 6270 12112 6276 12164
rect 6328 12152 6334 12164
rect 7576 12152 7604 12183
rect 8018 12180 8024 12192
rect 8076 12180 8082 12232
rect 9674 12180 9680 12232
rect 9732 12220 9738 12232
rect 10137 12223 10195 12229
rect 10137 12220 10149 12223
rect 9732 12192 10149 12220
rect 9732 12180 9738 12192
rect 10137 12189 10149 12192
rect 10183 12189 10195 12223
rect 10137 12183 10195 12189
rect 10321 12223 10379 12229
rect 10321 12189 10333 12223
rect 10367 12220 10379 12223
rect 10778 12220 10784 12232
rect 10367 12192 10784 12220
rect 10367 12189 10379 12192
rect 10321 12183 10379 12189
rect 6328 12124 7604 12152
rect 9493 12155 9551 12161
rect 6328 12112 6334 12124
rect 9493 12121 9505 12155
rect 9539 12152 9551 12155
rect 10336 12152 10364 12183
rect 10778 12180 10784 12192
rect 10836 12180 10842 12232
rect 11054 12180 11060 12232
rect 11112 12220 11118 12232
rect 11238 12220 11244 12232
rect 11112 12192 11244 12220
rect 11112 12180 11118 12192
rect 11238 12180 11244 12192
rect 11296 12220 11302 12232
rect 11793 12223 11851 12229
rect 11793 12220 11805 12223
rect 11296 12192 11805 12220
rect 11296 12180 11302 12192
rect 11793 12189 11805 12192
rect 11839 12189 11851 12223
rect 11974 12220 11980 12232
rect 11935 12192 11980 12220
rect 11793 12183 11851 12189
rect 11974 12180 11980 12192
rect 12032 12180 12038 12232
rect 13081 12223 13139 12229
rect 13081 12189 13093 12223
rect 13127 12220 13139 12223
rect 13265 12223 13323 12229
rect 13265 12220 13277 12223
rect 13127 12192 13277 12220
rect 13127 12189 13139 12192
rect 13081 12183 13139 12189
rect 13265 12189 13277 12192
rect 13311 12189 13323 12223
rect 13265 12183 13323 12189
rect 14093 12223 14151 12229
rect 14093 12189 14105 12223
rect 14139 12189 14151 12223
rect 14274 12220 14280 12232
rect 14235 12192 14280 12220
rect 14093 12183 14151 12189
rect 9539 12124 10364 12152
rect 12437 12155 12495 12161
rect 9539 12121 9551 12124
rect 9493 12115 9551 12121
rect 12437 12121 12449 12155
rect 12483 12152 12495 12155
rect 14108 12152 14136 12183
rect 14274 12180 14280 12192
rect 14332 12180 14338 12232
rect 14366 12180 14372 12232
rect 14424 12180 14430 12232
rect 14734 12180 14740 12232
rect 14792 12220 14798 12232
rect 15289 12223 15347 12229
rect 15289 12220 15301 12223
rect 14792 12192 15301 12220
rect 14792 12180 14798 12192
rect 15289 12189 15301 12192
rect 15335 12189 15347 12223
rect 15289 12183 15347 12189
rect 12483 12124 14872 12152
rect 12483 12121 12495 12124
rect 12437 12115 12495 12121
rect 14844 12096 14872 12124
rect 3510 12084 3516 12096
rect 3423 12056 3516 12084
rect 3510 12044 3516 12056
rect 3568 12084 3574 12096
rect 5074 12084 5080 12096
rect 3568 12056 5080 12084
rect 3568 12044 3574 12056
rect 5074 12044 5080 12056
rect 5132 12044 5138 12096
rect 6546 12044 6552 12096
rect 6604 12084 6610 12096
rect 6825 12087 6883 12093
rect 6825 12084 6837 12087
rect 6604 12056 6837 12084
rect 6604 12044 6610 12056
rect 6825 12053 6837 12056
rect 6871 12053 6883 12087
rect 6825 12047 6883 12053
rect 7834 12044 7840 12096
rect 7892 12084 7898 12096
rect 8021 12087 8079 12093
rect 8021 12084 8033 12087
rect 7892 12056 8033 12084
rect 7892 12044 7898 12056
rect 8021 12053 8033 12056
rect 8067 12053 8079 12087
rect 8021 12047 8079 12053
rect 8110 12044 8116 12096
rect 8168 12084 8174 12096
rect 8386 12084 8392 12096
rect 8168 12056 8392 12084
rect 8168 12044 8174 12056
rect 8386 12044 8392 12056
rect 8444 12084 8450 12096
rect 8757 12087 8815 12093
rect 8757 12084 8769 12087
rect 8444 12056 8769 12084
rect 8444 12044 8450 12056
rect 8757 12053 8769 12056
rect 8803 12053 8815 12087
rect 10870 12084 10876 12096
rect 10831 12056 10876 12084
rect 8757 12047 8815 12053
rect 10870 12044 10876 12056
rect 10928 12044 10934 12096
rect 13170 12044 13176 12096
rect 13228 12084 13234 12096
rect 13265 12087 13323 12093
rect 13265 12084 13277 12087
rect 13228 12056 13277 12084
rect 13228 12044 13234 12056
rect 13265 12053 13277 12056
rect 13311 12084 13323 12087
rect 13541 12087 13599 12093
rect 13541 12084 13553 12087
rect 13311 12056 13553 12084
rect 13311 12053 13323 12056
rect 13265 12047 13323 12053
rect 13541 12053 13553 12056
rect 13587 12084 13599 12087
rect 14642 12084 14648 12096
rect 13587 12056 14648 12084
rect 13587 12053 13599 12056
rect 13541 12047 13599 12053
rect 14642 12044 14648 12056
rect 14700 12044 14706 12096
rect 14826 12044 14832 12096
rect 14884 12044 14890 12096
rect 16209 12087 16267 12093
rect 16209 12053 16221 12087
rect 16255 12084 16267 12087
rect 16298 12084 16304 12096
rect 16255 12056 16304 12084
rect 16255 12053 16267 12056
rect 16209 12047 16267 12053
rect 16298 12044 16304 12056
rect 16356 12044 16362 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 3421 11883 3479 11889
rect 3421 11849 3433 11883
rect 3467 11880 3479 11883
rect 3510 11880 3516 11892
rect 3467 11852 3516 11880
rect 3467 11849 3479 11852
rect 3421 11843 3479 11849
rect 3510 11840 3516 11852
rect 3568 11840 3574 11892
rect 4430 11840 4436 11892
rect 4488 11880 4494 11892
rect 4525 11883 4583 11889
rect 4525 11880 4537 11883
rect 4488 11852 4537 11880
rect 4488 11840 4494 11852
rect 4525 11849 4537 11852
rect 4571 11849 4583 11883
rect 6270 11880 6276 11892
rect 6231 11852 6276 11880
rect 4525 11843 4583 11849
rect 6270 11840 6276 11852
rect 6328 11840 6334 11892
rect 6641 11883 6699 11889
rect 6641 11849 6653 11883
rect 6687 11880 6699 11883
rect 7374 11880 7380 11892
rect 6687 11852 7380 11880
rect 6687 11849 6699 11852
rect 6641 11843 6699 11849
rect 7374 11840 7380 11852
rect 7432 11840 7438 11892
rect 8110 11840 8116 11892
rect 8168 11880 8174 11892
rect 8570 11880 8576 11892
rect 8168 11852 8576 11880
rect 8168 11840 8174 11852
rect 8570 11840 8576 11852
rect 8628 11880 8634 11892
rect 8849 11883 8907 11889
rect 8849 11880 8861 11883
rect 8628 11852 8861 11880
rect 8628 11840 8634 11852
rect 8849 11849 8861 11852
rect 8895 11849 8907 11883
rect 9674 11880 9680 11892
rect 9635 11852 9680 11880
rect 8849 11843 8907 11849
rect 9674 11840 9680 11852
rect 9732 11840 9738 11892
rect 11974 11840 11980 11892
rect 12032 11880 12038 11892
rect 12069 11883 12127 11889
rect 12069 11880 12081 11883
rect 12032 11852 12081 11880
rect 12032 11840 12038 11852
rect 12069 11849 12081 11852
rect 12115 11849 12127 11883
rect 12069 11843 12127 11849
rect 13173 11883 13231 11889
rect 13173 11849 13185 11883
rect 13219 11880 13231 11883
rect 14274 11880 14280 11892
rect 13219 11852 14280 11880
rect 13219 11849 13231 11852
rect 13173 11843 13231 11849
rect 14274 11840 14280 11852
rect 14332 11840 14338 11892
rect 14642 11880 14648 11892
rect 14603 11852 14648 11880
rect 14642 11840 14648 11852
rect 14700 11840 14706 11892
rect 14826 11840 14832 11892
rect 14884 11880 14890 11892
rect 15197 11883 15255 11889
rect 15197 11880 15209 11883
rect 14884 11852 15209 11880
rect 14884 11840 14890 11852
rect 15197 11849 15209 11852
rect 15243 11849 15255 11883
rect 16114 11880 16120 11892
rect 16075 11852 16120 11880
rect 15197 11843 15255 11849
rect 16114 11840 16120 11852
rect 16172 11840 16178 11892
rect 18506 11880 18512 11892
rect 18467 11852 18512 11880
rect 18506 11840 18512 11852
rect 18564 11840 18570 11892
rect 4982 11772 4988 11824
rect 5040 11812 5046 11824
rect 7009 11815 7067 11821
rect 7009 11812 7021 11815
rect 5040 11784 7021 11812
rect 5040 11772 5046 11784
rect 7009 11781 7021 11784
rect 7055 11812 7067 11815
rect 7190 11812 7196 11824
rect 7055 11784 7196 11812
rect 7055 11781 7067 11784
rect 7009 11775 7067 11781
rect 7190 11772 7196 11784
rect 7248 11772 7254 11824
rect 14292 11812 14320 11840
rect 15286 11812 15292 11824
rect 14292 11784 15292 11812
rect 15286 11772 15292 11784
rect 15344 11772 15350 11824
rect 4338 11704 4344 11756
rect 4396 11744 4402 11756
rect 4433 11747 4491 11753
rect 4433 11744 4445 11747
rect 4396 11716 4445 11744
rect 4396 11704 4402 11716
rect 4433 11713 4445 11716
rect 4479 11744 4491 11747
rect 4614 11744 4620 11756
rect 4479 11716 4620 11744
rect 4479 11713 4491 11716
rect 4433 11707 4491 11713
rect 4614 11704 4620 11716
rect 4672 11704 4678 11756
rect 5074 11744 5080 11756
rect 5035 11716 5080 11744
rect 5074 11704 5080 11716
rect 5132 11744 5138 11756
rect 5537 11747 5595 11753
rect 5537 11744 5549 11747
rect 5132 11716 5549 11744
rect 5132 11704 5138 11716
rect 5537 11713 5549 11716
rect 5583 11713 5595 11747
rect 5537 11707 5595 11713
rect 9490 11704 9496 11756
rect 9548 11744 9554 11756
rect 10505 11747 10563 11753
rect 10505 11744 10517 11747
rect 9548 11716 10517 11744
rect 9548 11704 9554 11716
rect 10505 11713 10517 11716
rect 10551 11713 10563 11747
rect 10505 11707 10563 11713
rect 13262 11704 13268 11756
rect 13320 11753 13326 11756
rect 13320 11744 13330 11753
rect 15657 11747 15715 11753
rect 13320 11716 13365 11744
rect 13320 11707 13330 11716
rect 15657 11713 15669 11747
rect 15703 11744 15715 11747
rect 16669 11747 16727 11753
rect 16669 11744 16681 11747
rect 15703 11716 16681 11744
rect 15703 11713 15715 11716
rect 15657 11707 15715 11713
rect 16669 11713 16681 11716
rect 16715 11744 16727 11747
rect 16850 11744 16856 11756
rect 16715 11716 16856 11744
rect 16715 11713 16727 11716
rect 16669 11707 16727 11713
rect 13320 11704 13326 11707
rect 16850 11704 16856 11716
rect 16908 11744 16914 11756
rect 17129 11747 17187 11753
rect 17129 11744 17141 11747
rect 16908 11716 17141 11744
rect 16908 11704 16914 11716
rect 17129 11713 17141 11716
rect 17175 11713 17187 11747
rect 17129 11707 17187 11713
rect 2038 11676 2044 11688
rect 1999 11648 2044 11676
rect 2038 11636 2044 11648
rect 2096 11636 2102 11688
rect 4065 11679 4123 11685
rect 4065 11645 4077 11679
rect 4111 11676 4123 11679
rect 4890 11676 4896 11688
rect 4111 11648 4896 11676
rect 4111 11645 4123 11648
rect 4065 11639 4123 11645
rect 4890 11636 4896 11648
rect 4948 11636 4954 11688
rect 7374 11636 7380 11688
rect 7432 11676 7438 11688
rect 7469 11679 7527 11685
rect 7469 11676 7481 11679
rect 7432 11648 7481 11676
rect 7432 11636 7438 11648
rect 7469 11645 7481 11648
rect 7515 11645 7527 11679
rect 7469 11639 7527 11645
rect 10042 11636 10048 11688
rect 10100 11676 10106 11688
rect 10965 11679 11023 11685
rect 10965 11676 10977 11679
rect 10100 11648 10977 11676
rect 10100 11636 10106 11648
rect 10965 11645 10977 11648
rect 11011 11645 11023 11679
rect 10965 11639 11023 11645
rect 11425 11679 11483 11685
rect 11425 11645 11437 11679
rect 11471 11676 11483 11679
rect 12066 11676 12072 11688
rect 11471 11648 12072 11676
rect 11471 11645 11483 11648
rect 11425 11639 11483 11645
rect 12066 11636 12072 11648
rect 12124 11636 12130 11688
rect 1949 11611 2007 11617
rect 1949 11577 1961 11611
rect 1995 11608 2007 11611
rect 2308 11611 2366 11617
rect 2308 11608 2320 11611
rect 1995 11580 2320 11608
rect 1995 11577 2007 11580
rect 1949 11571 2007 11577
rect 2308 11577 2320 11580
rect 2354 11608 2366 11611
rect 2406 11608 2412 11620
rect 2354 11580 2412 11608
rect 2354 11577 2366 11580
rect 2308 11571 2366 11577
rect 2406 11568 2412 11580
rect 2464 11568 2470 11620
rect 4614 11568 4620 11620
rect 4672 11608 4678 11620
rect 4985 11611 5043 11617
rect 4985 11608 4997 11611
rect 4672 11580 4997 11608
rect 4672 11568 4678 11580
rect 4985 11577 4997 11580
rect 5031 11577 5043 11611
rect 4985 11571 5043 11577
rect 7736 11611 7794 11617
rect 7736 11577 7748 11611
rect 7782 11608 7794 11611
rect 7834 11608 7840 11620
rect 7782 11580 7840 11608
rect 7782 11577 7794 11580
rect 7736 11571 7794 11577
rect 7834 11568 7840 11580
rect 7892 11568 7898 11620
rect 9858 11568 9864 11620
rect 9916 11608 9922 11620
rect 10413 11611 10471 11617
rect 10413 11608 10425 11611
rect 9916 11580 10425 11608
rect 9916 11568 9922 11580
rect 10413 11577 10425 11580
rect 10459 11608 10471 11611
rect 10459 11580 11836 11608
rect 10459 11577 10471 11580
rect 10413 11571 10471 11577
rect 1394 11500 1400 11552
rect 1452 11540 1458 11552
rect 7282 11540 7288 11552
rect 1452 11512 7288 11540
rect 1452 11500 1458 11512
rect 7282 11500 7288 11512
rect 7340 11500 7346 11552
rect 9306 11500 9312 11552
rect 9364 11540 9370 11552
rect 9953 11543 10011 11549
rect 9953 11540 9965 11543
rect 9364 11512 9965 11540
rect 9364 11500 9370 11512
rect 9953 11509 9965 11512
rect 9999 11509 10011 11543
rect 9953 11503 10011 11509
rect 10321 11543 10379 11549
rect 10321 11509 10333 11543
rect 10367 11540 10379 11543
rect 10686 11540 10692 11552
rect 10367 11512 10692 11540
rect 10367 11509 10379 11512
rect 10321 11503 10379 11509
rect 10686 11500 10692 11512
rect 10744 11500 10750 11552
rect 11808 11549 11836 11580
rect 12342 11568 12348 11620
rect 12400 11608 12406 11620
rect 13538 11617 13544 11620
rect 12805 11611 12863 11617
rect 12805 11608 12817 11611
rect 12400 11580 12817 11608
rect 12400 11568 12406 11580
rect 12805 11577 12817 11580
rect 12851 11608 12863 11611
rect 13532 11608 13544 11617
rect 12851 11580 13544 11608
rect 12851 11577 12863 11580
rect 12805 11571 12863 11577
rect 13532 11571 13544 11580
rect 13538 11568 13544 11571
rect 13596 11568 13602 11620
rect 15930 11608 15936 11620
rect 15891 11580 15936 11608
rect 15930 11568 15936 11580
rect 15988 11608 15994 11620
rect 16390 11608 16396 11620
rect 15988 11580 16396 11608
rect 15988 11568 15994 11580
rect 16390 11568 16396 11580
rect 16448 11608 16454 11620
rect 16485 11611 16543 11617
rect 16485 11608 16497 11611
rect 16448 11580 16497 11608
rect 16448 11568 16454 11580
rect 16485 11577 16497 11580
rect 16531 11577 16543 11611
rect 16485 11571 16543 11577
rect 17681 11611 17739 11617
rect 17681 11577 17693 11611
rect 17727 11608 17739 11611
rect 17954 11608 17960 11620
rect 17727 11580 17960 11608
rect 17727 11577 17739 11580
rect 17681 11571 17739 11577
rect 17954 11568 17960 11580
rect 18012 11568 18018 11620
rect 11793 11543 11851 11549
rect 11793 11509 11805 11543
rect 11839 11540 11851 11543
rect 11882 11540 11888 11552
rect 11839 11512 11888 11540
rect 11839 11509 11851 11512
rect 11793 11503 11851 11509
rect 11882 11500 11888 11512
rect 11940 11500 11946 11552
rect 13630 11500 13636 11552
rect 13688 11540 13694 11552
rect 13906 11540 13912 11552
rect 13688 11512 13912 11540
rect 13688 11500 13694 11512
rect 13906 11500 13912 11512
rect 13964 11500 13970 11552
rect 16298 11500 16304 11552
rect 16356 11540 16362 11552
rect 16577 11543 16635 11549
rect 16577 11540 16589 11543
rect 16356 11512 16589 11540
rect 16356 11500 16362 11512
rect 16577 11509 16589 11512
rect 16623 11509 16635 11543
rect 18046 11540 18052 11552
rect 18007 11512 18052 11540
rect 16577 11503 16635 11509
rect 18046 11500 18052 11512
rect 18104 11500 18110 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1762 11296 1768 11348
rect 1820 11336 1826 11348
rect 1949 11339 2007 11345
rect 1949 11336 1961 11339
rect 1820 11308 1961 11336
rect 1820 11296 1826 11308
rect 1949 11305 1961 11308
rect 1995 11336 2007 11339
rect 3786 11336 3792 11348
rect 1995 11308 3792 11336
rect 1995 11305 2007 11308
rect 1949 11299 2007 11305
rect 3786 11296 3792 11308
rect 3844 11296 3850 11348
rect 4065 11339 4123 11345
rect 4065 11305 4077 11339
rect 4111 11336 4123 11339
rect 4522 11336 4528 11348
rect 4111 11308 4528 11336
rect 4111 11305 4123 11308
rect 4065 11299 4123 11305
rect 4522 11296 4528 11308
rect 4580 11336 4586 11348
rect 5077 11339 5135 11345
rect 5077 11336 5089 11339
rect 4580 11308 5089 11336
rect 4580 11296 4586 11308
rect 5077 11305 5089 11308
rect 5123 11305 5135 11339
rect 6086 11336 6092 11348
rect 6047 11308 6092 11336
rect 5077 11299 5135 11305
rect 6086 11296 6092 11308
rect 6144 11296 6150 11348
rect 7834 11336 7840 11348
rect 7747 11308 7840 11336
rect 7834 11296 7840 11308
rect 7892 11336 7898 11348
rect 9490 11336 9496 11348
rect 7892 11308 9496 11336
rect 7892 11296 7898 11308
rect 9490 11296 9496 11308
rect 9548 11296 9554 11348
rect 11238 11336 11244 11348
rect 11199 11308 11244 11336
rect 11238 11296 11244 11308
rect 11296 11296 11302 11348
rect 12710 11336 12716 11348
rect 12671 11308 12716 11336
rect 12710 11296 12716 11308
rect 12768 11296 12774 11348
rect 13170 11336 13176 11348
rect 13131 11308 13176 11336
rect 13170 11296 13176 11308
rect 13228 11296 13234 11348
rect 13265 11339 13323 11345
rect 13265 11305 13277 11339
rect 13311 11336 13323 11339
rect 13998 11336 14004 11348
rect 13311 11308 14004 11336
rect 13311 11305 13323 11308
rect 13265 11299 13323 11305
rect 13998 11296 14004 11308
rect 14056 11336 14062 11348
rect 15013 11339 15071 11345
rect 15013 11336 15025 11339
rect 14056 11308 15025 11336
rect 14056 11296 14062 11308
rect 15013 11305 15025 11308
rect 15059 11305 15071 11339
rect 15013 11299 15071 11305
rect 15473 11339 15531 11345
rect 15473 11305 15485 11339
rect 15519 11336 15531 11339
rect 15746 11336 15752 11348
rect 15519 11308 15752 11336
rect 15519 11305 15531 11308
rect 15473 11299 15531 11305
rect 15746 11296 15752 11308
rect 15804 11296 15810 11348
rect 16390 11336 16396 11348
rect 16351 11308 16396 11336
rect 16390 11296 16396 11308
rect 16448 11296 16454 11348
rect 16666 11296 16672 11348
rect 16724 11336 16730 11348
rect 17129 11339 17187 11345
rect 17129 11336 17141 11339
rect 16724 11308 17141 11336
rect 16724 11296 16730 11308
rect 17129 11305 17141 11308
rect 17175 11336 17187 11339
rect 18046 11336 18052 11348
rect 17175 11308 18052 11336
rect 17175 11305 17187 11308
rect 17129 11299 17187 11305
rect 18046 11296 18052 11308
rect 18104 11296 18110 11348
rect 1673 11271 1731 11277
rect 1673 11237 1685 11271
rect 1719 11268 1731 11271
rect 3510 11268 3516 11280
rect 1719 11240 3516 11268
rect 1719 11237 1731 11240
rect 1673 11231 1731 11237
rect 3510 11228 3516 11240
rect 3568 11228 3574 11280
rect 6638 11228 6644 11280
rect 6696 11277 6702 11280
rect 6696 11271 6760 11277
rect 6696 11237 6714 11271
rect 6748 11237 6760 11271
rect 6696 11231 6760 11237
rect 6696 11228 6702 11231
rect 7374 11228 7380 11280
rect 7432 11228 7438 11280
rect 9122 11228 9128 11280
rect 9180 11268 9186 11280
rect 9858 11268 9864 11280
rect 9180 11240 9864 11268
rect 9180 11228 9186 11240
rect 9858 11228 9864 11240
rect 9916 11268 9922 11280
rect 10137 11271 10195 11277
rect 10137 11268 10149 11271
rect 9916 11240 10149 11268
rect 9916 11228 9922 11240
rect 10137 11237 10149 11240
rect 10183 11237 10195 11271
rect 10137 11231 10195 11237
rect 10686 11228 10692 11280
rect 10744 11268 10750 11280
rect 10781 11271 10839 11277
rect 10781 11268 10793 11271
rect 10744 11240 10793 11268
rect 10744 11228 10750 11240
rect 10781 11237 10793 11240
rect 10827 11268 10839 11271
rect 10870 11268 10876 11280
rect 10827 11240 10876 11268
rect 10827 11237 10839 11240
rect 10781 11231 10839 11237
rect 10870 11228 10876 11240
rect 10928 11268 10934 11280
rect 12526 11268 12532 11280
rect 10928 11240 12532 11268
rect 10928 11228 10934 11240
rect 12526 11228 12532 11240
rect 12584 11228 12590 11280
rect 13354 11228 13360 11280
rect 13412 11268 13418 11280
rect 14366 11268 14372 11280
rect 13412 11240 14228 11268
rect 14327 11240 14372 11268
rect 13412 11228 13418 11240
rect 1486 11160 1492 11212
rect 1544 11200 1550 11212
rect 1854 11200 1860 11212
rect 1544 11172 1860 11200
rect 1544 11160 1550 11172
rect 1854 11160 1860 11172
rect 1912 11160 1918 11212
rect 2777 11203 2835 11209
rect 2777 11169 2789 11203
rect 2823 11200 2835 11203
rect 3234 11200 3240 11212
rect 2823 11172 3240 11200
rect 2823 11169 2835 11172
rect 2777 11163 2835 11169
rect 3234 11160 3240 11172
rect 3292 11200 3298 11212
rect 4433 11203 4491 11209
rect 4433 11200 4445 11203
rect 3292 11172 4445 11200
rect 3292 11160 3298 11172
rect 4433 11169 4445 11172
rect 4479 11200 4491 11203
rect 4798 11200 4804 11212
rect 4479 11172 4804 11200
rect 4479 11169 4491 11172
rect 4433 11163 4491 11169
rect 4798 11160 4804 11172
rect 4856 11200 4862 11212
rect 5442 11200 5448 11212
rect 4856 11172 5448 11200
rect 4856 11160 4862 11172
rect 5442 11160 5448 11172
rect 5500 11160 5506 11212
rect 6457 11203 6515 11209
rect 6457 11169 6469 11203
rect 6503 11200 6515 11203
rect 6546 11200 6552 11212
rect 6503 11172 6552 11200
rect 6503 11169 6515 11172
rect 6457 11163 6515 11169
rect 6546 11160 6552 11172
rect 6604 11200 6610 11212
rect 7392 11200 7420 11228
rect 8386 11200 8392 11212
rect 6604 11172 8392 11200
rect 6604 11160 6610 11172
rect 8386 11160 8392 11172
rect 8444 11200 8450 11212
rect 8757 11203 8815 11209
rect 8757 11200 8769 11203
rect 8444 11172 8769 11200
rect 8444 11160 8450 11172
rect 8757 11169 8769 11172
rect 8803 11169 8815 11203
rect 10042 11200 10048 11212
rect 10003 11172 10048 11200
rect 8757 11163 8815 11169
rect 10042 11160 10048 11172
rect 10100 11160 10106 11212
rect 11606 11160 11612 11212
rect 11664 11200 11670 11212
rect 12069 11203 12127 11209
rect 12069 11200 12081 11203
rect 11664 11172 12081 11200
rect 11664 11160 11670 11172
rect 12069 11169 12081 11172
rect 12115 11169 12127 11203
rect 12069 11163 12127 11169
rect 13633 11203 13691 11209
rect 13633 11169 13645 11203
rect 13679 11200 13691 11203
rect 13998 11200 14004 11212
rect 13679 11172 14004 11200
rect 13679 11169 13691 11172
rect 13633 11163 13691 11169
rect 13998 11160 14004 11172
rect 14056 11160 14062 11212
rect 14200 11200 14228 11240
rect 14366 11228 14372 11240
rect 14424 11228 14430 11280
rect 15562 11228 15568 11280
rect 15620 11268 15626 11280
rect 15620 11240 17356 11268
rect 15620 11228 15626 11240
rect 17126 11200 17132 11212
rect 14200 11172 17132 11200
rect 17126 11160 17132 11172
rect 17184 11160 17190 11212
rect 17328 11200 17356 11240
rect 17402 11228 17408 11280
rect 17460 11268 17466 11280
rect 17460 11240 18184 11268
rect 17460 11228 17466 11240
rect 17678 11200 17684 11212
rect 17328 11172 17684 11200
rect 17678 11160 17684 11172
rect 17736 11200 17742 11212
rect 17957 11203 18015 11209
rect 17957 11200 17969 11203
rect 17736 11172 17969 11200
rect 17736 11160 17742 11172
rect 17957 11169 17969 11172
rect 18003 11169 18015 11203
rect 17957 11163 18015 11169
rect 2869 11135 2927 11141
rect 2869 11101 2881 11135
rect 2915 11101 2927 11135
rect 2869 11095 2927 11101
rect 3053 11135 3111 11141
rect 3053 11101 3065 11135
rect 3099 11132 3111 11135
rect 4525 11135 4583 11141
rect 3099 11104 3556 11132
rect 3099 11101 3111 11104
rect 3053 11095 3111 11101
rect 2130 11024 2136 11076
rect 2188 11064 2194 11076
rect 2409 11067 2467 11073
rect 2409 11064 2421 11067
rect 2188 11036 2421 11064
rect 2188 11024 2194 11036
rect 2409 11033 2421 11036
rect 2455 11033 2467 11067
rect 2409 11027 2467 11033
rect 2774 11024 2780 11076
rect 2832 11064 2838 11076
rect 2884 11064 2912 11095
rect 3528 11073 3556 11104
rect 4525 11101 4537 11135
rect 4571 11101 4583 11135
rect 4525 11095 4583 11101
rect 4709 11135 4767 11141
rect 4709 11101 4721 11135
rect 4755 11132 4767 11135
rect 5074 11132 5080 11144
rect 4755 11104 5080 11132
rect 4755 11101 4767 11104
rect 4709 11095 4767 11101
rect 3513 11067 3571 11073
rect 2832 11036 3464 11064
rect 2832 11024 2838 11036
rect 3436 10996 3464 11036
rect 3513 11033 3525 11067
rect 3559 11064 3571 11067
rect 3878 11064 3884 11076
rect 3559 11036 3884 11064
rect 3559 11033 3571 11036
rect 3513 11027 3571 11033
rect 3878 11024 3884 11036
rect 3936 11024 3942 11076
rect 4540 11064 4568 11095
rect 5074 11092 5080 11104
rect 5132 11092 5138 11144
rect 10318 11132 10324 11144
rect 10279 11104 10324 11132
rect 10318 11092 10324 11104
rect 10376 11092 10382 11144
rect 12158 11132 12164 11144
rect 12119 11104 12164 11132
rect 12158 11092 12164 11104
rect 12216 11092 12222 11144
rect 12342 11132 12348 11144
rect 12303 11104 12348 11132
rect 12342 11092 12348 11104
rect 12400 11092 12406 11144
rect 13722 11132 13728 11144
rect 13096 11104 13728 11132
rect 4890 11064 4896 11076
rect 3988 11036 4896 11064
rect 3988 10996 4016 11036
rect 4890 11024 4896 11036
rect 4948 11064 4954 11076
rect 5166 11064 5172 11076
rect 4948 11036 5172 11064
rect 4948 11024 4954 11036
rect 5166 11024 5172 11036
rect 5224 11024 5230 11076
rect 8202 11024 8208 11076
rect 8260 11064 8266 11076
rect 9677 11067 9735 11073
rect 9677 11064 9689 11067
rect 8260 11036 9689 11064
rect 8260 11024 8266 11036
rect 9677 11033 9689 11036
rect 9723 11033 9735 11067
rect 9677 11027 9735 11033
rect 11609 11067 11667 11073
rect 11609 11033 11621 11067
rect 11655 11064 11667 11067
rect 12360 11064 12388 11092
rect 11655 11036 12388 11064
rect 11655 11033 11667 11036
rect 11609 11027 11667 11033
rect 3436 10968 4016 10996
rect 5534 10956 5540 11008
rect 5592 10996 5598 11008
rect 5629 10999 5687 11005
rect 5629 10996 5641 10999
rect 5592 10968 5641 10996
rect 5592 10956 5598 10968
rect 5629 10965 5641 10968
rect 5675 10965 5687 10999
rect 5629 10959 5687 10965
rect 6086 10956 6092 11008
rect 6144 10996 6150 11008
rect 8386 10996 8392 11008
rect 6144 10968 8392 10996
rect 6144 10956 6150 10968
rect 8386 10956 8392 10968
rect 8444 10956 8450 11008
rect 11701 10999 11759 11005
rect 11701 10965 11713 10999
rect 11747 10996 11759 10999
rect 13096 10996 13124 11104
rect 13722 11092 13728 11104
rect 13780 11092 13786 11144
rect 13817 11135 13875 11141
rect 13817 11101 13829 11135
rect 13863 11101 13875 11135
rect 13817 11095 13875 11101
rect 13170 11024 13176 11076
rect 13228 11064 13234 11076
rect 13832 11064 13860 11095
rect 15286 11092 15292 11144
rect 15344 11132 15350 11144
rect 16298 11132 16304 11144
rect 15344 11104 16304 11132
rect 15344 11092 15350 11104
rect 16298 11092 16304 11104
rect 16356 11132 16362 11144
rect 16485 11135 16543 11141
rect 16485 11132 16497 11135
rect 16356 11104 16497 11132
rect 16356 11092 16362 11104
rect 16485 11101 16497 11104
rect 16531 11101 16543 11135
rect 16485 11095 16543 11101
rect 16577 11135 16635 11141
rect 16577 11101 16589 11135
rect 16623 11101 16635 11135
rect 18046 11132 18052 11144
rect 18007 11104 18052 11132
rect 16577 11095 16635 11101
rect 13228 11036 13860 11064
rect 13228 11024 13234 11036
rect 15562 11024 15568 11076
rect 15620 11064 15626 11076
rect 16025 11067 16083 11073
rect 16025 11064 16037 11067
rect 15620 11036 16037 11064
rect 15620 11024 15626 11036
rect 16025 11033 16037 11036
rect 16071 11033 16083 11067
rect 16592 11064 16620 11095
rect 18046 11092 18052 11104
rect 18104 11092 18110 11144
rect 18156 11141 18184 11240
rect 18141 11135 18199 11141
rect 18141 11101 18153 11135
rect 18187 11132 18199 11135
rect 18598 11132 18604 11144
rect 18187 11104 18604 11132
rect 18187 11101 18199 11104
rect 18141 11095 18199 11101
rect 18598 11092 18604 11104
rect 18656 11092 18662 11144
rect 17402 11064 17408 11076
rect 16025 11027 16083 11033
rect 16500 11036 16620 11064
rect 17363 11036 17408 11064
rect 14642 10996 14648 11008
rect 11747 10968 13124 10996
rect 14603 10968 14648 10996
rect 11747 10965 11759 10968
rect 11701 10959 11759 10965
rect 14642 10956 14648 10968
rect 14700 10956 14706 11008
rect 15838 10996 15844 11008
rect 15799 10968 15844 10996
rect 15838 10956 15844 10968
rect 15896 10996 15902 11008
rect 16500 10996 16528 11036
rect 17402 11024 17408 11036
rect 17460 11024 17466 11076
rect 17589 11067 17647 11073
rect 17589 11033 17601 11067
rect 17635 11064 17647 11067
rect 17635 11036 17908 11064
rect 17635 11033 17647 11036
rect 17589 11027 17647 11033
rect 15896 10968 16528 10996
rect 17880 10996 17908 11036
rect 18506 10996 18512 11008
rect 17880 10968 18512 10996
rect 15896 10956 15902 10968
rect 18506 10956 18512 10968
rect 18564 10956 18570 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 2682 10792 2688 10804
rect 2643 10764 2688 10792
rect 2682 10752 2688 10764
rect 2740 10752 2746 10804
rect 5166 10792 5172 10804
rect 5127 10764 5172 10792
rect 5166 10752 5172 10764
rect 5224 10752 5230 10804
rect 5442 10752 5448 10804
rect 5500 10792 5506 10804
rect 5537 10795 5595 10801
rect 5537 10792 5549 10795
rect 5500 10764 5549 10792
rect 5500 10752 5506 10764
rect 5537 10761 5549 10764
rect 5583 10761 5595 10795
rect 5537 10755 5595 10761
rect 7558 10752 7564 10804
rect 7616 10792 7622 10804
rect 8021 10795 8079 10801
rect 8021 10792 8033 10795
rect 7616 10764 8033 10792
rect 7616 10752 7622 10764
rect 8021 10761 8033 10764
rect 8067 10761 8079 10795
rect 8021 10755 8079 10761
rect 9217 10795 9275 10801
rect 9217 10761 9229 10795
rect 9263 10792 9275 10795
rect 10318 10792 10324 10804
rect 9263 10764 10324 10792
rect 9263 10761 9275 10764
rect 9217 10755 9275 10761
rect 10318 10752 10324 10764
rect 10376 10792 10382 10804
rect 10686 10792 10692 10804
rect 10376 10764 10692 10792
rect 10376 10752 10382 10764
rect 10686 10752 10692 10764
rect 10744 10792 10750 10804
rect 11057 10795 11115 10801
rect 11057 10792 11069 10795
rect 10744 10764 11069 10792
rect 10744 10752 10750 10764
rect 11057 10761 11069 10764
rect 11103 10761 11115 10795
rect 11057 10755 11115 10761
rect 11606 10752 11612 10804
rect 11664 10792 11670 10804
rect 11701 10795 11759 10801
rect 11701 10792 11713 10795
rect 11664 10764 11713 10792
rect 11664 10752 11670 10764
rect 11701 10761 11713 10764
rect 11747 10761 11759 10795
rect 11701 10755 11759 10761
rect 11974 10752 11980 10804
rect 12032 10792 12038 10804
rect 12161 10795 12219 10801
rect 12161 10792 12173 10795
rect 12032 10764 12173 10792
rect 12032 10752 12038 10764
rect 12161 10761 12173 10764
rect 12207 10761 12219 10795
rect 13998 10792 14004 10804
rect 13911 10764 14004 10792
rect 12161 10755 12219 10761
rect 13998 10752 14004 10764
rect 14056 10792 14062 10804
rect 14642 10792 14648 10804
rect 14056 10764 14648 10792
rect 14056 10752 14062 10764
rect 14642 10752 14648 10764
rect 14700 10752 14706 10804
rect 16117 10795 16175 10801
rect 16117 10761 16129 10795
rect 16163 10792 16175 10795
rect 16390 10792 16396 10804
rect 16163 10764 16396 10792
rect 16163 10761 16175 10764
rect 16117 10755 16175 10761
rect 16390 10752 16396 10764
rect 16448 10752 16454 10804
rect 17678 10792 17684 10804
rect 17639 10764 17684 10792
rect 17678 10752 17684 10764
rect 17736 10752 17742 10804
rect 5810 10724 5816 10736
rect 5771 10696 5816 10724
rect 5810 10684 5816 10696
rect 5868 10684 5874 10736
rect 13906 10724 13912 10736
rect 13867 10696 13912 10724
rect 13906 10684 13912 10696
rect 13964 10684 13970 10736
rect 2222 10656 2228 10668
rect 2183 10628 2228 10656
rect 2222 10616 2228 10628
rect 2280 10616 2286 10668
rect 8570 10656 8576 10668
rect 8531 10628 8576 10656
rect 8570 10616 8576 10628
rect 8628 10616 8634 10668
rect 9585 10659 9643 10665
rect 9585 10625 9597 10659
rect 9631 10656 9643 10659
rect 9631 10628 9812 10656
rect 9631 10625 9643 10628
rect 9585 10619 9643 10625
rect 2038 10548 2044 10600
rect 2096 10588 2102 10600
rect 2774 10588 2780 10600
rect 2096 10560 2780 10588
rect 2096 10548 2102 10560
rect 2774 10548 2780 10560
rect 2832 10588 2838 10600
rect 3145 10591 3203 10597
rect 3145 10588 3157 10591
rect 2832 10560 3157 10588
rect 2832 10548 2838 10560
rect 3145 10557 3157 10560
rect 3191 10557 3203 10591
rect 3145 10551 3203 10557
rect 5534 10548 5540 10600
rect 5592 10588 5598 10600
rect 5629 10591 5687 10597
rect 5629 10588 5641 10591
rect 5592 10560 5641 10588
rect 5592 10548 5598 10560
rect 5629 10557 5641 10560
rect 5675 10557 5687 10591
rect 5629 10551 5687 10557
rect 7561 10591 7619 10597
rect 7561 10557 7573 10591
rect 7607 10588 7619 10591
rect 8481 10591 8539 10597
rect 8481 10588 8493 10591
rect 7607 10560 8493 10588
rect 7607 10557 7619 10560
rect 7561 10551 7619 10557
rect 8481 10557 8493 10560
rect 8527 10588 8539 10591
rect 9306 10588 9312 10600
rect 8527 10560 9312 10588
rect 8527 10557 8539 10560
rect 8481 10551 8539 10557
rect 9306 10548 9312 10560
rect 9364 10548 9370 10600
rect 9677 10591 9735 10597
rect 9677 10557 9689 10591
rect 9723 10557 9735 10591
rect 9784 10588 9812 10628
rect 12710 10616 12716 10668
rect 12768 10656 12774 10668
rect 12897 10659 12955 10665
rect 12897 10656 12909 10659
rect 12768 10628 12909 10656
rect 12768 10616 12774 10628
rect 12897 10625 12909 10628
rect 12943 10625 12955 10659
rect 12897 10619 12955 10625
rect 12986 10616 12992 10668
rect 13044 10656 13050 10668
rect 13538 10656 13544 10668
rect 13044 10628 13089 10656
rect 13451 10628 13544 10656
rect 13044 10616 13050 10628
rect 13538 10616 13544 10628
rect 13596 10656 13602 10668
rect 14550 10656 14556 10668
rect 13596 10628 14556 10656
rect 13596 10616 13602 10628
rect 14550 10616 14556 10628
rect 14608 10616 14614 10668
rect 15749 10659 15807 10665
rect 15749 10625 15761 10659
rect 15795 10656 15807 10659
rect 16758 10656 16764 10668
rect 15795 10628 16764 10656
rect 15795 10625 15807 10628
rect 15749 10619 15807 10625
rect 16758 10616 16764 10628
rect 16816 10616 16822 10668
rect 16942 10656 16948 10668
rect 16903 10628 16948 10656
rect 16942 10616 16948 10628
rect 17000 10616 17006 10668
rect 18598 10656 18604 10668
rect 18559 10628 18604 10656
rect 18598 10616 18604 10628
rect 18656 10616 18662 10668
rect 9950 10597 9956 10600
rect 9933 10591 9956 10597
rect 9933 10588 9945 10591
rect 9784 10560 9945 10588
rect 9677 10551 9735 10557
rect 9933 10557 9945 10560
rect 9933 10551 9956 10557
rect 2866 10480 2872 10532
rect 2924 10520 2930 10532
rect 3418 10529 3424 10532
rect 3390 10523 3424 10529
rect 3390 10520 3402 10523
rect 2924 10492 3402 10520
rect 2924 10480 2930 10492
rect 3390 10489 3402 10492
rect 3476 10520 3482 10532
rect 6822 10520 6828 10532
rect 3476 10492 3538 10520
rect 6783 10492 6828 10520
rect 3390 10483 3424 10489
rect 3418 10480 3424 10483
rect 3476 10480 3482 10492
rect 6822 10480 6828 10492
rect 6880 10480 6886 10532
rect 9692 10520 9720 10551
rect 9950 10548 9956 10551
rect 10008 10548 10014 10600
rect 14090 10548 14096 10600
rect 14148 10588 14154 10600
rect 14369 10591 14427 10597
rect 14369 10588 14381 10591
rect 14148 10560 14381 10588
rect 14148 10548 14154 10560
rect 14369 10557 14381 10560
rect 14415 10588 14427 10591
rect 14734 10588 14740 10600
rect 14415 10560 14740 10588
rect 14415 10557 14427 10560
rect 14369 10551 14427 10557
rect 14734 10548 14740 10560
rect 14792 10548 14798 10600
rect 16666 10588 16672 10600
rect 16627 10560 16672 10588
rect 16666 10548 16672 10560
rect 16724 10548 16730 10600
rect 18046 10548 18052 10600
rect 18104 10588 18110 10600
rect 18509 10591 18567 10597
rect 18509 10588 18521 10591
rect 18104 10560 18521 10588
rect 18104 10548 18110 10560
rect 18509 10557 18521 10560
rect 18555 10557 18567 10591
rect 18509 10551 18567 10557
rect 10134 10520 10140 10532
rect 9692 10492 10140 10520
rect 10134 10480 10140 10492
rect 10192 10480 10198 10532
rect 11974 10480 11980 10532
rect 12032 10520 12038 10532
rect 12805 10523 12863 10529
rect 12805 10520 12817 10523
rect 12032 10492 12817 10520
rect 12032 10480 12038 10492
rect 12805 10489 12817 10492
rect 12851 10489 12863 10523
rect 12805 10483 12863 10489
rect 13906 10480 13912 10532
rect 13964 10520 13970 10532
rect 14461 10523 14519 10529
rect 14461 10520 14473 10523
rect 13964 10492 14473 10520
rect 13964 10480 13970 10492
rect 14461 10489 14473 10492
rect 14507 10489 14519 10523
rect 15470 10520 15476 10532
rect 14461 10483 14519 10489
rect 14660 10492 15476 10520
rect 1578 10452 1584 10464
rect 1539 10424 1584 10452
rect 1578 10412 1584 10424
rect 1636 10412 1642 10464
rect 1854 10412 1860 10464
rect 1912 10452 1918 10464
rect 1949 10455 2007 10461
rect 1949 10452 1961 10455
rect 1912 10424 1961 10452
rect 1912 10412 1918 10424
rect 1949 10421 1961 10424
rect 1995 10421 2007 10455
rect 1949 10415 2007 10421
rect 2038 10412 2044 10464
rect 2096 10452 2102 10464
rect 3053 10455 3111 10461
rect 2096 10424 2141 10452
rect 2096 10412 2102 10424
rect 3053 10421 3065 10455
rect 3099 10452 3111 10455
rect 3234 10452 3240 10464
rect 3099 10424 3240 10452
rect 3099 10421 3111 10424
rect 3053 10415 3111 10421
rect 3234 10412 3240 10424
rect 3292 10412 3298 10464
rect 4430 10412 4436 10464
rect 4488 10452 4494 10464
rect 4525 10455 4583 10461
rect 4525 10452 4537 10455
rect 4488 10424 4537 10452
rect 4488 10412 4494 10424
rect 4525 10421 4537 10424
rect 4571 10421 4583 10455
rect 4525 10415 4583 10421
rect 6549 10455 6607 10461
rect 6549 10421 6561 10455
rect 6595 10452 6607 10455
rect 6638 10452 6644 10464
rect 6595 10424 6644 10452
rect 6595 10421 6607 10424
rect 6549 10415 6607 10421
rect 6638 10412 6644 10424
rect 6696 10452 6702 10464
rect 7098 10452 7104 10464
rect 6696 10424 7104 10452
rect 6696 10412 6702 10424
rect 7098 10412 7104 10424
rect 7156 10412 7162 10464
rect 7929 10455 7987 10461
rect 7929 10421 7941 10455
rect 7975 10452 7987 10455
rect 8389 10455 8447 10461
rect 8389 10452 8401 10455
rect 7975 10424 8401 10452
rect 7975 10421 7987 10424
rect 7929 10415 7987 10421
rect 8389 10421 8401 10424
rect 8435 10452 8447 10455
rect 8938 10452 8944 10464
rect 8435 10424 8944 10452
rect 8435 10421 8447 10424
rect 8389 10415 8447 10421
rect 8938 10412 8944 10424
rect 8996 10412 9002 10464
rect 12434 10412 12440 10464
rect 12492 10452 12498 10464
rect 12492 10424 12537 10452
rect 12492 10412 12498 10424
rect 12710 10412 12716 10464
rect 12768 10452 12774 10464
rect 14660 10452 14688 10492
rect 15470 10480 15476 10492
rect 15528 10480 15534 10532
rect 18414 10520 18420 10532
rect 18375 10492 18420 10520
rect 18414 10480 18420 10492
rect 18472 10520 18478 10532
rect 19061 10523 19119 10529
rect 19061 10520 19073 10523
rect 18472 10492 19073 10520
rect 18472 10480 18478 10492
rect 19061 10489 19073 10492
rect 19107 10489 19119 10523
rect 19061 10483 19119 10489
rect 12768 10424 14688 10452
rect 12768 10412 12774 10424
rect 14734 10412 14740 10464
rect 14792 10452 14798 10464
rect 15286 10452 15292 10464
rect 14792 10424 15292 10452
rect 14792 10412 14798 10424
rect 15286 10412 15292 10424
rect 15344 10412 15350 10464
rect 16298 10452 16304 10464
rect 16259 10424 16304 10452
rect 16298 10412 16304 10424
rect 16356 10412 16362 10464
rect 17954 10412 17960 10464
rect 18012 10452 18018 10464
rect 18049 10455 18107 10461
rect 18049 10452 18061 10455
rect 18012 10424 18061 10452
rect 18012 10412 18018 10424
rect 18049 10421 18061 10424
rect 18095 10421 18107 10455
rect 18049 10415 18107 10421
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 3418 10248 3424 10260
rect 3379 10220 3424 10248
rect 3418 10208 3424 10220
rect 3476 10208 3482 10260
rect 3510 10208 3516 10260
rect 3568 10248 3574 10260
rect 3789 10251 3847 10257
rect 3789 10248 3801 10251
rect 3568 10220 3801 10248
rect 3568 10208 3574 10220
rect 3789 10217 3801 10220
rect 3835 10217 3847 10251
rect 3789 10211 3847 10217
rect 5537 10251 5595 10257
rect 5537 10217 5549 10251
rect 5583 10248 5595 10251
rect 5626 10248 5632 10260
rect 5583 10220 5632 10248
rect 5583 10217 5595 10220
rect 5537 10211 5595 10217
rect 5626 10208 5632 10220
rect 5684 10208 5690 10260
rect 7745 10251 7803 10257
rect 7745 10217 7757 10251
rect 7791 10248 7803 10251
rect 8202 10248 8208 10260
rect 7791 10220 8208 10248
rect 7791 10217 7803 10220
rect 7745 10211 7803 10217
rect 8202 10208 8208 10220
rect 8260 10208 8266 10260
rect 9858 10248 9864 10260
rect 9819 10220 9864 10248
rect 9858 10208 9864 10220
rect 9916 10208 9922 10260
rect 10042 10208 10048 10260
rect 10100 10248 10106 10260
rect 10229 10251 10287 10257
rect 10229 10248 10241 10251
rect 10100 10220 10241 10248
rect 10100 10208 10106 10220
rect 10229 10217 10241 10220
rect 10275 10217 10287 10251
rect 10229 10211 10287 10217
rect 12434 10208 12440 10260
rect 12492 10248 12498 10260
rect 13078 10248 13084 10260
rect 12492 10220 13084 10248
rect 12492 10208 12498 10220
rect 13078 10208 13084 10220
rect 13136 10248 13142 10260
rect 13449 10251 13507 10257
rect 13449 10248 13461 10251
rect 13136 10220 13461 10248
rect 13136 10208 13142 10220
rect 13449 10217 13461 10220
rect 13495 10217 13507 10251
rect 13449 10211 13507 10217
rect 13722 10208 13728 10260
rect 13780 10208 13786 10260
rect 14090 10248 14096 10260
rect 14051 10220 14096 10248
rect 14090 10208 14096 10220
rect 14148 10208 14154 10260
rect 14829 10251 14887 10257
rect 14829 10217 14841 10251
rect 14875 10248 14887 10251
rect 15286 10248 15292 10260
rect 14875 10220 15292 10248
rect 14875 10217 14887 10220
rect 14829 10211 14887 10217
rect 15286 10208 15292 10220
rect 15344 10248 15350 10260
rect 15746 10248 15752 10260
rect 15344 10220 15752 10248
rect 15344 10208 15350 10220
rect 15746 10208 15752 10220
rect 15804 10208 15810 10260
rect 17954 10208 17960 10260
rect 18012 10248 18018 10260
rect 18785 10251 18843 10257
rect 18785 10248 18797 10251
rect 18012 10220 18797 10248
rect 18012 10208 18018 10220
rect 18785 10217 18797 10220
rect 18831 10217 18843 10251
rect 18785 10211 18843 10217
rect 2590 10140 2596 10192
rect 2648 10180 2654 10192
rect 2869 10183 2927 10189
rect 2869 10180 2881 10183
rect 2648 10152 2881 10180
rect 2648 10140 2654 10152
rect 2869 10149 2881 10152
rect 2915 10180 2927 10183
rect 3326 10180 3332 10192
rect 2915 10152 3332 10180
rect 2915 10149 2927 10152
rect 2869 10143 2927 10149
rect 3326 10140 3332 10152
rect 3384 10140 3390 10192
rect 5988 10183 6046 10189
rect 5988 10149 6000 10183
rect 6034 10180 6046 10183
rect 6086 10180 6092 10192
rect 6034 10152 6092 10180
rect 6034 10149 6046 10152
rect 5988 10143 6046 10149
rect 6086 10140 6092 10152
rect 6144 10140 6150 10192
rect 8113 10183 8171 10189
rect 8113 10149 8125 10183
rect 8159 10180 8171 10183
rect 8570 10180 8576 10192
rect 8159 10152 8576 10180
rect 8159 10149 8171 10152
rect 8113 10143 8171 10149
rect 8570 10140 8576 10152
rect 8628 10140 8634 10192
rect 9217 10183 9275 10189
rect 9217 10149 9229 10183
rect 9263 10180 9275 10183
rect 9950 10180 9956 10192
rect 9263 10152 9956 10180
rect 9263 10149 9275 10152
rect 9217 10143 9275 10149
rect 9950 10140 9956 10152
rect 10008 10140 10014 10192
rect 10686 10140 10692 10192
rect 10744 10189 10750 10192
rect 10744 10183 10808 10189
rect 10744 10149 10762 10183
rect 10796 10149 10808 10183
rect 13740 10180 13768 10208
rect 14369 10183 14427 10189
rect 14369 10180 14381 10183
rect 13740 10152 14381 10180
rect 10744 10143 10808 10149
rect 14369 10149 14381 10152
rect 14415 10149 14427 10183
rect 14369 10143 14427 10149
rect 10744 10140 10750 10143
rect 17126 10140 17132 10192
rect 17184 10180 17190 10192
rect 18046 10180 18052 10192
rect 17184 10152 18052 10180
rect 17184 10140 17190 10152
rect 18046 10140 18052 10152
rect 18104 10140 18110 10192
rect 18506 10140 18512 10192
rect 18564 10180 18570 10192
rect 18877 10183 18935 10189
rect 18877 10180 18889 10183
rect 18564 10152 18889 10180
rect 18564 10140 18570 10152
rect 18877 10149 18889 10152
rect 18923 10180 18935 10183
rect 19334 10180 19340 10192
rect 18923 10152 19340 10180
rect 18923 10149 18935 10152
rect 18877 10143 18935 10149
rect 19334 10140 19340 10152
rect 19392 10140 19398 10192
rect 2317 10115 2375 10121
rect 2317 10081 2329 10115
rect 2363 10112 2375 10115
rect 2777 10115 2835 10121
rect 2777 10112 2789 10115
rect 2363 10084 2789 10112
rect 2363 10081 2375 10084
rect 2317 10075 2375 10081
rect 2777 10081 2789 10084
rect 2823 10112 2835 10115
rect 3694 10112 3700 10124
rect 2823 10084 3700 10112
rect 2823 10081 2835 10084
rect 2777 10075 2835 10081
rect 3694 10072 3700 10084
rect 3752 10072 3758 10124
rect 4433 10115 4491 10121
rect 4433 10081 4445 10115
rect 4479 10112 4491 10115
rect 5442 10112 5448 10124
rect 4479 10084 5448 10112
rect 4479 10081 4491 10084
rect 4433 10075 4491 10081
rect 5442 10072 5448 10084
rect 5500 10072 5506 10124
rect 10134 10072 10140 10124
rect 10192 10112 10198 10124
rect 10505 10115 10563 10121
rect 10505 10112 10517 10115
rect 10192 10084 10517 10112
rect 10192 10072 10198 10084
rect 10505 10081 10517 10084
rect 10551 10112 10563 10115
rect 11054 10112 11060 10124
rect 10551 10084 11060 10112
rect 10551 10081 10563 10084
rect 10505 10075 10563 10081
rect 11054 10072 11060 10084
rect 11112 10072 11118 10124
rect 13354 10112 13360 10124
rect 13315 10084 13360 10112
rect 13354 10072 13360 10084
rect 13412 10072 13418 10124
rect 15838 10112 15844 10124
rect 15751 10084 15844 10112
rect 2961 10047 3019 10053
rect 2961 10013 2973 10047
rect 3007 10013 3019 10047
rect 4522 10044 4528 10056
rect 4483 10016 4528 10044
rect 2961 10007 3019 10013
rect 1673 9979 1731 9985
rect 1673 9945 1685 9979
rect 1719 9976 1731 9979
rect 2222 9976 2228 9988
rect 1719 9948 2228 9976
rect 1719 9945 1731 9948
rect 1673 9939 1731 9945
rect 2222 9936 2228 9948
rect 2280 9976 2286 9988
rect 2682 9976 2688 9988
rect 2280 9948 2688 9976
rect 2280 9936 2286 9948
rect 2682 9936 2688 9948
rect 2740 9936 2746 9988
rect 2976 9976 3004 10007
rect 4522 10004 4528 10016
rect 4580 10004 4586 10056
rect 4706 10044 4712 10056
rect 4667 10016 4712 10044
rect 4706 10004 4712 10016
rect 4764 10004 4770 10056
rect 5166 10004 5172 10056
rect 5224 10044 5230 10056
rect 5721 10047 5779 10053
rect 5721 10044 5733 10047
rect 5224 10016 5733 10044
rect 5224 10004 5230 10016
rect 5721 10013 5733 10016
rect 5767 10013 5779 10047
rect 5721 10007 5779 10013
rect 13633 10047 13691 10053
rect 13633 10013 13645 10047
rect 13679 10044 13691 10047
rect 13722 10044 13728 10056
rect 13679 10016 13728 10044
rect 13679 10013 13691 10016
rect 13633 10007 13691 10013
rect 13722 10004 13728 10016
rect 13780 10004 13786 10056
rect 3050 9976 3056 9988
rect 2976 9948 3056 9976
rect 3050 9936 3056 9948
rect 3108 9976 3114 9988
rect 4430 9976 4436 9988
rect 3108 9948 4436 9976
rect 3108 9936 3114 9948
rect 4430 9936 4436 9948
rect 4488 9936 4494 9988
rect 7098 9976 7104 9988
rect 7059 9948 7104 9976
rect 7098 9936 7104 9948
rect 7156 9936 7162 9988
rect 12894 9976 12900 9988
rect 12855 9948 12900 9976
rect 12894 9936 12900 9948
rect 12952 9936 12958 9988
rect 1946 9868 1952 9920
rect 2004 9908 2010 9920
rect 2409 9911 2467 9917
rect 2409 9908 2421 9911
rect 2004 9880 2421 9908
rect 2004 9868 2010 9880
rect 2409 9877 2421 9880
rect 2455 9877 2467 9911
rect 2409 9871 2467 9877
rect 3142 9868 3148 9920
rect 3200 9908 3206 9920
rect 4065 9911 4123 9917
rect 4065 9908 4077 9911
rect 3200 9880 4077 9908
rect 3200 9868 3206 9880
rect 4065 9877 4077 9880
rect 4111 9877 4123 9911
rect 4065 9871 4123 9877
rect 4154 9868 4160 9920
rect 4212 9908 4218 9920
rect 5077 9911 5135 9917
rect 5077 9908 5089 9911
rect 4212 9880 5089 9908
rect 4212 9868 4218 9880
rect 5077 9877 5089 9880
rect 5123 9877 5135 9911
rect 5077 9871 5135 9877
rect 8386 9868 8392 9920
rect 8444 9908 8450 9920
rect 8481 9911 8539 9917
rect 8481 9908 8493 9911
rect 8444 9880 8493 9908
rect 8444 9868 8450 9880
rect 8481 9877 8493 9880
rect 8527 9908 8539 9911
rect 8849 9911 8907 9917
rect 8849 9908 8861 9911
rect 8527 9880 8861 9908
rect 8527 9877 8539 9880
rect 8481 9871 8539 9877
rect 8849 9877 8861 9880
rect 8895 9908 8907 9911
rect 9398 9908 9404 9920
rect 8895 9880 9404 9908
rect 8895 9877 8907 9880
rect 8849 9871 8907 9877
rect 9398 9868 9404 9880
rect 9456 9868 9462 9920
rect 11422 9868 11428 9920
rect 11480 9908 11486 9920
rect 11885 9911 11943 9917
rect 11885 9908 11897 9911
rect 11480 9880 11897 9908
rect 11480 9868 11486 9880
rect 11885 9877 11897 9880
rect 11931 9877 11943 9911
rect 11885 9871 11943 9877
rect 12158 9868 12164 9920
rect 12216 9908 12222 9920
rect 12434 9908 12440 9920
rect 12216 9880 12440 9908
rect 12216 9868 12222 9880
rect 12434 9868 12440 9880
rect 12492 9908 12498 9920
rect 12986 9908 12992 9920
rect 12492 9880 12585 9908
rect 12947 9880 12992 9908
rect 12492 9868 12498 9880
rect 12986 9868 12992 9880
rect 13044 9868 13050 9920
rect 15470 9868 15476 9920
rect 15528 9908 15534 9920
rect 15764 9917 15792 10084
rect 15838 10072 15844 10084
rect 15896 10112 15902 10124
rect 16189 10115 16247 10121
rect 16189 10112 16201 10115
rect 15896 10084 16201 10112
rect 15896 10072 15902 10084
rect 16189 10081 16201 10084
rect 16235 10112 16247 10115
rect 16942 10112 16948 10124
rect 16235 10084 16948 10112
rect 16235 10081 16247 10084
rect 16189 10075 16247 10081
rect 16942 10072 16948 10084
rect 17000 10072 17006 10124
rect 15930 10044 15936 10056
rect 15891 10016 15936 10044
rect 15930 10004 15936 10016
rect 15988 10004 15994 10056
rect 18966 10044 18972 10056
rect 18927 10016 18972 10044
rect 18966 10004 18972 10016
rect 19024 10004 19030 10056
rect 18138 9936 18144 9988
rect 18196 9976 18202 9988
rect 18417 9979 18475 9985
rect 18417 9976 18429 9979
rect 18196 9948 18429 9976
rect 18196 9936 18202 9948
rect 18417 9945 18429 9948
rect 18463 9945 18475 9979
rect 18417 9939 18475 9945
rect 15749 9911 15807 9917
rect 15749 9908 15761 9911
rect 15528 9880 15761 9908
rect 15528 9868 15534 9880
rect 15749 9877 15761 9880
rect 15795 9877 15807 9911
rect 15749 9871 15807 9877
rect 16574 9868 16580 9920
rect 16632 9908 16638 9920
rect 17313 9911 17371 9917
rect 17313 9908 17325 9911
rect 16632 9880 17325 9908
rect 16632 9868 16638 9880
rect 17313 9877 17325 9880
rect 17359 9877 17371 9911
rect 19426 9908 19432 9920
rect 19387 9880 19432 9908
rect 17313 9871 17371 9877
rect 19426 9868 19432 9880
rect 19484 9908 19490 9920
rect 19797 9911 19855 9917
rect 19797 9908 19809 9911
rect 19484 9880 19809 9908
rect 19484 9868 19490 9880
rect 19797 9877 19809 9880
rect 19843 9877 19855 9911
rect 19797 9871 19855 9877
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 2501 9707 2559 9713
rect 2501 9673 2513 9707
rect 2547 9704 2559 9707
rect 2590 9704 2596 9716
rect 2547 9676 2596 9704
rect 2547 9673 2559 9676
rect 2501 9667 2559 9673
rect 2590 9664 2596 9676
rect 2648 9664 2654 9716
rect 4246 9664 4252 9716
rect 4304 9704 4310 9716
rect 4706 9704 4712 9716
rect 4304 9676 4712 9704
rect 4304 9664 4310 9676
rect 4706 9664 4712 9676
rect 4764 9664 4770 9716
rect 4798 9664 4804 9716
rect 4856 9704 4862 9716
rect 6086 9704 6092 9716
rect 4856 9676 5488 9704
rect 6047 9676 6092 9704
rect 4856 9664 4862 9676
rect 5460 9636 5488 9676
rect 6086 9664 6092 9676
rect 6144 9664 6150 9716
rect 15378 9704 15384 9716
rect 10704 9676 15384 9704
rect 6365 9639 6423 9645
rect 6365 9636 6377 9639
rect 5460 9608 6377 9636
rect 6365 9605 6377 9608
rect 6411 9605 6423 9639
rect 6365 9599 6423 9605
rect 7101 9639 7159 9645
rect 7101 9605 7113 9639
rect 7147 9636 7159 9639
rect 7190 9636 7196 9648
rect 7147 9608 7196 9636
rect 7147 9605 7159 9608
rect 7101 9599 7159 9605
rect 7190 9596 7196 9608
rect 7248 9596 7254 9648
rect 7561 9639 7619 9645
rect 7561 9605 7573 9639
rect 7607 9636 7619 9639
rect 7742 9636 7748 9648
rect 7607 9608 7748 9636
rect 7607 9605 7619 9608
rect 7561 9599 7619 9605
rect 7742 9596 7748 9608
rect 7800 9596 7806 9648
rect 9122 9636 9128 9648
rect 9083 9608 9128 9636
rect 9122 9596 9128 9608
rect 9180 9596 9186 9648
rect 10704 9636 10732 9676
rect 15378 9664 15384 9676
rect 15436 9664 15442 9716
rect 15930 9664 15936 9716
rect 15988 9704 15994 9716
rect 15988 9676 16620 9704
rect 15988 9664 15994 9676
rect 9600 9608 10732 9636
rect 2038 9528 2044 9580
rect 2096 9568 2102 9580
rect 2774 9568 2780 9580
rect 2096 9540 2780 9568
rect 2096 9528 2102 9540
rect 2774 9528 2780 9540
rect 2832 9528 2838 9580
rect 5074 9568 5080 9580
rect 5035 9540 5080 9568
rect 5074 9528 5080 9540
rect 5132 9528 5138 9580
rect 5534 9568 5540 9580
rect 5495 9540 5540 9568
rect 5534 9528 5540 9540
rect 5592 9528 5598 9580
rect 7469 9571 7527 9577
rect 7469 9537 7481 9571
rect 7515 9568 7527 9571
rect 8110 9568 8116 9580
rect 7515 9540 8116 9568
rect 7515 9537 7527 9540
rect 7469 9531 7527 9537
rect 8110 9528 8116 9540
rect 8168 9528 8174 9580
rect 9214 9528 9220 9580
rect 9272 9568 9278 9580
rect 9600 9577 9628 9608
rect 10778 9596 10784 9648
rect 10836 9636 10842 9648
rect 11146 9636 11152 9648
rect 10836 9608 11152 9636
rect 10836 9596 10842 9608
rect 11146 9596 11152 9608
rect 11204 9596 11210 9648
rect 15562 9636 15568 9648
rect 15523 9608 15568 9636
rect 15562 9596 15568 9608
rect 15620 9636 15626 9648
rect 16592 9636 16620 9676
rect 17034 9636 17040 9648
rect 15620 9608 16528 9636
rect 16592 9608 17040 9636
rect 15620 9596 15626 9608
rect 9585 9571 9643 9577
rect 9585 9568 9597 9571
rect 9272 9540 9597 9568
rect 9272 9528 9278 9540
rect 9585 9537 9597 9540
rect 9631 9537 9643 9571
rect 9585 9531 9643 9537
rect 9769 9571 9827 9577
rect 9769 9537 9781 9571
rect 9815 9568 9827 9571
rect 9950 9568 9956 9580
rect 9815 9540 9956 9568
rect 9815 9537 9827 9540
rect 9769 9531 9827 9537
rect 9950 9528 9956 9540
rect 10008 9568 10014 9580
rect 10229 9571 10287 9577
rect 10229 9568 10241 9571
rect 10008 9540 10241 9568
rect 10008 9528 10014 9540
rect 10229 9537 10241 9540
rect 10275 9568 10287 9571
rect 11241 9571 11299 9577
rect 11241 9568 11253 9571
rect 10275 9540 11253 9568
rect 10275 9537 10287 9540
rect 10229 9531 10287 9537
rect 11241 9537 11253 9540
rect 11287 9537 11299 9571
rect 11241 9531 11299 9537
rect 14274 9528 14280 9580
rect 14332 9568 14338 9580
rect 14550 9568 14556 9580
rect 14332 9540 14556 9568
rect 14332 9528 14338 9540
rect 14550 9528 14556 9540
rect 14608 9528 14614 9580
rect 16500 9577 16528 9608
rect 17034 9596 17040 9608
rect 17092 9596 17098 9648
rect 17497 9639 17555 9645
rect 17497 9605 17509 9639
rect 17543 9636 17555 9639
rect 17862 9636 17868 9648
rect 17543 9608 17868 9636
rect 17543 9605 17555 9608
rect 17497 9599 17555 9605
rect 17862 9596 17868 9608
rect 17920 9596 17926 9648
rect 19334 9596 19340 9648
rect 19392 9636 19398 9648
rect 19981 9639 20039 9645
rect 19981 9636 19993 9639
rect 19392 9608 19993 9636
rect 19392 9596 19398 9608
rect 19981 9605 19993 9608
rect 20027 9605 20039 9639
rect 19981 9599 20039 9605
rect 16485 9571 16543 9577
rect 16485 9537 16497 9571
rect 16531 9537 16543 9571
rect 16485 9531 16543 9537
rect 16574 9528 16580 9580
rect 16632 9568 16638 9580
rect 17773 9571 17831 9577
rect 17773 9568 17785 9571
rect 16632 9540 17785 9568
rect 16632 9528 16638 9540
rect 17773 9537 17785 9540
rect 17819 9568 17831 9571
rect 17819 9540 18184 9568
rect 17819 9537 17831 9540
rect 17773 9531 17831 9537
rect 1394 9500 1400 9512
rect 1355 9472 1400 9500
rect 1394 9460 1400 9472
rect 1452 9460 1458 9512
rect 1673 9503 1731 9509
rect 1673 9469 1685 9503
rect 1719 9500 1731 9503
rect 2498 9500 2504 9512
rect 1719 9472 2504 9500
rect 1719 9469 1731 9472
rect 1673 9463 1731 9469
rect 2498 9460 2504 9472
rect 2556 9460 2562 9512
rect 2792 9432 2820 9528
rect 3050 9509 3056 9512
rect 3044 9500 3056 9509
rect 3011 9472 3056 9500
rect 3044 9463 3056 9472
rect 3050 9460 3056 9463
rect 3108 9460 3114 9512
rect 3602 9460 3608 9512
rect 3660 9500 3666 9512
rect 4985 9503 5043 9509
rect 4985 9500 4997 9503
rect 3660 9472 4997 9500
rect 3660 9460 3666 9472
rect 4985 9469 4997 9472
rect 5031 9469 5043 9503
rect 5092 9500 5120 9528
rect 5261 9503 5319 9509
rect 5261 9500 5273 9503
rect 5092 9472 5273 9500
rect 4985 9463 5043 9469
rect 5261 9469 5273 9472
rect 5307 9469 5319 9503
rect 5261 9463 5319 9469
rect 8021 9503 8079 9509
rect 8021 9469 8033 9503
rect 8067 9500 8079 9503
rect 8202 9500 8208 9512
rect 8067 9472 8208 9500
rect 8067 9469 8079 9472
rect 8021 9463 8079 9469
rect 8202 9460 8208 9472
rect 8260 9460 8266 9512
rect 10134 9460 10140 9512
rect 10192 9500 10198 9512
rect 10594 9500 10600 9512
rect 10192 9472 10600 9500
rect 10192 9460 10198 9472
rect 10594 9460 10600 9472
rect 10652 9460 10658 9512
rect 10686 9460 10692 9512
rect 10744 9500 10750 9512
rect 11701 9503 11759 9509
rect 11701 9500 11713 9503
rect 10744 9472 11713 9500
rect 10744 9460 10750 9472
rect 11701 9469 11713 9472
rect 11747 9469 11759 9503
rect 11701 9463 11759 9469
rect 12526 9460 12532 9512
rect 12584 9500 12590 9512
rect 13262 9500 13268 9512
rect 12584 9472 13268 9500
rect 12584 9460 12590 9472
rect 13262 9460 13268 9472
rect 13320 9460 13326 9512
rect 16298 9460 16304 9512
rect 16356 9500 16362 9512
rect 16393 9503 16451 9509
rect 16393 9500 16405 9503
rect 16356 9472 16405 9500
rect 16356 9460 16362 9472
rect 16393 9469 16405 9472
rect 16439 9469 16451 9503
rect 16393 9463 16451 9469
rect 17034 9460 17040 9512
rect 17092 9500 17098 9512
rect 18049 9503 18107 9509
rect 18049 9500 18061 9503
rect 17092 9472 18061 9500
rect 17092 9460 17098 9472
rect 18049 9469 18061 9472
rect 18095 9469 18107 9503
rect 18156 9500 18184 9540
rect 18305 9503 18363 9509
rect 18305 9500 18317 9503
rect 18156 9472 18317 9500
rect 18049 9463 18107 9469
rect 18305 9469 18317 9472
rect 18351 9469 18363 9503
rect 18305 9463 18363 9469
rect 5074 9432 5080 9444
rect 2792 9404 5080 9432
rect 5074 9392 5080 9404
rect 5132 9392 5138 9444
rect 7929 9435 7987 9441
rect 7929 9401 7941 9435
rect 7975 9432 7987 9435
rect 8665 9435 8723 9441
rect 8665 9432 8677 9435
rect 7975 9404 8677 9432
rect 7975 9401 7987 9404
rect 7929 9395 7987 9401
rect 8665 9401 8677 9404
rect 8711 9432 8723 9435
rect 9950 9432 9956 9444
rect 8711 9404 9956 9432
rect 8711 9401 8723 9404
rect 8665 9395 8723 9401
rect 9950 9392 9956 9404
rect 10008 9392 10014 9444
rect 10042 9392 10048 9444
rect 10100 9432 10106 9444
rect 10100 9404 10732 9432
rect 10100 9392 10106 9404
rect 4154 9364 4160 9376
rect 4115 9336 4160 9364
rect 4154 9324 4160 9336
rect 4212 9324 4218 9376
rect 4985 9367 5043 9373
rect 4985 9333 4997 9367
rect 5031 9364 5043 9367
rect 8941 9367 8999 9373
rect 8941 9364 8953 9367
rect 5031 9336 8953 9364
rect 5031 9333 5043 9336
rect 4985 9327 5043 9333
rect 8941 9333 8953 9336
rect 8987 9364 8999 9367
rect 9490 9364 9496 9376
rect 8987 9336 9496 9364
rect 8987 9333 8999 9336
rect 8941 9327 8999 9333
rect 9490 9324 9496 9336
rect 9548 9324 9554 9376
rect 10704 9373 10732 9404
rect 10778 9392 10784 9444
rect 10836 9432 10842 9444
rect 10962 9432 10968 9444
rect 10836 9404 10968 9432
rect 10836 9392 10842 9404
rect 10962 9392 10968 9404
rect 11020 9432 11026 9444
rect 11149 9435 11207 9441
rect 11149 9432 11161 9435
rect 11020 9404 11161 9432
rect 11020 9392 11026 9404
rect 11149 9401 11161 9404
rect 11195 9401 11207 9435
rect 11149 9395 11207 9401
rect 12253 9435 12311 9441
rect 12253 9401 12265 9435
rect 12299 9432 12311 9435
rect 13354 9432 13360 9444
rect 12299 9404 13360 9432
rect 12299 9401 12311 9404
rect 12253 9395 12311 9401
rect 13354 9392 13360 9404
rect 13412 9392 13418 9444
rect 13532 9435 13590 9441
rect 13532 9432 13544 9435
rect 13464 9404 13544 9432
rect 10689 9367 10747 9373
rect 10689 9333 10701 9367
rect 10735 9333 10747 9367
rect 10689 9327 10747 9333
rect 11057 9367 11115 9373
rect 11057 9333 11069 9367
rect 11103 9364 11115 9367
rect 11238 9364 11244 9376
rect 11103 9336 11244 9364
rect 11103 9333 11115 9336
rect 11057 9327 11115 9333
rect 11238 9324 11244 9336
rect 11296 9324 11302 9376
rect 12802 9364 12808 9376
rect 12763 9336 12808 9364
rect 12802 9324 12808 9336
rect 12860 9324 12866 9376
rect 12894 9324 12900 9376
rect 12952 9364 12958 9376
rect 13173 9367 13231 9373
rect 13173 9364 13185 9367
rect 12952 9336 13185 9364
rect 12952 9324 12958 9336
rect 13173 9333 13185 9336
rect 13219 9364 13231 9367
rect 13464 9364 13492 9404
rect 13532 9401 13544 9404
rect 13578 9432 13590 9435
rect 14274 9432 14280 9444
rect 13578 9404 14280 9432
rect 13578 9401 13590 9404
rect 13532 9395 13590 9401
rect 14274 9392 14280 9404
rect 14332 9392 14338 9444
rect 18064 9432 18092 9463
rect 19334 9432 19340 9444
rect 18064 9404 19340 9432
rect 19334 9392 19340 9404
rect 19392 9392 19398 9444
rect 13219 9336 13492 9364
rect 13219 9333 13231 9336
rect 13173 9327 13231 9333
rect 13722 9324 13728 9376
rect 13780 9364 13786 9376
rect 14645 9367 14703 9373
rect 14645 9364 14657 9367
rect 13780 9336 14657 9364
rect 13780 9324 13786 9336
rect 14645 9333 14657 9336
rect 14691 9333 14703 9367
rect 14645 9327 14703 9333
rect 15470 9324 15476 9376
rect 15528 9364 15534 9376
rect 15841 9367 15899 9373
rect 15841 9364 15853 9367
rect 15528 9336 15853 9364
rect 15528 9324 15534 9336
rect 15841 9333 15853 9336
rect 15887 9333 15899 9367
rect 16022 9364 16028 9376
rect 15983 9336 16028 9364
rect 15841 9327 15899 9333
rect 16022 9324 16028 9336
rect 16080 9324 16086 9376
rect 17129 9367 17187 9373
rect 17129 9333 17141 9367
rect 17175 9364 17187 9367
rect 17218 9364 17224 9376
rect 17175 9336 17224 9364
rect 17175 9333 17187 9336
rect 17129 9327 17187 9333
rect 17218 9324 17224 9336
rect 17276 9324 17282 9376
rect 19426 9364 19432 9376
rect 19387 9336 19432 9364
rect 19426 9324 19432 9336
rect 19484 9324 19490 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 2774 9120 2780 9172
rect 2832 9160 2838 9172
rect 2832 9132 2877 9160
rect 2832 9120 2838 9132
rect 5074 9120 5080 9172
rect 5132 9160 5138 9172
rect 5629 9163 5687 9169
rect 5629 9160 5641 9163
rect 5132 9132 5641 9160
rect 5132 9120 5138 9132
rect 5629 9129 5641 9132
rect 5675 9129 5687 9163
rect 8478 9160 8484 9172
rect 8439 9132 8484 9160
rect 5629 9123 5687 9129
rect 8478 9120 8484 9132
rect 8536 9120 8542 9172
rect 9214 9160 9220 9172
rect 9175 9132 9220 9160
rect 9214 9120 9220 9132
rect 9272 9120 9278 9172
rect 9398 9120 9404 9172
rect 9456 9160 9462 9172
rect 9861 9163 9919 9169
rect 9861 9160 9873 9163
rect 9456 9132 9873 9160
rect 9456 9120 9462 9132
rect 9861 9129 9873 9132
rect 9907 9160 9919 9163
rect 10962 9160 10968 9172
rect 9907 9132 10968 9160
rect 9907 9129 9919 9132
rect 9861 9123 9919 9129
rect 10962 9120 10968 9132
rect 11020 9120 11026 9172
rect 13078 9160 13084 9172
rect 13039 9132 13084 9160
rect 13078 9120 13084 9132
rect 13136 9120 13142 9172
rect 13354 9120 13360 9172
rect 13412 9160 13418 9172
rect 13633 9163 13691 9169
rect 13633 9160 13645 9163
rect 13412 9132 13645 9160
rect 13412 9120 13418 9132
rect 13633 9129 13645 9132
rect 13679 9129 13691 9163
rect 13633 9123 13691 9129
rect 16298 9120 16304 9172
rect 16356 9160 16362 9172
rect 16393 9163 16451 9169
rect 16393 9160 16405 9163
rect 16356 9132 16405 9160
rect 16356 9120 16362 9132
rect 16393 9129 16405 9132
rect 16439 9129 16451 9163
rect 17218 9160 17224 9172
rect 16393 9123 16451 9129
rect 16684 9132 17224 9160
rect 1664 9095 1722 9101
rect 1664 9061 1676 9095
rect 1710 9092 1722 9095
rect 2222 9092 2228 9104
rect 1710 9064 2228 9092
rect 1710 9061 1722 9064
rect 1664 9055 1722 9061
rect 2222 9052 2228 9064
rect 2280 9052 2286 9104
rect 4525 9095 4583 9101
rect 4525 9061 4537 9095
rect 4571 9092 4583 9095
rect 4614 9092 4620 9104
rect 4571 9064 4620 9092
rect 4571 9061 4583 9064
rect 4525 9055 4583 9061
rect 4614 9052 4620 9064
rect 4672 9052 4678 9104
rect 11330 9052 11336 9104
rect 11388 9101 11394 9104
rect 11388 9095 11452 9101
rect 11388 9061 11406 9095
rect 11440 9061 11452 9095
rect 11388 9055 11452 9061
rect 11388 9052 11394 9055
rect 15286 9052 15292 9104
rect 15344 9092 15350 9104
rect 15565 9095 15623 9101
rect 15565 9092 15577 9095
rect 15344 9064 15577 9092
rect 15344 9052 15350 9064
rect 15565 9061 15577 9064
rect 15611 9092 15623 9095
rect 16684 9092 16712 9132
rect 17218 9120 17224 9132
rect 17276 9120 17282 9172
rect 17954 9160 17960 9172
rect 17915 9132 17960 9160
rect 17954 9120 17960 9132
rect 18012 9120 18018 9172
rect 18601 9163 18659 9169
rect 18601 9129 18613 9163
rect 18647 9160 18659 9163
rect 18966 9160 18972 9172
rect 18647 9132 18972 9160
rect 18647 9129 18659 9132
rect 18601 9123 18659 9129
rect 18966 9120 18972 9132
rect 19024 9120 19030 9172
rect 16850 9101 16856 9104
rect 16844 9092 16856 9101
rect 15611 9064 16712 9092
rect 16811 9064 16856 9092
rect 15611 9061 15623 9064
rect 15565 9055 15623 9061
rect 16844 9055 16856 9064
rect 16850 9052 16856 9055
rect 16908 9052 16914 9104
rect 17034 9052 17040 9104
rect 17092 9052 17098 9104
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 9024 1455 9027
rect 2038 9024 2044 9036
rect 1443 8996 2044 9024
rect 1443 8993 1455 8996
rect 1397 8987 1455 8993
rect 2038 8984 2044 8996
rect 2096 8984 2102 9036
rect 4433 9027 4491 9033
rect 4433 8993 4445 9027
rect 4479 9024 4491 9027
rect 4798 9024 4804 9036
rect 4479 8996 4804 9024
rect 4479 8993 4491 8996
rect 4433 8987 4491 8993
rect 4798 8984 4804 8996
rect 4856 8984 4862 9036
rect 5813 9027 5871 9033
rect 5813 8993 5825 9027
rect 5859 9024 5871 9027
rect 6638 9024 6644 9036
rect 5859 8996 6644 9024
rect 5859 8993 5871 8996
rect 5813 8987 5871 8993
rect 6638 8984 6644 8996
rect 6696 8984 6702 9036
rect 7368 9027 7426 9033
rect 7368 8993 7380 9027
rect 7414 9024 7426 9027
rect 8202 9024 8208 9036
rect 7414 8996 8208 9024
rect 7414 8993 7426 8996
rect 7368 8987 7426 8993
rect 8202 8984 8208 8996
rect 8260 8984 8266 9036
rect 13262 8984 13268 9036
rect 13320 9024 13326 9036
rect 14001 9027 14059 9033
rect 14001 9024 14013 9027
rect 13320 8996 14013 9024
rect 13320 8984 13326 8996
rect 14001 8993 14013 8996
rect 14047 8993 14059 9027
rect 14001 8987 14059 8993
rect 16577 9027 16635 9033
rect 16577 8993 16589 9027
rect 16623 9024 16635 9027
rect 17052 9024 17080 9052
rect 19426 9024 19432 9036
rect 16623 8996 17080 9024
rect 19387 8996 19432 9024
rect 16623 8993 16635 8996
rect 16577 8987 16635 8993
rect 19426 8984 19432 8996
rect 19484 8984 19490 9036
rect 4617 8959 4675 8965
rect 4617 8925 4629 8959
rect 4663 8925 4675 8959
rect 4617 8919 4675 8925
rect 3418 8888 3424 8900
rect 3331 8860 3424 8888
rect 3418 8848 3424 8860
rect 3476 8888 3482 8900
rect 4430 8888 4436 8900
rect 3476 8860 4436 8888
rect 3476 8848 3482 8860
rect 4430 8848 4436 8860
rect 4488 8888 4494 8900
rect 4632 8888 4660 8919
rect 5534 8916 5540 8968
rect 5592 8956 5598 8968
rect 5592 8928 6224 8956
rect 5592 8916 5598 8928
rect 5077 8891 5135 8897
rect 5077 8888 5089 8891
rect 4488 8860 5089 8888
rect 4488 8848 4494 8860
rect 5077 8857 5089 8860
rect 5123 8888 5135 8891
rect 5166 8888 5172 8900
rect 5123 8860 5172 8888
rect 5123 8857 5135 8860
rect 5077 8851 5135 8857
rect 5166 8848 5172 8860
rect 5224 8848 5230 8900
rect 3510 8780 3516 8832
rect 3568 8820 3574 8832
rect 3789 8823 3847 8829
rect 3789 8820 3801 8823
rect 3568 8792 3801 8820
rect 3568 8780 3574 8792
rect 3789 8789 3801 8792
rect 3835 8820 3847 8823
rect 4065 8823 4123 8829
rect 4065 8820 4077 8823
rect 3835 8792 4077 8820
rect 3835 8789 3847 8792
rect 3789 8783 3847 8789
rect 4065 8789 4077 8792
rect 4111 8789 4123 8823
rect 5534 8820 5540 8832
rect 5495 8792 5540 8820
rect 4065 8783 4123 8789
rect 5534 8780 5540 8792
rect 5592 8780 5598 8832
rect 6196 8829 6224 8928
rect 6546 8916 6552 8968
rect 6604 8956 6610 8968
rect 6822 8956 6828 8968
rect 6604 8928 6828 8956
rect 6604 8916 6610 8928
rect 6822 8916 6828 8928
rect 6880 8956 6886 8968
rect 7101 8959 7159 8965
rect 7101 8956 7113 8959
rect 6880 8928 7113 8956
rect 6880 8916 6886 8928
rect 7101 8925 7113 8928
rect 7147 8925 7159 8959
rect 7101 8919 7159 8925
rect 9858 8916 9864 8968
rect 9916 8956 9922 8968
rect 10045 8959 10103 8965
rect 10045 8956 10057 8959
rect 9916 8928 10057 8956
rect 9916 8916 9922 8928
rect 10045 8925 10057 8928
rect 10091 8925 10103 8959
rect 10045 8919 10103 8925
rect 11054 8916 11060 8968
rect 11112 8956 11118 8968
rect 11149 8959 11207 8965
rect 11149 8956 11161 8959
rect 11112 8928 11161 8956
rect 11112 8916 11118 8928
rect 11149 8925 11161 8928
rect 11195 8925 11207 8959
rect 11149 8919 11207 8925
rect 13538 8916 13544 8968
rect 13596 8956 13602 8968
rect 14093 8959 14151 8965
rect 14093 8956 14105 8959
rect 13596 8928 14105 8956
rect 13596 8916 13602 8928
rect 14093 8925 14105 8928
rect 14139 8925 14151 8959
rect 14274 8956 14280 8968
rect 14235 8928 14280 8956
rect 14093 8919 14151 8925
rect 14274 8916 14280 8928
rect 14332 8916 14338 8968
rect 19334 8916 19340 8968
rect 19392 8956 19398 8968
rect 19521 8959 19579 8965
rect 19521 8956 19533 8959
rect 19392 8928 19533 8956
rect 19392 8916 19398 8928
rect 19521 8925 19533 8928
rect 19567 8925 19579 8959
rect 19521 8919 19579 8925
rect 19613 8959 19671 8965
rect 19613 8925 19625 8959
rect 19659 8925 19671 8959
rect 19613 8919 19671 8925
rect 12894 8848 12900 8900
rect 12952 8888 12958 8900
rect 12952 8860 14780 8888
rect 12952 8848 12958 8860
rect 6181 8823 6239 8829
rect 6181 8789 6193 8823
rect 6227 8820 6239 8823
rect 6270 8820 6276 8832
rect 6227 8792 6276 8820
rect 6227 8789 6239 8792
rect 6181 8783 6239 8789
rect 6270 8780 6276 8792
rect 6328 8780 6334 8832
rect 6546 8820 6552 8832
rect 6507 8792 6552 8820
rect 6546 8780 6552 8792
rect 6604 8780 6610 8832
rect 6914 8820 6920 8832
rect 6875 8792 6920 8820
rect 6914 8780 6920 8792
rect 6972 8780 6978 8832
rect 10778 8820 10784 8832
rect 10739 8792 10784 8820
rect 10778 8780 10784 8792
rect 10836 8780 10842 8832
rect 12434 8780 12440 8832
rect 12492 8820 12498 8832
rect 12529 8823 12587 8829
rect 12529 8820 12541 8823
rect 12492 8792 12541 8820
rect 12492 8780 12498 8792
rect 12529 8789 12541 8792
rect 12575 8789 12587 8823
rect 12529 8783 12587 8789
rect 12802 8780 12808 8832
rect 12860 8820 12866 8832
rect 13541 8823 13599 8829
rect 13541 8820 13553 8823
rect 12860 8792 13553 8820
rect 12860 8780 12866 8792
rect 13541 8789 13553 8792
rect 13587 8820 13599 8823
rect 13722 8820 13728 8832
rect 13587 8792 13728 8820
rect 13587 8789 13599 8792
rect 13541 8783 13599 8789
rect 13722 8780 13728 8792
rect 13780 8780 13786 8832
rect 14752 8829 14780 8860
rect 18598 8848 18604 8900
rect 18656 8888 18662 8900
rect 19628 8888 19656 8919
rect 20070 8888 20076 8900
rect 18656 8860 19656 8888
rect 20031 8860 20076 8888
rect 18656 8848 18662 8860
rect 19536 8832 19564 8860
rect 20070 8848 20076 8860
rect 20128 8848 20134 8900
rect 14737 8823 14795 8829
rect 14737 8789 14749 8823
rect 14783 8820 14795 8823
rect 15013 8823 15071 8829
rect 15013 8820 15025 8823
rect 14783 8792 15025 8820
rect 14783 8789 14795 8792
rect 14737 8783 14795 8789
rect 15013 8789 15025 8792
rect 15059 8820 15071 8823
rect 15378 8820 15384 8832
rect 15059 8792 15384 8820
rect 15059 8789 15071 8792
rect 15013 8783 15071 8789
rect 15378 8780 15384 8792
rect 15436 8780 15442 8832
rect 15562 8780 15568 8832
rect 15620 8820 15626 8832
rect 16025 8823 16083 8829
rect 16025 8820 16037 8823
rect 15620 8792 16037 8820
rect 15620 8780 15626 8792
rect 16025 8789 16037 8792
rect 16071 8820 16083 8823
rect 16574 8820 16580 8832
rect 16071 8792 16580 8820
rect 16071 8789 16083 8792
rect 16025 8783 16083 8789
rect 16574 8780 16580 8792
rect 16632 8780 16638 8832
rect 18782 8780 18788 8832
rect 18840 8820 18846 8832
rect 18877 8823 18935 8829
rect 18877 8820 18889 8823
rect 18840 8792 18889 8820
rect 18840 8780 18846 8792
rect 18877 8789 18889 8792
rect 18923 8789 18935 8823
rect 19058 8820 19064 8832
rect 19019 8792 19064 8820
rect 18877 8783 18935 8789
rect 19058 8780 19064 8792
rect 19116 8780 19122 8832
rect 19518 8780 19524 8832
rect 19576 8780 19582 8832
rect 20438 8820 20444 8832
rect 20399 8792 20444 8820
rect 20438 8780 20444 8792
rect 20496 8780 20502 8832
rect 21174 8820 21180 8832
rect 21135 8792 21180 8820
rect 21174 8780 21180 8792
rect 21232 8780 21238 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 1489 8619 1547 8625
rect 1489 8585 1501 8619
rect 1535 8616 1547 8619
rect 1854 8616 1860 8628
rect 1535 8588 1860 8616
rect 1535 8585 1547 8588
rect 1489 8579 1547 8585
rect 1854 8576 1860 8588
rect 1912 8576 1918 8628
rect 3053 8619 3111 8625
rect 3053 8585 3065 8619
rect 3099 8616 3111 8619
rect 4062 8616 4068 8628
rect 3099 8588 4068 8616
rect 3099 8585 3111 8588
rect 3053 8579 3111 8585
rect 4062 8576 4068 8588
rect 4120 8576 4126 8628
rect 9858 8616 9864 8628
rect 9819 8588 9864 8616
rect 9858 8576 9864 8588
rect 9916 8576 9922 8628
rect 9950 8576 9956 8628
rect 10008 8616 10014 8628
rect 11241 8619 11299 8625
rect 10008 8588 10053 8616
rect 10008 8576 10014 8588
rect 11241 8585 11253 8619
rect 11287 8616 11299 8619
rect 11330 8616 11336 8628
rect 11287 8588 11336 8616
rect 11287 8585 11299 8588
rect 11241 8579 11299 8585
rect 11330 8576 11336 8588
rect 11388 8576 11394 8628
rect 11422 8576 11428 8628
rect 11480 8616 11486 8628
rect 11609 8619 11667 8625
rect 11609 8616 11621 8619
rect 11480 8588 11621 8616
rect 11480 8576 11486 8588
rect 11609 8585 11621 8588
rect 11655 8616 11667 8619
rect 12894 8616 12900 8628
rect 11655 8588 12900 8616
rect 11655 8585 11667 8588
rect 11609 8579 11667 8585
rect 12894 8576 12900 8588
rect 12952 8576 12958 8628
rect 13262 8616 13268 8628
rect 13223 8588 13268 8616
rect 13262 8576 13268 8588
rect 13320 8576 13326 8628
rect 13538 8616 13544 8628
rect 13499 8588 13544 8616
rect 13538 8576 13544 8588
rect 13596 8576 13602 8628
rect 14090 8616 14096 8628
rect 13648 8588 14096 8616
rect 2593 8551 2651 8557
rect 2593 8517 2605 8551
rect 2639 8548 2651 8551
rect 2958 8548 2964 8560
rect 2639 8520 2964 8548
rect 2639 8517 2651 8520
rect 2593 8511 2651 8517
rect 2958 8508 2964 8520
rect 3016 8548 3022 8560
rect 3418 8548 3424 8560
rect 3016 8520 3424 8548
rect 3016 8508 3022 8520
rect 3418 8508 3424 8520
rect 3476 8508 3482 8560
rect 3878 8508 3884 8560
rect 3936 8548 3942 8560
rect 4617 8551 4675 8557
rect 4617 8548 4629 8551
rect 3936 8520 4629 8548
rect 3936 8508 3942 8520
rect 4617 8517 4629 8520
rect 4663 8517 4675 8551
rect 5994 8548 6000 8560
rect 5955 8520 6000 8548
rect 4617 8511 4675 8517
rect 5994 8508 6000 8520
rect 6052 8508 6058 8560
rect 6457 8551 6515 8557
rect 6457 8517 6469 8551
rect 6503 8548 6515 8551
rect 6822 8548 6828 8560
rect 6503 8520 6828 8548
rect 6503 8517 6515 8520
rect 6457 8511 6515 8517
rect 6822 8508 6828 8520
rect 6880 8508 6886 8560
rect 8202 8548 8208 8560
rect 8163 8520 8208 8548
rect 8202 8508 8208 8520
rect 8260 8508 8266 8560
rect 8846 8548 8852 8560
rect 8759 8520 8852 8548
rect 8846 8508 8852 8520
rect 8904 8548 8910 8560
rect 8904 8520 12020 8548
rect 8904 8508 8910 8520
rect 1946 8480 1952 8492
rect 1907 8452 1952 8480
rect 1946 8440 1952 8452
rect 2004 8440 2010 8492
rect 2133 8483 2191 8489
rect 2133 8449 2145 8483
rect 2179 8480 2191 8483
rect 2222 8480 2228 8492
rect 2179 8452 2228 8480
rect 2179 8449 2191 8452
rect 2133 8443 2191 8449
rect 2222 8440 2228 8452
rect 2280 8440 2286 8492
rect 3510 8480 3516 8492
rect 3471 8452 3516 8480
rect 3510 8440 3516 8452
rect 3568 8440 3574 8492
rect 3602 8440 3608 8492
rect 3660 8480 3666 8492
rect 3697 8483 3755 8489
rect 3697 8480 3709 8483
rect 3660 8452 3709 8480
rect 3660 8440 3666 8452
rect 3697 8449 3709 8452
rect 3743 8480 3755 8483
rect 4154 8480 4160 8492
rect 3743 8452 4160 8480
rect 3743 8449 3755 8452
rect 3697 8443 3755 8449
rect 4154 8440 4160 8452
rect 4212 8440 4218 8492
rect 5166 8480 5172 8492
rect 5127 8452 5172 8480
rect 5166 8440 5172 8452
rect 5224 8480 5230 8492
rect 5629 8483 5687 8489
rect 5629 8480 5641 8483
rect 5224 8452 5641 8480
rect 5224 8440 5230 8452
rect 5629 8449 5641 8452
rect 5675 8449 5687 8483
rect 5629 8443 5687 8449
rect 2240 8412 2268 8440
rect 2961 8415 3019 8421
rect 2961 8412 2973 8415
rect 2240 8384 2973 8412
rect 2961 8381 2973 8384
rect 3007 8412 3019 8415
rect 3620 8412 3648 8440
rect 3007 8384 3648 8412
rect 4525 8415 4583 8421
rect 3007 8381 3019 8384
rect 2961 8375 3019 8381
rect 4525 8381 4537 8415
rect 4571 8412 4583 8415
rect 6638 8412 6644 8424
rect 4571 8384 5120 8412
rect 6599 8384 6644 8412
rect 4571 8381 4583 8384
rect 4525 8375 4583 8381
rect 1857 8347 1915 8353
rect 1857 8313 1869 8347
rect 1903 8344 1915 8347
rect 2406 8344 2412 8356
rect 1903 8316 2412 8344
rect 1903 8313 1915 8316
rect 1857 8307 1915 8313
rect 2406 8304 2412 8316
rect 2464 8304 2470 8356
rect 4157 8347 4215 8353
rect 4157 8313 4169 8347
rect 4203 8344 4215 8347
rect 4798 8344 4804 8356
rect 4203 8316 4804 8344
rect 4203 8313 4215 8316
rect 4157 8307 4215 8313
rect 4798 8304 4804 8316
rect 4856 8304 4862 8356
rect 3421 8279 3479 8285
rect 3421 8245 3433 8279
rect 3467 8276 3479 8279
rect 3878 8276 3884 8288
rect 3467 8248 3884 8276
rect 3467 8245 3479 8248
rect 3421 8239 3479 8245
rect 3878 8236 3884 8248
rect 3936 8236 3942 8288
rect 4706 8236 4712 8288
rect 4764 8276 4770 8288
rect 4982 8276 4988 8288
rect 4764 8248 4988 8276
rect 4764 8236 4770 8248
rect 4982 8236 4988 8248
rect 5040 8236 5046 8288
rect 5092 8285 5120 8384
rect 6638 8372 6644 8384
rect 6696 8372 6702 8424
rect 6840 8421 6868 8508
rect 9493 8483 9551 8489
rect 9493 8449 9505 8483
rect 9539 8480 9551 8483
rect 10505 8483 10563 8489
rect 10505 8480 10517 8483
rect 9539 8452 10517 8480
rect 9539 8449 9551 8452
rect 9493 8443 9551 8449
rect 10505 8449 10517 8452
rect 10551 8480 10563 8483
rect 10686 8480 10692 8492
rect 10551 8452 10692 8480
rect 10551 8449 10563 8452
rect 10505 8443 10563 8449
rect 10686 8440 10692 8452
rect 10744 8440 10750 8492
rect 6825 8415 6883 8421
rect 6825 8381 6837 8415
rect 6871 8412 6883 8415
rect 8570 8412 8576 8424
rect 6871 8384 8576 8412
rect 6871 8381 6883 8384
rect 6825 8375 6883 8381
rect 8570 8372 8576 8384
rect 8628 8372 8634 8424
rect 9858 8372 9864 8424
rect 9916 8412 9922 8424
rect 11992 8421 12020 8520
rect 12713 8483 12771 8489
rect 12713 8449 12725 8483
rect 12759 8480 12771 8483
rect 13280 8480 13308 8576
rect 13449 8551 13507 8557
rect 13449 8517 13461 8551
rect 13495 8548 13507 8551
rect 13648 8548 13676 8588
rect 14090 8576 14096 8588
rect 14148 8576 14154 8628
rect 15749 8619 15807 8625
rect 15749 8585 15761 8619
rect 15795 8616 15807 8619
rect 16022 8616 16028 8628
rect 15795 8588 16028 8616
rect 15795 8585 15807 8588
rect 15749 8579 15807 8585
rect 16022 8576 16028 8588
rect 16080 8576 16086 8628
rect 16117 8619 16175 8625
rect 16117 8585 16129 8619
rect 16163 8616 16175 8619
rect 16850 8616 16856 8628
rect 16163 8588 16856 8616
rect 16163 8585 16175 8588
rect 16117 8579 16175 8585
rect 16850 8576 16856 8588
rect 16908 8616 16914 8628
rect 17221 8619 17279 8625
rect 17221 8616 17233 8619
rect 16908 8588 17233 8616
rect 16908 8576 16914 8588
rect 17221 8585 17233 8588
rect 17267 8585 17279 8619
rect 17221 8579 17279 8585
rect 20714 8576 20720 8628
rect 20772 8616 20778 8628
rect 21177 8619 21235 8625
rect 21177 8616 21189 8619
rect 20772 8588 21189 8616
rect 20772 8576 20778 8588
rect 21177 8585 21189 8588
rect 21223 8585 21235 8619
rect 21177 8579 21235 8585
rect 13495 8520 13676 8548
rect 13495 8517 13507 8520
rect 13449 8511 13507 8517
rect 12759 8452 13308 8480
rect 12759 8449 12771 8452
rect 12713 8443 12771 8449
rect 13354 8440 13360 8492
rect 13412 8480 13418 8492
rect 16868 8489 16896 8576
rect 17954 8508 17960 8560
rect 18012 8548 18018 8560
rect 19061 8551 19119 8557
rect 19061 8548 19073 8551
rect 18012 8520 19073 8548
rect 18012 8508 18018 8520
rect 19061 8517 19073 8520
rect 19107 8548 19119 8551
rect 19334 8548 19340 8560
rect 19107 8520 19340 8548
rect 19107 8517 19119 8520
rect 19061 8511 19119 8517
rect 19334 8508 19340 8520
rect 19392 8508 19398 8560
rect 19610 8548 19616 8560
rect 19571 8520 19616 8548
rect 19610 8508 19616 8520
rect 19668 8508 19674 8560
rect 20070 8508 20076 8560
rect 20128 8548 20134 8560
rect 20990 8548 20996 8560
rect 20128 8520 20208 8548
rect 20951 8520 20996 8548
rect 20128 8508 20134 8520
rect 16853 8483 16911 8489
rect 13412 8452 13860 8480
rect 13412 8440 13418 8452
rect 10321 8415 10379 8421
rect 10321 8412 10333 8415
rect 9916 8384 10333 8412
rect 9916 8372 9922 8384
rect 10321 8381 10333 8384
rect 10367 8381 10379 8415
rect 10321 8375 10379 8381
rect 11977 8415 12035 8421
rect 11977 8381 11989 8415
rect 12023 8412 12035 8415
rect 12253 8415 12311 8421
rect 12253 8412 12265 8415
rect 12023 8384 12265 8412
rect 12023 8381 12035 8384
rect 11977 8375 12035 8381
rect 12253 8381 12265 8384
rect 12299 8412 12311 8415
rect 13449 8415 13507 8421
rect 13449 8412 13461 8415
rect 12299 8384 13461 8412
rect 12299 8381 12311 8384
rect 12253 8375 12311 8381
rect 13449 8381 13461 8384
rect 13495 8381 13507 8415
rect 13449 8375 13507 8381
rect 13538 8372 13544 8424
rect 13596 8412 13602 8424
rect 13725 8415 13783 8421
rect 13725 8412 13737 8415
rect 13596 8384 13737 8412
rect 13596 8372 13602 8384
rect 13725 8381 13737 8384
rect 13771 8381 13783 8415
rect 13832 8412 13860 8452
rect 16853 8449 16865 8483
rect 16899 8449 16911 8483
rect 18598 8480 18604 8492
rect 16853 8443 16911 8449
rect 17788 8452 18604 8480
rect 13832 8384 14780 8412
rect 13725 8375 13783 8381
rect 6914 8344 6920 8356
rect 6827 8316 6920 8344
rect 5077 8279 5135 8285
rect 5077 8245 5089 8279
rect 5123 8276 5135 8279
rect 6362 8276 6368 8288
rect 5123 8248 6368 8276
rect 5123 8245 5135 8248
rect 5077 8239 5135 8245
rect 6362 8236 6368 8248
rect 6420 8236 6426 8288
rect 6638 8236 6644 8288
rect 6696 8276 6702 8288
rect 6840 8276 6868 8316
rect 6914 8304 6920 8316
rect 6972 8344 6978 8356
rect 7070 8347 7128 8353
rect 7070 8344 7082 8347
rect 6972 8316 7082 8344
rect 6972 8304 6978 8316
rect 7070 8313 7082 8316
rect 7116 8313 7128 8347
rect 7070 8307 7128 8313
rect 9122 8304 9128 8356
rect 9180 8344 9186 8356
rect 10134 8344 10140 8356
rect 9180 8316 10140 8344
rect 9180 8304 9186 8316
rect 10134 8304 10140 8316
rect 10192 8344 10198 8356
rect 10413 8347 10471 8353
rect 10413 8344 10425 8347
rect 10192 8316 10425 8344
rect 10192 8304 10198 8316
rect 10413 8313 10425 8316
rect 10459 8313 10471 8347
rect 10413 8307 10471 8313
rect 13970 8347 14028 8353
rect 13970 8313 13982 8347
rect 14016 8313 14028 8347
rect 14752 8344 14780 8384
rect 16022 8372 16028 8424
rect 16080 8412 16086 8424
rect 16577 8415 16635 8421
rect 16577 8412 16589 8415
rect 16080 8384 16589 8412
rect 16080 8372 16086 8384
rect 16577 8381 16589 8384
rect 16623 8381 16635 8415
rect 16577 8375 16635 8381
rect 16666 8344 16672 8356
rect 14752 8316 16344 8344
rect 16627 8316 16672 8344
rect 13970 8307 14028 8313
rect 6696 8248 6868 8276
rect 6696 8236 6702 8248
rect 8570 8236 8576 8288
rect 8628 8276 8634 8288
rect 9398 8276 9404 8288
rect 8628 8248 9404 8276
rect 8628 8236 8634 8248
rect 9398 8236 9404 8248
rect 9456 8276 9462 8288
rect 10686 8276 10692 8288
rect 9456 8248 10692 8276
rect 9456 8236 9462 8248
rect 10686 8236 10692 8248
rect 10744 8236 10750 8288
rect 11054 8236 11060 8288
rect 11112 8276 11118 8288
rect 11238 8276 11244 8288
rect 11112 8248 11244 8276
rect 11112 8236 11118 8248
rect 11238 8236 11244 8248
rect 11296 8276 11302 8288
rect 12069 8279 12127 8285
rect 12069 8276 12081 8279
rect 11296 8248 12081 8276
rect 11296 8236 11302 8248
rect 12069 8245 12081 8248
rect 12115 8276 12127 8279
rect 12526 8276 12532 8288
rect 12115 8248 12532 8276
rect 12115 8245 12127 8248
rect 12069 8239 12127 8245
rect 12526 8236 12532 8248
rect 12584 8276 12590 8288
rect 13538 8276 13544 8288
rect 12584 8248 13544 8276
rect 12584 8236 12590 8248
rect 13538 8236 13544 8248
rect 13596 8236 13602 8288
rect 13722 8236 13728 8288
rect 13780 8276 13786 8288
rect 13985 8276 14013 8307
rect 13780 8248 14013 8276
rect 13780 8236 13786 8248
rect 14642 8236 14648 8288
rect 14700 8276 14706 8288
rect 15105 8279 15163 8285
rect 15105 8276 15117 8279
rect 14700 8248 15117 8276
rect 14700 8236 14706 8248
rect 15105 8245 15117 8248
rect 15151 8245 15163 8279
rect 16206 8276 16212 8288
rect 16167 8248 16212 8276
rect 15105 8239 15163 8245
rect 16206 8236 16212 8248
rect 16264 8236 16270 8288
rect 16316 8276 16344 8316
rect 16666 8304 16672 8316
rect 16724 8304 16730 8356
rect 17788 8285 17816 8452
rect 18598 8440 18604 8452
rect 18656 8440 18662 8492
rect 19426 8480 19432 8492
rect 19387 8452 19432 8480
rect 19426 8440 19432 8452
rect 19484 8440 19490 8492
rect 20180 8489 20208 8520
rect 20990 8508 20996 8520
rect 21048 8508 21054 8560
rect 20165 8483 20223 8489
rect 20165 8449 20177 8483
rect 20211 8449 20223 8483
rect 20165 8443 20223 8449
rect 19058 8372 19064 8424
rect 19116 8412 19122 8424
rect 19981 8415 20039 8421
rect 19981 8412 19993 8415
rect 19116 8384 19993 8412
rect 19116 8372 19122 8384
rect 19981 8381 19993 8384
rect 20027 8381 20039 8415
rect 19981 8375 20039 8381
rect 20073 8415 20131 8421
rect 20073 8381 20085 8415
rect 20119 8412 20131 8415
rect 20438 8412 20444 8424
rect 20119 8384 20444 8412
rect 20119 8381 20131 8384
rect 20073 8375 20131 8381
rect 18417 8347 18475 8353
rect 18417 8313 18429 8347
rect 18463 8344 18475 8347
rect 18782 8344 18788 8356
rect 18463 8316 18788 8344
rect 18463 8313 18475 8316
rect 18417 8307 18475 8313
rect 18782 8304 18788 8316
rect 18840 8304 18846 8356
rect 19334 8304 19340 8356
rect 19392 8344 19398 8356
rect 20088 8344 20116 8375
rect 20438 8372 20444 8384
rect 20496 8372 20502 8424
rect 21008 8412 21036 8508
rect 21174 8440 21180 8492
rect 21232 8480 21238 8492
rect 21729 8483 21787 8489
rect 21729 8480 21741 8483
rect 21232 8452 21741 8480
rect 21232 8440 21238 8452
rect 21729 8449 21741 8452
rect 21775 8449 21787 8483
rect 21729 8443 21787 8449
rect 21545 8415 21603 8421
rect 21545 8412 21557 8415
rect 21008 8384 21557 8412
rect 21545 8381 21557 8384
rect 21591 8381 21603 8415
rect 21545 8375 21603 8381
rect 19392 8316 20116 8344
rect 19392 8304 19398 8316
rect 17773 8279 17831 8285
rect 17773 8276 17785 8279
rect 16316 8248 17785 8276
rect 17773 8245 17785 8248
rect 17819 8245 17831 8279
rect 18046 8276 18052 8288
rect 18007 8248 18052 8276
rect 17773 8239 17831 8245
rect 18046 8236 18052 8248
rect 18104 8236 18110 8288
rect 18509 8279 18567 8285
rect 18509 8245 18521 8279
rect 18555 8276 18567 8279
rect 18690 8276 18696 8288
rect 18555 8248 18696 8276
rect 18555 8245 18567 8248
rect 18509 8239 18567 8245
rect 18690 8236 18696 8248
rect 18748 8236 18754 8288
rect 19518 8236 19524 8288
rect 19576 8276 19582 8288
rect 20625 8279 20683 8285
rect 20625 8276 20637 8279
rect 19576 8248 20637 8276
rect 19576 8236 19582 8248
rect 20625 8245 20637 8248
rect 20671 8245 20683 8279
rect 21634 8276 21640 8288
rect 21595 8248 21640 8276
rect 20625 8239 20683 8245
rect 21634 8236 21640 8248
rect 21692 8236 21698 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1673 8075 1731 8081
rect 1673 8041 1685 8075
rect 1719 8072 1731 8075
rect 2222 8072 2228 8084
rect 1719 8044 2228 8072
rect 1719 8041 1731 8044
rect 1673 8035 1731 8041
rect 2222 8032 2228 8044
rect 2280 8032 2286 8084
rect 2406 8072 2412 8084
rect 2367 8044 2412 8072
rect 2406 8032 2412 8044
rect 2464 8032 2470 8084
rect 3513 8075 3571 8081
rect 3513 8041 3525 8075
rect 3559 8072 3571 8075
rect 3602 8072 3608 8084
rect 3559 8044 3608 8072
rect 3559 8041 3571 8044
rect 3513 8035 3571 8041
rect 3602 8032 3608 8044
rect 3660 8032 3666 8084
rect 3878 8072 3884 8084
rect 3839 8044 3884 8072
rect 3878 8032 3884 8044
rect 3936 8032 3942 8084
rect 4614 8072 4620 8084
rect 4575 8044 4620 8072
rect 4614 8032 4620 8044
rect 4672 8032 4678 8084
rect 7285 8075 7343 8081
rect 7285 8041 7297 8075
rect 7331 8072 7343 8075
rect 8202 8072 8208 8084
rect 7331 8044 8208 8072
rect 7331 8041 7343 8044
rect 7285 8035 7343 8041
rect 8202 8032 8208 8044
rect 8260 8032 8266 8084
rect 8846 8072 8852 8084
rect 8807 8044 8852 8072
rect 8846 8032 8852 8044
rect 8904 8032 8910 8084
rect 10134 8072 10140 8084
rect 10095 8044 10140 8072
rect 10134 8032 10140 8044
rect 10192 8032 10198 8084
rect 11057 8075 11115 8081
rect 11057 8041 11069 8075
rect 11103 8072 11115 8075
rect 12342 8072 12348 8084
rect 11103 8044 12348 8072
rect 11103 8041 11115 8044
rect 11057 8035 11115 8041
rect 12342 8032 12348 8044
rect 12400 8032 12406 8084
rect 13541 8075 13599 8081
rect 13541 8041 13553 8075
rect 13587 8072 13599 8075
rect 14274 8072 14280 8084
rect 13587 8044 14280 8072
rect 13587 8041 13599 8044
rect 13541 8035 13599 8041
rect 14274 8032 14280 8044
rect 14332 8032 14338 8084
rect 15102 8072 15108 8084
rect 15063 8044 15108 8072
rect 15102 8032 15108 8044
rect 15160 8032 15166 8084
rect 19058 8072 19064 8084
rect 16132 8044 17172 8072
rect 19019 8044 19064 8072
rect 2866 8004 2872 8016
rect 2827 7976 2872 8004
rect 2866 7964 2872 7976
rect 2924 7964 2930 8016
rect 6822 8004 6828 8016
rect 5276 7976 6828 8004
rect 2774 7896 2780 7948
rect 2832 7936 2838 7948
rect 5276 7945 5304 7976
rect 6822 7964 6828 7976
rect 6880 7964 6886 8016
rect 13814 7964 13820 8016
rect 13872 8004 13878 8016
rect 14001 8007 14059 8013
rect 14001 8004 14013 8007
rect 13872 7976 14013 8004
rect 13872 7964 13878 7976
rect 14001 7973 14013 7976
rect 14047 7973 14059 8007
rect 14001 7967 14059 7973
rect 14921 8007 14979 8013
rect 14921 7973 14933 8007
rect 14967 8004 14979 8007
rect 16132 8004 16160 8044
rect 17034 8004 17040 8016
rect 14967 7976 16160 8004
rect 16684 7976 17040 8004
rect 14967 7973 14979 7976
rect 14921 7967 14979 7973
rect 5534 7945 5540 7948
rect 4065 7939 4123 7945
rect 4065 7936 4077 7939
rect 2832 7908 4077 7936
rect 2832 7896 2838 7908
rect 4065 7905 4077 7908
rect 4111 7905 4123 7939
rect 4065 7899 4123 7905
rect 5261 7939 5319 7945
rect 5261 7905 5273 7939
rect 5307 7905 5319 7939
rect 5528 7936 5540 7945
rect 5495 7908 5540 7936
rect 5261 7899 5319 7905
rect 5528 7899 5540 7908
rect 5534 7896 5540 7899
rect 5592 7896 5598 7948
rect 8110 7936 8116 7948
rect 8071 7908 8116 7936
rect 8110 7896 8116 7908
rect 8168 7896 8174 7948
rect 9674 7936 9680 7948
rect 9635 7908 9680 7936
rect 9674 7896 9680 7908
rect 9732 7896 9738 7948
rect 11149 7939 11207 7945
rect 11149 7905 11161 7939
rect 11195 7936 11207 7939
rect 11238 7936 11244 7948
rect 11195 7908 11244 7936
rect 11195 7905 11207 7908
rect 11149 7899 11207 7905
rect 11238 7896 11244 7908
rect 11296 7896 11302 7948
rect 11416 7939 11474 7945
rect 11416 7905 11428 7939
rect 11462 7936 11474 7939
rect 12342 7936 12348 7948
rect 11462 7908 12348 7936
rect 11462 7905 11474 7908
rect 11416 7899 11474 7905
rect 12342 7896 12348 7908
rect 12400 7936 12406 7948
rect 12434 7936 12440 7948
rect 12400 7908 12440 7936
rect 12400 7896 12406 7908
rect 12434 7896 12440 7908
rect 12492 7896 12498 7948
rect 14734 7896 14740 7948
rect 14792 7936 14798 7948
rect 15289 7939 15347 7945
rect 15289 7936 15301 7939
rect 14792 7908 15301 7936
rect 14792 7896 14798 7908
rect 15289 7905 15301 7908
rect 15335 7936 15347 7939
rect 15746 7936 15752 7948
rect 15335 7908 15752 7936
rect 15335 7905 15347 7908
rect 15289 7899 15347 7905
rect 15746 7896 15752 7908
rect 15804 7896 15810 7948
rect 16684 7945 16712 7976
rect 17034 7964 17040 7976
rect 17092 7964 17098 8016
rect 16669 7939 16727 7945
rect 16669 7905 16681 7939
rect 16715 7905 16727 7939
rect 16669 7899 16727 7905
rect 16758 7896 16764 7948
rect 16816 7936 16822 7948
rect 16925 7939 16983 7945
rect 16925 7936 16937 7939
rect 16816 7908 16937 7936
rect 16816 7896 16822 7908
rect 16925 7905 16937 7908
rect 16971 7905 16983 7939
rect 17144 7936 17172 8044
rect 19058 8032 19064 8044
rect 19116 8032 19122 8084
rect 19153 8075 19211 8081
rect 19153 8041 19165 8075
rect 19199 8072 19211 8075
rect 19242 8072 19248 8084
rect 19199 8044 19248 8072
rect 19199 8041 19211 8044
rect 19153 8035 19211 8041
rect 19242 8032 19248 8044
rect 19300 8032 19306 8084
rect 19521 8075 19579 8081
rect 19521 8041 19533 8075
rect 19567 8072 19579 8075
rect 19978 8072 19984 8084
rect 19567 8044 19984 8072
rect 19567 8041 19579 8044
rect 19521 8035 19579 8041
rect 19978 8032 19984 8044
rect 20036 8032 20042 8084
rect 18874 7964 18880 8016
rect 18932 8004 18938 8016
rect 19613 8007 19671 8013
rect 19613 8004 19625 8007
rect 18932 7976 19625 8004
rect 18932 7964 18938 7976
rect 19613 7973 19625 7976
rect 19659 7973 19671 8007
rect 19613 7967 19671 7973
rect 21177 7939 21235 7945
rect 21177 7936 21189 7939
rect 17144 7908 21189 7936
rect 16925 7899 16983 7905
rect 21177 7905 21189 7908
rect 21223 7936 21235 7939
rect 21634 7936 21640 7948
rect 21223 7908 21640 7936
rect 21223 7905 21235 7908
rect 21177 7899 21235 7905
rect 21634 7896 21640 7908
rect 21692 7896 21698 7948
rect 2958 7868 2964 7880
rect 2919 7840 2964 7868
rect 2958 7828 2964 7840
rect 3016 7828 3022 7880
rect 7834 7828 7840 7880
rect 7892 7868 7898 7880
rect 8205 7871 8263 7877
rect 8205 7868 8217 7871
rect 7892 7840 8217 7868
rect 7892 7828 7898 7840
rect 8205 7837 8217 7840
rect 8251 7837 8263 7871
rect 8205 7831 8263 7837
rect 8389 7871 8447 7877
rect 8389 7837 8401 7871
rect 8435 7868 8447 7871
rect 8662 7868 8668 7880
rect 8435 7840 8668 7868
rect 8435 7837 8447 7840
rect 8389 7831 8447 7837
rect 8662 7828 8668 7840
rect 8720 7828 8726 7880
rect 13354 7868 13360 7880
rect 12544 7840 13360 7868
rect 1302 7760 1308 7812
rect 1360 7800 1366 7812
rect 4706 7800 4712 7812
rect 1360 7772 4712 7800
rect 1360 7760 1366 7772
rect 4706 7760 4712 7772
rect 4764 7800 4770 7812
rect 4893 7803 4951 7809
rect 4893 7800 4905 7803
rect 4764 7772 4905 7800
rect 4764 7760 4770 7772
rect 4893 7769 4905 7772
rect 4939 7769 4951 7803
rect 4893 7763 4951 7769
rect 7006 7760 7012 7812
rect 7064 7800 7070 7812
rect 7745 7803 7803 7809
rect 7745 7800 7757 7803
rect 7064 7772 7757 7800
rect 7064 7760 7070 7772
rect 7745 7769 7757 7772
rect 7791 7769 7803 7803
rect 9306 7800 9312 7812
rect 9267 7772 9312 7800
rect 7745 7763 7803 7769
rect 9306 7760 9312 7772
rect 9364 7760 9370 7812
rect 2314 7732 2320 7744
rect 2275 7704 2320 7732
rect 2314 7692 2320 7704
rect 2372 7732 2378 7744
rect 2682 7732 2688 7744
rect 2372 7704 2688 7732
rect 2372 7692 2378 7704
rect 2682 7692 2688 7704
rect 2740 7692 2746 7744
rect 6638 7732 6644 7744
rect 6599 7704 6644 7732
rect 6638 7692 6644 7704
rect 6696 7692 6702 7744
rect 7558 7732 7564 7744
rect 7519 7704 7564 7732
rect 7558 7692 7564 7704
rect 7616 7692 7622 7744
rect 10686 7692 10692 7744
rect 10744 7732 10750 7744
rect 10781 7735 10839 7741
rect 10781 7732 10793 7735
rect 10744 7704 10793 7732
rect 10744 7692 10750 7704
rect 10781 7701 10793 7704
rect 10827 7732 10839 7735
rect 11057 7735 11115 7741
rect 11057 7732 11069 7735
rect 10827 7704 11069 7732
rect 10827 7701 10839 7704
rect 10781 7695 10839 7701
rect 11057 7701 11069 7704
rect 11103 7701 11115 7735
rect 11057 7695 11115 7701
rect 12066 7692 12072 7744
rect 12124 7732 12130 7744
rect 12544 7741 12572 7840
rect 13354 7828 13360 7840
rect 13412 7828 13418 7880
rect 14093 7871 14151 7877
rect 14093 7837 14105 7871
rect 14139 7837 14151 7871
rect 14274 7868 14280 7880
rect 14235 7840 14280 7868
rect 14093 7831 14151 7837
rect 13173 7803 13231 7809
rect 13173 7769 13185 7803
rect 13219 7800 13231 7803
rect 13630 7800 13636 7812
rect 13219 7772 13636 7800
rect 13219 7769 13231 7772
rect 13173 7763 13231 7769
rect 13630 7760 13636 7772
rect 13688 7760 13694 7812
rect 14108 7800 14136 7831
rect 14274 7828 14280 7840
rect 14332 7828 14338 7880
rect 14645 7871 14703 7877
rect 14645 7837 14657 7871
rect 14691 7868 14703 7871
rect 15378 7868 15384 7880
rect 14691 7840 15384 7868
rect 14691 7837 14703 7840
rect 14645 7831 14703 7837
rect 15378 7828 15384 7840
rect 15436 7828 15442 7880
rect 19705 7871 19763 7877
rect 19705 7837 19717 7871
rect 19751 7837 19763 7871
rect 19705 7831 19763 7837
rect 14921 7803 14979 7809
rect 14921 7800 14933 7803
rect 14108 7772 14933 7800
rect 12529 7735 12587 7741
rect 12529 7732 12541 7735
rect 12124 7704 12541 7732
rect 12124 7692 12130 7704
rect 12529 7701 12541 7704
rect 12575 7701 12587 7735
rect 12529 7695 12587 7701
rect 13262 7692 13268 7744
rect 13320 7732 13326 7744
rect 14108 7732 14136 7772
rect 14921 7769 14933 7772
rect 14967 7769 14979 7803
rect 14921 7763 14979 7769
rect 15473 7803 15531 7809
rect 15473 7769 15485 7803
rect 15519 7800 15531 7803
rect 16390 7800 16396 7812
rect 15519 7772 16396 7800
rect 15519 7769 15531 7772
rect 15473 7763 15531 7769
rect 16390 7760 16396 7772
rect 16448 7760 16454 7812
rect 19518 7760 19524 7812
rect 19576 7800 19582 7812
rect 19720 7800 19748 7831
rect 19576 7772 19748 7800
rect 19576 7760 19582 7772
rect 13320 7704 14136 7732
rect 13320 7692 13326 7704
rect 15286 7692 15292 7744
rect 15344 7732 15350 7744
rect 15841 7735 15899 7741
rect 15841 7732 15853 7735
rect 15344 7704 15853 7732
rect 15344 7692 15350 7704
rect 15841 7701 15853 7704
rect 15887 7701 15899 7735
rect 15841 7695 15899 7701
rect 16022 7692 16028 7744
rect 16080 7732 16086 7744
rect 16209 7735 16267 7741
rect 16209 7732 16221 7735
rect 16080 7704 16221 7732
rect 16080 7692 16086 7704
rect 16209 7701 16221 7704
rect 16255 7732 16267 7735
rect 16666 7732 16672 7744
rect 16255 7704 16672 7732
rect 16255 7701 16267 7704
rect 16209 7695 16267 7701
rect 16666 7692 16672 7704
rect 16724 7692 16730 7744
rect 18049 7735 18107 7741
rect 18049 7701 18061 7735
rect 18095 7732 18107 7735
rect 18138 7732 18144 7744
rect 18095 7704 18144 7732
rect 18095 7701 18107 7704
rect 18049 7695 18107 7701
rect 18138 7692 18144 7704
rect 18196 7692 18202 7744
rect 18690 7732 18696 7744
rect 18651 7704 18696 7732
rect 18690 7692 18696 7704
rect 18748 7692 18754 7744
rect 20070 7692 20076 7744
rect 20128 7732 20134 7744
rect 20165 7735 20223 7741
rect 20165 7732 20177 7735
rect 20128 7704 20177 7732
rect 20128 7692 20134 7704
rect 20165 7701 20177 7704
rect 20211 7701 20223 7735
rect 20530 7732 20536 7744
rect 20491 7704 20536 7732
rect 20165 7695 20223 7701
rect 20530 7692 20536 7704
rect 20588 7692 20594 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 1670 7528 1676 7540
rect 1631 7500 1676 7528
rect 1670 7488 1676 7500
rect 1728 7488 1734 7540
rect 2958 7488 2964 7540
rect 3016 7528 3022 7540
rect 4157 7531 4215 7537
rect 4157 7528 4169 7531
rect 3016 7500 4169 7528
rect 3016 7488 3022 7500
rect 4157 7497 4169 7500
rect 4203 7497 4215 7531
rect 4157 7491 4215 7497
rect 6273 7531 6331 7537
rect 6273 7497 6285 7531
rect 6319 7528 6331 7531
rect 6454 7528 6460 7540
rect 6319 7500 6460 7528
rect 6319 7497 6331 7500
rect 6273 7491 6331 7497
rect 6454 7488 6460 7500
rect 6512 7488 6518 7540
rect 6641 7531 6699 7537
rect 6641 7497 6653 7531
rect 6687 7528 6699 7531
rect 6730 7528 6736 7540
rect 6687 7500 6736 7528
rect 6687 7497 6699 7500
rect 6641 7491 6699 7497
rect 6730 7488 6736 7500
rect 6788 7488 6794 7540
rect 7834 7528 7840 7540
rect 7795 7500 7840 7528
rect 7834 7488 7840 7500
rect 7892 7488 7898 7540
rect 8662 7528 8668 7540
rect 8623 7500 8668 7528
rect 8662 7488 8668 7500
rect 8720 7488 8726 7540
rect 11885 7531 11943 7537
rect 11885 7497 11897 7531
rect 11931 7528 11943 7531
rect 12342 7528 12348 7540
rect 11931 7500 12348 7528
rect 11931 7497 11943 7500
rect 11885 7491 11943 7497
rect 12342 7488 12348 7500
rect 12400 7488 12406 7540
rect 13081 7531 13139 7537
rect 13081 7497 13093 7531
rect 13127 7528 13139 7531
rect 13170 7528 13176 7540
rect 13127 7500 13176 7528
rect 13127 7497 13139 7500
rect 13081 7491 13139 7497
rect 13170 7488 13176 7500
rect 13228 7488 13234 7540
rect 13814 7488 13820 7540
rect 13872 7528 13878 7540
rect 14185 7531 14243 7537
rect 14185 7528 14197 7531
rect 13872 7500 14197 7528
rect 13872 7488 13878 7500
rect 14185 7497 14197 7500
rect 14231 7528 14243 7531
rect 16666 7528 16672 7540
rect 14231 7500 16672 7528
rect 14231 7497 14243 7500
rect 14185 7491 14243 7497
rect 16666 7488 16672 7500
rect 16724 7488 16730 7540
rect 18874 7488 18880 7540
rect 18932 7528 18938 7540
rect 19061 7531 19119 7537
rect 19061 7528 19073 7531
rect 18932 7500 19073 7528
rect 18932 7488 18938 7500
rect 19061 7497 19073 7500
rect 19107 7497 19119 7531
rect 19610 7528 19616 7540
rect 19571 7500 19616 7528
rect 19061 7491 19119 7497
rect 19610 7488 19616 7500
rect 19668 7488 19674 7540
rect 20714 7488 20720 7540
rect 20772 7528 20778 7540
rect 21177 7531 21235 7537
rect 21177 7528 21189 7531
rect 20772 7500 21189 7528
rect 20772 7488 20778 7500
rect 21177 7497 21189 7500
rect 21223 7497 21235 7531
rect 21177 7491 21235 7497
rect 3605 7463 3663 7469
rect 3605 7460 3617 7463
rect 3232 7432 3617 7460
rect 1578 7352 1584 7404
rect 1636 7392 1642 7404
rect 2038 7392 2044 7404
rect 1636 7364 2044 7392
rect 1636 7352 1642 7364
rect 2038 7352 2044 7364
rect 2096 7392 2102 7404
rect 2225 7395 2283 7401
rect 2225 7392 2237 7395
rect 2096 7364 2237 7392
rect 2096 7352 2102 7364
rect 2225 7361 2237 7364
rect 2271 7361 2283 7395
rect 2225 7355 2283 7361
rect 2314 7284 2320 7336
rect 2372 7324 2378 7336
rect 2481 7327 2539 7333
rect 2481 7324 2493 7327
rect 2372 7296 2493 7324
rect 2372 7284 2378 7296
rect 2481 7293 2493 7296
rect 2527 7293 2539 7327
rect 2481 7287 2539 7293
rect 2958 7284 2964 7336
rect 3016 7324 3022 7336
rect 3232 7324 3260 7432
rect 3605 7429 3617 7432
rect 3651 7460 3663 7463
rect 3970 7460 3976 7472
rect 3651 7432 3976 7460
rect 3651 7429 3663 7432
rect 3605 7423 3663 7429
rect 3970 7420 3976 7432
rect 4028 7420 4034 7472
rect 5166 7460 5172 7472
rect 5127 7432 5172 7460
rect 5166 7420 5172 7432
rect 5224 7420 5230 7472
rect 11146 7460 11152 7472
rect 9876 7432 11152 7460
rect 5813 7395 5871 7401
rect 5813 7361 5825 7395
rect 5859 7392 5871 7395
rect 6086 7392 6092 7404
rect 5859 7364 6092 7392
rect 5859 7361 5871 7364
rect 5813 7355 5871 7361
rect 6086 7352 6092 7364
rect 6144 7352 6150 7404
rect 7374 7392 7380 7404
rect 7335 7364 7380 7392
rect 7374 7352 7380 7364
rect 7432 7352 7438 7404
rect 8662 7352 8668 7404
rect 8720 7392 8726 7404
rect 9876 7401 9904 7432
rect 11146 7420 11152 7432
rect 11204 7420 11210 7472
rect 9125 7395 9183 7401
rect 9125 7392 9137 7395
rect 8720 7364 9137 7392
rect 8720 7352 8726 7364
rect 9125 7361 9137 7364
rect 9171 7392 9183 7395
rect 9861 7395 9919 7401
rect 9861 7392 9873 7395
rect 9171 7364 9873 7392
rect 9171 7361 9183 7364
rect 9125 7355 9183 7361
rect 9861 7361 9873 7364
rect 9907 7361 9919 7395
rect 9861 7355 9919 7361
rect 10321 7395 10379 7401
rect 10321 7361 10333 7395
rect 10367 7392 10379 7395
rect 11333 7395 11391 7401
rect 11333 7392 11345 7395
rect 10367 7364 11345 7392
rect 10367 7361 10379 7364
rect 10321 7355 10379 7361
rect 11333 7361 11345 7364
rect 11379 7392 11391 7395
rect 12802 7392 12808 7404
rect 11379 7364 12808 7392
rect 11379 7361 11391 7364
rect 11333 7355 11391 7361
rect 12802 7352 12808 7364
rect 12860 7352 12866 7404
rect 13630 7392 13636 7404
rect 13591 7364 13636 7392
rect 13630 7352 13636 7364
rect 13688 7352 13694 7404
rect 13817 7395 13875 7401
rect 13817 7361 13829 7395
rect 13863 7361 13875 7395
rect 13817 7355 13875 7361
rect 17865 7395 17923 7401
rect 17865 7361 17877 7395
rect 17911 7392 17923 7395
rect 18414 7392 18420 7404
rect 17911 7364 18420 7392
rect 17911 7361 17923 7364
rect 17865 7355 17923 7361
rect 3016 7296 3260 7324
rect 3016 7284 3022 7296
rect 3418 7284 3424 7336
rect 3476 7324 3482 7336
rect 4338 7324 4344 7336
rect 3476 7296 4344 7324
rect 3476 7284 3482 7296
rect 4338 7284 4344 7296
rect 4396 7324 4402 7336
rect 4985 7327 5043 7333
rect 4985 7324 4997 7327
rect 4396 7296 4997 7324
rect 4396 7284 4402 7296
rect 4985 7293 4997 7296
rect 5031 7324 5043 7327
rect 5629 7327 5687 7333
rect 5629 7324 5641 7327
rect 5031 7296 5641 7324
rect 5031 7293 5043 7296
rect 4985 7287 5043 7293
rect 5629 7293 5641 7296
rect 5675 7293 5687 7327
rect 5629 7287 5687 7293
rect 6730 7284 6736 7336
rect 6788 7324 6794 7336
rect 7193 7327 7251 7333
rect 7193 7324 7205 7327
rect 6788 7296 7205 7324
rect 6788 7284 6794 7296
rect 7193 7293 7205 7296
rect 7239 7293 7251 7327
rect 7193 7287 7251 7293
rect 9582 7284 9588 7336
rect 9640 7324 9646 7336
rect 9677 7327 9735 7333
rect 9677 7324 9689 7327
rect 9640 7296 9689 7324
rect 9640 7284 9646 7296
rect 9677 7293 9689 7296
rect 9723 7293 9735 7327
rect 9677 7287 9735 7293
rect 10505 7327 10563 7333
rect 10505 7293 10517 7327
rect 10551 7324 10563 7327
rect 11241 7327 11299 7333
rect 11241 7324 11253 7327
rect 10551 7296 11253 7324
rect 10551 7293 10563 7296
rect 10505 7287 10563 7293
rect 11241 7293 11253 7296
rect 11287 7293 11299 7327
rect 11241 7287 11299 7293
rect 12713 7327 12771 7333
rect 12713 7293 12725 7327
rect 12759 7324 12771 7327
rect 13722 7324 13728 7336
rect 12759 7296 13728 7324
rect 12759 7293 12771 7296
rect 12713 7287 12771 7293
rect 13722 7284 13728 7296
rect 13780 7324 13786 7336
rect 13832 7324 13860 7355
rect 18414 7352 18420 7364
rect 18472 7392 18478 7404
rect 18601 7395 18659 7401
rect 18601 7392 18613 7395
rect 18472 7364 18613 7392
rect 18472 7352 18478 7364
rect 18601 7361 18613 7364
rect 18647 7361 18659 7395
rect 18601 7355 18659 7361
rect 19518 7352 19524 7404
rect 19576 7392 19582 7404
rect 20165 7395 20223 7401
rect 20165 7392 20177 7395
rect 19576 7364 20177 7392
rect 19576 7352 19582 7364
rect 20165 7361 20177 7364
rect 20211 7392 20223 7395
rect 20625 7395 20683 7401
rect 20625 7392 20637 7395
rect 20211 7364 20637 7392
rect 20211 7361 20223 7364
rect 20165 7355 20223 7361
rect 20625 7361 20637 7364
rect 20671 7361 20683 7395
rect 20990 7392 20996 7404
rect 20951 7364 20996 7392
rect 20625 7355 20683 7361
rect 20990 7352 20996 7364
rect 21048 7392 21054 7404
rect 21729 7395 21787 7401
rect 21729 7392 21741 7395
rect 21048 7364 21741 7392
rect 21048 7352 21054 7364
rect 21729 7361 21741 7364
rect 21775 7361 21787 7395
rect 21729 7355 21787 7361
rect 14642 7324 14648 7336
rect 13780 7296 13860 7324
rect 14603 7296 14648 7324
rect 13780 7284 13786 7296
rect 14642 7284 14648 7296
rect 14700 7284 14706 7336
rect 14737 7327 14795 7333
rect 14737 7293 14749 7327
rect 14783 7324 14795 7327
rect 17034 7324 17040 7336
rect 14783 7296 17040 7324
rect 14783 7293 14795 7296
rect 14737 7287 14795 7293
rect 17034 7284 17040 7296
rect 17092 7284 17098 7336
rect 17402 7324 17408 7336
rect 17363 7296 17408 7324
rect 17402 7284 17408 7296
rect 17460 7284 17466 7336
rect 5537 7259 5595 7265
rect 5537 7256 5549 7259
rect 4632 7228 5549 7256
rect 1118 7148 1124 7200
rect 1176 7188 1182 7200
rect 2041 7191 2099 7197
rect 2041 7188 2053 7191
rect 1176 7160 2053 7188
rect 1176 7148 1182 7160
rect 2041 7157 2053 7160
rect 2087 7188 2099 7191
rect 2866 7188 2872 7200
rect 2087 7160 2872 7188
rect 2087 7157 2099 7160
rect 2041 7151 2099 7157
rect 2866 7148 2872 7160
rect 2924 7148 2930 7200
rect 3694 7148 3700 7200
rect 3752 7188 3758 7200
rect 4632 7197 4660 7228
rect 5537 7225 5549 7228
rect 5583 7256 5595 7259
rect 5994 7256 6000 7268
rect 5583 7228 6000 7256
rect 5583 7225 5595 7228
rect 5537 7219 5595 7225
rect 5994 7216 6000 7228
rect 6052 7216 6058 7268
rect 6454 7216 6460 7268
rect 6512 7256 6518 7268
rect 7285 7259 7343 7265
rect 7285 7256 7297 7259
rect 6512 7228 7297 7256
rect 6512 7216 6518 7228
rect 7285 7225 7297 7228
rect 7331 7225 7343 7259
rect 7285 7219 7343 7225
rect 9306 7216 9312 7268
rect 9364 7256 9370 7268
rect 9364 7228 9628 7256
rect 9364 7216 9370 7228
rect 4617 7191 4675 7197
rect 4617 7188 4629 7191
rect 3752 7160 4629 7188
rect 3752 7148 3758 7160
rect 4617 7157 4629 7160
rect 4663 7157 4675 7191
rect 6822 7188 6828 7200
rect 6783 7160 6828 7188
rect 4617 7151 4675 7157
rect 6822 7148 6828 7160
rect 6880 7148 6886 7200
rect 8202 7188 8208 7200
rect 8163 7160 8208 7188
rect 8202 7148 8208 7160
rect 8260 7148 8266 7200
rect 9217 7191 9275 7197
rect 9217 7157 9229 7191
rect 9263 7188 9275 7191
rect 9490 7188 9496 7200
rect 9263 7160 9496 7188
rect 9263 7157 9275 7160
rect 9217 7151 9275 7157
rect 9490 7148 9496 7160
rect 9548 7148 9554 7200
rect 9600 7197 9628 7228
rect 10134 7216 10140 7268
rect 10192 7256 10198 7268
rect 10686 7256 10692 7268
rect 10192 7228 10692 7256
rect 10192 7216 10198 7228
rect 10686 7216 10692 7228
rect 10744 7256 10750 7268
rect 11149 7259 11207 7265
rect 11149 7256 11161 7259
rect 10744 7228 11161 7256
rect 10744 7216 10750 7228
rect 11149 7225 11161 7228
rect 11195 7225 11207 7259
rect 11149 7219 11207 7225
rect 14090 7216 14096 7268
rect 14148 7256 14154 7268
rect 14660 7256 14688 7284
rect 14982 7259 15040 7265
rect 14982 7256 14994 7259
rect 14148 7228 14994 7256
rect 14148 7216 14154 7228
rect 14982 7225 14994 7228
rect 15028 7225 15040 7259
rect 14982 7219 15040 7225
rect 16574 7216 16580 7268
rect 16632 7256 16638 7268
rect 17129 7259 17187 7265
rect 17129 7256 17141 7259
rect 16632 7228 17141 7256
rect 16632 7216 16638 7228
rect 17129 7225 17141 7228
rect 17175 7256 17187 7259
rect 18417 7259 18475 7265
rect 18417 7256 18429 7259
rect 17175 7228 18429 7256
rect 17175 7225 17187 7228
rect 17129 7219 17187 7225
rect 18417 7225 18429 7228
rect 18463 7225 18475 7259
rect 18417 7219 18475 7225
rect 19521 7259 19579 7265
rect 19521 7225 19533 7259
rect 19567 7256 19579 7259
rect 19981 7259 20039 7265
rect 19981 7256 19993 7259
rect 19567 7228 19993 7256
rect 19567 7225 19579 7228
rect 19521 7219 19579 7225
rect 19981 7225 19993 7228
rect 20027 7256 20039 7259
rect 20162 7256 20168 7268
rect 20027 7228 20168 7256
rect 20027 7225 20039 7228
rect 19981 7219 20039 7225
rect 20162 7216 20168 7228
rect 20220 7216 20226 7268
rect 21174 7216 21180 7268
rect 21232 7256 21238 7268
rect 21637 7259 21695 7265
rect 21637 7256 21649 7259
rect 21232 7228 21649 7256
rect 21232 7216 21238 7228
rect 21637 7225 21649 7228
rect 21683 7225 21695 7259
rect 21637 7219 21695 7225
rect 9585 7191 9643 7197
rect 9585 7157 9597 7191
rect 9631 7157 9643 7191
rect 9585 7151 9643 7157
rect 9858 7148 9864 7200
rect 9916 7188 9922 7200
rect 10505 7191 10563 7197
rect 10505 7188 10517 7191
rect 9916 7160 10517 7188
rect 9916 7148 9922 7160
rect 10505 7157 10517 7160
rect 10551 7188 10563 7191
rect 10597 7191 10655 7197
rect 10597 7188 10609 7191
rect 10551 7160 10609 7188
rect 10551 7157 10563 7160
rect 10505 7151 10563 7157
rect 10597 7157 10609 7160
rect 10643 7157 10655 7191
rect 10597 7151 10655 7157
rect 10781 7191 10839 7197
rect 10781 7157 10793 7191
rect 10827 7188 10839 7191
rect 10962 7188 10968 7200
rect 10827 7160 10968 7188
rect 10827 7157 10839 7160
rect 10781 7151 10839 7157
rect 10962 7148 10968 7160
rect 11020 7148 11026 7200
rect 11974 7148 11980 7200
rect 12032 7188 12038 7200
rect 12161 7191 12219 7197
rect 12161 7188 12173 7191
rect 12032 7160 12173 7188
rect 12032 7148 12038 7160
rect 12161 7157 12173 7160
rect 12207 7157 12219 7191
rect 13170 7188 13176 7200
rect 13131 7160 13176 7188
rect 12161 7151 12219 7157
rect 13170 7148 13176 7160
rect 13228 7148 13234 7200
rect 13538 7188 13544 7200
rect 13499 7160 13544 7188
rect 13538 7148 13544 7160
rect 13596 7148 13602 7200
rect 15378 7148 15384 7200
rect 15436 7188 15442 7200
rect 16117 7191 16175 7197
rect 16117 7188 16129 7191
rect 15436 7160 16129 7188
rect 15436 7148 15442 7160
rect 16117 7157 16129 7160
rect 16163 7188 16175 7191
rect 16669 7191 16727 7197
rect 16669 7188 16681 7191
rect 16163 7160 16681 7188
rect 16163 7157 16175 7160
rect 16117 7151 16175 7157
rect 16669 7157 16681 7160
rect 16715 7188 16727 7191
rect 16758 7188 16764 7200
rect 16715 7160 16764 7188
rect 16715 7157 16727 7160
rect 16669 7151 16727 7157
rect 16758 7148 16764 7160
rect 16816 7148 16822 7200
rect 17034 7148 17040 7200
rect 17092 7188 17098 7200
rect 17221 7191 17279 7197
rect 17221 7188 17233 7191
rect 17092 7160 17233 7188
rect 17092 7148 17098 7160
rect 17221 7157 17233 7160
rect 17267 7157 17279 7191
rect 18046 7188 18052 7200
rect 18007 7160 18052 7188
rect 17221 7151 17279 7157
rect 18046 7148 18052 7160
rect 18104 7148 18110 7200
rect 18506 7188 18512 7200
rect 18467 7160 18512 7188
rect 18506 7148 18512 7160
rect 18564 7148 18570 7200
rect 20070 7188 20076 7200
rect 20031 7160 20076 7188
rect 20070 7148 20076 7160
rect 20128 7148 20134 7200
rect 21542 7188 21548 7200
rect 21503 7160 21548 7188
rect 21542 7148 21548 7160
rect 21600 7148 21606 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 1670 6944 1676 6996
rect 1728 6984 1734 6996
rect 1765 6987 1823 6993
rect 1765 6984 1777 6987
rect 1728 6956 1777 6984
rect 1728 6944 1734 6956
rect 1765 6953 1777 6956
rect 1811 6953 1823 6987
rect 1765 6947 1823 6953
rect 2774 6944 2780 6996
rect 2832 6984 2838 6996
rect 7101 6987 7159 6993
rect 2832 6956 2877 6984
rect 2832 6944 2838 6956
rect 7101 6953 7113 6987
rect 7147 6984 7159 6987
rect 7374 6984 7380 6996
rect 7147 6956 7380 6984
rect 7147 6953 7159 6956
rect 7101 6947 7159 6953
rect 7374 6944 7380 6956
rect 7432 6944 7438 6996
rect 8662 6984 8668 6996
rect 8623 6956 8668 6984
rect 8662 6944 8668 6956
rect 8720 6944 8726 6996
rect 9309 6987 9367 6993
rect 9309 6953 9321 6987
rect 9355 6984 9367 6987
rect 9582 6984 9588 6996
rect 9355 6956 9588 6984
rect 9355 6953 9367 6956
rect 9309 6947 9367 6953
rect 9582 6944 9588 6956
rect 9640 6944 9646 6996
rect 11054 6944 11060 6996
rect 11112 6984 11118 6996
rect 11609 6987 11667 6993
rect 11609 6984 11621 6987
rect 11112 6956 11621 6984
rect 11112 6944 11118 6956
rect 11609 6953 11621 6956
rect 11655 6984 11667 6987
rect 11974 6984 11980 6996
rect 11655 6956 11980 6984
rect 11655 6953 11667 6956
rect 11609 6947 11667 6953
rect 11974 6944 11980 6956
rect 12032 6944 12038 6996
rect 12805 6987 12863 6993
rect 12805 6953 12817 6987
rect 12851 6984 12863 6987
rect 12897 6987 12955 6993
rect 12897 6984 12909 6987
rect 12851 6956 12909 6984
rect 12851 6953 12863 6956
rect 12805 6947 12863 6953
rect 12897 6953 12909 6956
rect 12943 6984 12955 6987
rect 13538 6984 13544 6996
rect 12943 6956 13544 6984
rect 12943 6953 12955 6956
rect 12897 6947 12955 6953
rect 13538 6944 13544 6956
rect 13596 6944 13602 6996
rect 14001 6987 14059 6993
rect 14001 6953 14013 6987
rect 14047 6984 14059 6987
rect 14274 6984 14280 6996
rect 14047 6956 14280 6984
rect 14047 6953 14059 6956
rect 14001 6947 14059 6953
rect 1486 6876 1492 6928
rect 1544 6916 1550 6928
rect 1857 6919 1915 6925
rect 1857 6916 1869 6919
rect 1544 6888 1869 6916
rect 1544 6876 1550 6888
rect 1857 6885 1869 6888
rect 1903 6916 1915 6919
rect 2409 6919 2467 6925
rect 2409 6916 2421 6919
rect 1903 6888 2421 6916
rect 1903 6885 1915 6888
rect 1857 6879 1915 6885
rect 2409 6885 2421 6888
rect 2455 6885 2467 6919
rect 2409 6879 2467 6885
rect 4706 6876 4712 6928
rect 4764 6916 4770 6928
rect 7929 6919 7987 6925
rect 7929 6916 7941 6919
rect 4764 6888 7941 6916
rect 4764 6876 4770 6888
rect 7929 6885 7941 6888
rect 7975 6916 7987 6919
rect 8294 6916 8300 6928
rect 7975 6888 8300 6916
rect 7975 6885 7987 6888
rect 7929 6879 7987 6885
rect 8294 6876 8300 6888
rect 8352 6876 8358 6928
rect 4982 6848 4988 6860
rect 4895 6820 4988 6848
rect 4982 6808 4988 6820
rect 5040 6848 5046 6860
rect 5344 6851 5402 6857
rect 5344 6848 5356 6851
rect 5040 6820 5356 6848
rect 5040 6808 5046 6820
rect 5344 6817 5356 6820
rect 5390 6848 5402 6851
rect 6086 6848 6092 6860
rect 5390 6820 6092 6848
rect 5390 6817 5402 6820
rect 5344 6811 5402 6817
rect 6086 6808 6092 6820
rect 6144 6808 6150 6860
rect 8018 6808 8024 6860
rect 8076 6848 8082 6860
rect 9944 6851 10002 6857
rect 8076 6820 8121 6848
rect 8076 6808 8082 6820
rect 9944 6817 9956 6851
rect 9990 6848 10002 6851
rect 10318 6848 10324 6860
rect 9990 6820 10324 6848
rect 9990 6817 10002 6820
rect 9944 6811 10002 6817
rect 10318 6808 10324 6820
rect 10376 6848 10382 6860
rect 12066 6848 12072 6860
rect 10376 6820 12072 6848
rect 10376 6808 10382 6820
rect 12066 6808 12072 6820
rect 12124 6808 12130 6860
rect 12437 6851 12495 6857
rect 12437 6817 12449 6851
rect 12483 6848 12495 6851
rect 12986 6848 12992 6860
rect 12483 6820 12992 6848
rect 12483 6817 12495 6820
rect 12437 6811 12495 6817
rect 12986 6808 12992 6820
rect 13044 6808 13050 6860
rect 13262 6848 13268 6860
rect 13223 6820 13268 6848
rect 13262 6808 13268 6820
rect 13320 6808 13326 6860
rect 1949 6783 2007 6789
rect 1949 6749 1961 6783
rect 1995 6749 2007 6783
rect 1949 6743 2007 6749
rect 1762 6672 1768 6724
rect 1820 6712 1826 6724
rect 1964 6712 1992 6743
rect 2498 6740 2504 6792
rect 2556 6780 2562 6792
rect 2961 6783 3019 6789
rect 2961 6780 2973 6783
rect 2556 6752 2973 6780
rect 2556 6740 2562 6752
rect 2961 6749 2973 6752
rect 3007 6749 3019 6783
rect 5074 6780 5080 6792
rect 5035 6752 5080 6780
rect 2961 6743 3019 6749
rect 5074 6740 5080 6752
rect 5132 6740 5138 6792
rect 7650 6740 7656 6792
rect 7708 6780 7714 6792
rect 8113 6783 8171 6789
rect 8113 6780 8125 6783
rect 7708 6752 8125 6780
rect 7708 6740 7714 6752
rect 8113 6749 8125 6752
rect 8159 6749 8171 6783
rect 8113 6743 8171 6749
rect 9677 6783 9735 6789
rect 9677 6749 9689 6783
rect 9723 6749 9735 6783
rect 9677 6743 9735 6749
rect 1820 6684 1992 6712
rect 1820 6672 1826 6684
rect 6546 6672 6552 6724
rect 6604 6712 6610 6724
rect 7561 6715 7619 6721
rect 7561 6712 7573 6715
rect 6604 6684 7573 6712
rect 6604 6672 6610 6684
rect 7561 6681 7573 6684
rect 7607 6681 7619 6715
rect 7561 6675 7619 6681
rect 9398 6672 9404 6724
rect 9456 6712 9462 6724
rect 9692 6712 9720 6743
rect 12526 6740 12532 6792
rect 12584 6780 12590 6792
rect 13357 6783 13415 6789
rect 13357 6780 13369 6783
rect 12584 6752 13369 6780
rect 12584 6740 12590 6752
rect 13357 6749 13369 6752
rect 13403 6749 13415 6783
rect 13357 6743 13415 6749
rect 13541 6783 13599 6789
rect 13541 6749 13553 6783
rect 13587 6780 13599 6783
rect 13630 6780 13636 6792
rect 13587 6752 13636 6780
rect 13587 6749 13599 6752
rect 13541 6743 13599 6749
rect 13630 6740 13636 6752
rect 13688 6780 13694 6792
rect 14016 6780 14044 6947
rect 14274 6944 14280 6956
rect 14332 6944 14338 6996
rect 15746 6984 15752 6996
rect 15707 6956 15752 6984
rect 15746 6944 15752 6956
rect 15804 6944 15810 6996
rect 18414 6944 18420 6996
rect 18472 6984 18478 6996
rect 19245 6987 19303 6993
rect 19245 6984 19257 6987
rect 18472 6956 19257 6984
rect 18472 6944 18478 6956
rect 19245 6953 19257 6956
rect 19291 6953 19303 6987
rect 19245 6947 19303 6953
rect 19518 6944 19524 6996
rect 19576 6984 19582 6996
rect 20165 6987 20223 6993
rect 20165 6984 20177 6987
rect 19576 6956 20177 6984
rect 19576 6944 19582 6956
rect 20165 6953 20177 6956
rect 20211 6953 20223 6987
rect 20165 6947 20223 6953
rect 16669 6919 16727 6925
rect 16669 6916 16681 6919
rect 16500 6888 16681 6916
rect 16114 6848 16120 6860
rect 16075 6820 16120 6848
rect 16114 6808 16120 6820
rect 16172 6808 16178 6860
rect 16500 6848 16528 6888
rect 16669 6885 16681 6888
rect 16715 6885 16727 6919
rect 18506 6916 18512 6928
rect 16669 6879 16727 6885
rect 17880 6888 18512 6916
rect 16224 6820 16528 6848
rect 16224 6792 16252 6820
rect 16942 6808 16948 6860
rect 17000 6848 17006 6860
rect 17773 6851 17831 6857
rect 17773 6848 17785 6851
rect 17000 6820 17785 6848
rect 17000 6808 17006 6820
rect 17773 6817 17785 6820
rect 17819 6848 17831 6851
rect 17880 6848 17908 6888
rect 18506 6876 18512 6888
rect 18564 6876 18570 6928
rect 19889 6919 19947 6925
rect 19889 6885 19901 6919
rect 19935 6916 19947 6919
rect 19978 6916 19984 6928
rect 19935 6888 19984 6916
rect 19935 6885 19947 6888
rect 19889 6879 19947 6885
rect 19978 6876 19984 6888
rect 20036 6876 20042 6928
rect 18138 6857 18144 6860
rect 18132 6848 18144 6857
rect 17819 6820 17908 6848
rect 18099 6820 18144 6848
rect 17819 6817 17831 6820
rect 17773 6811 17831 6817
rect 18132 6811 18144 6820
rect 18138 6808 18144 6811
rect 18196 6808 18202 6860
rect 13688 6752 14044 6780
rect 15289 6783 15347 6789
rect 13688 6740 13694 6752
rect 15289 6749 15301 6783
rect 15335 6780 15347 6783
rect 16206 6780 16212 6792
rect 15335 6752 16212 6780
rect 15335 6749 15347 6752
rect 15289 6743 15347 6749
rect 16206 6740 16212 6752
rect 16264 6740 16270 6792
rect 16761 6783 16819 6789
rect 16761 6749 16773 6783
rect 16807 6749 16819 6783
rect 16761 6743 16819 6749
rect 9456 6684 9720 6712
rect 11057 6715 11115 6721
rect 9456 6672 9462 6684
rect 11057 6681 11069 6715
rect 11103 6712 11115 6715
rect 11146 6712 11152 6724
rect 11103 6684 11152 6712
rect 11103 6681 11115 6684
rect 11057 6675 11115 6681
rect 11146 6672 11152 6684
rect 11204 6672 11210 6724
rect 14553 6715 14611 6721
rect 14553 6681 14565 6715
rect 14599 6712 14611 6715
rect 15930 6712 15936 6724
rect 14599 6684 15936 6712
rect 14599 6681 14611 6684
rect 14553 6675 14611 6681
rect 15930 6672 15936 6684
rect 15988 6672 15994 6724
rect 16301 6715 16359 6721
rect 16301 6681 16313 6715
rect 16347 6712 16359 6715
rect 16482 6712 16488 6724
rect 16347 6684 16488 6712
rect 16347 6681 16359 6684
rect 16301 6675 16359 6681
rect 16482 6672 16488 6684
rect 16540 6672 16546 6724
rect 1397 6647 1455 6653
rect 1397 6613 1409 6647
rect 1443 6644 1455 6647
rect 1854 6644 1860 6656
rect 1443 6616 1860 6644
rect 1443 6613 1455 6616
rect 1397 6607 1455 6613
rect 1854 6604 1860 6616
rect 1912 6604 1918 6656
rect 2590 6604 2596 6656
rect 2648 6644 2654 6656
rect 3510 6644 3516 6656
rect 2648 6616 3516 6644
rect 2648 6604 2654 6616
rect 3510 6604 3516 6616
rect 3568 6604 3574 6656
rect 3878 6644 3884 6656
rect 3839 6616 3884 6644
rect 3878 6604 3884 6616
rect 3936 6604 3942 6656
rect 4614 6644 4620 6656
rect 4575 6616 4620 6644
rect 4614 6604 4620 6616
rect 4672 6604 4678 6656
rect 6270 6604 6276 6656
rect 6328 6644 6334 6656
rect 6457 6647 6515 6653
rect 6457 6644 6469 6647
rect 6328 6616 6469 6644
rect 6328 6604 6334 6616
rect 6457 6613 6469 6616
rect 6503 6613 6515 6647
rect 7374 6644 7380 6656
rect 7335 6616 7380 6644
rect 6457 6607 6515 6613
rect 7374 6604 7380 6616
rect 7432 6604 7438 6656
rect 14826 6644 14832 6656
rect 14787 6616 14832 6644
rect 14826 6604 14832 6616
rect 14884 6604 14890 6656
rect 16114 6604 16120 6656
rect 16172 6644 16178 6656
rect 16776 6644 16804 6743
rect 16850 6740 16856 6792
rect 16908 6780 16914 6792
rect 17310 6780 17316 6792
rect 16908 6752 16953 6780
rect 17271 6752 17316 6780
rect 16908 6740 16914 6752
rect 17310 6740 17316 6752
rect 17368 6740 17374 6792
rect 17865 6783 17923 6789
rect 17865 6749 17877 6783
rect 17911 6749 17923 6783
rect 21174 6780 21180 6792
rect 21135 6752 21180 6780
rect 17865 6743 17923 6749
rect 17034 6672 17040 6724
rect 17092 6712 17098 6724
rect 17880 6712 17908 6743
rect 21174 6740 21180 6752
rect 21232 6740 21238 6792
rect 17092 6684 17908 6712
rect 17092 6672 17098 6684
rect 20530 6644 20536 6656
rect 16172 6616 16804 6644
rect 20491 6616 20536 6644
rect 16172 6604 16178 6616
rect 20530 6604 20536 6616
rect 20588 6604 20594 6656
rect 21542 6644 21548 6656
rect 21503 6616 21548 6644
rect 21542 6604 21548 6616
rect 21600 6604 21606 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 2682 6400 2688 6452
rect 2740 6440 2746 6452
rect 2961 6443 3019 6449
rect 2961 6440 2973 6443
rect 2740 6412 2973 6440
rect 2740 6400 2746 6412
rect 2961 6409 2973 6412
rect 3007 6440 3019 6443
rect 4154 6440 4160 6452
rect 3007 6412 4160 6440
rect 3007 6409 3019 6412
rect 2961 6403 3019 6409
rect 4154 6400 4160 6412
rect 4212 6400 4218 6452
rect 4982 6440 4988 6452
rect 4943 6412 4988 6440
rect 4982 6400 4988 6412
rect 5040 6400 5046 6452
rect 7929 6443 7987 6449
rect 7929 6409 7941 6443
rect 7975 6440 7987 6443
rect 8018 6440 8024 6452
rect 7975 6412 8024 6440
rect 7975 6409 7987 6412
rect 7929 6403 7987 6409
rect 8018 6400 8024 6412
rect 8076 6400 8082 6452
rect 8294 6440 8300 6452
rect 8255 6412 8300 6440
rect 8294 6400 8300 6412
rect 8352 6400 8358 6452
rect 8570 6440 8576 6452
rect 8404 6412 8576 6440
rect 2866 6332 2872 6384
rect 2924 6372 2930 6384
rect 6549 6375 6607 6381
rect 6549 6372 6561 6375
rect 2924 6344 6561 6372
rect 2924 6332 2930 6344
rect 6549 6341 6561 6344
rect 6595 6341 6607 6375
rect 6822 6372 6828 6384
rect 6783 6344 6828 6372
rect 6549 6335 6607 6341
rect 1578 6304 1584 6316
rect 1539 6276 1584 6304
rect 1578 6264 1584 6276
rect 1636 6264 1642 6316
rect 4614 6304 4620 6316
rect 4527 6276 4620 6304
rect 4614 6264 4620 6276
rect 4672 6304 4678 6316
rect 5534 6304 5540 6316
rect 4672 6276 5540 6304
rect 4672 6264 4678 6276
rect 5534 6264 5540 6276
rect 5592 6304 5598 6316
rect 5721 6307 5779 6313
rect 5721 6304 5733 6307
rect 5592 6276 5733 6304
rect 5592 6264 5598 6276
rect 5721 6273 5733 6276
rect 5767 6304 5779 6307
rect 6270 6304 6276 6316
rect 5767 6276 6276 6304
rect 5767 6273 5779 6276
rect 5721 6267 5779 6273
rect 6270 6264 6276 6276
rect 6328 6264 6334 6316
rect 6564 6304 6592 6335
rect 6822 6332 6828 6344
rect 6880 6332 6886 6384
rect 7285 6307 7343 6313
rect 7285 6304 7297 6307
rect 6564 6276 7297 6304
rect 7285 6273 7297 6276
rect 7331 6273 7343 6307
rect 7285 6267 7343 6273
rect 7469 6307 7527 6313
rect 7469 6273 7481 6307
rect 7515 6304 7527 6307
rect 7650 6304 7656 6316
rect 7515 6276 7656 6304
rect 7515 6273 7527 6276
rect 7469 6267 7527 6273
rect 6086 6196 6092 6248
rect 6144 6236 6150 6248
rect 6181 6239 6239 6245
rect 6181 6236 6193 6239
rect 6144 6208 6193 6236
rect 6144 6196 6150 6208
rect 6181 6205 6193 6208
rect 6227 6236 6239 6239
rect 6362 6236 6368 6248
rect 6227 6208 6368 6236
rect 6227 6205 6239 6208
rect 6181 6199 6239 6205
rect 6362 6196 6368 6208
rect 6420 6236 6426 6248
rect 7484 6236 7512 6267
rect 7650 6264 7656 6276
rect 7708 6264 7714 6316
rect 8404 6313 8432 6412
rect 8570 6400 8576 6412
rect 8628 6440 8634 6452
rect 9398 6440 9404 6452
rect 8628 6412 9404 6440
rect 8628 6400 8634 6412
rect 9398 6400 9404 6412
rect 9456 6400 9462 6452
rect 10318 6440 10324 6452
rect 10279 6412 10324 6440
rect 10318 6400 10324 6412
rect 10376 6400 10382 6452
rect 11054 6440 11060 6452
rect 11015 6412 11060 6440
rect 11054 6400 11060 6412
rect 11112 6440 11118 6452
rect 11425 6443 11483 6449
rect 11425 6440 11437 6443
rect 11112 6412 11437 6440
rect 11112 6400 11118 6412
rect 11425 6409 11437 6412
rect 11471 6440 11483 6443
rect 11793 6443 11851 6449
rect 11793 6440 11805 6443
rect 11471 6412 11805 6440
rect 11471 6409 11483 6412
rect 11425 6403 11483 6409
rect 11793 6409 11805 6412
rect 11839 6409 11851 6443
rect 11793 6403 11851 6409
rect 12253 6443 12311 6449
rect 12253 6409 12265 6443
rect 12299 6440 12311 6443
rect 13630 6440 13636 6452
rect 12299 6412 13636 6440
rect 12299 6409 12311 6412
rect 12253 6403 12311 6409
rect 13630 6400 13636 6412
rect 13688 6400 13694 6452
rect 14090 6400 14096 6452
rect 14148 6440 14154 6452
rect 14277 6443 14335 6449
rect 14277 6440 14289 6443
rect 14148 6412 14289 6440
rect 14148 6400 14154 6412
rect 14277 6409 14289 6412
rect 14323 6409 14335 6443
rect 16206 6440 16212 6452
rect 16167 6412 16212 6440
rect 14277 6403 14335 6409
rect 16206 6400 16212 6412
rect 16264 6400 16270 6452
rect 16393 6443 16451 6449
rect 16393 6409 16405 6443
rect 16439 6440 16451 6443
rect 16942 6440 16948 6452
rect 16439 6412 16948 6440
rect 16439 6409 16451 6412
rect 16393 6403 16451 6409
rect 16942 6400 16948 6412
rect 17000 6400 17006 6452
rect 17865 6443 17923 6449
rect 17865 6409 17877 6443
rect 17911 6440 17923 6443
rect 18138 6440 18144 6452
rect 17911 6412 18144 6440
rect 17911 6409 17923 6412
rect 17865 6403 17923 6409
rect 8389 6307 8447 6313
rect 8389 6273 8401 6307
rect 8435 6273 8447 6307
rect 10686 6304 10692 6316
rect 10647 6276 10692 6304
rect 8389 6267 8447 6273
rect 10686 6264 10692 6276
rect 10744 6264 10750 6316
rect 13170 6264 13176 6316
rect 13228 6304 13234 6316
rect 13722 6304 13728 6316
rect 13228 6276 13728 6304
rect 13228 6264 13234 6276
rect 13722 6264 13728 6276
rect 13780 6264 13786 6316
rect 13909 6307 13967 6313
rect 13909 6273 13921 6307
rect 13955 6304 13967 6307
rect 14108 6304 14136 6400
rect 14734 6372 14740 6384
rect 14695 6344 14740 6372
rect 14734 6332 14740 6344
rect 14792 6332 14798 6384
rect 13955 6276 14136 6304
rect 13955 6273 13967 6276
rect 13909 6267 13967 6273
rect 8662 6245 8668 6248
rect 8656 6236 8668 6245
rect 6420 6208 7512 6236
rect 8623 6208 8668 6236
rect 6420 6196 6426 6208
rect 8656 6199 8668 6208
rect 8662 6196 8668 6199
rect 8720 6196 8726 6248
rect 12986 6196 12992 6248
rect 13044 6236 13050 6248
rect 13633 6239 13691 6245
rect 13633 6236 13645 6239
rect 13044 6208 13645 6236
rect 13044 6196 13050 6208
rect 13633 6205 13645 6208
rect 13679 6205 13691 6239
rect 14752 6236 14780 6332
rect 14826 6264 14832 6316
rect 14884 6304 14890 6316
rect 15378 6304 15384 6316
rect 14884 6276 15384 6304
rect 14884 6264 14890 6276
rect 15378 6264 15384 6276
rect 15436 6264 15442 6316
rect 15933 6307 15991 6313
rect 15933 6273 15945 6307
rect 15979 6304 15991 6307
rect 16574 6304 16580 6316
rect 15979 6276 16580 6304
rect 15979 6273 15991 6276
rect 15933 6267 15991 6273
rect 16574 6264 16580 6276
rect 16632 6304 16638 6316
rect 16850 6304 16856 6316
rect 16632 6276 16856 6304
rect 16632 6264 16638 6276
rect 16850 6264 16856 6276
rect 16908 6304 16914 6316
rect 16945 6307 17003 6313
rect 16945 6304 16957 6307
rect 16908 6276 16957 6304
rect 16908 6264 16914 6276
rect 16945 6273 16957 6276
rect 16991 6304 17003 6307
rect 17880 6304 17908 6403
rect 18138 6400 18144 6412
rect 18196 6400 18202 6452
rect 18414 6440 18420 6452
rect 18375 6412 18420 6440
rect 18414 6400 18420 6412
rect 18472 6400 18478 6452
rect 20438 6440 20444 6452
rect 20399 6412 20444 6440
rect 20438 6400 20444 6412
rect 20496 6440 20502 6452
rect 20496 6412 21496 6440
rect 20496 6400 20502 6412
rect 16991 6276 17908 6304
rect 18432 6304 18460 6400
rect 20806 6372 20812 6384
rect 20767 6344 20812 6372
rect 20806 6332 20812 6344
rect 20864 6332 20870 6384
rect 20990 6372 20996 6384
rect 20951 6344 20996 6372
rect 20990 6332 20996 6344
rect 21048 6332 21054 6384
rect 18432 6276 18644 6304
rect 16991 6273 17003 6276
rect 16945 6267 17003 6273
rect 15197 6239 15255 6245
rect 15197 6236 15209 6239
rect 14752 6208 15209 6236
rect 13633 6199 13691 6205
rect 15197 6205 15209 6208
rect 15243 6236 15255 6239
rect 16206 6236 16212 6248
rect 15243 6208 16212 6236
rect 15243 6205 15255 6208
rect 15197 6199 15255 6205
rect 16206 6196 16212 6208
rect 16264 6196 16270 6248
rect 17034 6196 17040 6248
rect 17092 6236 17098 6248
rect 18506 6236 18512 6248
rect 17092 6208 18512 6236
rect 17092 6196 17098 6208
rect 18506 6196 18512 6208
rect 18564 6196 18570 6248
rect 18616 6236 18644 6276
rect 18765 6239 18823 6245
rect 18765 6236 18777 6239
rect 18616 6208 18777 6236
rect 18765 6205 18777 6208
rect 18811 6205 18823 6239
rect 20824 6236 20852 6332
rect 21468 6313 21496 6412
rect 21453 6307 21511 6313
rect 21453 6273 21465 6307
rect 21499 6273 21511 6307
rect 21634 6304 21640 6316
rect 21595 6276 21640 6304
rect 21453 6267 21511 6273
rect 21634 6264 21640 6276
rect 21692 6264 21698 6316
rect 21361 6239 21419 6245
rect 21361 6236 21373 6239
rect 20824 6208 21373 6236
rect 18765 6199 18823 6205
rect 21361 6205 21373 6208
rect 21407 6236 21419 6239
rect 22002 6236 22008 6248
rect 21407 6208 22008 6236
rect 21407 6205 21419 6208
rect 21361 6199 21419 6205
rect 22002 6196 22008 6208
rect 22060 6196 22066 6248
rect 1848 6171 1906 6177
rect 1848 6137 1860 6171
rect 1894 6168 1906 6171
rect 1946 6168 1952 6180
rect 1894 6140 1952 6168
rect 1894 6137 1906 6140
rect 1848 6131 1906 6137
rect 1946 6128 1952 6140
rect 2004 6168 2010 6180
rect 2866 6168 2872 6180
rect 2004 6140 2872 6168
rect 2004 6128 2010 6140
rect 2866 6128 2872 6140
rect 2924 6168 2930 6180
rect 3881 6171 3939 6177
rect 3881 6168 3893 6171
rect 2924 6140 3893 6168
rect 2924 6128 2930 6140
rect 3881 6137 3893 6140
rect 3927 6137 3939 6171
rect 3881 6131 3939 6137
rect 5166 6128 5172 6180
rect 5224 6168 5230 6180
rect 5537 6171 5595 6177
rect 5537 6168 5549 6171
rect 5224 6140 5549 6168
rect 5224 6128 5230 6140
rect 5537 6137 5549 6140
rect 5583 6137 5595 6171
rect 16850 6168 16856 6180
rect 5537 6131 5595 6137
rect 14844 6140 16856 6168
rect 3602 6100 3608 6112
rect 3563 6072 3608 6100
rect 3602 6060 3608 6072
rect 3660 6060 3666 6112
rect 4062 6100 4068 6112
rect 4023 6072 4068 6100
rect 4062 6060 4068 6072
rect 4120 6060 4126 6112
rect 5074 6100 5080 6112
rect 5035 6072 5080 6100
rect 5074 6060 5080 6072
rect 5132 6060 5138 6112
rect 5445 6103 5503 6109
rect 5445 6069 5457 6103
rect 5491 6100 5503 6103
rect 6822 6100 6828 6112
rect 5491 6072 6828 6100
rect 5491 6069 5503 6072
rect 5445 6063 5503 6069
rect 6822 6060 6828 6072
rect 6880 6060 6886 6112
rect 6914 6060 6920 6112
rect 6972 6100 6978 6112
rect 7193 6103 7251 6109
rect 7193 6100 7205 6103
rect 6972 6072 7205 6100
rect 6972 6060 6978 6072
rect 7193 6069 7205 6072
rect 7239 6069 7251 6103
rect 7193 6063 7251 6069
rect 9769 6103 9827 6109
rect 9769 6069 9781 6103
rect 9815 6100 9827 6103
rect 10134 6100 10140 6112
rect 9815 6072 10140 6100
rect 9815 6069 9827 6072
rect 9769 6063 9827 6069
rect 10134 6060 10140 6072
rect 10192 6060 10198 6112
rect 12526 6060 12532 6112
rect 12584 6100 12590 6112
rect 12897 6103 12955 6109
rect 12897 6100 12909 6103
rect 12584 6072 12909 6100
rect 12584 6060 12590 6072
rect 12897 6069 12909 6072
rect 12943 6069 12955 6103
rect 12897 6063 12955 6069
rect 13078 6060 13084 6112
rect 13136 6100 13142 6112
rect 14844 6109 14872 6140
rect 16850 6128 16856 6140
rect 16908 6128 16914 6180
rect 13265 6103 13323 6109
rect 13265 6100 13277 6103
rect 13136 6072 13277 6100
rect 13136 6060 13142 6072
rect 13265 6069 13277 6072
rect 13311 6069 13323 6103
rect 13265 6063 13323 6069
rect 14829 6103 14887 6109
rect 14829 6069 14841 6103
rect 14875 6069 14887 6103
rect 15286 6100 15292 6112
rect 15247 6072 15292 6100
rect 14829 6063 14887 6069
rect 15286 6060 15292 6072
rect 15344 6060 15350 6112
rect 16758 6100 16764 6112
rect 16719 6072 16764 6100
rect 16758 6060 16764 6072
rect 16816 6100 16822 6112
rect 17405 6103 17463 6109
rect 17405 6100 17417 6103
rect 16816 6072 17417 6100
rect 16816 6060 16822 6072
rect 17405 6069 17417 6072
rect 17451 6069 17463 6103
rect 17405 6063 17463 6069
rect 19334 6060 19340 6112
rect 19392 6100 19398 6112
rect 19889 6103 19947 6109
rect 19889 6100 19901 6103
rect 19392 6072 19901 6100
rect 19392 6060 19398 6072
rect 19889 6069 19901 6072
rect 19935 6069 19947 6103
rect 19889 6063 19947 6069
rect 22094 6060 22100 6112
rect 22152 6100 22158 6112
rect 22152 6072 22197 6100
rect 22152 6060 22158 6072
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 2866 5896 2872 5908
rect 2827 5868 2872 5896
rect 2866 5856 2872 5868
rect 2924 5856 2930 5908
rect 3510 5856 3516 5908
rect 3568 5896 3574 5908
rect 4433 5899 4491 5905
rect 4433 5896 4445 5899
rect 3568 5868 4445 5896
rect 3568 5856 3574 5868
rect 4433 5865 4445 5868
rect 4479 5865 4491 5899
rect 4433 5859 4491 5865
rect 5629 5899 5687 5905
rect 5629 5865 5641 5899
rect 5675 5896 5687 5899
rect 5902 5896 5908 5908
rect 5675 5868 5908 5896
rect 5675 5865 5687 5868
rect 5629 5859 5687 5865
rect 5902 5856 5908 5868
rect 5960 5856 5966 5908
rect 5997 5899 6055 5905
rect 5997 5865 6009 5899
rect 6043 5896 6055 5899
rect 6546 5896 6552 5908
rect 6043 5868 6552 5896
rect 6043 5865 6055 5868
rect 5997 5859 6055 5865
rect 6546 5856 6552 5868
rect 6604 5856 6610 5908
rect 6914 5896 6920 5908
rect 6875 5868 6920 5896
rect 6914 5856 6920 5868
rect 6972 5856 6978 5908
rect 7561 5899 7619 5905
rect 7561 5865 7573 5899
rect 7607 5896 7619 5899
rect 7650 5896 7656 5908
rect 7607 5868 7656 5896
rect 7607 5865 7619 5868
rect 7561 5859 7619 5865
rect 7650 5856 7656 5868
rect 7708 5856 7714 5908
rect 8018 5896 8024 5908
rect 7979 5868 8024 5896
rect 8018 5856 8024 5868
rect 8076 5856 8082 5908
rect 9674 5856 9680 5908
rect 9732 5896 9738 5908
rect 10137 5899 10195 5905
rect 10137 5896 10149 5899
rect 9732 5868 10149 5896
rect 9732 5856 9738 5868
rect 10137 5865 10149 5868
rect 10183 5865 10195 5899
rect 10137 5859 10195 5865
rect 11054 5856 11060 5908
rect 11112 5896 11118 5908
rect 11333 5899 11391 5905
rect 11333 5896 11345 5899
rect 11112 5868 11345 5896
rect 11112 5856 11118 5868
rect 11333 5865 11345 5868
rect 11379 5865 11391 5899
rect 11514 5896 11520 5908
rect 11475 5868 11520 5896
rect 11333 5859 11391 5865
rect 1762 5837 1768 5840
rect 1756 5828 1768 5837
rect 1723 5800 1768 5828
rect 1756 5791 1768 5800
rect 1762 5788 1768 5791
rect 1820 5788 1826 5840
rect 1854 5788 1860 5840
rect 1912 5828 1918 5840
rect 3789 5831 3847 5837
rect 3789 5828 3801 5831
rect 1912 5800 3801 5828
rect 1912 5788 1918 5800
rect 3789 5797 3801 5800
rect 3835 5797 3847 5831
rect 3789 5791 3847 5797
rect 9493 5831 9551 5837
rect 9493 5797 9505 5831
rect 9539 5828 9551 5831
rect 10042 5828 10048 5840
rect 9539 5800 10048 5828
rect 9539 5797 9551 5800
rect 9493 5791 9551 5797
rect 10042 5788 10048 5800
rect 10100 5788 10106 5840
rect 10686 5828 10692 5840
rect 10647 5800 10692 5828
rect 10686 5788 10692 5800
rect 10744 5788 10750 5840
rect 11348 5828 11376 5859
rect 11514 5856 11520 5868
rect 11572 5856 11578 5908
rect 12986 5896 12992 5908
rect 12899 5868 12992 5896
rect 12986 5856 12992 5868
rect 13044 5896 13050 5908
rect 13262 5896 13268 5908
rect 13044 5868 13268 5896
rect 13044 5856 13050 5868
rect 13262 5856 13268 5868
rect 13320 5856 13326 5908
rect 13446 5856 13452 5908
rect 13504 5896 13510 5908
rect 13541 5899 13599 5905
rect 13541 5896 13553 5899
rect 13504 5868 13553 5896
rect 13504 5856 13510 5868
rect 13541 5865 13553 5868
rect 13587 5865 13599 5899
rect 13541 5859 13599 5865
rect 13722 5856 13728 5908
rect 13780 5896 13786 5908
rect 14093 5899 14151 5905
rect 14093 5896 14105 5899
rect 13780 5868 14105 5896
rect 13780 5856 13786 5868
rect 14093 5865 14105 5868
rect 14139 5865 14151 5899
rect 14093 5859 14151 5865
rect 15378 5856 15384 5908
rect 15436 5896 15442 5908
rect 15841 5899 15899 5905
rect 15841 5896 15853 5899
rect 15436 5868 15853 5896
rect 15436 5856 15442 5868
rect 15841 5865 15853 5868
rect 15887 5865 15899 5899
rect 15841 5859 15899 5865
rect 15930 5856 15936 5908
rect 15988 5896 15994 5908
rect 16574 5896 16580 5908
rect 15988 5868 16033 5896
rect 16535 5868 16580 5896
rect 15988 5856 15994 5868
rect 16574 5856 16580 5868
rect 16632 5856 16638 5908
rect 16850 5896 16856 5908
rect 16811 5868 16856 5896
rect 16850 5856 16856 5868
rect 16908 5856 16914 5908
rect 18506 5856 18512 5908
rect 18564 5896 18570 5908
rect 19337 5899 19395 5905
rect 19337 5896 19349 5899
rect 18564 5868 19349 5896
rect 18564 5856 18570 5868
rect 19337 5865 19349 5868
rect 19383 5896 19395 5899
rect 20441 5899 20499 5905
rect 20441 5896 20453 5899
rect 19383 5868 20453 5896
rect 19383 5865 19395 5868
rect 19337 5859 19395 5865
rect 20441 5865 20453 5868
rect 20487 5896 20499 5899
rect 20530 5896 20536 5908
rect 20487 5868 20536 5896
rect 20487 5865 20499 5868
rect 20441 5859 20499 5865
rect 20530 5856 20536 5868
rect 20588 5856 20594 5908
rect 12434 5828 12440 5840
rect 11348 5800 12440 5828
rect 12434 5788 12440 5800
rect 12492 5788 12498 5840
rect 17218 5788 17224 5840
rect 17276 5837 17282 5840
rect 17276 5831 17340 5837
rect 17276 5797 17294 5831
rect 17328 5797 17340 5831
rect 17276 5791 17340 5797
rect 17276 5788 17282 5791
rect 1489 5763 1547 5769
rect 1489 5729 1501 5763
rect 1535 5760 1547 5763
rect 1578 5760 1584 5772
rect 1535 5732 1584 5760
rect 1535 5729 1547 5732
rect 1489 5723 1547 5729
rect 1578 5720 1584 5732
rect 1636 5720 1642 5772
rect 2682 5720 2688 5772
rect 2740 5760 2746 5772
rect 3878 5760 3884 5772
rect 2740 5732 3884 5760
rect 2740 5720 2746 5732
rect 3878 5720 3884 5732
rect 3936 5760 3942 5772
rect 4525 5763 4583 5769
rect 4525 5760 4537 5763
rect 3936 5732 4537 5760
rect 3936 5720 3942 5732
rect 4525 5729 4537 5732
rect 4571 5729 4583 5763
rect 4525 5723 4583 5729
rect 5442 5720 5448 5772
rect 5500 5760 5506 5772
rect 6086 5760 6092 5772
rect 5500 5732 6092 5760
rect 5500 5720 5506 5732
rect 6086 5720 6092 5732
rect 6144 5720 6150 5772
rect 8386 5760 8392 5772
rect 8347 5732 8392 5760
rect 8386 5720 8392 5732
rect 8444 5720 8450 5772
rect 11882 5760 11888 5772
rect 8496 5732 11888 5760
rect 4154 5652 4160 5704
rect 4212 5692 4218 5704
rect 4617 5695 4675 5701
rect 4617 5692 4629 5695
rect 4212 5664 4629 5692
rect 4212 5652 4218 5664
rect 4617 5661 4629 5664
rect 4663 5661 4675 5695
rect 6270 5692 6276 5704
rect 6231 5664 6276 5692
rect 4617 5655 4675 5661
rect 6270 5652 6276 5664
rect 6328 5652 6334 5704
rect 8294 5652 8300 5704
rect 8352 5692 8358 5704
rect 8496 5701 8524 5732
rect 11882 5720 11888 5732
rect 11940 5720 11946 5772
rect 13449 5763 13507 5769
rect 13449 5729 13461 5763
rect 13495 5760 13507 5763
rect 13722 5760 13728 5772
rect 13495 5732 13728 5760
rect 13495 5729 13507 5732
rect 13449 5723 13507 5729
rect 13722 5720 13728 5732
rect 13780 5720 13786 5772
rect 14550 5720 14556 5772
rect 14608 5760 14614 5772
rect 14829 5763 14887 5769
rect 14829 5760 14841 5763
rect 14608 5732 14841 5760
rect 14608 5720 14614 5732
rect 14829 5729 14841 5732
rect 14875 5760 14887 5763
rect 15286 5760 15292 5772
rect 14875 5732 15292 5760
rect 14875 5729 14887 5732
rect 14829 5723 14887 5729
rect 15286 5720 15292 5732
rect 15344 5760 15350 5772
rect 15838 5760 15844 5772
rect 15344 5732 15844 5760
rect 15344 5720 15350 5732
rect 15838 5720 15844 5732
rect 15896 5720 15902 5772
rect 19518 5760 19524 5772
rect 19479 5732 19524 5760
rect 19518 5720 19524 5732
rect 19576 5760 19582 5772
rect 20073 5763 20131 5769
rect 20073 5760 20085 5763
rect 19576 5732 20085 5760
rect 19576 5720 19582 5732
rect 20073 5729 20085 5732
rect 20119 5729 20131 5763
rect 20073 5723 20131 5729
rect 8481 5695 8539 5701
rect 8481 5692 8493 5695
rect 8352 5664 8493 5692
rect 8352 5652 8358 5664
rect 8481 5661 8493 5664
rect 8527 5661 8539 5695
rect 8481 5655 8539 5661
rect 8573 5695 8631 5701
rect 8573 5661 8585 5695
rect 8619 5661 8631 5695
rect 10226 5692 10232 5704
rect 10187 5664 10232 5692
rect 8573 5655 8631 5661
rect 4062 5624 4068 5636
rect 4023 5596 4068 5624
rect 4062 5584 4068 5596
rect 4120 5584 4126 5636
rect 8588 5624 8616 5655
rect 10226 5652 10232 5664
rect 10284 5652 10290 5704
rect 11974 5692 11980 5704
rect 11935 5664 11980 5692
rect 11974 5652 11980 5664
rect 12032 5652 12038 5704
rect 12066 5652 12072 5704
rect 12124 5692 12130 5704
rect 12124 5664 12217 5692
rect 12124 5652 12130 5664
rect 12802 5652 12808 5704
rect 12860 5692 12866 5704
rect 13633 5695 13691 5701
rect 13633 5692 13645 5695
rect 12860 5664 13645 5692
rect 12860 5652 12866 5664
rect 13633 5661 13645 5664
rect 13679 5661 13691 5695
rect 13633 5655 13691 5661
rect 9030 5624 9036 5636
rect 7852 5596 8616 5624
rect 8991 5596 9036 5624
rect 7852 5568 7880 5596
rect 9030 5584 9036 5596
rect 9088 5584 9094 5636
rect 11146 5584 11152 5636
rect 11204 5624 11210 5636
rect 12084 5624 12112 5652
rect 11204 5596 12112 5624
rect 12621 5627 12679 5633
rect 11204 5584 11210 5596
rect 12621 5593 12633 5627
rect 12667 5624 12679 5627
rect 13262 5624 13268 5636
rect 12667 5596 13268 5624
rect 12667 5593 12679 5596
rect 12621 5587 12679 5593
rect 13262 5584 13268 5596
rect 13320 5584 13326 5636
rect 13648 5624 13676 5655
rect 15562 5652 15568 5704
rect 15620 5692 15626 5704
rect 16114 5692 16120 5704
rect 15620 5664 16120 5692
rect 15620 5652 15626 5664
rect 16114 5652 16120 5664
rect 16172 5652 16178 5704
rect 16574 5652 16580 5704
rect 16632 5692 16638 5704
rect 17034 5692 17040 5704
rect 16632 5664 17040 5692
rect 16632 5652 16638 5664
rect 17034 5652 17040 5664
rect 17092 5652 17098 5704
rect 13722 5624 13728 5636
rect 13648 5596 13728 5624
rect 13722 5584 13728 5596
rect 13780 5584 13786 5636
rect 2958 5516 2964 5568
rect 3016 5556 3022 5568
rect 3421 5559 3479 5565
rect 3421 5556 3433 5559
rect 3016 5528 3433 5556
rect 3016 5516 3022 5528
rect 3421 5525 3433 5528
rect 3467 5525 3479 5559
rect 3421 5519 3479 5525
rect 5261 5559 5319 5565
rect 5261 5525 5273 5559
rect 5307 5556 5319 5559
rect 5350 5556 5356 5568
rect 5307 5528 5356 5556
rect 5307 5525 5319 5528
rect 5261 5519 5319 5525
rect 5350 5516 5356 5528
rect 5408 5516 5414 5568
rect 7834 5556 7840 5568
rect 7795 5528 7840 5556
rect 7834 5516 7840 5528
rect 7892 5516 7898 5568
rect 9677 5559 9735 5565
rect 9677 5525 9689 5559
rect 9723 5556 9735 5559
rect 10134 5556 10140 5568
rect 9723 5528 10140 5556
rect 9723 5525 9735 5528
rect 9677 5519 9735 5525
rect 10134 5516 10140 5528
rect 10192 5516 10198 5568
rect 13081 5559 13139 5565
rect 13081 5525 13093 5559
rect 13127 5556 13139 5559
rect 13630 5556 13636 5568
rect 13127 5528 13636 5556
rect 13127 5525 13139 5528
rect 13081 5519 13139 5525
rect 13630 5516 13636 5528
rect 13688 5516 13694 5568
rect 14553 5559 14611 5565
rect 14553 5525 14565 5559
rect 14599 5556 14611 5559
rect 14642 5556 14648 5568
rect 14599 5528 14648 5556
rect 14599 5525 14611 5528
rect 14553 5519 14611 5525
rect 14642 5516 14648 5528
rect 14700 5516 14706 5568
rect 15473 5559 15531 5565
rect 15473 5525 15485 5559
rect 15519 5556 15531 5559
rect 16022 5556 16028 5568
rect 15519 5528 16028 5556
rect 15519 5525 15531 5528
rect 15473 5519 15531 5525
rect 16022 5516 16028 5528
rect 16080 5516 16086 5568
rect 18322 5516 18328 5568
rect 18380 5556 18386 5568
rect 18417 5559 18475 5565
rect 18417 5556 18429 5559
rect 18380 5528 18429 5556
rect 18380 5516 18386 5528
rect 18417 5525 18429 5528
rect 18463 5525 18475 5559
rect 18417 5519 18475 5525
rect 18506 5516 18512 5568
rect 18564 5556 18570 5568
rect 18969 5559 19027 5565
rect 18969 5556 18981 5559
rect 18564 5528 18981 5556
rect 18564 5516 18570 5528
rect 18969 5525 18981 5528
rect 19015 5525 19027 5559
rect 18969 5519 19027 5525
rect 19426 5516 19432 5568
rect 19484 5556 19490 5568
rect 19705 5559 19763 5565
rect 19705 5556 19717 5559
rect 19484 5528 19717 5556
rect 19484 5516 19490 5528
rect 19705 5525 19717 5528
rect 19751 5525 19763 5559
rect 19705 5519 19763 5525
rect 20714 5516 20720 5568
rect 20772 5556 20778 5568
rect 21085 5559 21143 5565
rect 21085 5556 21097 5559
rect 20772 5528 21097 5556
rect 20772 5516 20778 5528
rect 21085 5525 21097 5528
rect 21131 5556 21143 5559
rect 21634 5556 21640 5568
rect 21131 5528 21640 5556
rect 21131 5525 21143 5528
rect 21085 5519 21143 5525
rect 21634 5516 21640 5528
rect 21692 5516 21698 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 1397 5355 1455 5361
rect 1397 5321 1409 5355
rect 1443 5352 1455 5355
rect 2590 5352 2596 5364
rect 1443 5324 2596 5352
rect 1443 5321 1455 5324
rect 1397 5315 1455 5321
rect 2590 5312 2596 5324
rect 2648 5312 2654 5364
rect 2958 5352 2964 5364
rect 2919 5324 2964 5352
rect 2958 5312 2964 5324
rect 3016 5312 3022 5364
rect 4154 5352 4160 5364
rect 4115 5324 4160 5352
rect 4154 5312 4160 5324
rect 4212 5312 4218 5364
rect 5169 5355 5227 5361
rect 5169 5321 5181 5355
rect 5215 5352 5227 5355
rect 5442 5352 5448 5364
rect 5215 5324 5448 5352
rect 5215 5321 5227 5324
rect 5169 5315 5227 5321
rect 5442 5312 5448 5324
rect 5500 5312 5506 5364
rect 6641 5355 6699 5361
rect 6641 5321 6653 5355
rect 6687 5352 6699 5355
rect 7282 5352 7288 5364
rect 6687 5324 7288 5352
rect 6687 5321 6699 5324
rect 6641 5315 6699 5321
rect 7282 5312 7288 5324
rect 7340 5312 7346 5364
rect 9950 5312 9956 5364
rect 10008 5352 10014 5364
rect 10962 5352 10968 5364
rect 10008 5324 10968 5352
rect 10008 5312 10014 5324
rect 10962 5312 10968 5324
rect 11020 5312 11026 5364
rect 11146 5352 11152 5364
rect 11107 5324 11152 5352
rect 11146 5312 11152 5324
rect 11204 5312 11210 5364
rect 11882 5312 11888 5364
rect 11940 5352 11946 5364
rect 12161 5355 12219 5361
rect 12161 5352 12173 5355
rect 11940 5324 12173 5352
rect 11940 5312 11946 5324
rect 12161 5321 12173 5324
rect 12207 5321 12219 5355
rect 13446 5352 13452 5364
rect 13407 5324 13452 5352
rect 12161 5315 12219 5321
rect 13446 5312 13452 5324
rect 13504 5312 13510 5364
rect 13906 5352 13912 5364
rect 13867 5324 13912 5352
rect 13906 5312 13912 5324
rect 13964 5312 13970 5364
rect 14921 5355 14979 5361
rect 14921 5321 14933 5355
rect 14967 5352 14979 5355
rect 15378 5352 15384 5364
rect 14967 5324 15384 5352
rect 14967 5321 14979 5324
rect 14921 5315 14979 5321
rect 15378 5312 15384 5324
rect 15436 5312 15442 5364
rect 16114 5312 16120 5364
rect 16172 5352 16178 5364
rect 16301 5355 16359 5361
rect 16301 5352 16313 5355
rect 16172 5324 16313 5352
rect 16172 5312 16178 5324
rect 16301 5321 16313 5324
rect 16347 5321 16359 5355
rect 18046 5352 18052 5364
rect 18007 5324 18052 5352
rect 16301 5315 16359 5321
rect 18046 5312 18052 5324
rect 18104 5312 18110 5364
rect 19613 5355 19671 5361
rect 19613 5321 19625 5355
rect 19659 5352 19671 5355
rect 20070 5352 20076 5364
rect 19659 5324 20076 5352
rect 19659 5321 19671 5324
rect 19613 5315 19671 5321
rect 20070 5312 20076 5324
rect 20128 5312 20134 5364
rect 20530 5312 20536 5364
rect 20588 5352 20594 5364
rect 20625 5355 20683 5361
rect 20625 5352 20637 5355
rect 20588 5324 20637 5352
rect 20588 5312 20594 5324
rect 20625 5321 20637 5324
rect 20671 5321 20683 5355
rect 20625 5315 20683 5321
rect 1762 5244 1768 5296
rect 1820 5284 1826 5296
rect 1820 5256 2176 5284
rect 1820 5244 1826 5256
rect 1946 5216 1952 5228
rect 1907 5188 1952 5216
rect 1946 5176 1952 5188
rect 2004 5176 2010 5228
rect 2148 5216 2176 5256
rect 13814 5244 13820 5296
rect 13872 5284 13878 5296
rect 14185 5287 14243 5293
rect 14185 5284 14197 5287
rect 13872 5256 14197 5284
rect 13872 5244 13878 5256
rect 14185 5253 14197 5256
rect 14231 5253 14243 5287
rect 14185 5247 14243 5253
rect 15470 5244 15476 5296
rect 15528 5284 15534 5296
rect 16025 5287 16083 5293
rect 16025 5284 16037 5287
rect 15528 5256 16037 5284
rect 15528 5244 15534 5256
rect 2222 5216 2228 5228
rect 2135 5188 2228 5216
rect 2222 5176 2228 5188
rect 2280 5216 2286 5228
rect 2409 5219 2467 5225
rect 2409 5216 2421 5219
rect 2280 5188 2421 5216
rect 2280 5176 2286 5188
rect 2409 5185 2421 5188
rect 2455 5216 2467 5219
rect 3602 5216 3608 5228
rect 2455 5188 3608 5216
rect 2455 5185 2467 5188
rect 2409 5179 2467 5185
rect 3602 5176 3608 5188
rect 3660 5176 3666 5228
rect 4709 5219 4767 5225
rect 4709 5185 4721 5219
rect 4755 5216 4767 5219
rect 5626 5216 5632 5228
rect 4755 5188 5632 5216
rect 4755 5185 4767 5188
rect 4709 5179 4767 5185
rect 5626 5176 5632 5188
rect 5684 5216 5690 5228
rect 5813 5219 5871 5225
rect 5813 5216 5825 5219
rect 5684 5188 5825 5216
rect 5684 5176 5690 5188
rect 5813 5185 5825 5188
rect 5859 5216 5871 5219
rect 6362 5216 6368 5228
rect 5859 5188 6368 5216
rect 5859 5185 5871 5188
rect 5813 5179 5871 5185
rect 6362 5176 6368 5188
rect 6420 5176 6426 5228
rect 7377 5219 7435 5225
rect 7377 5216 7389 5219
rect 7300 5188 7389 5216
rect 1854 5148 1860 5160
rect 1815 5120 1860 5148
rect 1854 5108 1860 5120
rect 1912 5108 1918 5160
rect 5077 5151 5135 5157
rect 5077 5117 5089 5151
rect 5123 5148 5135 5151
rect 5537 5151 5595 5157
rect 5537 5148 5549 5151
rect 5123 5120 5549 5148
rect 5123 5117 5135 5120
rect 5077 5111 5135 5117
rect 5537 5117 5549 5120
rect 5583 5148 5595 5151
rect 6546 5148 6552 5160
rect 5583 5120 6552 5148
rect 5583 5117 5595 5120
rect 5537 5111 5595 5117
rect 6546 5108 6552 5120
rect 6604 5108 6610 5160
rect 7190 5148 7196 5160
rect 7151 5120 7196 5148
rect 7190 5108 7196 5120
rect 7248 5108 7254 5160
rect 1670 5040 1676 5092
rect 1728 5080 1734 5092
rect 1765 5083 1823 5089
rect 1765 5080 1777 5083
rect 1728 5052 1777 5080
rect 1728 5040 1734 5052
rect 1765 5049 1777 5052
rect 1811 5080 1823 5083
rect 2498 5080 2504 5092
rect 1811 5052 2504 5080
rect 1811 5049 1823 5052
rect 1765 5043 1823 5049
rect 2498 5040 2504 5052
rect 2556 5040 2562 5092
rect 7300 5080 7328 5188
rect 7377 5185 7389 5188
rect 7423 5185 7435 5219
rect 8570 5216 8576 5228
rect 8531 5188 8576 5216
rect 7377 5179 7435 5185
rect 8570 5176 8576 5188
rect 8628 5176 8634 5228
rect 12894 5216 12900 5228
rect 12855 5188 12900 5216
rect 12894 5176 12900 5188
rect 12952 5176 12958 5228
rect 13081 5219 13139 5225
rect 13081 5185 13093 5219
rect 13127 5216 13139 5219
rect 13262 5216 13268 5228
rect 13127 5188 13268 5216
rect 13127 5185 13139 5188
rect 13081 5179 13139 5185
rect 13262 5176 13268 5188
rect 13320 5176 13326 5228
rect 15580 5225 15608 5256
rect 16025 5253 16037 5256
rect 16071 5284 16083 5287
rect 16071 5256 18368 5284
rect 16071 5253 16083 5256
rect 16025 5247 16083 5253
rect 18340 5228 18368 5256
rect 15565 5219 15623 5225
rect 15565 5185 15577 5219
rect 15611 5185 15623 5219
rect 16758 5216 16764 5228
rect 16719 5188 16764 5216
rect 15565 5179 15623 5185
rect 16758 5176 16764 5188
rect 16816 5176 16822 5228
rect 18322 5176 18328 5228
rect 18380 5216 18386 5228
rect 18601 5219 18659 5225
rect 18601 5216 18613 5219
rect 18380 5188 18613 5216
rect 18380 5176 18386 5188
rect 18601 5185 18613 5188
rect 18647 5185 18659 5219
rect 18601 5179 18659 5185
rect 18966 5176 18972 5228
rect 19024 5216 19030 5228
rect 20165 5219 20223 5225
rect 20165 5216 20177 5219
rect 19024 5188 20177 5216
rect 19024 5176 19030 5188
rect 20165 5185 20177 5188
rect 20211 5216 20223 5219
rect 20714 5216 20720 5228
rect 20211 5188 20720 5216
rect 20211 5185 20223 5188
rect 20165 5179 20223 5185
rect 20714 5176 20720 5188
rect 20772 5176 20778 5228
rect 11146 5108 11152 5160
rect 11204 5148 11210 5160
rect 11241 5151 11299 5157
rect 11241 5148 11253 5151
rect 11204 5120 11253 5148
rect 11204 5108 11210 5120
rect 11241 5117 11253 5120
rect 11287 5117 11299 5151
rect 11241 5111 11299 5117
rect 12434 5108 12440 5160
rect 12492 5148 12498 5160
rect 12805 5151 12863 5157
rect 12805 5148 12817 5151
rect 12492 5120 12817 5148
rect 12492 5108 12498 5120
rect 12805 5117 12817 5120
rect 12851 5117 12863 5151
rect 12805 5111 12863 5117
rect 16298 5108 16304 5160
rect 16356 5148 16362 5160
rect 16485 5151 16543 5157
rect 16485 5148 16497 5151
rect 16356 5120 16497 5148
rect 16356 5108 16362 5120
rect 16485 5117 16497 5120
rect 16531 5117 16543 5151
rect 16485 5111 16543 5117
rect 17865 5151 17923 5157
rect 17865 5117 17877 5151
rect 17911 5148 17923 5151
rect 18417 5151 18475 5157
rect 18417 5148 18429 5151
rect 17911 5120 18429 5148
rect 17911 5117 17923 5120
rect 17865 5111 17923 5117
rect 18417 5117 18429 5120
rect 18463 5148 18475 5151
rect 19242 5148 19248 5160
rect 18463 5120 19248 5148
rect 18463 5117 18475 5120
rect 18417 5111 18475 5117
rect 19242 5108 19248 5120
rect 19300 5108 19306 5160
rect 21174 5148 21180 5160
rect 21135 5120 21180 5148
rect 21174 5108 21180 5120
rect 21232 5148 21238 5160
rect 21913 5151 21971 5157
rect 21913 5148 21925 5151
rect 21232 5120 21925 5148
rect 21232 5108 21238 5120
rect 21913 5117 21925 5120
rect 21959 5117 21971 5151
rect 21913 5111 21971 5117
rect 6380 5052 7328 5080
rect 6380 5024 6408 5052
rect 8662 5040 8668 5092
rect 8720 5080 8726 5092
rect 8818 5083 8876 5089
rect 8818 5080 8830 5083
rect 8720 5052 8830 5080
rect 8720 5040 8726 5052
rect 8818 5049 8830 5052
rect 8864 5080 8876 5083
rect 10226 5080 10232 5092
rect 8864 5052 10232 5080
rect 8864 5049 8876 5052
rect 8818 5043 8876 5049
rect 10226 5040 10232 5052
rect 10284 5080 10290 5092
rect 10505 5083 10563 5089
rect 10505 5080 10517 5083
rect 10284 5052 10517 5080
rect 10284 5040 10290 5052
rect 10505 5049 10517 5052
rect 10551 5049 10563 5083
rect 10505 5043 10563 5049
rect 11330 5040 11336 5092
rect 11388 5080 11394 5092
rect 11793 5083 11851 5089
rect 11793 5080 11805 5083
rect 11388 5052 11805 5080
rect 11388 5040 11394 5052
rect 11793 5049 11805 5052
rect 11839 5080 11851 5083
rect 11974 5080 11980 5092
rect 11839 5052 11980 5080
rect 11839 5049 11851 5052
rect 11793 5043 11851 5049
rect 11974 5040 11980 5052
rect 12032 5040 12038 5092
rect 14550 5040 14556 5092
rect 14608 5080 14614 5092
rect 14737 5083 14795 5089
rect 14737 5080 14749 5083
rect 14608 5052 14749 5080
rect 14608 5040 14614 5052
rect 14737 5049 14749 5052
rect 14783 5080 14795 5083
rect 15378 5080 15384 5092
rect 14783 5052 15384 5080
rect 14783 5049 14795 5052
rect 14737 5043 14795 5049
rect 15378 5040 15384 5052
rect 15436 5040 15442 5092
rect 19981 5083 20039 5089
rect 19981 5080 19993 5083
rect 19076 5052 19993 5080
rect 19076 5024 19104 5052
rect 19981 5049 19993 5052
rect 20027 5049 20039 5083
rect 21450 5080 21456 5092
rect 21411 5052 21456 5080
rect 19981 5043 20039 5049
rect 21450 5040 21456 5052
rect 21508 5040 21514 5092
rect 2590 4972 2596 5024
rect 2648 5012 2654 5024
rect 2869 5015 2927 5021
rect 2869 5012 2881 5015
rect 2648 4984 2881 5012
rect 2648 4972 2654 4984
rect 2869 4981 2881 4984
rect 2915 5012 2927 5015
rect 3329 5015 3387 5021
rect 3329 5012 3341 5015
rect 2915 4984 3341 5012
rect 2915 4981 2927 4984
rect 2869 4975 2927 4981
rect 3329 4981 3341 4984
rect 3375 4981 3387 5015
rect 3329 4975 3387 4981
rect 3421 5015 3479 5021
rect 3421 4981 3433 5015
rect 3467 5012 3479 5015
rect 3878 5012 3884 5024
rect 3467 4984 3884 5012
rect 3467 4981 3479 4984
rect 3421 4975 3479 4981
rect 3878 4972 3884 4984
rect 3936 4972 3942 5024
rect 5350 4972 5356 5024
rect 5408 5012 5414 5024
rect 5629 5015 5687 5021
rect 5629 5012 5641 5015
rect 5408 4984 5641 5012
rect 5408 4972 5414 4984
rect 5629 4981 5641 4984
rect 5675 5012 5687 5015
rect 5994 5012 6000 5024
rect 5675 4984 6000 5012
rect 5675 4981 5687 4984
rect 5629 4975 5687 4981
rect 5994 4972 6000 4984
rect 6052 4972 6058 5024
rect 6273 5015 6331 5021
rect 6273 4981 6285 5015
rect 6319 5012 6331 5015
rect 6362 5012 6368 5024
rect 6319 4984 6368 5012
rect 6319 4981 6331 4984
rect 6273 4975 6331 4981
rect 6362 4972 6368 4984
rect 6420 4972 6426 5024
rect 6822 5012 6828 5024
rect 6783 4984 6828 5012
rect 6822 4972 6828 4984
rect 6880 4972 6886 5024
rect 7282 4972 7288 5024
rect 7340 5012 7346 5024
rect 7340 4984 7385 5012
rect 7340 4972 7346 4984
rect 7926 4972 7932 5024
rect 7984 5012 7990 5024
rect 8021 5015 8079 5021
rect 8021 5012 8033 5015
rect 7984 4984 8033 5012
rect 7984 4972 7990 4984
rect 8021 4981 8033 4984
rect 8067 5012 8079 5015
rect 8202 5012 8208 5024
rect 8067 4984 8208 5012
rect 8067 4981 8079 4984
rect 8021 4975 8079 4981
rect 8202 4972 8208 4984
rect 8260 4972 8266 5024
rect 8386 5012 8392 5024
rect 8347 4984 8392 5012
rect 8386 4972 8392 4984
rect 8444 4972 8450 5024
rect 9950 5012 9956 5024
rect 9911 4984 9956 5012
rect 9950 4972 9956 4984
rect 10008 4972 10014 5024
rect 11425 5015 11483 5021
rect 11425 4981 11437 5015
rect 11471 5012 11483 5015
rect 11606 5012 11612 5024
rect 11471 4984 11612 5012
rect 11471 4981 11483 4984
rect 11425 4975 11483 4981
rect 11606 4972 11612 4984
rect 11664 4972 11670 5024
rect 12434 4972 12440 5024
rect 12492 5012 12498 5024
rect 12492 4984 12537 5012
rect 12492 4972 12498 4984
rect 14918 4972 14924 5024
rect 14976 5012 14982 5024
rect 15289 5015 15347 5021
rect 15289 5012 15301 5015
rect 14976 4984 15301 5012
rect 14976 4972 14982 4984
rect 15289 4981 15301 4984
rect 15335 4981 15347 5015
rect 15289 4975 15347 4981
rect 16390 4972 16396 5024
rect 16448 5012 16454 5024
rect 16850 5012 16856 5024
rect 16448 4984 16856 5012
rect 16448 4972 16454 4984
rect 16850 4972 16856 4984
rect 16908 4972 16914 5024
rect 17218 5012 17224 5024
rect 17179 4984 17224 5012
rect 17218 4972 17224 4984
rect 17276 4972 17282 5024
rect 18506 4972 18512 5024
rect 18564 5012 18570 5024
rect 19058 5012 19064 5024
rect 18564 4984 18609 5012
rect 19019 4984 19064 5012
rect 18564 4972 18570 4984
rect 19058 4972 19064 4984
rect 19116 4972 19122 5024
rect 19334 4972 19340 5024
rect 19392 5012 19398 5024
rect 19429 5015 19487 5021
rect 19429 5012 19441 5015
rect 19392 4984 19441 5012
rect 19392 4972 19398 4984
rect 19429 4981 19441 4984
rect 19475 5012 19487 5015
rect 20073 5015 20131 5021
rect 20073 5012 20085 5015
rect 19475 4984 20085 5012
rect 19475 4981 19487 4984
rect 19429 4975 19487 4981
rect 20073 4981 20085 4984
rect 20119 4981 20131 5015
rect 20073 4975 20131 4981
rect 21358 4972 21364 5024
rect 21416 5012 21422 5024
rect 22094 5012 22100 5024
rect 21416 4984 22100 5012
rect 21416 4972 21422 4984
rect 22094 4972 22100 4984
rect 22152 4972 22158 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1670 4808 1676 4820
rect 1631 4780 1676 4808
rect 1670 4768 1676 4780
rect 1728 4768 1734 4820
rect 2317 4811 2375 4817
rect 2317 4777 2329 4811
rect 2363 4808 2375 4811
rect 2958 4808 2964 4820
rect 2363 4780 2964 4808
rect 2363 4777 2375 4780
rect 2317 4771 2375 4777
rect 2958 4768 2964 4780
rect 3016 4768 3022 4820
rect 3421 4811 3479 4817
rect 3421 4777 3433 4811
rect 3467 4808 3479 4811
rect 3602 4808 3608 4820
rect 3467 4780 3608 4808
rect 3467 4777 3479 4780
rect 3421 4771 3479 4777
rect 3602 4768 3608 4780
rect 3660 4768 3666 4820
rect 3789 4811 3847 4817
rect 3789 4777 3801 4811
rect 3835 4808 3847 4811
rect 4062 4808 4068 4820
rect 3835 4780 4068 4808
rect 3835 4777 3847 4780
rect 3789 4771 3847 4777
rect 4062 4768 4068 4780
rect 4120 4768 4126 4820
rect 5626 4808 5632 4820
rect 5587 4780 5632 4808
rect 5626 4768 5632 4780
rect 5684 4768 5690 4820
rect 6270 4808 6276 4820
rect 6231 4780 6276 4808
rect 6270 4768 6276 4780
rect 6328 4768 6334 4820
rect 6822 4768 6828 4820
rect 6880 4808 6886 4820
rect 7193 4811 7251 4817
rect 7193 4808 7205 4811
rect 6880 4780 7205 4808
rect 6880 4768 6886 4780
rect 7193 4777 7205 4780
rect 7239 4808 7251 4811
rect 7282 4808 7288 4820
rect 7239 4780 7288 4808
rect 7239 4777 7251 4780
rect 7193 4771 7251 4777
rect 7282 4768 7288 4780
rect 7340 4768 7346 4820
rect 8662 4808 8668 4820
rect 8623 4780 8668 4808
rect 8662 4768 8668 4780
rect 8720 4768 8726 4820
rect 9490 4808 9496 4820
rect 9451 4780 9496 4808
rect 9490 4768 9496 4780
rect 9548 4768 9554 4820
rect 9766 4768 9772 4820
rect 9824 4808 9830 4820
rect 10042 4808 10048 4820
rect 9824 4780 10048 4808
rect 9824 4768 9830 4780
rect 10042 4768 10048 4780
rect 10100 4768 10106 4820
rect 10137 4811 10195 4817
rect 10137 4777 10149 4811
rect 10183 4808 10195 4811
rect 10962 4808 10968 4820
rect 10183 4780 10968 4808
rect 10183 4777 10195 4780
rect 10137 4771 10195 4777
rect 10962 4768 10968 4780
rect 11020 4768 11026 4820
rect 12894 4768 12900 4820
rect 12952 4808 12958 4820
rect 12989 4811 13047 4817
rect 12989 4808 13001 4811
rect 12952 4780 13001 4808
rect 12952 4768 12958 4780
rect 12989 4777 13001 4780
rect 13035 4777 13047 4811
rect 13630 4808 13636 4820
rect 13591 4780 13636 4808
rect 12989 4771 13047 4777
rect 13630 4768 13636 4780
rect 13688 4808 13694 4820
rect 14553 4811 14611 4817
rect 14553 4808 14565 4811
rect 13688 4780 14565 4808
rect 13688 4768 13694 4780
rect 14553 4777 14565 4780
rect 14599 4777 14611 4811
rect 14553 4771 14611 4777
rect 17218 4768 17224 4820
rect 17276 4808 17282 4820
rect 17681 4811 17739 4817
rect 17681 4808 17693 4811
rect 17276 4780 17693 4808
rect 17276 4768 17282 4780
rect 17681 4777 17693 4780
rect 17727 4777 17739 4811
rect 18322 4808 18328 4820
rect 18283 4780 18328 4808
rect 17681 4771 17739 4777
rect 18322 4768 18328 4780
rect 18380 4768 18386 4820
rect 18598 4808 18604 4820
rect 18559 4780 18604 4808
rect 18598 4768 18604 4780
rect 18656 4768 18662 4820
rect 18782 4808 18788 4820
rect 18743 4780 18788 4808
rect 18782 4768 18788 4780
rect 18840 4768 18846 4820
rect 20530 4808 20536 4820
rect 20491 4780 20536 4808
rect 20530 4768 20536 4780
rect 20588 4808 20594 4820
rect 21358 4808 21364 4820
rect 20588 4780 21364 4808
rect 20588 4768 20594 4780
rect 21358 4768 21364 4780
rect 21416 4768 21422 4820
rect 3053 4743 3111 4749
rect 3053 4709 3065 4743
rect 3099 4740 3111 4743
rect 3878 4740 3884 4752
rect 3099 4712 3884 4740
rect 3099 4709 3111 4712
rect 3053 4703 3111 4709
rect 3878 4700 3884 4712
rect 3936 4700 3942 4752
rect 4430 4700 4436 4752
rect 4488 4749 4494 4752
rect 4488 4743 4552 4749
rect 4488 4709 4506 4743
rect 4540 4709 4552 4743
rect 4488 4703 4552 4709
rect 4488 4700 4494 4703
rect 9950 4700 9956 4752
rect 10008 4740 10014 4752
rect 10008 4712 10272 4740
rect 10008 4700 10014 4712
rect 2130 4632 2136 4684
rect 2188 4672 2194 4684
rect 2225 4675 2283 4681
rect 2225 4672 2237 4675
rect 2188 4644 2237 4672
rect 2188 4632 2194 4644
rect 2225 4641 2237 4644
rect 2271 4641 2283 4675
rect 2225 4635 2283 4641
rect 4062 4632 4068 4684
rect 4120 4672 4126 4684
rect 4249 4675 4307 4681
rect 4249 4672 4261 4675
rect 4120 4644 4261 4672
rect 4120 4632 4126 4644
rect 4249 4641 4261 4644
rect 4295 4672 4307 4675
rect 4982 4672 4988 4684
rect 4295 4644 4988 4672
rect 4295 4641 4307 4644
rect 4249 4635 4307 4641
rect 4982 4632 4988 4644
rect 5040 4632 5046 4684
rect 6917 4675 6975 4681
rect 6917 4641 6929 4675
rect 6963 4672 6975 4675
rect 7190 4672 7196 4684
rect 6963 4644 7196 4672
rect 6963 4641 6975 4644
rect 6917 4635 6975 4641
rect 7190 4632 7196 4644
rect 7248 4632 7254 4684
rect 7926 4672 7932 4684
rect 7887 4644 7932 4672
rect 7926 4632 7932 4644
rect 7984 4632 7990 4684
rect 8021 4675 8079 4681
rect 8021 4641 8033 4675
rect 8067 4672 8079 4675
rect 8202 4672 8208 4684
rect 8067 4644 8208 4672
rect 8067 4641 8079 4644
rect 8021 4635 8079 4641
rect 8202 4632 8208 4644
rect 8260 4632 8266 4684
rect 10244 4616 10272 4712
rect 14458 4700 14464 4752
rect 14516 4740 14522 4752
rect 14918 4740 14924 4752
rect 14516 4712 14924 4740
rect 14516 4700 14522 4712
rect 14918 4700 14924 4712
rect 14976 4740 14982 4752
rect 16298 4740 16304 4752
rect 14976 4712 16304 4740
rect 14976 4700 14982 4712
rect 16298 4700 16304 4712
rect 16356 4700 16362 4752
rect 11977 4675 12035 4681
rect 11977 4641 11989 4675
rect 12023 4672 12035 4675
rect 12342 4672 12348 4684
rect 12023 4644 12348 4672
rect 12023 4641 12035 4644
rect 11977 4635 12035 4641
rect 12342 4632 12348 4644
rect 12400 4632 12406 4684
rect 13446 4632 13452 4684
rect 13504 4672 13510 4684
rect 13541 4675 13599 4681
rect 13541 4672 13553 4675
rect 13504 4644 13553 4672
rect 13504 4632 13510 4644
rect 13541 4641 13553 4644
rect 13587 4672 13599 4675
rect 15289 4675 15347 4681
rect 15289 4672 15301 4675
rect 13587 4644 15301 4672
rect 13587 4641 13599 4644
rect 13541 4635 13599 4641
rect 15289 4641 15301 4644
rect 15335 4641 15347 4675
rect 15289 4635 15347 4641
rect 16206 4632 16212 4684
rect 16264 4672 16270 4684
rect 16557 4675 16615 4681
rect 16557 4672 16569 4675
rect 16264 4644 16569 4672
rect 16264 4632 16270 4644
rect 16557 4641 16569 4644
rect 16603 4641 16615 4675
rect 19150 4672 19156 4684
rect 19111 4644 19156 4672
rect 16557 4635 16615 4641
rect 19150 4632 19156 4644
rect 19208 4632 19214 4684
rect 20901 4675 20959 4681
rect 20901 4641 20913 4675
rect 20947 4672 20959 4675
rect 21450 4672 21456 4684
rect 20947 4644 21456 4672
rect 20947 4641 20959 4644
rect 20901 4635 20959 4641
rect 21450 4632 21456 4644
rect 21508 4632 21514 4684
rect 22370 4672 22376 4684
rect 22331 4644 22376 4672
rect 22370 4632 22376 4644
rect 22428 4632 22434 4684
rect 1946 4564 1952 4616
rect 2004 4604 2010 4616
rect 2409 4607 2467 4613
rect 2409 4604 2421 4607
rect 2004 4576 2421 4604
rect 2004 4564 2010 4576
rect 2409 4573 2421 4576
rect 2455 4604 2467 4607
rect 2774 4604 2780 4616
rect 2455 4576 2780 4604
rect 2455 4573 2467 4576
rect 2409 4567 2467 4573
rect 2774 4564 2780 4576
rect 2832 4564 2838 4616
rect 8110 4604 8116 4616
rect 8071 4576 8116 4604
rect 8110 4564 8116 4576
rect 8168 4564 8174 4616
rect 10226 4564 10232 4616
rect 10284 4604 10290 4616
rect 12069 4607 12127 4613
rect 10284 4576 10329 4604
rect 10284 4564 10290 4576
rect 12069 4573 12081 4607
rect 12115 4604 12127 4607
rect 12253 4607 12311 4613
rect 12115 4576 12149 4604
rect 12115 4573 12127 4576
rect 12069 4567 12127 4573
rect 12253 4573 12265 4607
rect 12299 4604 12311 4607
rect 13262 4604 13268 4616
rect 12299 4576 13268 4604
rect 12299 4573 12311 4576
rect 12253 4567 12311 4573
rect 1857 4539 1915 4545
rect 1857 4505 1869 4539
rect 1903 4536 1915 4539
rect 2682 4536 2688 4548
rect 1903 4508 2688 4536
rect 1903 4505 1915 4508
rect 1857 4499 1915 4505
rect 2682 4496 2688 4508
rect 2740 4496 2746 4548
rect 9766 4536 9772 4548
rect 9048 4508 9772 4536
rect 9048 4477 9076 4508
rect 9766 4496 9772 4508
rect 9824 4496 9830 4548
rect 11974 4496 11980 4548
rect 12032 4536 12038 4548
rect 12084 4536 12112 4567
rect 13262 4564 13268 4576
rect 13320 4564 13326 4616
rect 13817 4607 13875 4613
rect 13817 4573 13829 4607
rect 13863 4604 13875 4607
rect 16301 4607 16359 4613
rect 13863 4576 14136 4604
rect 13863 4573 13875 4576
rect 13817 4567 13875 4573
rect 12621 4539 12679 4545
rect 12621 4536 12633 4539
rect 12032 4508 12633 4536
rect 12032 4496 12038 4508
rect 12621 4505 12633 4508
rect 12667 4505 12679 4539
rect 12621 4499 12679 4505
rect 14108 4480 14136 4576
rect 16301 4573 16313 4607
rect 16347 4573 16359 4607
rect 19242 4604 19248 4616
rect 19203 4576 19248 4604
rect 16301 4567 16359 4573
rect 15286 4496 15292 4548
rect 15344 4536 15350 4548
rect 16316 4536 16344 4567
rect 19242 4564 19248 4576
rect 19300 4564 19306 4616
rect 19337 4607 19395 4613
rect 19337 4573 19349 4607
rect 19383 4604 19395 4607
rect 19797 4607 19855 4613
rect 19797 4604 19809 4607
rect 19383 4576 19809 4604
rect 19383 4573 19395 4576
rect 19337 4567 19395 4573
rect 19797 4573 19809 4576
rect 19843 4573 19855 4607
rect 19797 4567 19855 4573
rect 22649 4607 22707 4613
rect 22649 4573 22661 4607
rect 22695 4604 22707 4607
rect 23474 4604 23480 4616
rect 22695 4576 23480 4604
rect 22695 4573 22707 4576
rect 22649 4567 22707 4573
rect 15344 4508 16344 4536
rect 15344 4496 15350 4508
rect 7561 4471 7619 4477
rect 7561 4437 7573 4471
rect 7607 4468 7619 4471
rect 9033 4471 9091 4477
rect 9033 4468 9045 4471
rect 7607 4440 9045 4468
rect 7607 4437 7619 4440
rect 7561 4431 7619 4437
rect 9033 4437 9045 4440
rect 9079 4437 9091 4471
rect 9674 4468 9680 4480
rect 9635 4440 9680 4468
rect 9033 4431 9091 4437
rect 9674 4428 9680 4440
rect 9732 4428 9738 4480
rect 10686 4468 10692 4480
rect 10647 4440 10692 4468
rect 10686 4428 10692 4440
rect 10744 4428 10750 4480
rect 11146 4428 11152 4480
rect 11204 4468 11210 4480
rect 11241 4471 11299 4477
rect 11241 4468 11253 4471
rect 11204 4440 11253 4468
rect 11204 4428 11210 4440
rect 11241 4437 11253 4440
rect 11287 4437 11299 4471
rect 11241 4431 11299 4437
rect 11609 4471 11667 4477
rect 11609 4437 11621 4471
rect 11655 4468 11667 4471
rect 12066 4468 12072 4480
rect 11655 4440 12072 4468
rect 11655 4437 11667 4440
rect 11609 4431 11667 4437
rect 12066 4428 12072 4440
rect 12124 4428 12130 4480
rect 13170 4468 13176 4480
rect 13131 4440 13176 4468
rect 13170 4428 13176 4440
rect 13228 4428 13234 4480
rect 14090 4428 14096 4480
rect 14148 4468 14154 4480
rect 14185 4471 14243 4477
rect 14185 4468 14197 4471
rect 14148 4440 14197 4468
rect 14148 4428 14154 4440
rect 14185 4437 14197 4440
rect 14231 4437 14243 4471
rect 15838 4468 15844 4480
rect 15799 4440 15844 4468
rect 14185 4431 14243 4437
rect 15838 4428 15844 4440
rect 15896 4428 15902 4480
rect 16206 4468 16212 4480
rect 16167 4440 16212 4468
rect 16206 4428 16212 4440
rect 16264 4428 16270 4480
rect 16316 4468 16344 4508
rect 18966 4496 18972 4548
rect 19024 4536 19030 4548
rect 19352 4536 19380 4567
rect 23474 4564 23480 4576
rect 23532 4564 23538 4616
rect 19024 4508 19380 4536
rect 19024 4496 19030 4508
rect 16574 4468 16580 4480
rect 16316 4440 16580 4468
rect 16574 4428 16580 4440
rect 16632 4428 16638 4480
rect 20254 4468 20260 4480
rect 20167 4440 20260 4468
rect 20254 4428 20260 4440
rect 20312 4468 20318 4480
rect 20622 4468 20628 4480
rect 20312 4440 20628 4468
rect 20312 4428 20318 4440
rect 20622 4428 20628 4440
rect 20680 4428 20686 4480
rect 21085 4471 21143 4477
rect 21085 4437 21097 4471
rect 21131 4468 21143 4471
rect 23106 4468 23112 4480
rect 21131 4440 23112 4468
rect 21131 4437 21143 4440
rect 21085 4431 21143 4437
rect 23106 4428 23112 4440
rect 23164 4428 23170 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 6273 4267 6331 4273
rect 6273 4233 6285 4267
rect 6319 4264 6331 4267
rect 6362 4264 6368 4276
rect 6319 4236 6368 4264
rect 6319 4233 6331 4236
rect 6273 4227 6331 4233
rect 2222 4088 2228 4140
rect 2280 4128 2286 4140
rect 2409 4131 2467 4137
rect 2409 4128 2421 4131
rect 2280 4100 2421 4128
rect 2280 4088 2286 4100
rect 2409 4097 2421 4100
rect 2455 4097 2467 4131
rect 2409 4091 2467 4097
rect 2774 4088 2780 4140
rect 2832 4128 2838 4140
rect 2869 4131 2927 4137
rect 2869 4128 2881 4131
rect 2832 4100 2881 4128
rect 2832 4088 2838 4100
rect 2869 4097 2881 4100
rect 2915 4128 2927 4131
rect 3237 4131 3295 4137
rect 3237 4128 3249 4131
rect 2915 4100 3249 4128
rect 2915 4097 2927 4100
rect 2869 4091 2927 4097
rect 3237 4097 3249 4100
rect 3283 4097 3295 4131
rect 3237 4091 3295 4097
rect 4065 4131 4123 4137
rect 4065 4097 4077 4131
rect 4111 4128 4123 4131
rect 4154 4128 4160 4140
rect 4111 4100 4160 4128
rect 4111 4097 4123 4100
rect 4065 4091 4123 4097
rect 4154 4088 4160 4100
rect 4212 4088 4218 4140
rect 5077 4131 5135 4137
rect 5077 4097 5089 4131
rect 5123 4128 5135 4131
rect 5258 4128 5264 4140
rect 5123 4100 5264 4128
rect 5123 4097 5135 4100
rect 5077 4091 5135 4097
rect 5258 4088 5264 4100
rect 5316 4128 5322 4140
rect 5629 4131 5687 4137
rect 5629 4128 5641 4131
rect 5316 4100 5641 4128
rect 5316 4088 5322 4100
rect 5629 4097 5641 4100
rect 5675 4097 5687 4131
rect 5629 4091 5687 4097
rect 5813 4131 5871 4137
rect 5813 4097 5825 4131
rect 5859 4128 5871 4131
rect 6288 4128 6316 4227
rect 6362 4224 6368 4236
rect 6420 4224 6426 4276
rect 10042 4224 10048 4276
rect 10100 4264 10106 4276
rect 10689 4267 10747 4273
rect 10689 4264 10701 4267
rect 10100 4236 10701 4264
rect 10100 4224 10106 4236
rect 10689 4233 10701 4236
rect 10735 4264 10747 4267
rect 12989 4267 13047 4273
rect 12989 4264 13001 4267
rect 10735 4236 13001 4264
rect 10735 4233 10747 4236
rect 10689 4227 10747 4233
rect 7282 4128 7288 4140
rect 5859 4100 6316 4128
rect 7243 4100 7288 4128
rect 5859 4097 5871 4100
rect 5813 4091 5871 4097
rect 7282 4088 7288 4100
rect 7340 4088 7346 4140
rect 7377 4131 7435 4137
rect 7377 4097 7389 4131
rect 7423 4097 7435 4131
rect 7377 4091 7435 4097
rect 1765 4063 1823 4069
rect 1765 4029 1777 4063
rect 1811 4060 1823 4063
rect 2314 4060 2320 4072
rect 1811 4032 2320 4060
rect 1811 4029 1823 4032
rect 1765 4023 1823 4029
rect 2314 4020 2320 4032
rect 2372 4020 2378 4072
rect 3050 4020 3056 4072
rect 3108 4060 3114 4072
rect 3418 4060 3424 4072
rect 3108 4032 3424 4060
rect 3108 4020 3114 4032
rect 3418 4020 3424 4032
rect 3476 4020 3482 4072
rect 7392 4060 7420 4091
rect 8570 4088 8576 4140
rect 8628 4128 8634 4140
rect 8757 4131 8815 4137
rect 8757 4128 8769 4131
rect 8628 4100 8769 4128
rect 8628 4088 8634 4100
rect 8757 4097 8769 4100
rect 8803 4097 8815 4131
rect 8757 4091 8815 4097
rect 7837 4063 7895 4069
rect 7837 4060 7849 4063
rect 6656 4032 7849 4060
rect 2130 3992 2136 4004
rect 1872 3964 2136 3992
rect 1872 3933 1900 3964
rect 2130 3952 2136 3964
rect 2188 3992 2194 4004
rect 2958 3992 2964 4004
rect 2188 3964 2964 3992
rect 2188 3952 2194 3964
rect 2958 3952 2964 3964
rect 3016 3952 3022 4004
rect 3786 3992 3792 4004
rect 3747 3964 3792 3992
rect 3786 3952 3792 3964
rect 3844 3952 3850 4004
rect 4709 3995 4767 4001
rect 4709 3961 4721 3995
rect 4755 3992 4767 3995
rect 5534 3992 5540 4004
rect 4755 3964 5540 3992
rect 4755 3961 4767 3964
rect 4709 3955 4767 3961
rect 5534 3952 5540 3964
rect 5592 3952 5598 4004
rect 6656 3936 6684 4032
rect 7837 4029 7849 4032
rect 7883 4060 7895 4063
rect 8110 4060 8116 4072
rect 7883 4032 8116 4060
rect 7883 4029 7895 4032
rect 7837 4023 7895 4029
rect 8110 4020 8116 4032
rect 8168 4020 8174 4072
rect 11238 4060 11244 4072
rect 11199 4032 11244 4060
rect 11238 4020 11244 4032
rect 11296 4060 11302 4072
rect 12452 4069 12480 4236
rect 12989 4233 13001 4236
rect 13035 4233 13047 4267
rect 13446 4264 13452 4276
rect 13407 4236 13452 4264
rect 12989 4227 13047 4233
rect 13446 4224 13452 4236
rect 13504 4224 13510 4276
rect 16390 4264 16396 4276
rect 16351 4236 16396 4264
rect 16390 4224 16396 4236
rect 16448 4224 16454 4276
rect 19150 4264 19156 4276
rect 19111 4236 19156 4264
rect 19150 4224 19156 4236
rect 19208 4224 19214 4276
rect 21450 4224 21456 4276
rect 21508 4264 21514 4276
rect 21637 4267 21695 4273
rect 21637 4264 21649 4267
rect 21508 4236 21649 4264
rect 21508 4224 21514 4236
rect 21637 4233 21649 4236
rect 21683 4233 21695 4267
rect 22370 4264 22376 4276
rect 22331 4236 22376 4264
rect 21637 4227 21695 4233
rect 22370 4224 22376 4236
rect 22428 4224 22434 4276
rect 15838 4156 15844 4208
rect 15896 4196 15902 4208
rect 17218 4196 17224 4208
rect 15896 4168 17224 4196
rect 15896 4156 15902 4168
rect 15930 4088 15936 4140
rect 15988 4128 15994 4140
rect 16960 4137 16988 4168
rect 17218 4156 17224 4168
rect 17276 4156 17282 4208
rect 18598 4156 18604 4208
rect 18656 4196 18662 4208
rect 18656 4168 18736 4196
rect 18656 4156 18662 4168
rect 16117 4131 16175 4137
rect 16117 4128 16129 4131
rect 15988 4100 16129 4128
rect 15988 4088 15994 4100
rect 16117 4097 16129 4100
rect 16163 4128 16175 4131
rect 16209 4131 16267 4137
rect 16209 4128 16221 4131
rect 16163 4100 16221 4128
rect 16163 4097 16175 4100
rect 16117 4091 16175 4097
rect 16209 4097 16221 4100
rect 16255 4097 16267 4131
rect 16209 4091 16267 4097
rect 16945 4131 17003 4137
rect 16945 4097 16957 4131
rect 16991 4097 17003 4131
rect 16945 4091 17003 4097
rect 17126 4088 17132 4140
rect 17184 4128 17190 4140
rect 17405 4131 17463 4137
rect 17405 4128 17417 4131
rect 17184 4100 17417 4128
rect 17184 4088 17190 4100
rect 17405 4097 17417 4100
rect 17451 4128 17463 4131
rect 17681 4131 17739 4137
rect 17681 4128 17693 4131
rect 17451 4100 17693 4128
rect 17451 4097 17463 4100
rect 17405 4091 17463 4097
rect 17681 4097 17693 4100
rect 17727 4097 17739 4131
rect 17862 4128 17868 4140
rect 17775 4100 17868 4128
rect 17681 4091 17739 4097
rect 17862 4088 17868 4100
rect 17920 4128 17926 4140
rect 18414 4128 18420 4140
rect 17920 4100 18420 4128
rect 17920 4088 17926 4100
rect 18414 4088 18420 4100
rect 18472 4128 18478 4140
rect 18708 4137 18736 4168
rect 18509 4131 18567 4137
rect 18509 4128 18521 4131
rect 18472 4100 18521 4128
rect 18472 4088 18478 4100
rect 18509 4097 18521 4100
rect 18555 4097 18567 4131
rect 18509 4091 18567 4097
rect 18693 4131 18751 4137
rect 18693 4097 18705 4131
rect 18739 4097 18751 4131
rect 18693 4091 18751 4097
rect 19536 4100 20760 4128
rect 11793 4063 11851 4069
rect 11793 4060 11805 4063
rect 11296 4032 11805 4060
rect 11296 4020 11302 4032
rect 11793 4029 11805 4032
rect 11839 4029 11851 4063
rect 11793 4023 11851 4029
rect 12443 4063 12501 4069
rect 12443 4029 12455 4063
rect 12489 4029 12501 4063
rect 12443 4023 12501 4029
rect 13446 4020 13452 4072
rect 13504 4060 13510 4072
rect 13817 4063 13875 4069
rect 13817 4060 13829 4063
rect 13504 4032 13829 4060
rect 13504 4020 13510 4032
rect 13817 4029 13829 4032
rect 13863 4029 13875 4063
rect 13817 4023 13875 4029
rect 13906 4020 13912 4072
rect 13964 4060 13970 4072
rect 14366 4060 14372 4072
rect 13964 4032 14372 4060
rect 13964 4020 13970 4032
rect 14366 4020 14372 4032
rect 14424 4020 14430 4072
rect 15746 4020 15752 4072
rect 15804 4060 15810 4072
rect 15841 4063 15899 4069
rect 15841 4060 15853 4063
rect 15804 4032 15853 4060
rect 15804 4020 15810 4032
rect 15841 4029 15853 4032
rect 15887 4060 15899 4063
rect 16853 4063 16911 4069
rect 16853 4060 16865 4063
rect 15887 4032 16865 4060
rect 15887 4029 15899 4032
rect 15841 4023 15899 4029
rect 16853 4029 16865 4032
rect 16899 4060 16911 4063
rect 19536 4060 19564 4100
rect 16899 4032 19564 4060
rect 19613 4063 19671 4069
rect 16899 4029 16911 4032
rect 16853 4023 16911 4029
rect 19613 4029 19625 4063
rect 19659 4060 19671 4063
rect 19978 4060 19984 4072
rect 19659 4032 19984 4060
rect 19659 4029 19671 4032
rect 19613 4023 19671 4029
rect 19978 4020 19984 4032
rect 20036 4060 20042 4072
rect 20165 4063 20223 4069
rect 20165 4060 20177 4063
rect 20036 4032 20177 4060
rect 20036 4020 20042 4032
rect 20165 4029 20177 4032
rect 20211 4029 20223 4063
rect 20165 4023 20223 4029
rect 20346 4020 20352 4072
rect 20404 4060 20410 4072
rect 20732 4069 20760 4100
rect 20533 4063 20591 4069
rect 20533 4060 20545 4063
rect 20404 4032 20545 4060
rect 20404 4020 20410 4032
rect 20533 4029 20545 4032
rect 20579 4029 20591 4063
rect 20533 4023 20591 4029
rect 20717 4063 20775 4069
rect 20717 4029 20729 4063
rect 20763 4060 20775 4063
rect 21269 4063 21327 4069
rect 21269 4060 21281 4063
rect 20763 4032 21281 4060
rect 20763 4029 20775 4032
rect 20717 4023 20775 4029
rect 21269 4029 21281 4032
rect 21315 4029 21327 4063
rect 21818 4060 21824 4072
rect 21779 4032 21824 4060
rect 21269 4023 21327 4029
rect 21818 4020 21824 4032
rect 21876 4020 21882 4072
rect 23474 4020 23480 4072
rect 23532 4060 23538 4072
rect 23661 4063 23719 4069
rect 23661 4060 23673 4063
rect 23532 4032 23673 4060
rect 23532 4020 23538 4032
rect 23661 4029 23673 4032
rect 23707 4060 23719 4063
rect 24213 4063 24271 4069
rect 24213 4060 24225 4063
rect 23707 4032 24225 4060
rect 23707 4029 23719 4032
rect 23661 4023 23719 4029
rect 24213 4029 24225 4032
rect 24259 4029 24271 4063
rect 24213 4023 24271 4029
rect 8665 3995 8723 4001
rect 8665 3961 8677 3995
rect 8711 3992 8723 3995
rect 9024 3995 9082 4001
rect 9024 3992 9036 3995
rect 8711 3964 9036 3992
rect 8711 3961 8723 3964
rect 8665 3955 8723 3961
rect 9024 3961 9036 3964
rect 9070 3992 9082 3995
rect 9490 3992 9496 4004
rect 9070 3964 9496 3992
rect 9070 3961 9082 3964
rect 9024 3955 9082 3961
rect 9490 3952 9496 3964
rect 9548 3992 9554 4004
rect 10226 3992 10232 4004
rect 9548 3964 10232 3992
rect 9548 3952 9554 3964
rect 10226 3952 10232 3964
rect 10284 3952 10290 4004
rect 11054 3952 11060 4004
rect 11112 3992 11118 4004
rect 11149 3995 11207 4001
rect 11149 3992 11161 3995
rect 11112 3964 11161 3992
rect 11112 3952 11118 3964
rect 11149 3961 11161 3964
rect 11195 3992 11207 3995
rect 11882 3992 11888 4004
rect 11195 3964 11888 3992
rect 11195 3961 11207 3964
rect 11149 3955 11207 3961
rect 11882 3952 11888 3964
rect 11940 3952 11946 4004
rect 12253 3995 12311 4001
rect 12253 3961 12265 3995
rect 12299 3992 12311 3995
rect 13262 3992 13268 4004
rect 12299 3964 13268 3992
rect 12299 3961 12311 3964
rect 12253 3955 12311 3961
rect 13262 3952 13268 3964
rect 13320 3992 13326 4004
rect 14090 4001 14096 4004
rect 14062 3995 14096 4001
rect 14062 3992 14074 3995
rect 13320 3964 14074 3992
rect 13320 3952 13326 3964
rect 14062 3961 14074 3964
rect 14148 3992 14154 4004
rect 16117 3995 16175 4001
rect 14148 3964 14210 3992
rect 14062 3955 14096 3961
rect 14090 3952 14096 3955
rect 14148 3952 14154 3964
rect 16117 3961 16129 3995
rect 16163 3992 16175 3995
rect 16758 3992 16764 4004
rect 16163 3964 16764 3992
rect 16163 3961 16175 3964
rect 16117 3955 16175 3961
rect 16758 3952 16764 3964
rect 16816 3952 16822 4004
rect 17681 3995 17739 4001
rect 17681 3961 17693 3995
rect 17727 3992 17739 3995
rect 18417 3995 18475 4001
rect 18417 3992 18429 3995
rect 17727 3964 18429 3992
rect 17727 3961 17739 3964
rect 17681 3955 17739 3961
rect 18417 3961 18429 3964
rect 18463 3961 18475 3995
rect 18417 3955 18475 3961
rect 20254 3952 20260 4004
rect 20312 3992 20318 4004
rect 20312 3964 20944 3992
rect 20312 3952 20318 3964
rect 1857 3927 1915 3933
rect 1857 3893 1869 3927
rect 1903 3893 1915 3927
rect 1857 3887 1915 3893
rect 1946 3884 1952 3936
rect 2004 3924 2010 3936
rect 2225 3927 2283 3933
rect 2225 3924 2237 3927
rect 2004 3896 2237 3924
rect 2004 3884 2010 3896
rect 2225 3893 2237 3896
rect 2271 3893 2283 3927
rect 2225 3887 2283 3893
rect 2314 3884 2320 3936
rect 2372 3924 2378 3936
rect 3418 3924 3424 3936
rect 2372 3896 2417 3924
rect 3379 3896 3424 3924
rect 2372 3884 2378 3896
rect 3418 3884 3424 3896
rect 3476 3884 3482 3936
rect 3878 3924 3884 3936
rect 3839 3896 3884 3924
rect 3878 3884 3884 3896
rect 3936 3884 3942 3936
rect 5166 3924 5172 3936
rect 5127 3896 5172 3924
rect 5166 3884 5172 3896
rect 5224 3884 5230 3936
rect 6638 3924 6644 3936
rect 6599 3896 6644 3924
rect 6638 3884 6644 3896
rect 6696 3884 6702 3936
rect 6822 3924 6828 3936
rect 6783 3896 6828 3924
rect 6822 3884 6828 3896
rect 6880 3884 6886 3936
rect 7190 3924 7196 3936
rect 7151 3896 7196 3924
rect 7190 3884 7196 3896
rect 7248 3884 7254 3936
rect 8294 3924 8300 3936
rect 8255 3896 8300 3924
rect 8294 3884 8300 3896
rect 8352 3884 8358 3936
rect 10042 3884 10048 3936
rect 10100 3924 10106 3936
rect 10137 3927 10195 3933
rect 10137 3924 10149 3927
rect 10100 3896 10149 3924
rect 10100 3884 10106 3896
rect 10137 3893 10149 3896
rect 10183 3893 10195 3927
rect 11422 3924 11428 3936
rect 11383 3896 11428 3924
rect 10137 3887 10195 3893
rect 11422 3884 11428 3896
rect 11480 3884 11486 3936
rect 12621 3927 12679 3933
rect 12621 3893 12633 3927
rect 12667 3924 12679 3927
rect 13630 3924 13636 3936
rect 12667 3896 13636 3924
rect 12667 3893 12679 3896
rect 12621 3887 12679 3893
rect 13630 3884 13636 3896
rect 13688 3884 13694 3936
rect 13722 3884 13728 3936
rect 13780 3924 13786 3936
rect 15194 3924 15200 3936
rect 13780 3896 15200 3924
rect 13780 3884 13786 3896
rect 15194 3884 15200 3896
rect 15252 3884 15258 3936
rect 17954 3884 17960 3936
rect 18012 3924 18018 3936
rect 18049 3927 18107 3933
rect 18049 3924 18061 3927
rect 18012 3896 18061 3924
rect 18012 3884 18018 3896
rect 18049 3893 18061 3896
rect 18095 3893 18107 3927
rect 18049 3887 18107 3893
rect 19242 3884 19248 3936
rect 19300 3924 19306 3936
rect 19518 3924 19524 3936
rect 19300 3896 19524 3924
rect 19300 3884 19306 3896
rect 19518 3884 19524 3896
rect 19576 3884 19582 3936
rect 19797 3927 19855 3933
rect 19797 3893 19809 3927
rect 19843 3924 19855 3927
rect 20070 3924 20076 3936
rect 19843 3896 20076 3924
rect 19843 3893 19855 3896
rect 19797 3887 19855 3893
rect 20070 3884 20076 3896
rect 20128 3884 20134 3936
rect 20916 3933 20944 3964
rect 20901 3927 20959 3933
rect 20901 3893 20913 3927
rect 20947 3893 20959 3927
rect 22002 3924 22008 3936
rect 21963 3896 22008 3924
rect 20901 3887 20959 3893
rect 22002 3884 22008 3896
rect 22060 3884 22066 3936
rect 23845 3927 23903 3933
rect 23845 3893 23857 3927
rect 23891 3924 23903 3927
rect 25314 3924 25320 3936
rect 23891 3896 25320 3924
rect 23891 3893 23903 3896
rect 23845 3887 23903 3893
rect 25314 3884 25320 3896
rect 25372 3884 25378 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1946 3720 1952 3732
rect 1907 3692 1952 3720
rect 1946 3680 1952 3692
rect 2004 3680 2010 3732
rect 2222 3720 2228 3732
rect 2183 3692 2228 3720
rect 2222 3680 2228 3692
rect 2280 3680 2286 3732
rect 2406 3720 2412 3732
rect 2367 3692 2412 3720
rect 2406 3680 2412 3692
rect 2464 3680 2470 3732
rect 2777 3723 2835 3729
rect 2777 3689 2789 3723
rect 2823 3720 2835 3723
rect 3418 3720 3424 3732
rect 2823 3692 3424 3720
rect 2823 3689 2835 3692
rect 2777 3683 2835 3689
rect 3418 3680 3424 3692
rect 3476 3680 3482 3732
rect 5166 3680 5172 3732
rect 5224 3720 5230 3732
rect 6549 3723 6607 3729
rect 6549 3720 6561 3723
rect 5224 3692 6561 3720
rect 5224 3680 5230 3692
rect 6549 3689 6561 3692
rect 6595 3720 6607 3723
rect 7190 3720 7196 3732
rect 6595 3692 7196 3720
rect 6595 3689 6607 3692
rect 6549 3683 6607 3689
rect 7190 3680 7196 3692
rect 7248 3680 7254 3732
rect 7561 3723 7619 3729
rect 7561 3689 7573 3723
rect 7607 3720 7619 3723
rect 7926 3720 7932 3732
rect 7607 3692 7932 3720
rect 7607 3689 7619 3692
rect 7561 3683 7619 3689
rect 7926 3680 7932 3692
rect 7984 3720 7990 3732
rect 8021 3723 8079 3729
rect 8021 3720 8033 3723
rect 7984 3692 8033 3720
rect 7984 3680 7990 3692
rect 8021 3689 8033 3692
rect 8067 3689 8079 3723
rect 8021 3683 8079 3689
rect 8294 3680 8300 3732
rect 8352 3720 8358 3732
rect 9677 3723 9735 3729
rect 9677 3720 9689 3723
rect 8352 3692 9689 3720
rect 8352 3680 8358 3692
rect 9677 3689 9689 3692
rect 9723 3689 9735 3723
rect 9677 3683 9735 3689
rect 10045 3723 10103 3729
rect 10045 3689 10057 3723
rect 10091 3720 10103 3723
rect 11238 3720 11244 3732
rect 10091 3692 11244 3720
rect 10091 3689 10103 3692
rect 10045 3683 10103 3689
rect 11238 3680 11244 3692
rect 11296 3680 11302 3732
rect 11701 3723 11759 3729
rect 11701 3689 11713 3723
rect 11747 3720 11759 3723
rect 12526 3720 12532 3732
rect 11747 3692 12532 3720
rect 11747 3689 11759 3692
rect 11701 3683 11759 3689
rect 12526 3680 12532 3692
rect 12584 3680 12590 3732
rect 13170 3680 13176 3732
rect 13228 3720 13234 3732
rect 13725 3723 13783 3729
rect 13725 3720 13737 3723
rect 13228 3692 13737 3720
rect 13228 3680 13234 3692
rect 13725 3689 13737 3692
rect 13771 3720 13783 3723
rect 13814 3720 13820 3732
rect 13771 3692 13820 3720
rect 13771 3689 13783 3692
rect 13725 3683 13783 3689
rect 13814 3680 13820 3692
rect 13872 3680 13878 3732
rect 18141 3723 18199 3729
rect 18141 3689 18153 3723
rect 18187 3720 18199 3723
rect 18322 3720 18328 3732
rect 18187 3692 18328 3720
rect 18187 3689 18199 3692
rect 18141 3683 18199 3689
rect 18322 3680 18328 3692
rect 18380 3680 18386 3732
rect 18877 3723 18935 3729
rect 18877 3689 18889 3723
rect 18923 3720 18935 3723
rect 18966 3720 18972 3732
rect 18923 3692 18972 3720
rect 18923 3689 18935 3692
rect 18877 3683 18935 3689
rect 18966 3680 18972 3692
rect 19024 3680 19030 3732
rect 19981 3723 20039 3729
rect 19981 3689 19993 3723
rect 20027 3720 20039 3723
rect 20162 3720 20168 3732
rect 20027 3692 20168 3720
rect 20027 3689 20039 3692
rect 19981 3683 20039 3689
rect 20162 3680 20168 3692
rect 20220 3720 20226 3732
rect 20346 3720 20352 3732
rect 20220 3692 20352 3720
rect 20220 3680 20226 3692
rect 20346 3680 20352 3692
rect 20404 3680 20410 3732
rect 20714 3720 20720 3732
rect 20675 3692 20720 3720
rect 20714 3680 20720 3692
rect 20772 3680 20778 3732
rect 21358 3680 21364 3732
rect 21416 3720 21422 3732
rect 21453 3723 21511 3729
rect 21453 3720 21465 3723
rect 21416 3692 21465 3720
rect 21416 3680 21422 3692
rect 21453 3689 21465 3692
rect 21499 3689 21511 3723
rect 21453 3683 21511 3689
rect 2869 3655 2927 3661
rect 2869 3621 2881 3655
rect 2915 3652 2927 3655
rect 3142 3652 3148 3664
rect 2915 3624 3148 3652
rect 2915 3621 2927 3624
rect 2869 3615 2927 3621
rect 3142 3612 3148 3624
rect 3200 3612 3206 3664
rect 4154 3612 4160 3664
rect 4212 3652 4218 3664
rect 4310 3655 4368 3661
rect 4310 3652 4322 3655
rect 4212 3624 4322 3652
rect 4212 3612 4218 3624
rect 4310 3621 4322 3624
rect 4356 3621 4368 3655
rect 4310 3615 4368 3621
rect 6362 3612 6368 3664
rect 6420 3652 6426 3664
rect 7837 3655 7895 3661
rect 7837 3652 7849 3655
rect 6420 3624 7849 3652
rect 6420 3612 6426 3624
rect 7837 3621 7849 3624
rect 7883 3621 7895 3655
rect 7837 3615 7895 3621
rect 4062 3584 4068 3596
rect 4023 3556 4068 3584
rect 4062 3544 4068 3556
rect 4120 3544 4126 3596
rect 6730 3584 6736 3596
rect 6691 3556 6736 3584
rect 6730 3544 6736 3556
rect 6788 3544 6794 3596
rect 7009 3587 7067 3593
rect 7009 3553 7021 3587
rect 7055 3584 7067 3587
rect 7098 3584 7104 3596
rect 7055 3556 7104 3584
rect 7055 3553 7067 3556
rect 7009 3547 7067 3553
rect 7098 3544 7104 3556
rect 7156 3544 7162 3596
rect 3053 3519 3111 3525
rect 3053 3485 3065 3519
rect 3099 3516 3111 3519
rect 6086 3516 6092 3528
rect 3099 3488 3924 3516
rect 5999 3488 6092 3516
rect 3099 3485 3111 3488
rect 3053 3479 3111 3485
rect 2498 3408 2504 3460
rect 2556 3448 2562 3460
rect 3068 3448 3096 3479
rect 2556 3420 3096 3448
rect 2556 3408 2562 3420
rect 2866 3340 2872 3392
rect 2924 3380 2930 3392
rect 3050 3380 3056 3392
rect 2924 3352 3056 3380
rect 2924 3340 2930 3352
rect 3050 3340 3056 3352
rect 3108 3380 3114 3392
rect 3896 3389 3924 3488
rect 6086 3476 6092 3488
rect 6144 3516 6150 3528
rect 6822 3516 6828 3528
rect 6144 3488 6828 3516
rect 6144 3476 6150 3488
rect 6822 3476 6828 3488
rect 6880 3476 6886 3528
rect 7852 3516 7880 3615
rect 10134 3612 10140 3664
rect 10192 3652 10198 3664
rect 10870 3652 10876 3664
rect 10192 3624 10876 3652
rect 10192 3612 10198 3624
rect 10870 3612 10876 3624
rect 10928 3612 10934 3664
rect 15194 3612 15200 3664
rect 15252 3652 15258 3664
rect 15534 3655 15592 3661
rect 15534 3652 15546 3655
rect 15252 3624 15546 3652
rect 15252 3612 15258 3624
rect 15534 3621 15546 3624
rect 15580 3652 15592 3655
rect 15930 3652 15936 3664
rect 15580 3624 15936 3652
rect 15580 3621 15592 3624
rect 15534 3615 15592 3621
rect 15930 3612 15936 3624
rect 15988 3612 15994 3664
rect 8386 3584 8392 3596
rect 8347 3556 8392 3584
rect 8386 3544 8392 3556
rect 8444 3544 8450 3596
rect 8481 3587 8539 3593
rect 8481 3553 8493 3587
rect 8527 3584 8539 3587
rect 8754 3584 8760 3596
rect 8527 3556 8760 3584
rect 8527 3553 8539 3556
rect 8481 3547 8539 3553
rect 8754 3544 8760 3556
rect 8812 3544 8818 3596
rect 10042 3584 10048 3596
rect 9048 3556 10048 3584
rect 9048 3525 9076 3556
rect 10042 3544 10048 3556
rect 10100 3584 10106 3596
rect 10100 3556 10272 3584
rect 10100 3544 10106 3556
rect 8573 3519 8631 3525
rect 8573 3516 8585 3519
rect 7852 3488 8585 3516
rect 8573 3485 8585 3488
rect 8619 3516 8631 3519
rect 9033 3519 9091 3525
rect 9033 3516 9045 3519
rect 8619 3488 9045 3516
rect 8619 3485 8631 3488
rect 8573 3479 8631 3485
rect 9033 3485 9045 3488
rect 9079 3485 9091 3519
rect 9033 3479 9091 3485
rect 9674 3476 9680 3528
rect 9732 3516 9738 3528
rect 10244 3525 10272 3556
rect 11514 3544 11520 3596
rect 11572 3584 11578 3596
rect 11609 3587 11667 3593
rect 11609 3584 11621 3587
rect 11572 3556 11621 3584
rect 11572 3544 11578 3556
rect 11609 3553 11621 3556
rect 11655 3553 11667 3587
rect 11609 3547 11667 3553
rect 12434 3544 12440 3596
rect 12492 3584 12498 3596
rect 13630 3584 13636 3596
rect 12492 3556 13636 3584
rect 12492 3544 12498 3556
rect 13630 3544 13636 3556
rect 13688 3584 13694 3596
rect 13817 3587 13875 3593
rect 13817 3584 13829 3587
rect 13688 3556 13829 3584
rect 13688 3544 13694 3556
rect 13817 3553 13829 3556
rect 13863 3553 13875 3587
rect 15286 3584 15292 3596
rect 15247 3556 15292 3584
rect 13817 3547 13875 3553
rect 15286 3544 15292 3556
rect 15344 3544 15350 3596
rect 19150 3584 19156 3596
rect 17236 3556 18368 3584
rect 19111 3556 19156 3584
rect 10137 3519 10195 3525
rect 10137 3516 10149 3519
rect 9732 3488 10149 3516
rect 9732 3476 9738 3488
rect 10137 3485 10149 3488
rect 10183 3485 10195 3519
rect 10137 3479 10195 3485
rect 10229 3519 10287 3525
rect 10229 3485 10241 3519
rect 10275 3485 10287 3519
rect 11790 3516 11796 3528
rect 11751 3488 11796 3516
rect 10229 3479 10287 3485
rect 6454 3408 6460 3460
rect 6512 3448 6518 3460
rect 7098 3448 7104 3460
rect 6512 3420 7104 3448
rect 6512 3408 6518 3420
rect 7098 3408 7104 3420
rect 7156 3408 7162 3460
rect 10152 3448 10180 3479
rect 11790 3476 11796 3488
rect 11848 3476 11854 3528
rect 12529 3519 12587 3525
rect 12529 3485 12541 3519
rect 12575 3516 12587 3519
rect 12710 3516 12716 3528
rect 12575 3488 12716 3516
rect 12575 3485 12587 3488
rect 12529 3479 12587 3485
rect 12710 3476 12716 3488
rect 12768 3476 12774 3528
rect 13909 3519 13967 3525
rect 13909 3485 13921 3519
rect 13955 3485 13967 3519
rect 13909 3479 13967 3485
rect 11054 3448 11060 3460
rect 10152 3420 11060 3448
rect 11054 3408 11060 3420
rect 11112 3408 11118 3460
rect 12342 3408 12348 3460
rect 12400 3448 12406 3460
rect 12805 3451 12863 3457
rect 12805 3448 12817 3451
rect 12400 3420 12817 3448
rect 12400 3408 12406 3420
rect 12805 3417 12817 3420
rect 12851 3448 12863 3451
rect 12894 3448 12900 3460
rect 12851 3420 12900 3448
rect 12851 3417 12863 3420
rect 12805 3411 12863 3417
rect 12894 3408 12900 3420
rect 12952 3408 12958 3460
rect 13722 3408 13728 3460
rect 13780 3448 13786 3460
rect 13924 3448 13952 3479
rect 16298 3476 16304 3528
rect 16356 3516 16362 3528
rect 17236 3525 17264 3556
rect 18340 3525 18368 3556
rect 19150 3544 19156 3556
rect 19208 3544 19214 3596
rect 19334 3584 19340 3596
rect 19295 3556 19340 3584
rect 19334 3544 19340 3556
rect 19392 3544 19398 3596
rect 20898 3584 20904 3596
rect 20859 3556 20904 3584
rect 20898 3544 20904 3556
rect 20956 3544 20962 3596
rect 22005 3587 22063 3593
rect 22005 3553 22017 3587
rect 22051 3553 22063 3587
rect 22005 3547 22063 3553
rect 17221 3519 17279 3525
rect 17221 3516 17233 3519
rect 16356 3488 17233 3516
rect 16356 3476 16362 3488
rect 17221 3485 17233 3488
rect 17267 3485 17279 3519
rect 17221 3479 17279 3485
rect 18233 3519 18291 3525
rect 18233 3485 18245 3519
rect 18279 3485 18291 3519
rect 18233 3479 18291 3485
rect 18325 3519 18383 3525
rect 18325 3485 18337 3519
rect 18371 3516 18383 3519
rect 18598 3516 18604 3528
rect 18371 3488 18604 3516
rect 18371 3485 18383 3488
rect 18325 3479 18383 3485
rect 13780 3420 13952 3448
rect 13780 3408 13786 3420
rect 16574 3408 16580 3460
rect 16632 3448 16638 3460
rect 17773 3451 17831 3457
rect 17773 3448 17785 3451
rect 16632 3420 17785 3448
rect 16632 3408 16638 3420
rect 17773 3417 17785 3420
rect 17819 3417 17831 3451
rect 17773 3411 17831 3417
rect 18248 3448 18276 3479
rect 18598 3476 18604 3488
rect 18656 3476 18662 3528
rect 22020 3516 22048 3547
rect 22020 3488 22140 3516
rect 22112 3460 22140 3488
rect 22094 3448 22100 3460
rect 18248 3420 22100 3448
rect 3421 3383 3479 3389
rect 3421 3380 3433 3383
rect 3108 3352 3433 3380
rect 3108 3340 3114 3352
rect 3421 3349 3433 3352
rect 3467 3349 3479 3383
rect 3421 3343 3479 3349
rect 3881 3383 3939 3389
rect 3881 3349 3893 3383
rect 3927 3380 3939 3383
rect 4430 3380 4436 3392
rect 3927 3352 4436 3380
rect 3927 3349 3939 3352
rect 3881 3343 3939 3349
rect 4430 3340 4436 3352
rect 4488 3380 4494 3392
rect 5445 3383 5503 3389
rect 5445 3380 5457 3383
rect 4488 3352 5457 3380
rect 4488 3340 4494 3352
rect 5445 3349 5457 3352
rect 5491 3349 5503 3383
rect 9490 3380 9496 3392
rect 9451 3352 9496 3380
rect 5445 3343 5503 3349
rect 9490 3340 9496 3352
rect 9548 3340 9554 3392
rect 12434 3340 12440 3392
rect 12492 3380 12498 3392
rect 12710 3380 12716 3392
rect 12492 3352 12716 3380
rect 12492 3340 12498 3352
rect 12710 3340 12716 3352
rect 12768 3340 12774 3392
rect 13262 3380 13268 3392
rect 13223 3352 13268 3380
rect 13262 3340 13268 3352
rect 13320 3340 13326 3392
rect 13357 3383 13415 3389
rect 13357 3349 13369 3383
rect 13403 3380 13415 3383
rect 14550 3380 14556 3392
rect 13403 3352 14556 3380
rect 13403 3349 13415 3352
rect 13357 3343 13415 3349
rect 14550 3340 14556 3352
rect 14608 3340 14614 3392
rect 14826 3340 14832 3392
rect 14884 3380 14890 3392
rect 14921 3383 14979 3389
rect 14921 3380 14933 3383
rect 14884 3352 14933 3380
rect 14884 3340 14890 3352
rect 14921 3349 14933 3352
rect 14967 3349 14979 3383
rect 14921 3343 14979 3349
rect 15470 3340 15476 3392
rect 15528 3380 15534 3392
rect 16206 3380 16212 3392
rect 15528 3352 16212 3380
rect 15528 3340 15534 3352
rect 16206 3340 16212 3352
rect 16264 3380 16270 3392
rect 16669 3383 16727 3389
rect 16669 3380 16681 3383
rect 16264 3352 16681 3380
rect 16264 3340 16270 3352
rect 16669 3349 16681 3352
rect 16715 3349 16727 3383
rect 17586 3380 17592 3392
rect 17547 3352 17592 3380
rect 16669 3343 16727 3349
rect 17586 3340 17592 3352
rect 17644 3380 17650 3392
rect 18248 3380 18276 3420
rect 22094 3408 22100 3420
rect 22152 3408 22158 3460
rect 19518 3380 19524 3392
rect 17644 3352 18276 3380
rect 19479 3352 19524 3380
rect 17644 3340 17650 3352
rect 19518 3340 19524 3352
rect 19576 3340 19582 3392
rect 20806 3340 20812 3392
rect 20864 3380 20870 3392
rect 21085 3383 21143 3389
rect 21085 3380 21097 3383
rect 20864 3352 21097 3380
rect 20864 3340 20870 3352
rect 21085 3349 21097 3352
rect 21131 3349 21143 3383
rect 21818 3380 21824 3392
rect 21779 3352 21824 3380
rect 21085 3343 21143 3349
rect 21818 3340 21824 3352
rect 21876 3340 21882 3392
rect 22186 3380 22192 3392
rect 22147 3352 22192 3380
rect 22186 3340 22192 3352
rect 22244 3340 22250 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 2498 3176 2504 3188
rect 2459 3148 2504 3176
rect 2498 3136 2504 3148
rect 2556 3136 2562 3188
rect 3878 3136 3884 3188
rect 3936 3176 3942 3188
rect 5169 3179 5227 3185
rect 5169 3176 5181 3179
rect 3936 3148 5181 3176
rect 3936 3136 3942 3148
rect 5169 3145 5181 3148
rect 5215 3145 5227 3179
rect 5169 3139 5227 3145
rect 6273 3179 6331 3185
rect 6273 3145 6285 3179
rect 6319 3176 6331 3179
rect 6730 3176 6736 3188
rect 6319 3148 6736 3176
rect 6319 3145 6331 3148
rect 6273 3139 6331 3145
rect 6730 3136 6736 3148
rect 6788 3136 6794 3188
rect 8386 3136 8392 3188
rect 8444 3176 8450 3188
rect 9125 3179 9183 3185
rect 9125 3176 9137 3179
rect 8444 3148 9137 3176
rect 8444 3136 8450 3148
rect 9125 3145 9137 3148
rect 9171 3145 9183 3179
rect 9306 3176 9312 3188
rect 9267 3148 9312 3176
rect 9125 3139 9183 3145
rect 9306 3136 9312 3148
rect 9364 3136 9370 3188
rect 9490 3136 9496 3188
rect 9548 3176 9554 3188
rect 10781 3179 10839 3185
rect 10781 3176 10793 3179
rect 9548 3148 10793 3176
rect 9548 3136 9554 3148
rect 10781 3145 10793 3148
rect 10827 3176 10839 3179
rect 11790 3176 11796 3188
rect 10827 3148 11796 3176
rect 10827 3145 10839 3148
rect 10781 3139 10839 3145
rect 11790 3136 11796 3148
rect 11848 3136 11854 3188
rect 15930 3176 15936 3188
rect 15891 3148 15936 3176
rect 15930 3136 15936 3148
rect 15988 3136 15994 3188
rect 16298 3176 16304 3188
rect 16259 3148 16304 3176
rect 16298 3136 16304 3148
rect 16356 3136 16362 3188
rect 18322 3136 18328 3188
rect 18380 3176 18386 3188
rect 19058 3176 19064 3188
rect 18380 3148 19064 3176
rect 18380 3136 18386 3148
rect 19058 3136 19064 3148
rect 19116 3136 19122 3188
rect 19334 3136 19340 3188
rect 19392 3176 19398 3188
rect 19429 3179 19487 3185
rect 19429 3176 19441 3179
rect 19392 3148 19441 3176
rect 19392 3136 19398 3148
rect 19429 3145 19441 3148
rect 19475 3145 19487 3179
rect 20809 3179 20867 3185
rect 20809 3176 20821 3179
rect 19429 3139 19487 3145
rect 19904 3148 20821 3176
rect 1486 3068 1492 3120
rect 1544 3108 1550 3120
rect 1544 3080 1716 3108
rect 1544 3068 1550 3080
rect 1688 3049 1716 3080
rect 4154 3068 4160 3120
rect 4212 3108 4218 3120
rect 4249 3111 4307 3117
rect 4249 3108 4261 3111
rect 4212 3080 4261 3108
rect 4212 3068 4218 3080
rect 4249 3077 4261 3080
rect 4295 3108 4307 3111
rect 4801 3111 4859 3117
rect 4801 3108 4813 3111
rect 4295 3080 4813 3108
rect 4295 3077 4307 3080
rect 4249 3071 4307 3077
rect 4801 3077 4813 3080
rect 4847 3077 4859 3111
rect 5626 3108 5632 3120
rect 5587 3080 5632 3108
rect 4801 3071 4859 3077
rect 5626 3068 5632 3080
rect 5684 3068 5690 3120
rect 6362 3068 6368 3120
rect 6420 3108 6426 3120
rect 6549 3111 6607 3117
rect 6549 3108 6561 3111
rect 6420 3080 6561 3108
rect 6420 3068 6426 3080
rect 6549 3077 6561 3080
rect 6595 3077 6607 3111
rect 6549 3071 6607 3077
rect 1673 3043 1731 3049
rect 1673 3009 1685 3043
rect 1719 3009 1731 3043
rect 1673 3003 1731 3009
rect 5534 3000 5540 3052
rect 5592 3040 5598 3052
rect 5721 3043 5779 3049
rect 5721 3040 5733 3043
rect 5592 3012 5733 3040
rect 5592 3000 5598 3012
rect 5721 3009 5733 3012
rect 5767 3009 5779 3043
rect 6564 3040 6592 3071
rect 11514 3068 11520 3120
rect 11572 3108 11578 3120
rect 11977 3111 12035 3117
rect 11977 3108 11989 3111
rect 11572 3080 11989 3108
rect 11572 3068 11578 3080
rect 11977 3077 11989 3080
rect 12023 3077 12035 3111
rect 11977 3071 12035 3077
rect 14921 3111 14979 3117
rect 14921 3077 14933 3111
rect 14967 3108 14979 3111
rect 14967 3080 16528 3108
rect 14967 3077 14979 3080
rect 14921 3071 14979 3077
rect 9766 3040 9772 3052
rect 6564 3012 6960 3040
rect 9727 3012 9772 3040
rect 5721 3003 5779 3009
rect 1489 2975 1547 2981
rect 1489 2941 1501 2975
rect 1535 2972 1547 2975
rect 2406 2972 2412 2984
rect 1535 2944 2412 2972
rect 1535 2941 1547 2944
rect 1489 2935 1547 2941
rect 2406 2932 2412 2944
rect 2464 2932 2470 2984
rect 2869 2975 2927 2981
rect 2869 2941 2881 2975
rect 2915 2972 2927 2975
rect 4062 2972 4068 2984
rect 2915 2944 4068 2972
rect 2915 2941 2927 2944
rect 2869 2935 2927 2941
rect 4062 2932 4068 2944
rect 4120 2932 4126 2984
rect 6822 2972 6828 2984
rect 6783 2944 6828 2972
rect 6822 2932 6828 2944
rect 6880 2932 6886 2984
rect 6932 2972 6960 3012
rect 9766 3000 9772 3012
rect 9824 3000 9830 3052
rect 9858 3000 9864 3052
rect 9916 3040 9922 3052
rect 9953 3043 10011 3049
rect 9953 3040 9965 3043
rect 9916 3012 9965 3040
rect 9916 3000 9922 3012
rect 9953 3009 9965 3012
rect 9999 3040 10011 3043
rect 10321 3043 10379 3049
rect 10321 3040 10333 3043
rect 9999 3012 10333 3040
rect 9999 3009 10011 3012
rect 9953 3003 10011 3009
rect 10321 3009 10333 3012
rect 10367 3009 10379 3043
rect 11146 3040 11152 3052
rect 11107 3012 11152 3040
rect 10321 3003 10379 3009
rect 11146 3000 11152 3012
rect 11204 3000 11210 3052
rect 14829 3043 14887 3049
rect 14829 3009 14841 3043
rect 14875 3040 14887 3043
rect 15470 3040 15476 3052
rect 14875 3012 15476 3040
rect 14875 3009 14887 3012
rect 14829 3003 14887 3009
rect 15470 3000 15476 3012
rect 15528 3000 15534 3052
rect 7081 2975 7139 2981
rect 7081 2972 7093 2975
rect 6932 2944 7093 2972
rect 7081 2941 7093 2944
rect 7127 2941 7139 2975
rect 7081 2935 7139 2941
rect 9677 2975 9735 2981
rect 9677 2941 9689 2975
rect 9723 2972 9735 2975
rect 10686 2972 10692 2984
rect 9723 2944 10692 2972
rect 9723 2941 9735 2944
rect 9677 2935 9735 2941
rect 10686 2932 10692 2944
rect 10744 2932 10750 2984
rect 10870 2972 10876 2984
rect 10831 2944 10876 2972
rect 10870 2932 10876 2944
rect 10928 2932 10934 2984
rect 12437 2975 12495 2981
rect 12437 2941 12449 2975
rect 12483 2972 12495 2975
rect 13446 2972 13452 2984
rect 12483 2944 13452 2972
rect 12483 2941 12495 2944
rect 12437 2935 12495 2941
rect 13446 2932 13452 2944
rect 13504 2932 13510 2984
rect 13722 2932 13728 2984
rect 13780 2972 13786 2984
rect 14369 2975 14427 2981
rect 14369 2972 14381 2975
rect 13780 2944 14381 2972
rect 13780 2932 13786 2944
rect 14369 2941 14381 2944
rect 14415 2941 14427 2975
rect 14369 2935 14427 2941
rect 14550 2932 14556 2984
rect 14608 2972 14614 2984
rect 16500 2981 16528 3080
rect 16758 3040 16764 3052
rect 16719 3012 16764 3040
rect 16758 3000 16764 3012
rect 16816 3000 16822 3052
rect 18598 3040 18604 3052
rect 18559 3012 18604 3040
rect 18598 3000 18604 3012
rect 18656 3000 18662 3052
rect 19904 3049 19932 3148
rect 20809 3145 20821 3148
rect 20855 3176 20867 3179
rect 20898 3176 20904 3188
rect 20855 3148 20904 3176
rect 20855 3145 20867 3148
rect 20809 3139 20867 3145
rect 20898 3136 20904 3148
rect 20956 3136 20962 3188
rect 21726 3136 21732 3188
rect 21784 3176 21790 3188
rect 21821 3179 21879 3185
rect 21821 3176 21833 3179
rect 21784 3148 21833 3176
rect 21784 3136 21790 3148
rect 21821 3145 21833 3148
rect 21867 3145 21879 3179
rect 21821 3139 21879 3145
rect 22094 3136 22100 3188
rect 22152 3176 22158 3188
rect 22557 3179 22615 3185
rect 22557 3176 22569 3179
rect 22152 3148 22569 3176
rect 22152 3136 22158 3148
rect 22557 3145 22569 3148
rect 22603 3145 22615 3179
rect 22557 3139 22615 3145
rect 21358 3068 21364 3120
rect 21416 3108 21422 3120
rect 22189 3111 22247 3117
rect 22189 3108 22201 3111
rect 21416 3080 22201 3108
rect 21416 3068 21422 3080
rect 22189 3077 22201 3080
rect 22235 3077 22247 3111
rect 22189 3071 22247 3077
rect 19889 3043 19947 3049
rect 19889 3009 19901 3043
rect 19935 3009 19947 3043
rect 19889 3003 19947 3009
rect 15289 2975 15347 2981
rect 15289 2972 15301 2975
rect 14608 2944 15301 2972
rect 14608 2932 14614 2944
rect 15289 2941 15301 2944
rect 15335 2941 15347 2975
rect 15289 2935 15347 2941
rect 16485 2975 16543 2981
rect 16485 2941 16497 2975
rect 16531 2941 16543 2975
rect 16485 2935 16543 2941
rect 17497 2975 17555 2981
rect 17497 2941 17509 2975
rect 17543 2972 17555 2975
rect 18509 2975 18567 2981
rect 18509 2972 18521 2975
rect 17543 2944 18521 2972
rect 17543 2941 17555 2944
rect 17497 2935 17555 2941
rect 18509 2941 18521 2944
rect 18555 2972 18567 2975
rect 19242 2972 19248 2984
rect 18555 2944 19248 2972
rect 18555 2941 18567 2944
rect 18509 2935 18567 2941
rect 3050 2864 3056 2916
rect 3108 2913 3114 2916
rect 3108 2907 3172 2913
rect 3108 2873 3126 2907
rect 3160 2873 3172 2907
rect 3108 2867 3172 2873
rect 11624 2876 12112 2904
rect 3108 2864 3114 2867
rect 11624 2848 11652 2876
rect 8202 2836 8208 2848
rect 8163 2808 8208 2836
rect 8202 2796 8208 2808
rect 8260 2796 8266 2848
rect 8754 2836 8760 2848
rect 8715 2808 8760 2836
rect 8754 2796 8760 2808
rect 8812 2796 8818 2848
rect 11606 2836 11612 2848
rect 11567 2808 11612 2836
rect 11606 2796 11612 2808
rect 11664 2796 11670 2848
rect 12084 2836 12112 2876
rect 12342 2864 12348 2916
rect 12400 2904 12406 2916
rect 12682 2907 12740 2913
rect 12682 2904 12694 2907
rect 12400 2876 12694 2904
rect 12400 2864 12406 2876
rect 12682 2873 12694 2876
rect 12728 2873 12740 2907
rect 12682 2867 12740 2873
rect 13170 2864 13176 2916
rect 13228 2904 13234 2916
rect 14826 2904 14832 2916
rect 13228 2876 14832 2904
rect 13228 2864 13234 2876
rect 14826 2864 14832 2876
rect 14884 2904 14890 2916
rect 15381 2907 15439 2913
rect 15381 2904 15393 2907
rect 14884 2876 15393 2904
rect 14884 2864 14890 2876
rect 15381 2873 15393 2876
rect 15427 2873 15439 2907
rect 15381 2867 15439 2873
rect 12434 2836 12440 2848
rect 12084 2808 12440 2836
rect 12434 2796 12440 2808
rect 12492 2796 12498 2848
rect 13262 2796 13268 2848
rect 13320 2836 13326 2848
rect 13817 2839 13875 2845
rect 13817 2836 13829 2839
rect 13320 2808 13829 2836
rect 13320 2796 13326 2808
rect 13817 2805 13829 2808
rect 13863 2836 13875 2839
rect 15102 2836 15108 2848
rect 13863 2808 15108 2836
rect 13863 2805 13875 2808
rect 13817 2799 13875 2805
rect 15102 2796 15108 2808
rect 15160 2796 15166 2848
rect 16500 2836 16528 2935
rect 19242 2932 19248 2944
rect 19300 2932 19306 2984
rect 19334 2932 19340 2984
rect 19392 2972 19398 2984
rect 19613 2975 19671 2981
rect 19613 2972 19625 2975
rect 19392 2944 19625 2972
rect 19392 2932 19398 2944
rect 19613 2941 19625 2944
rect 19659 2972 19671 2975
rect 20349 2975 20407 2981
rect 20349 2972 20361 2975
rect 19659 2944 20361 2972
rect 19659 2941 19671 2944
rect 19613 2935 19671 2941
rect 20349 2941 20361 2944
rect 20395 2941 20407 2975
rect 20349 2935 20407 2941
rect 20714 2932 20720 2984
rect 20772 2972 20778 2984
rect 20901 2975 20959 2981
rect 20901 2972 20913 2975
rect 20772 2944 20913 2972
rect 20772 2932 20778 2944
rect 20901 2941 20913 2944
rect 20947 2972 20959 2975
rect 21453 2975 21511 2981
rect 21453 2972 21465 2975
rect 20947 2944 21465 2972
rect 20947 2941 20959 2944
rect 20901 2935 20959 2941
rect 21453 2941 21465 2944
rect 21499 2941 21511 2975
rect 21453 2935 21511 2941
rect 21726 2932 21732 2984
rect 21784 2972 21790 2984
rect 22005 2975 22063 2981
rect 22005 2972 22017 2975
rect 21784 2944 22017 2972
rect 21784 2932 21790 2944
rect 22005 2941 22017 2944
rect 22051 2941 22063 2975
rect 22005 2935 22063 2941
rect 17862 2904 17868 2916
rect 17775 2876 17868 2904
rect 17862 2864 17868 2876
rect 17920 2904 17926 2916
rect 18417 2907 18475 2913
rect 18417 2904 18429 2907
rect 17920 2876 18429 2904
rect 17920 2864 17926 2876
rect 18417 2873 18429 2876
rect 18463 2873 18475 2907
rect 22462 2904 22468 2916
rect 18417 2867 18475 2873
rect 21100 2876 22468 2904
rect 16574 2836 16580 2848
rect 16500 2808 16580 2836
rect 16574 2796 16580 2808
rect 16632 2796 16638 2848
rect 18046 2836 18052 2848
rect 18007 2808 18052 2836
rect 18046 2796 18052 2808
rect 18104 2796 18110 2848
rect 21100 2845 21128 2876
rect 22462 2864 22468 2876
rect 22520 2864 22526 2916
rect 21085 2839 21143 2845
rect 21085 2805 21097 2839
rect 21131 2805 21143 2839
rect 21085 2799 21143 2805
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 1670 2592 1676 2644
rect 1728 2632 1734 2644
rect 2409 2635 2467 2641
rect 2409 2632 2421 2635
rect 1728 2604 2421 2632
rect 1728 2592 1734 2604
rect 2409 2601 2421 2604
rect 2455 2601 2467 2635
rect 2866 2632 2872 2644
rect 2827 2604 2872 2632
rect 2409 2595 2467 2601
rect 2866 2592 2872 2604
rect 2924 2592 2930 2644
rect 2958 2592 2964 2644
rect 3016 2632 3022 2644
rect 3789 2635 3847 2641
rect 3789 2632 3801 2635
rect 3016 2604 3801 2632
rect 3016 2592 3022 2604
rect 3789 2601 3801 2604
rect 3835 2601 3847 2635
rect 3789 2595 3847 2601
rect 3970 2592 3976 2644
rect 4028 2632 4034 2644
rect 4065 2635 4123 2641
rect 4065 2632 4077 2635
rect 4028 2604 4077 2632
rect 4028 2592 4034 2604
rect 4065 2601 4077 2604
rect 4111 2601 4123 2635
rect 4706 2632 4712 2644
rect 4667 2604 4712 2632
rect 4065 2595 4123 2601
rect 4706 2592 4712 2604
rect 4764 2632 4770 2644
rect 5629 2635 5687 2641
rect 5629 2632 5641 2635
rect 4764 2604 5641 2632
rect 4764 2592 4770 2604
rect 5629 2601 5641 2604
rect 5675 2601 5687 2635
rect 5629 2595 5687 2601
rect 6638 2592 6644 2644
rect 6696 2632 6702 2644
rect 6733 2635 6791 2641
rect 6733 2632 6745 2635
rect 6696 2604 6745 2632
rect 6696 2592 6702 2604
rect 6733 2601 6745 2604
rect 6779 2632 6791 2635
rect 8202 2632 8208 2644
rect 6779 2604 8208 2632
rect 6779 2601 6791 2604
rect 6733 2595 6791 2601
rect 1949 2567 2007 2573
rect 1949 2533 1961 2567
rect 1995 2564 2007 2567
rect 2884 2564 2912 2592
rect 7484 2573 7512 2604
rect 8202 2592 8208 2604
rect 8260 2592 8266 2644
rect 9950 2592 9956 2644
rect 10008 2632 10014 2644
rect 10962 2632 10968 2644
rect 10008 2604 10968 2632
rect 10008 2592 10014 2604
rect 10962 2592 10968 2604
rect 11020 2592 11026 2644
rect 11054 2592 11060 2644
rect 11112 2632 11118 2644
rect 11793 2635 11851 2641
rect 11793 2632 11805 2635
rect 11112 2604 11805 2632
rect 11112 2592 11118 2604
rect 11793 2601 11805 2604
rect 11839 2601 11851 2635
rect 13170 2632 13176 2644
rect 13131 2604 13176 2632
rect 11793 2595 11851 2601
rect 13170 2592 13176 2604
rect 13228 2592 13234 2644
rect 13814 2592 13820 2644
rect 13872 2632 13878 2644
rect 14185 2635 14243 2641
rect 14185 2632 14197 2635
rect 13872 2604 14197 2632
rect 13872 2592 13878 2604
rect 14185 2601 14197 2604
rect 14231 2601 14243 2635
rect 15194 2632 15200 2644
rect 15155 2604 15200 2632
rect 14185 2595 14243 2601
rect 15194 2592 15200 2604
rect 15252 2632 15258 2644
rect 16574 2632 16580 2644
rect 15252 2604 16068 2632
rect 16535 2604 16580 2632
rect 15252 2592 15258 2604
rect 1995 2536 2912 2564
rect 7460 2567 7518 2573
rect 1995 2533 2007 2536
rect 1949 2527 2007 2533
rect 7460 2533 7472 2567
rect 7506 2533 7518 2567
rect 7460 2527 7518 2533
rect 11238 2524 11244 2576
rect 11296 2564 11302 2576
rect 12161 2567 12219 2573
rect 12161 2564 12173 2567
rect 11296 2536 12173 2564
rect 11296 2524 11302 2536
rect 12161 2533 12173 2536
rect 12207 2533 12219 2567
rect 12161 2527 12219 2533
rect 2317 2499 2375 2505
rect 2317 2465 2329 2499
rect 2363 2496 2375 2499
rect 2777 2499 2835 2505
rect 2777 2496 2789 2499
rect 2363 2468 2789 2496
rect 2363 2465 2375 2468
rect 2317 2459 2375 2465
rect 2777 2465 2789 2468
rect 2823 2496 2835 2499
rect 3602 2496 3608 2508
rect 2823 2468 3608 2496
rect 2823 2465 2835 2468
rect 2777 2459 2835 2465
rect 3602 2456 3608 2468
rect 3660 2456 3666 2508
rect 5166 2496 5172 2508
rect 5079 2468 5172 2496
rect 5166 2456 5172 2468
rect 5224 2496 5230 2508
rect 5721 2499 5779 2505
rect 5721 2496 5733 2499
rect 5224 2468 5733 2496
rect 5224 2456 5230 2468
rect 5721 2465 5733 2468
rect 5767 2496 5779 2499
rect 6086 2496 6092 2508
rect 5767 2468 6092 2496
rect 5767 2465 5779 2468
rect 5721 2459 5779 2465
rect 6086 2456 6092 2468
rect 6144 2456 6150 2508
rect 6822 2456 6828 2508
rect 6880 2496 6886 2508
rect 7193 2499 7251 2505
rect 7193 2496 7205 2499
rect 6880 2468 7205 2496
rect 6880 2456 6886 2468
rect 7193 2465 7205 2468
rect 7239 2496 7251 2499
rect 8570 2496 8576 2508
rect 7239 2468 8576 2496
rect 7239 2465 7251 2468
rect 7193 2459 7251 2465
rect 8570 2456 8576 2468
rect 8628 2496 8634 2508
rect 9861 2499 9919 2505
rect 9861 2496 9873 2499
rect 8628 2468 9873 2496
rect 8628 2456 8634 2468
rect 9861 2465 9873 2468
rect 9907 2465 9919 2499
rect 10117 2499 10175 2505
rect 10117 2496 10129 2499
rect 9861 2459 9919 2465
rect 9968 2468 10129 2496
rect 3050 2428 3056 2440
rect 3011 2400 3056 2428
rect 3050 2388 3056 2400
rect 3108 2428 3114 2440
rect 3421 2431 3479 2437
rect 3421 2428 3433 2431
rect 3108 2400 3433 2428
rect 3108 2388 3114 2400
rect 3421 2397 3433 2400
rect 3467 2397 3479 2431
rect 3421 2391 3479 2397
rect 5905 2431 5963 2437
rect 5905 2397 5917 2431
rect 5951 2428 5963 2431
rect 6362 2428 6368 2440
rect 5951 2400 6368 2428
rect 5951 2397 5963 2400
rect 5905 2391 5963 2397
rect 6362 2388 6368 2400
rect 6420 2388 6426 2440
rect 9968 2428 9996 2468
rect 10117 2465 10129 2468
rect 10163 2465 10175 2499
rect 10117 2459 10175 2465
rect 12066 2456 12072 2508
rect 12124 2496 12130 2508
rect 13538 2496 13544 2508
rect 12124 2468 13544 2496
rect 12124 2456 12130 2468
rect 13538 2456 13544 2468
rect 13596 2456 13602 2508
rect 13633 2499 13691 2505
rect 13633 2465 13645 2499
rect 13679 2496 13691 2499
rect 15838 2496 15844 2508
rect 13679 2468 14688 2496
rect 15799 2468 15844 2496
rect 13679 2465 13691 2468
rect 13633 2459 13691 2465
rect 9324 2400 9996 2428
rect 5258 2360 5264 2372
rect 5219 2332 5264 2360
rect 5258 2320 5264 2332
rect 5316 2320 5322 2372
rect 9324 2369 9352 2400
rect 9876 2372 9904 2400
rect 13722 2388 13728 2440
rect 13780 2428 13786 2440
rect 13780 2400 13825 2428
rect 13780 2388 13786 2400
rect 8573 2363 8631 2369
rect 8573 2329 8585 2363
rect 8619 2360 8631 2363
rect 9309 2363 9367 2369
rect 9309 2360 9321 2363
rect 8619 2332 9321 2360
rect 8619 2329 8631 2332
rect 8573 2323 8631 2329
rect 9309 2329 9321 2332
rect 9355 2329 9367 2363
rect 9309 2323 9367 2329
rect 9858 2320 9864 2372
rect 9916 2320 9922 2372
rect 11238 2360 11244 2372
rect 11151 2332 11244 2360
rect 11238 2320 11244 2332
rect 11296 2360 11302 2372
rect 12342 2360 12348 2372
rect 11296 2332 12348 2360
rect 11296 2320 11302 2332
rect 12342 2320 12348 2332
rect 12400 2320 12406 2372
rect 13081 2363 13139 2369
rect 13081 2329 13093 2363
rect 13127 2360 13139 2363
rect 13740 2360 13768 2388
rect 14660 2372 14688 2468
rect 15838 2456 15844 2468
rect 15896 2456 15902 2508
rect 16040 2437 16068 2604
rect 16574 2592 16580 2604
rect 16632 2592 16638 2644
rect 18138 2632 18144 2644
rect 18099 2604 18144 2632
rect 18138 2592 18144 2604
rect 18196 2632 18202 2644
rect 18785 2635 18843 2641
rect 18785 2632 18797 2635
rect 18196 2604 18797 2632
rect 18196 2592 18202 2604
rect 18785 2601 18797 2604
rect 18831 2601 18843 2635
rect 18785 2595 18843 2601
rect 21361 2635 21419 2641
rect 21361 2601 21373 2635
rect 21407 2632 21419 2635
rect 22002 2632 22008 2644
rect 21407 2604 22008 2632
rect 21407 2601 21419 2604
rect 21361 2595 21419 2601
rect 22002 2592 22008 2604
rect 22060 2592 22066 2644
rect 22094 2592 22100 2644
rect 22152 2632 22158 2644
rect 22152 2604 22197 2632
rect 22152 2592 22158 2604
rect 16114 2524 16120 2576
rect 16172 2564 16178 2576
rect 16945 2567 17003 2573
rect 16945 2564 16957 2567
rect 16172 2536 16957 2564
rect 16172 2524 16178 2536
rect 16945 2533 16957 2536
rect 16991 2533 17003 2567
rect 16945 2527 17003 2533
rect 16960 2496 16988 2527
rect 18046 2524 18052 2576
rect 18104 2564 18110 2576
rect 19705 2567 19763 2573
rect 19705 2564 19717 2567
rect 18104 2536 19717 2564
rect 18104 2524 18110 2536
rect 19705 2533 19717 2536
rect 19751 2533 19763 2567
rect 19705 2527 19763 2533
rect 17129 2499 17187 2505
rect 17129 2496 17141 2499
rect 16960 2468 17141 2496
rect 17129 2465 17141 2468
rect 17175 2465 17187 2499
rect 17129 2459 17187 2465
rect 18693 2499 18751 2505
rect 18693 2465 18705 2499
rect 18739 2465 18751 2499
rect 19886 2496 19892 2508
rect 19847 2468 19892 2496
rect 18693 2459 18751 2465
rect 14921 2431 14979 2437
rect 14921 2397 14933 2431
rect 14967 2428 14979 2431
rect 15933 2431 15991 2437
rect 15933 2428 15945 2431
rect 14967 2400 15945 2428
rect 14967 2397 14979 2400
rect 14921 2391 14979 2397
rect 15933 2397 15945 2400
rect 15979 2397 15991 2431
rect 15933 2391 15991 2397
rect 16025 2431 16083 2437
rect 16025 2397 16037 2431
rect 16071 2397 16083 2431
rect 16025 2391 16083 2397
rect 13127 2332 13768 2360
rect 13127 2329 13139 2332
rect 13081 2323 13139 2329
rect 14642 2320 14648 2372
rect 14700 2360 14706 2372
rect 15473 2363 15531 2369
rect 15473 2360 15485 2363
rect 14700 2332 15485 2360
rect 14700 2320 14706 2332
rect 15473 2329 15485 2332
rect 15519 2329 15531 2363
rect 15948 2360 15976 2391
rect 17034 2388 17040 2440
rect 17092 2428 17098 2440
rect 17681 2431 17739 2437
rect 17681 2428 17693 2431
rect 17092 2400 17693 2428
rect 17092 2388 17098 2400
rect 17681 2397 17693 2400
rect 17727 2428 17739 2431
rect 18708 2428 18736 2459
rect 19886 2456 19892 2468
rect 19944 2496 19950 2508
rect 20441 2499 20499 2505
rect 20441 2496 20453 2499
rect 19944 2468 20453 2496
rect 19944 2456 19950 2468
rect 20441 2465 20453 2468
rect 20487 2465 20499 2499
rect 21174 2496 21180 2508
rect 21135 2468 21180 2496
rect 20441 2459 20499 2465
rect 21174 2456 21180 2468
rect 21232 2496 21238 2508
rect 21729 2499 21787 2505
rect 21729 2496 21741 2499
rect 21232 2468 21741 2496
rect 21232 2456 21238 2468
rect 21729 2465 21741 2468
rect 21775 2465 21787 2499
rect 22278 2496 22284 2508
rect 22239 2468 22284 2496
rect 21729 2459 21787 2465
rect 22278 2456 22284 2468
rect 22336 2496 22342 2508
rect 22833 2499 22891 2505
rect 22833 2496 22845 2499
rect 22336 2468 22845 2496
rect 22336 2456 22342 2468
rect 22833 2465 22845 2468
rect 22879 2465 22891 2499
rect 24026 2496 24032 2508
rect 23987 2468 24032 2496
rect 22833 2459 22891 2465
rect 24026 2456 24032 2468
rect 24084 2496 24090 2508
rect 24581 2499 24639 2505
rect 24581 2496 24593 2499
rect 24084 2468 24593 2496
rect 24084 2456 24090 2468
rect 24581 2465 24593 2468
rect 24627 2465 24639 2499
rect 24581 2459 24639 2465
rect 17727 2400 18736 2428
rect 18877 2431 18935 2437
rect 17727 2397 17739 2400
rect 17681 2391 17739 2397
rect 18877 2397 18889 2431
rect 18923 2428 18935 2431
rect 19337 2431 19395 2437
rect 19337 2428 19349 2431
rect 18923 2400 19349 2428
rect 18923 2397 18935 2400
rect 18877 2391 18935 2397
rect 19337 2397 19349 2400
rect 19383 2397 19395 2431
rect 19337 2391 19395 2397
rect 16482 2360 16488 2372
rect 15948 2332 16488 2360
rect 15473 2323 15531 2329
rect 16482 2320 16488 2332
rect 16540 2320 16546 2372
rect 17310 2360 17316 2372
rect 17271 2332 17316 2360
rect 17310 2320 17316 2332
rect 17368 2320 17374 2372
rect 18598 2320 18604 2372
rect 18656 2360 18662 2372
rect 18892 2360 18920 2391
rect 18656 2332 18920 2360
rect 20073 2363 20131 2369
rect 18656 2320 18662 2332
rect 20073 2329 20085 2363
rect 20119 2360 20131 2363
rect 21910 2360 21916 2372
rect 20119 2332 21916 2360
rect 20119 2329 20131 2332
rect 20073 2323 20131 2329
rect 21910 2320 21916 2332
rect 21968 2320 21974 2372
rect 22465 2363 22523 2369
rect 22465 2329 22477 2363
rect 22511 2360 22523 2363
rect 23658 2360 23664 2372
rect 22511 2332 23664 2360
rect 22511 2329 22523 2332
rect 22465 2323 22523 2329
rect 23658 2320 23664 2332
rect 23716 2320 23722 2372
rect 18322 2292 18328 2304
rect 18283 2264 18328 2292
rect 18322 2252 18328 2264
rect 18380 2252 18386 2304
rect 20714 2252 20720 2304
rect 20772 2292 20778 2304
rect 20809 2295 20867 2301
rect 20809 2292 20821 2295
rect 20772 2264 20821 2292
rect 20772 2252 20778 2264
rect 20809 2261 20821 2264
rect 20855 2261 20867 2295
rect 20809 2255 20867 2261
rect 23474 2252 23480 2304
rect 23532 2292 23538 2304
rect 24213 2295 24271 2301
rect 24213 2292 24225 2295
rect 23532 2264 24225 2292
rect 23532 2252 23538 2264
rect 24213 2261 24225 2264
rect 24259 2261 24271 2295
rect 24213 2255 24271 2261
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 5994 552 6000 604
rect 6052 592 6058 604
rect 6178 592 6184 604
rect 6052 564 6184 592
rect 6052 552 6058 564
rect 6178 552 6184 564
rect 6236 552 6242 604
<< via1 >>
rect 5264 27412 5316 27464
rect 5356 27412 5408 27464
rect 8944 27412 8996 27464
rect 9404 27412 9456 27464
rect 3516 27208 3568 27260
rect 7012 27208 7064 27260
rect 4068 26528 4120 26580
rect 8116 26528 8168 26580
rect 3516 26256 3568 26308
rect 7196 26256 7248 26308
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 3056 25440 3108 25492
rect 4068 25440 4120 25492
rect 7196 25440 7248 25492
rect 2044 25372 2096 25424
rect 9496 25372 9548 25424
rect 1584 25304 1636 25356
rect 2596 25304 2648 25356
rect 4436 25304 4488 25356
rect 6920 25347 6972 25356
rect 2872 25236 2924 25288
rect 6920 25313 6929 25347
rect 6929 25313 6963 25347
rect 6963 25313 6972 25347
rect 6920 25304 6972 25313
rect 7748 25304 7800 25356
rect 15660 25304 15712 25356
rect 12624 25236 12676 25288
rect 4068 25168 4120 25220
rect 7012 25168 7064 25220
rect 2136 25100 2188 25152
rect 3516 25100 3568 25152
rect 26516 25100 26568 25152
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 3332 24896 3384 24948
rect 8116 24939 8168 24948
rect 8116 24905 8125 24939
rect 8125 24905 8159 24939
rect 8159 24905 8168 24939
rect 8116 24896 8168 24905
rect 6920 24828 6972 24880
rect 2136 24760 2188 24812
rect 6276 24760 6328 24812
rect 1584 24692 1636 24744
rect 2688 24692 2740 24744
rect 2964 24692 3016 24744
rect 12624 24803 12676 24812
rect 12624 24769 12633 24803
rect 12633 24769 12667 24803
rect 12667 24769 12676 24803
rect 12624 24760 12676 24769
rect 1768 24667 1820 24676
rect 1768 24633 1777 24667
rect 1777 24633 1811 24667
rect 1811 24633 1820 24667
rect 1768 24624 1820 24633
rect 2504 24624 2556 24676
rect 7840 24692 7892 24744
rect 9496 24735 9548 24744
rect 9496 24701 9505 24735
rect 9505 24701 9539 24735
rect 9539 24701 9548 24735
rect 9496 24692 9548 24701
rect 9956 24692 10008 24744
rect 2596 24599 2648 24608
rect 2596 24565 2605 24599
rect 2605 24565 2639 24599
rect 2639 24565 2648 24599
rect 2596 24556 2648 24565
rect 3240 24556 3292 24608
rect 4068 24599 4120 24608
rect 4068 24565 4077 24599
rect 4077 24565 4111 24599
rect 4111 24565 4120 24599
rect 4068 24556 4120 24565
rect 4436 24599 4488 24608
rect 4436 24565 4445 24599
rect 4445 24565 4479 24599
rect 4479 24565 4488 24599
rect 4436 24556 4488 24565
rect 5172 24599 5224 24608
rect 5172 24565 5181 24599
rect 5181 24565 5215 24599
rect 5215 24565 5224 24599
rect 5172 24556 5224 24565
rect 5540 24599 5592 24608
rect 5540 24565 5549 24599
rect 5549 24565 5583 24599
rect 5583 24565 5592 24599
rect 5540 24556 5592 24565
rect 6276 24599 6328 24608
rect 6276 24565 6285 24599
rect 6285 24565 6319 24599
rect 6319 24565 6328 24599
rect 6276 24556 6328 24565
rect 16120 24692 16172 24744
rect 18144 24692 18196 24744
rect 15384 24624 15436 24676
rect 6828 24556 6880 24608
rect 8852 24599 8904 24608
rect 8852 24565 8861 24599
rect 8861 24565 8895 24599
rect 8895 24565 8904 24599
rect 8852 24556 8904 24565
rect 13084 24556 13136 24608
rect 13636 24599 13688 24608
rect 13636 24565 13645 24599
rect 13645 24565 13679 24599
rect 13679 24565 13688 24599
rect 13636 24556 13688 24565
rect 16488 24624 16540 24676
rect 15660 24599 15712 24608
rect 15660 24565 15669 24599
rect 15669 24565 15703 24599
rect 15703 24565 15712 24599
rect 15660 24556 15712 24565
rect 16396 24599 16448 24608
rect 16396 24565 16405 24599
rect 16405 24565 16439 24599
rect 16439 24565 16448 24599
rect 16396 24556 16448 24565
rect 18236 24599 18288 24608
rect 18236 24565 18245 24599
rect 18245 24565 18279 24599
rect 18279 24565 18288 24599
rect 18236 24556 18288 24565
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 2872 24352 2924 24404
rect 3148 24352 3200 24404
rect 4896 24352 4948 24404
rect 9312 24352 9364 24404
rect 12072 24352 12124 24404
rect 13084 24395 13136 24404
rect 13084 24361 13093 24395
rect 13093 24361 13127 24395
rect 13127 24361 13136 24395
rect 13084 24352 13136 24361
rect 16212 24352 16264 24404
rect 18512 24352 18564 24404
rect 18788 24395 18840 24404
rect 18788 24361 18797 24395
rect 18797 24361 18831 24395
rect 18831 24361 18840 24395
rect 18788 24352 18840 24361
rect 23112 24352 23164 24404
rect 23296 24395 23348 24404
rect 23296 24361 23305 24395
rect 23305 24361 23339 24395
rect 23339 24361 23348 24395
rect 23296 24352 23348 24361
rect 1952 24327 2004 24336
rect 1952 24293 1961 24327
rect 1961 24293 1995 24327
rect 1995 24293 2004 24327
rect 1952 24284 2004 24293
rect 1676 24259 1728 24268
rect 1676 24225 1685 24259
rect 1685 24225 1719 24259
rect 1719 24225 1728 24259
rect 1676 24216 1728 24225
rect 2228 24216 2280 24268
rect 6276 24216 6328 24268
rect 9036 24216 9088 24268
rect 10324 24259 10376 24268
rect 10324 24225 10333 24259
rect 10333 24225 10367 24259
rect 10367 24225 10376 24259
rect 10324 24216 10376 24225
rect 12256 24216 12308 24268
rect 13360 24216 13412 24268
rect 15292 24259 15344 24268
rect 15292 24225 15301 24259
rect 15301 24225 15335 24259
rect 15335 24225 15344 24259
rect 15292 24216 15344 24225
rect 16396 24259 16448 24268
rect 16396 24225 16405 24259
rect 16405 24225 16439 24259
rect 16439 24225 16448 24259
rect 16396 24216 16448 24225
rect 17500 24259 17552 24268
rect 17500 24225 17509 24259
rect 17509 24225 17543 24259
rect 17543 24225 17552 24259
rect 17500 24216 17552 24225
rect 18512 24216 18564 24268
rect 20812 24216 20864 24268
rect 22008 24259 22060 24268
rect 22008 24225 22017 24259
rect 22017 24225 22051 24259
rect 22051 24225 22060 24259
rect 22008 24216 22060 24225
rect 23296 24216 23348 24268
rect 3332 24148 3384 24200
rect 8668 24191 8720 24200
rect 8668 24157 8677 24191
rect 8677 24157 8711 24191
rect 8711 24157 8720 24191
rect 8668 24148 8720 24157
rect 10140 24148 10192 24200
rect 12348 24148 12400 24200
rect 13544 24191 13596 24200
rect 13544 24157 13553 24191
rect 13553 24157 13587 24191
rect 13587 24157 13596 24191
rect 13544 24148 13596 24157
rect 13728 24191 13780 24200
rect 13728 24157 13737 24191
rect 13737 24157 13771 24191
rect 13771 24157 13780 24191
rect 13728 24148 13780 24157
rect 9956 24123 10008 24132
rect 9956 24089 9965 24123
rect 9965 24089 9999 24123
rect 9999 24089 10008 24123
rect 9956 24080 10008 24089
rect 12992 24123 13044 24132
rect 12992 24089 13001 24123
rect 13001 24089 13035 24123
rect 13035 24089 13044 24123
rect 12992 24080 13044 24089
rect 17868 24080 17920 24132
rect 22468 24080 22520 24132
rect 3976 24012 4028 24064
rect 6644 24055 6696 24064
rect 6644 24021 6653 24055
rect 6653 24021 6687 24055
rect 6687 24021 6696 24055
rect 6644 24012 6696 24021
rect 7012 24012 7064 24064
rect 8116 24012 8168 24064
rect 13820 24012 13872 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 1768 23715 1820 23724
rect 1768 23681 1777 23715
rect 1777 23681 1811 23715
rect 1811 23681 1820 23715
rect 1768 23672 1820 23681
rect 2412 23808 2464 23860
rect 3332 23808 3384 23860
rect 6276 23808 6328 23860
rect 9036 23851 9088 23860
rect 9036 23817 9045 23851
rect 9045 23817 9079 23851
rect 9079 23817 9088 23851
rect 9036 23808 9088 23817
rect 9312 23851 9364 23860
rect 9312 23817 9321 23851
rect 9321 23817 9355 23851
rect 9355 23817 9364 23851
rect 9312 23808 9364 23817
rect 11244 23851 11296 23860
rect 11244 23817 11253 23851
rect 11253 23817 11287 23851
rect 11287 23817 11296 23851
rect 11244 23808 11296 23817
rect 12072 23808 12124 23860
rect 13728 23808 13780 23860
rect 16396 23808 16448 23860
rect 19064 23808 19116 23860
rect 19524 23808 19576 23860
rect 21364 23808 21416 23860
rect 21916 23808 21968 23860
rect 23664 23808 23716 23860
rect 25320 23808 25372 23860
rect 12624 23783 12676 23792
rect 12624 23749 12633 23783
rect 12633 23749 12667 23783
rect 12667 23749 12676 23783
rect 12624 23740 12676 23749
rect 7012 23715 7064 23724
rect 7012 23681 7021 23715
rect 7021 23681 7055 23715
rect 7055 23681 7064 23715
rect 7012 23672 7064 23681
rect 15384 23672 15436 23724
rect 9956 23604 10008 23656
rect 12072 23604 12124 23656
rect 13636 23604 13688 23656
rect 18052 23647 18104 23656
rect 7564 23536 7616 23588
rect 10140 23579 10192 23588
rect 10140 23545 10174 23579
rect 10174 23545 10192 23579
rect 10140 23536 10192 23545
rect 10324 23536 10376 23588
rect 13912 23536 13964 23588
rect 2688 23511 2740 23520
rect 2688 23477 2697 23511
rect 2697 23477 2731 23511
rect 2731 23477 2740 23511
rect 2688 23468 2740 23477
rect 4068 23468 4120 23520
rect 4344 23468 4396 23520
rect 5816 23511 5868 23520
rect 5816 23477 5825 23511
rect 5825 23477 5859 23511
rect 5859 23477 5868 23511
rect 5816 23468 5868 23477
rect 6092 23468 6144 23520
rect 10968 23468 11020 23520
rect 12256 23511 12308 23520
rect 12256 23477 12265 23511
rect 12265 23477 12299 23511
rect 12299 23477 12308 23511
rect 12256 23468 12308 23477
rect 13360 23511 13412 23520
rect 13360 23477 13369 23511
rect 13369 23477 13403 23511
rect 13403 23477 13412 23511
rect 13360 23468 13412 23477
rect 13452 23468 13504 23520
rect 18052 23613 18061 23647
rect 18061 23613 18095 23647
rect 18095 23613 18104 23647
rect 18052 23604 18104 23613
rect 18420 23604 18472 23656
rect 18512 23536 18564 23588
rect 21364 23647 21416 23656
rect 21364 23613 21373 23647
rect 21373 23613 21407 23647
rect 21407 23613 21416 23647
rect 21364 23604 21416 23613
rect 22376 23604 22428 23656
rect 23480 23604 23532 23656
rect 15200 23468 15252 23520
rect 17132 23468 17184 23520
rect 17500 23511 17552 23520
rect 17500 23477 17509 23511
rect 17509 23477 17543 23511
rect 17543 23477 17552 23511
rect 17500 23468 17552 23477
rect 20076 23511 20128 23520
rect 20076 23477 20085 23511
rect 20085 23477 20119 23511
rect 20119 23477 20128 23511
rect 20076 23468 20128 23477
rect 20812 23468 20864 23520
rect 21180 23468 21232 23520
rect 22008 23468 22060 23520
rect 23296 23468 23348 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 1676 23264 1728 23316
rect 7012 23307 7064 23316
rect 7012 23273 7021 23307
rect 7021 23273 7055 23307
rect 7055 23273 7064 23307
rect 7012 23264 7064 23273
rect 7564 23264 7616 23316
rect 10140 23264 10192 23316
rect 2412 23128 2464 23180
rect 4344 23171 4396 23180
rect 2872 23103 2924 23112
rect 2872 23069 2881 23103
rect 2881 23069 2915 23103
rect 2915 23069 2924 23103
rect 2872 23060 2924 23069
rect 4344 23137 4367 23171
rect 4367 23137 4396 23171
rect 4344 23128 4396 23137
rect 6552 23128 6604 23180
rect 10508 23239 10560 23248
rect 10508 23205 10542 23239
rect 10542 23205 10560 23239
rect 12348 23264 12400 23316
rect 14740 23264 14792 23316
rect 20628 23264 20680 23316
rect 10508 23196 10560 23205
rect 13544 23196 13596 23248
rect 17132 23239 17184 23248
rect 17132 23205 17141 23239
rect 17141 23205 17175 23239
rect 17175 23205 17184 23239
rect 17132 23196 17184 23205
rect 21180 23239 21232 23248
rect 21180 23205 21189 23239
rect 21189 23205 21223 23239
rect 21223 23205 21232 23239
rect 21180 23196 21232 23205
rect 23388 23196 23440 23248
rect 7656 23128 7708 23180
rect 12992 23171 13044 23180
rect 12992 23137 13026 23171
rect 13026 23137 13044 23171
rect 12992 23128 13044 23137
rect 15568 23128 15620 23180
rect 16120 23128 16172 23180
rect 16764 23128 16816 23180
rect 18236 23128 18288 23180
rect 19432 23171 19484 23180
rect 19432 23137 19441 23171
rect 19441 23137 19475 23171
rect 19475 23137 19484 23171
rect 19432 23128 19484 23137
rect 20904 23171 20956 23180
rect 20904 23137 20913 23171
rect 20913 23137 20947 23171
rect 20947 23137 20956 23171
rect 20904 23128 20956 23137
rect 22468 23171 22520 23180
rect 22468 23137 22477 23171
rect 22477 23137 22511 23171
rect 22511 23137 22520 23171
rect 22468 23128 22520 23137
rect 2780 22992 2832 23044
rect 3332 23060 3384 23112
rect 3884 23060 3936 23112
rect 9036 23060 9088 23112
rect 9956 23060 10008 23112
rect 10232 23103 10284 23112
rect 10232 23069 10241 23103
rect 10241 23069 10275 23103
rect 10275 23069 10284 23103
rect 10232 23060 10284 23069
rect 12532 23060 12584 23112
rect 15936 23103 15988 23112
rect 15936 23069 15945 23103
rect 15945 23069 15979 23103
rect 15979 23069 15988 23103
rect 15936 23060 15988 23069
rect 3516 22967 3568 22976
rect 3516 22933 3525 22967
rect 3525 22933 3559 22967
rect 3559 22933 3568 22967
rect 3516 22924 3568 22933
rect 5448 22967 5500 22976
rect 5448 22933 5457 22967
rect 5457 22933 5491 22967
rect 5491 22933 5500 22967
rect 5448 22924 5500 22933
rect 15292 22967 15344 22976
rect 15292 22933 15301 22967
rect 15301 22933 15335 22967
rect 15335 22933 15344 22967
rect 15292 22924 15344 22933
rect 15476 22924 15528 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 2412 22763 2464 22772
rect 2412 22729 2421 22763
rect 2421 22729 2455 22763
rect 2455 22729 2464 22763
rect 2412 22720 2464 22729
rect 2688 22720 2740 22772
rect 2044 22584 2096 22636
rect 2872 22652 2924 22704
rect 3608 22627 3660 22636
rect 3608 22593 3617 22627
rect 3617 22593 3651 22627
rect 3651 22593 3660 22627
rect 3608 22584 3660 22593
rect 4160 22584 4212 22636
rect 6644 22720 6696 22772
rect 6828 22720 6880 22772
rect 8576 22720 8628 22772
rect 10508 22763 10560 22772
rect 10508 22729 10517 22763
rect 10517 22729 10551 22763
rect 10551 22729 10560 22763
rect 10508 22720 10560 22729
rect 12992 22720 13044 22772
rect 13544 22720 13596 22772
rect 14464 22720 14516 22772
rect 14740 22720 14792 22772
rect 19432 22763 19484 22772
rect 19432 22729 19441 22763
rect 19441 22729 19475 22763
rect 19475 22729 19484 22763
rect 19432 22720 19484 22729
rect 20904 22763 20956 22772
rect 20904 22729 20913 22763
rect 20913 22729 20947 22763
rect 20947 22729 20956 22763
rect 20904 22720 20956 22729
rect 16856 22695 16908 22704
rect 16856 22661 16865 22695
rect 16865 22661 16899 22695
rect 16899 22661 16908 22695
rect 16856 22652 16908 22661
rect 7564 22627 7616 22636
rect 7564 22593 7573 22627
rect 7573 22593 7607 22627
rect 7607 22593 7616 22627
rect 7564 22584 7616 22593
rect 13728 22627 13780 22636
rect 13728 22593 13737 22627
rect 13737 22593 13771 22627
rect 13771 22593 13780 22627
rect 13728 22584 13780 22593
rect 13912 22627 13964 22636
rect 13912 22593 13921 22627
rect 13921 22593 13955 22627
rect 13955 22593 13964 22627
rect 13912 22584 13964 22593
rect 15476 22627 15528 22636
rect 15476 22593 15485 22627
rect 15485 22593 15519 22627
rect 15519 22593 15528 22627
rect 15476 22584 15528 22593
rect 2688 22516 2740 22568
rect 2780 22516 2832 22568
rect 4988 22559 5040 22568
rect 4988 22525 4997 22559
rect 4997 22525 5031 22559
rect 5031 22525 5040 22559
rect 4988 22516 5040 22525
rect 7656 22516 7708 22568
rect 2872 22448 2924 22500
rect 3056 22448 3108 22500
rect 8668 22516 8720 22568
rect 13268 22516 13320 22568
rect 22468 22559 22520 22568
rect 22468 22525 22477 22559
rect 22477 22525 22511 22559
rect 22511 22525 22520 22559
rect 22468 22516 22520 22525
rect 3332 22423 3384 22432
rect 3332 22389 3341 22423
rect 3341 22389 3375 22423
rect 3375 22389 3384 22423
rect 3332 22380 3384 22389
rect 3516 22380 3568 22432
rect 4068 22380 4120 22432
rect 4528 22380 4580 22432
rect 7104 22380 7156 22432
rect 9036 22448 9088 22500
rect 10232 22448 10284 22500
rect 8760 22380 8812 22432
rect 9588 22380 9640 22432
rect 11060 22423 11112 22432
rect 11060 22389 11069 22423
rect 11069 22389 11103 22423
rect 11103 22389 11112 22423
rect 11060 22380 11112 22389
rect 15752 22491 15804 22500
rect 15752 22457 15764 22491
rect 15764 22457 15804 22491
rect 15752 22448 15804 22457
rect 16120 22448 16172 22500
rect 16764 22448 16816 22500
rect 12532 22380 12584 22432
rect 14188 22380 14240 22432
rect 15568 22380 15620 22432
rect 18236 22423 18288 22432
rect 18236 22389 18245 22423
rect 18245 22389 18279 22423
rect 18279 22389 18288 22423
rect 18236 22380 18288 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 10968 22176 11020 22228
rect 13360 22176 13412 22228
rect 13728 22219 13780 22228
rect 13728 22185 13737 22219
rect 13737 22185 13771 22219
rect 13771 22185 13780 22219
rect 13728 22176 13780 22185
rect 15476 22176 15528 22228
rect 3332 22108 3384 22160
rect 5448 22108 5500 22160
rect 7380 22108 7432 22160
rect 8024 22151 8076 22160
rect 8024 22117 8033 22151
rect 8033 22117 8067 22151
rect 8067 22117 8076 22151
rect 8024 22108 8076 22117
rect 1584 22083 1636 22092
rect 1584 22049 1593 22083
rect 1593 22049 1627 22083
rect 1627 22049 1636 22083
rect 1584 22040 1636 22049
rect 2412 22040 2464 22092
rect 2688 22040 2740 22092
rect 2780 22040 2832 22092
rect 7656 22040 7708 22092
rect 6644 21972 6696 22024
rect 8116 22015 8168 22024
rect 8116 21981 8125 22015
rect 8125 21981 8159 22015
rect 8159 21981 8168 22015
rect 8116 21972 8168 21981
rect 8392 22040 8444 22092
rect 9588 22040 9640 22092
rect 10048 22040 10100 22092
rect 13452 22040 13504 22092
rect 14832 22040 14884 22092
rect 9128 21972 9180 22024
rect 10232 22015 10284 22024
rect 10232 21981 10241 22015
rect 10241 21981 10275 22015
rect 10275 21981 10284 22015
rect 10232 21972 10284 21981
rect 10416 22015 10468 22024
rect 10416 21981 10425 22015
rect 10425 21981 10459 22015
rect 10459 21981 10468 22015
rect 10416 21972 10468 21981
rect 15936 22040 15988 22092
rect 6276 21947 6328 21956
rect 6276 21913 6285 21947
rect 6285 21913 6319 21947
rect 6319 21913 6328 21947
rect 6276 21904 6328 21913
rect 8024 21904 8076 21956
rect 10968 21904 11020 21956
rect 3056 21879 3108 21888
rect 3056 21845 3065 21879
rect 3065 21845 3099 21879
rect 3099 21845 3108 21879
rect 3056 21836 3108 21845
rect 3884 21879 3936 21888
rect 3884 21845 3893 21879
rect 3893 21845 3927 21879
rect 3927 21845 3936 21879
rect 3884 21836 3936 21845
rect 4528 21879 4580 21888
rect 4528 21845 4537 21879
rect 4537 21845 4571 21879
rect 4571 21845 4580 21879
rect 4528 21836 4580 21845
rect 7104 21879 7156 21888
rect 7104 21845 7113 21879
rect 7113 21845 7147 21879
rect 7147 21845 7156 21879
rect 7104 21836 7156 21845
rect 7656 21879 7708 21888
rect 7656 21845 7665 21879
rect 7665 21845 7699 21879
rect 7699 21845 7708 21879
rect 7656 21836 7708 21845
rect 9036 21879 9088 21888
rect 9036 21845 9045 21879
rect 9045 21845 9079 21879
rect 9079 21845 9088 21879
rect 9036 21836 9088 21845
rect 10692 21836 10744 21888
rect 12808 21836 12860 21888
rect 13268 21879 13320 21888
rect 13268 21845 13277 21879
rect 13277 21845 13311 21879
rect 13311 21845 13320 21879
rect 13268 21836 13320 21845
rect 15752 21836 15804 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 2780 21632 2832 21684
rect 4160 21675 4212 21684
rect 4160 21641 4169 21675
rect 4169 21641 4203 21675
rect 4203 21641 4212 21675
rect 4160 21632 4212 21641
rect 2228 21496 2280 21548
rect 3332 21496 3384 21548
rect 4344 21496 4396 21548
rect 5448 21632 5500 21684
rect 6644 21675 6696 21684
rect 6644 21641 6653 21675
rect 6653 21641 6687 21675
rect 6687 21641 6696 21675
rect 6644 21632 6696 21641
rect 7380 21675 7432 21684
rect 7380 21641 7389 21675
rect 7389 21641 7423 21675
rect 7423 21641 7432 21675
rect 7380 21632 7432 21641
rect 10140 21632 10192 21684
rect 10416 21632 10468 21684
rect 12164 21607 12216 21616
rect 12164 21573 12173 21607
rect 12173 21573 12207 21607
rect 12207 21573 12216 21607
rect 12164 21564 12216 21573
rect 5540 21496 5592 21548
rect 10692 21496 10744 21548
rect 11888 21496 11940 21548
rect 13636 21496 13688 21548
rect 13912 21496 13964 21548
rect 5172 21428 5224 21480
rect 9036 21428 9088 21480
rect 9772 21428 9824 21480
rect 1768 21335 1820 21344
rect 1768 21301 1777 21335
rect 1777 21301 1811 21335
rect 1811 21301 1820 21335
rect 1768 21292 1820 21301
rect 3424 21292 3476 21344
rect 6276 21360 6328 21412
rect 8024 21360 8076 21412
rect 9128 21360 9180 21412
rect 9680 21360 9732 21412
rect 12164 21360 12216 21412
rect 15476 21360 15528 21412
rect 5632 21335 5684 21344
rect 5632 21301 5641 21335
rect 5641 21301 5675 21335
rect 5675 21301 5684 21335
rect 5632 21292 5684 21301
rect 6552 21292 6604 21344
rect 9312 21292 9364 21344
rect 9772 21335 9824 21344
rect 9772 21301 9781 21335
rect 9781 21301 9815 21335
rect 9815 21301 9824 21335
rect 9772 21292 9824 21301
rect 9956 21335 10008 21344
rect 9956 21301 9965 21335
rect 9965 21301 9999 21335
rect 9999 21301 10008 21335
rect 9956 21292 10008 21301
rect 11888 21335 11940 21344
rect 11888 21301 11897 21335
rect 11897 21301 11931 21335
rect 11931 21301 11940 21335
rect 11888 21292 11940 21301
rect 12440 21335 12492 21344
rect 12440 21301 12449 21335
rect 12449 21301 12483 21335
rect 12483 21301 12492 21335
rect 12808 21335 12860 21344
rect 12440 21292 12492 21301
rect 12808 21301 12817 21335
rect 12817 21301 12851 21335
rect 12851 21301 12860 21335
rect 12808 21292 12860 21301
rect 13452 21335 13504 21344
rect 13452 21301 13461 21335
rect 13461 21301 13495 21335
rect 13495 21301 13504 21335
rect 13452 21292 13504 21301
rect 13820 21335 13872 21344
rect 13820 21301 13829 21335
rect 13829 21301 13863 21335
rect 13863 21301 13872 21335
rect 13820 21292 13872 21301
rect 15936 21335 15988 21344
rect 15936 21301 15945 21335
rect 15945 21301 15979 21335
rect 15979 21301 15988 21335
rect 15936 21292 15988 21301
rect 16396 21335 16448 21344
rect 16396 21301 16405 21335
rect 16405 21301 16439 21335
rect 16439 21301 16448 21335
rect 16396 21292 16448 21301
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 1584 21131 1636 21140
rect 1584 21097 1593 21131
rect 1593 21097 1627 21131
rect 1627 21097 1636 21131
rect 1584 21088 1636 21097
rect 4344 21131 4396 21140
rect 4344 21097 4353 21131
rect 4353 21097 4387 21131
rect 4387 21097 4396 21131
rect 4344 21088 4396 21097
rect 8392 21131 8444 21140
rect 8392 21097 8401 21131
rect 8401 21097 8435 21131
rect 8435 21097 8444 21131
rect 8392 21088 8444 21097
rect 12440 21088 12492 21140
rect 13912 21088 13964 21140
rect 15292 21088 15344 21140
rect 16028 21088 16080 21140
rect 2596 21020 2648 21072
rect 5080 21020 5132 21072
rect 10048 21020 10100 21072
rect 10876 21020 10928 21072
rect 1952 20995 2004 21004
rect 1952 20961 1961 20995
rect 1961 20961 1995 20995
rect 1995 20961 2004 20995
rect 1952 20952 2004 20961
rect 3884 20952 3936 21004
rect 5632 20952 5684 21004
rect 6276 20952 6328 21004
rect 8208 20952 8260 21004
rect 10692 20952 10744 21004
rect 12532 20952 12584 21004
rect 7104 20884 7156 20936
rect 7840 20927 7892 20936
rect 7840 20893 7849 20927
rect 7849 20893 7883 20927
rect 7883 20893 7892 20927
rect 7840 20884 7892 20893
rect 8024 20927 8076 20936
rect 8024 20893 8033 20927
rect 8033 20893 8067 20927
rect 8067 20893 8076 20927
rect 8024 20884 8076 20893
rect 12992 20927 13044 20936
rect 12992 20893 13001 20927
rect 13001 20893 13035 20927
rect 13035 20893 13044 20927
rect 12992 20884 13044 20893
rect 13820 20952 13872 21004
rect 15292 20952 15344 21004
rect 14556 20884 14608 20936
rect 15844 20927 15896 20936
rect 15844 20893 15853 20927
rect 15853 20893 15887 20927
rect 15887 20893 15896 20927
rect 15844 20884 15896 20893
rect 12532 20859 12584 20868
rect 12532 20825 12541 20859
rect 12541 20825 12575 20859
rect 12575 20825 12584 20859
rect 12532 20816 12584 20825
rect 15384 20816 15436 20868
rect 5540 20748 5592 20800
rect 6920 20748 6972 20800
rect 7380 20791 7432 20800
rect 7380 20757 7389 20791
rect 7389 20757 7423 20791
rect 7423 20757 7432 20791
rect 7380 20748 7432 20757
rect 9036 20791 9088 20800
rect 9036 20757 9045 20791
rect 9045 20757 9079 20791
rect 9079 20757 9088 20791
rect 9036 20748 9088 20757
rect 9404 20791 9456 20800
rect 9404 20757 9413 20791
rect 9413 20757 9447 20791
rect 9447 20757 9456 20791
rect 9404 20748 9456 20757
rect 11612 20748 11664 20800
rect 13360 20748 13412 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 1676 20587 1728 20596
rect 1676 20553 1685 20587
rect 1685 20553 1719 20587
rect 1719 20553 1728 20587
rect 1676 20544 1728 20553
rect 1952 20544 2004 20596
rect 2504 20587 2556 20596
rect 2504 20553 2513 20587
rect 2513 20553 2547 20587
rect 2547 20553 2556 20587
rect 2504 20544 2556 20553
rect 8208 20544 8260 20596
rect 11888 20587 11940 20596
rect 11888 20553 11897 20587
rect 11897 20553 11931 20587
rect 11931 20553 11940 20587
rect 11888 20544 11940 20553
rect 12348 20544 12400 20596
rect 13820 20544 13872 20596
rect 14556 20587 14608 20596
rect 14556 20553 14565 20587
rect 14565 20553 14599 20587
rect 14599 20553 14608 20587
rect 14556 20544 14608 20553
rect 15844 20544 15896 20596
rect 5080 20476 5132 20528
rect 7840 20476 7892 20528
rect 2044 20451 2096 20460
rect 2044 20417 2053 20451
rect 2053 20417 2087 20451
rect 2087 20417 2096 20451
rect 2044 20408 2096 20417
rect 5448 20408 5500 20460
rect 15292 20476 15344 20528
rect 15936 20408 15988 20460
rect 16672 20451 16724 20460
rect 16672 20417 16681 20451
rect 16681 20417 16715 20451
rect 16715 20417 16724 20451
rect 16672 20408 16724 20417
rect 1676 20340 1728 20392
rect 5908 20340 5960 20392
rect 6552 20383 6604 20392
rect 6552 20349 6561 20383
rect 6561 20349 6595 20383
rect 6595 20349 6604 20383
rect 6552 20340 6604 20349
rect 4344 20272 4396 20324
rect 6920 20340 6972 20392
rect 9036 20340 9088 20392
rect 11336 20340 11388 20392
rect 13360 20340 13412 20392
rect 14556 20340 14608 20392
rect 2872 20247 2924 20256
rect 2872 20213 2881 20247
rect 2881 20213 2915 20247
rect 2915 20213 2924 20247
rect 2872 20204 2924 20213
rect 3240 20247 3292 20256
rect 3240 20213 3249 20247
rect 3249 20213 3283 20247
rect 3283 20213 3292 20247
rect 3240 20204 3292 20213
rect 4804 20247 4856 20256
rect 4804 20213 4813 20247
rect 4813 20213 4847 20247
rect 4847 20213 4856 20247
rect 4804 20204 4856 20213
rect 6276 20204 6328 20256
rect 7748 20272 7800 20324
rect 9404 20272 9456 20324
rect 12716 20272 12768 20324
rect 8024 20204 8076 20256
rect 8576 20204 8628 20256
rect 9772 20204 9824 20256
rect 10692 20247 10744 20256
rect 10692 20213 10701 20247
rect 10701 20213 10735 20247
rect 10735 20213 10744 20247
rect 10692 20204 10744 20213
rect 15384 20204 15436 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 3884 20043 3936 20052
rect 3884 20009 3893 20043
rect 3893 20009 3927 20043
rect 3927 20009 3936 20043
rect 3884 20000 3936 20009
rect 4344 20043 4396 20052
rect 4344 20009 4353 20043
rect 4353 20009 4387 20043
rect 4387 20009 4396 20043
rect 4344 20000 4396 20009
rect 5908 20043 5960 20052
rect 5908 20009 5917 20043
rect 5917 20009 5951 20043
rect 5951 20009 5960 20043
rect 5908 20000 5960 20009
rect 6828 20000 6880 20052
rect 7380 20000 7432 20052
rect 9956 20000 10008 20052
rect 12716 20043 12768 20052
rect 12716 20009 12725 20043
rect 12725 20009 12759 20043
rect 12759 20009 12768 20043
rect 12716 20000 12768 20009
rect 13544 20000 13596 20052
rect 15292 20000 15344 20052
rect 16028 20043 16080 20052
rect 16028 20009 16037 20043
rect 16037 20009 16071 20043
rect 16071 20009 16080 20043
rect 16028 20000 16080 20009
rect 17408 20000 17460 20052
rect 2596 19932 2648 19984
rect 2964 19975 3016 19984
rect 2964 19941 2973 19975
rect 2973 19941 3007 19975
rect 3007 19941 3016 19975
rect 2964 19932 3016 19941
rect 3700 19932 3752 19984
rect 7288 19932 7340 19984
rect 10600 19932 10652 19984
rect 10876 19932 10928 19984
rect 14096 19975 14148 19984
rect 14096 19941 14105 19975
rect 14105 19941 14139 19975
rect 14139 19941 14148 19975
rect 14096 19932 14148 19941
rect 2688 19907 2740 19916
rect 2688 19873 2697 19907
rect 2697 19873 2731 19907
rect 2731 19873 2740 19907
rect 2688 19864 2740 19873
rect 2780 19864 2832 19916
rect 4712 19907 4764 19916
rect 4712 19873 4721 19907
rect 4721 19873 4755 19907
rect 4755 19873 4764 19907
rect 4712 19864 4764 19873
rect 2228 19839 2280 19848
rect 2228 19805 2237 19839
rect 2237 19805 2271 19839
rect 2271 19805 2280 19839
rect 2228 19796 2280 19805
rect 4344 19796 4396 19848
rect 4528 19796 4580 19848
rect 6644 19864 6696 19916
rect 8300 19864 8352 19916
rect 9128 19864 9180 19916
rect 11612 19907 11664 19916
rect 11612 19873 11635 19907
rect 11635 19873 11664 19907
rect 13820 19907 13872 19916
rect 11612 19864 11664 19873
rect 13820 19873 13829 19907
rect 13829 19873 13863 19907
rect 13863 19873 13872 19907
rect 13820 19864 13872 19873
rect 15292 19907 15344 19916
rect 15292 19873 15301 19907
rect 15301 19873 15335 19907
rect 15335 19873 15344 19907
rect 15292 19864 15344 19873
rect 16580 19907 16632 19916
rect 16580 19873 16589 19907
rect 16589 19873 16623 19907
rect 16623 19873 16632 19907
rect 16580 19864 16632 19873
rect 6552 19839 6604 19848
rect 4804 19728 4856 19780
rect 6552 19805 6561 19839
rect 6561 19805 6595 19839
rect 6595 19805 6604 19839
rect 6552 19796 6604 19805
rect 7748 19796 7800 19848
rect 10232 19839 10284 19848
rect 10232 19805 10241 19839
rect 10241 19805 10275 19839
rect 10275 19805 10284 19839
rect 10232 19796 10284 19805
rect 10324 19839 10376 19848
rect 10324 19805 10333 19839
rect 10333 19805 10367 19839
rect 10367 19805 10376 19839
rect 10324 19796 10376 19805
rect 5080 19728 5132 19780
rect 7012 19728 7064 19780
rect 10048 19728 10100 19780
rect 1952 19660 2004 19712
rect 2596 19660 2648 19712
rect 5264 19660 5316 19712
rect 7380 19703 7432 19712
rect 7380 19669 7389 19703
rect 7389 19669 7423 19703
rect 7423 19669 7432 19703
rect 7380 19660 7432 19669
rect 8576 19703 8628 19712
rect 8576 19669 8585 19703
rect 8585 19669 8619 19703
rect 8619 19669 8628 19703
rect 8576 19660 8628 19669
rect 9036 19703 9088 19712
rect 9036 19669 9045 19703
rect 9045 19669 9079 19703
rect 9079 19669 9088 19703
rect 9036 19660 9088 19669
rect 10876 19703 10928 19712
rect 10876 19669 10885 19703
rect 10885 19669 10919 19703
rect 10919 19669 10928 19703
rect 10876 19660 10928 19669
rect 11336 19660 11388 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 6644 19456 6696 19508
rect 10324 19456 10376 19508
rect 11612 19456 11664 19508
rect 12992 19499 13044 19508
rect 12992 19465 13001 19499
rect 13001 19465 13035 19499
rect 13035 19465 13044 19499
rect 12992 19456 13044 19465
rect 16580 19456 16632 19508
rect 10232 19388 10284 19440
rect 7288 19363 7340 19372
rect 1400 19252 1452 19304
rect 2504 19252 2556 19304
rect 1492 19159 1544 19168
rect 1492 19125 1501 19159
rect 1501 19125 1535 19159
rect 1535 19125 1544 19159
rect 1492 19116 1544 19125
rect 1952 19159 2004 19168
rect 1952 19125 1961 19159
rect 1961 19125 1995 19159
rect 1995 19125 2004 19159
rect 1952 19116 2004 19125
rect 7288 19329 7297 19363
rect 7297 19329 7331 19363
rect 7331 19329 7340 19363
rect 7288 19320 7340 19329
rect 8208 19320 8260 19372
rect 8576 19320 8628 19372
rect 10692 19320 10744 19372
rect 13544 19363 13596 19372
rect 13544 19329 13553 19363
rect 13553 19329 13587 19363
rect 13587 19329 13596 19363
rect 13544 19320 13596 19329
rect 3148 19252 3200 19304
rect 3884 19252 3936 19304
rect 5540 19295 5592 19304
rect 5540 19261 5549 19295
rect 5549 19261 5583 19295
rect 5583 19261 5592 19295
rect 5540 19252 5592 19261
rect 6828 19252 6880 19304
rect 8760 19295 8812 19304
rect 8760 19261 8769 19295
rect 8769 19261 8803 19295
rect 8803 19261 8812 19295
rect 8760 19252 8812 19261
rect 10232 19252 10284 19304
rect 11244 19295 11296 19304
rect 11244 19261 11253 19295
rect 11253 19261 11287 19295
rect 11287 19261 11296 19295
rect 11244 19252 11296 19261
rect 12440 19252 12492 19304
rect 13636 19252 13688 19304
rect 13728 19252 13780 19304
rect 15292 19320 15344 19372
rect 15476 19252 15528 19304
rect 11152 19227 11204 19236
rect 11152 19193 11161 19227
rect 11161 19193 11195 19227
rect 11195 19193 11204 19227
rect 11152 19184 11204 19193
rect 11336 19184 11388 19236
rect 13912 19184 13964 19236
rect 14280 19184 14332 19236
rect 16672 19184 16724 19236
rect 2688 19116 2740 19168
rect 3056 19116 3108 19168
rect 4528 19116 4580 19168
rect 4804 19116 4856 19168
rect 5356 19159 5408 19168
rect 5356 19125 5365 19159
rect 5365 19125 5399 19159
rect 5399 19125 5408 19159
rect 5356 19116 5408 19125
rect 5540 19116 5592 19168
rect 6828 19159 6880 19168
rect 6828 19125 6837 19159
rect 6837 19125 6871 19159
rect 6871 19125 6880 19159
rect 6828 19116 6880 19125
rect 7012 19116 7064 19168
rect 7380 19116 7432 19168
rect 7564 19116 7616 19168
rect 8300 19116 8352 19168
rect 8852 19159 8904 19168
rect 8852 19125 8861 19159
rect 8861 19125 8895 19159
rect 8895 19125 8904 19159
rect 8852 19116 8904 19125
rect 13544 19116 13596 19168
rect 13636 19116 13688 19168
rect 13820 19116 13872 19168
rect 15476 19116 15528 19168
rect 16764 19159 16816 19168
rect 16764 19125 16773 19159
rect 16773 19125 16807 19159
rect 16807 19125 16816 19159
rect 16764 19116 16816 19125
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 1400 18955 1452 18964
rect 1400 18921 1409 18955
rect 1409 18921 1443 18955
rect 1443 18921 1452 18955
rect 1400 18912 1452 18921
rect 2780 18955 2832 18964
rect 2780 18921 2789 18955
rect 2789 18921 2823 18955
rect 2823 18921 2832 18955
rect 2780 18912 2832 18921
rect 4712 18912 4764 18964
rect 5356 18912 5408 18964
rect 1400 18708 1452 18760
rect 4252 18844 4304 18896
rect 5080 18844 5132 18896
rect 1768 18819 1820 18828
rect 1768 18785 1777 18819
rect 1777 18785 1811 18819
rect 1811 18785 1820 18819
rect 1768 18776 1820 18785
rect 4160 18776 4212 18828
rect 6460 18912 6512 18964
rect 7748 18955 7800 18964
rect 7748 18921 7757 18955
rect 7757 18921 7791 18955
rect 7791 18921 7800 18955
rect 7748 18912 7800 18921
rect 8208 18912 8260 18964
rect 8300 18912 8352 18964
rect 9220 18955 9272 18964
rect 9220 18921 9229 18955
rect 9229 18921 9263 18955
rect 9263 18921 9272 18955
rect 9220 18912 9272 18921
rect 9956 18955 10008 18964
rect 9956 18921 9965 18955
rect 9965 18921 9999 18955
rect 9999 18921 10008 18955
rect 9956 18912 10008 18921
rect 10048 18912 10100 18964
rect 13636 18955 13688 18964
rect 13636 18921 13645 18955
rect 13645 18921 13679 18955
rect 13679 18921 13688 18955
rect 13636 18912 13688 18921
rect 14372 18912 14424 18964
rect 14648 18912 14700 18964
rect 16672 18955 16724 18964
rect 16672 18921 16681 18955
rect 16681 18921 16715 18955
rect 16715 18921 16724 18955
rect 16672 18912 16724 18921
rect 6184 18844 6236 18896
rect 10968 18844 11020 18896
rect 12624 18844 12676 18896
rect 18052 18844 18104 18896
rect 6276 18776 6328 18828
rect 8576 18776 8628 18828
rect 10140 18776 10192 18828
rect 11704 18776 11756 18828
rect 14004 18819 14056 18828
rect 14004 18785 14013 18819
rect 14013 18785 14047 18819
rect 14047 18785 14056 18819
rect 14004 18776 14056 18785
rect 14372 18776 14424 18828
rect 15936 18776 15988 18828
rect 4712 18751 4764 18760
rect 4712 18717 4721 18751
rect 4721 18717 4755 18751
rect 4755 18717 4764 18751
rect 4712 18708 4764 18717
rect 10600 18751 10652 18760
rect 10600 18717 10609 18751
rect 10609 18717 10643 18751
rect 10643 18717 10652 18751
rect 10600 18708 10652 18717
rect 12164 18751 12216 18760
rect 12164 18717 12173 18751
rect 12173 18717 12207 18751
rect 12207 18717 12216 18751
rect 12164 18708 12216 18717
rect 14280 18751 14332 18760
rect 14280 18717 14289 18751
rect 14289 18717 14323 18751
rect 14323 18717 14332 18751
rect 14280 18708 14332 18717
rect 4528 18640 4580 18692
rect 8392 18683 8444 18692
rect 8392 18649 8401 18683
rect 8401 18649 8435 18683
rect 8435 18649 8444 18683
rect 8392 18640 8444 18649
rect 2504 18615 2556 18624
rect 2504 18581 2513 18615
rect 2513 18581 2547 18615
rect 2547 18581 2556 18615
rect 2504 18572 2556 18581
rect 5080 18572 5132 18624
rect 5356 18572 5408 18624
rect 7012 18572 7064 18624
rect 10876 18572 10928 18624
rect 11152 18615 11204 18624
rect 11152 18581 11161 18615
rect 11161 18581 11195 18615
rect 11195 18581 11204 18615
rect 11152 18572 11204 18581
rect 12440 18572 12492 18624
rect 13544 18572 13596 18624
rect 13912 18572 13964 18624
rect 15476 18572 15528 18624
rect 16396 18572 16448 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 4160 18411 4212 18420
rect 4160 18377 4169 18411
rect 4169 18377 4203 18411
rect 4203 18377 4212 18411
rect 4160 18368 4212 18377
rect 4252 18368 4304 18420
rect 5172 18411 5224 18420
rect 5172 18377 5181 18411
rect 5181 18377 5215 18411
rect 5215 18377 5224 18411
rect 5172 18368 5224 18377
rect 8208 18368 8260 18420
rect 8668 18368 8720 18420
rect 10048 18368 10100 18420
rect 11888 18411 11940 18420
rect 11888 18377 11897 18411
rect 11897 18377 11931 18411
rect 11931 18377 11940 18411
rect 11888 18368 11940 18377
rect 12164 18368 12216 18420
rect 14004 18368 14056 18420
rect 5448 18300 5500 18352
rect 6276 18300 6328 18352
rect 10692 18300 10744 18352
rect 11244 18300 11296 18352
rect 14280 18300 14332 18352
rect 14740 18343 14792 18352
rect 14740 18309 14749 18343
rect 14749 18309 14783 18343
rect 14783 18309 14792 18343
rect 14740 18300 14792 18309
rect 7012 18232 7064 18284
rect 9680 18275 9732 18284
rect 1492 18164 1544 18216
rect 3148 18164 3200 18216
rect 5540 18164 5592 18216
rect 6276 18164 6328 18216
rect 9680 18241 9689 18275
rect 9689 18241 9723 18275
rect 9723 18241 9732 18275
rect 9680 18232 9732 18241
rect 10600 18232 10652 18284
rect 12164 18275 12216 18284
rect 12164 18241 12173 18275
rect 12173 18241 12207 18275
rect 12207 18241 12216 18275
rect 12164 18232 12216 18241
rect 11152 18207 11204 18216
rect 2688 18096 2740 18148
rect 1860 18028 1912 18080
rect 2964 18028 3016 18080
rect 3056 18028 3108 18080
rect 5264 18028 5316 18080
rect 6920 18096 6972 18148
rect 11152 18173 11161 18207
rect 11161 18173 11195 18207
rect 11195 18173 11204 18207
rect 11152 18164 11204 18173
rect 12440 18207 12492 18216
rect 12440 18173 12449 18207
rect 12449 18173 12483 18207
rect 12483 18173 12492 18207
rect 12440 18164 12492 18173
rect 15936 18232 15988 18284
rect 7840 18096 7892 18148
rect 10600 18139 10652 18148
rect 10600 18105 10609 18139
rect 10609 18105 10643 18139
rect 10643 18105 10652 18139
rect 10600 18096 10652 18105
rect 15108 18096 15160 18148
rect 6184 18071 6236 18080
rect 6184 18037 6193 18071
rect 6193 18037 6227 18071
rect 6227 18037 6236 18071
rect 6184 18028 6236 18037
rect 7012 18028 7064 18080
rect 7288 18028 7340 18080
rect 8576 18028 8628 18080
rect 9956 18028 10008 18080
rect 10784 18071 10836 18080
rect 10784 18037 10793 18071
rect 10793 18037 10827 18071
rect 10827 18037 10836 18071
rect 10784 18028 10836 18037
rect 11060 18028 11112 18080
rect 13820 18071 13872 18080
rect 13820 18037 13829 18071
rect 13829 18037 13863 18071
rect 13863 18037 13872 18071
rect 13820 18028 13872 18037
rect 15936 18071 15988 18080
rect 15936 18037 15945 18071
rect 15945 18037 15979 18071
rect 15979 18037 15988 18071
rect 15936 18028 15988 18037
rect 16396 18071 16448 18080
rect 16396 18037 16405 18071
rect 16405 18037 16439 18071
rect 16439 18037 16448 18071
rect 16396 18028 16448 18037
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 2964 17824 3016 17876
rect 3148 17824 3200 17876
rect 6920 17867 6972 17876
rect 6920 17833 6929 17867
rect 6929 17833 6963 17867
rect 6963 17833 6972 17867
rect 6920 17824 6972 17833
rect 9772 17824 9824 17876
rect 10968 17824 11020 17876
rect 12164 17867 12216 17876
rect 12164 17833 12173 17867
rect 12173 17833 12207 17867
rect 12207 17833 12216 17867
rect 12164 17824 12216 17833
rect 12716 17867 12768 17876
rect 12716 17833 12725 17867
rect 12725 17833 12759 17867
rect 12759 17833 12768 17867
rect 12716 17824 12768 17833
rect 15108 17824 15160 17876
rect 4620 17756 4672 17808
rect 10876 17756 10928 17808
rect 11888 17756 11940 17808
rect 12440 17756 12492 17808
rect 15660 17799 15712 17808
rect 848 17688 900 17740
rect 2412 17688 2464 17740
rect 2964 17688 3016 17740
rect 5448 17688 5500 17740
rect 7288 17731 7340 17740
rect 7288 17697 7297 17731
rect 7297 17697 7331 17731
rect 7331 17697 7340 17731
rect 7288 17688 7340 17697
rect 1860 17620 1912 17672
rect 3056 17663 3108 17672
rect 3056 17629 3065 17663
rect 3065 17629 3099 17663
rect 3099 17629 3108 17663
rect 3056 17620 3108 17629
rect 7380 17663 7432 17672
rect 7380 17629 7389 17663
rect 7389 17629 7423 17663
rect 7423 17629 7432 17663
rect 7380 17620 7432 17629
rect 8484 17663 8536 17672
rect 2044 17552 2096 17604
rect 5540 17552 5592 17604
rect 8484 17629 8493 17663
rect 8493 17629 8527 17663
rect 8527 17629 8536 17663
rect 8484 17620 8536 17629
rect 11336 17688 11388 17740
rect 12624 17688 12676 17740
rect 14004 17688 14056 17740
rect 14832 17688 14884 17740
rect 15660 17765 15669 17799
rect 15669 17765 15703 17799
rect 15703 17765 15712 17799
rect 15660 17756 15712 17765
rect 17408 17688 17460 17740
rect 13176 17663 13228 17672
rect 1676 17484 1728 17536
rect 3608 17484 3660 17536
rect 4620 17484 4672 17536
rect 5448 17484 5500 17536
rect 6184 17484 6236 17536
rect 6368 17527 6420 17536
rect 6368 17493 6377 17527
rect 6377 17493 6411 17527
rect 6411 17493 6420 17527
rect 6368 17484 6420 17493
rect 6644 17484 6696 17536
rect 8760 17552 8812 17604
rect 9036 17552 9088 17604
rect 13176 17629 13185 17663
rect 13185 17629 13219 17663
rect 13219 17629 13228 17663
rect 13820 17663 13872 17672
rect 13176 17620 13228 17629
rect 13820 17629 13829 17663
rect 13829 17629 13863 17663
rect 13863 17629 13872 17663
rect 13820 17620 13872 17629
rect 15752 17663 15804 17672
rect 15752 17629 15761 17663
rect 15761 17629 15795 17663
rect 15795 17629 15804 17663
rect 15752 17620 15804 17629
rect 13728 17552 13780 17604
rect 14832 17552 14884 17604
rect 16764 17620 16816 17672
rect 17500 17663 17552 17672
rect 17500 17629 17509 17663
rect 17509 17629 17543 17663
rect 17543 17629 17552 17663
rect 17500 17620 17552 17629
rect 7840 17484 7892 17536
rect 8392 17527 8444 17536
rect 8392 17493 8401 17527
rect 8401 17493 8435 17527
rect 8435 17493 8444 17527
rect 8392 17484 8444 17493
rect 9680 17484 9732 17536
rect 10140 17527 10192 17536
rect 10140 17493 10149 17527
rect 10149 17493 10183 17527
rect 10183 17493 10192 17527
rect 10140 17484 10192 17493
rect 14372 17527 14424 17536
rect 14372 17493 14381 17527
rect 14381 17493 14415 17527
rect 14415 17493 14424 17527
rect 14372 17484 14424 17493
rect 15292 17527 15344 17536
rect 15292 17493 15301 17527
rect 15301 17493 15335 17527
rect 15335 17493 15344 17527
rect 15292 17484 15344 17493
rect 16396 17484 16448 17536
rect 16672 17527 16724 17536
rect 16672 17493 16681 17527
rect 16681 17493 16715 17527
rect 16715 17493 16724 17527
rect 16672 17484 16724 17493
rect 16856 17527 16908 17536
rect 16856 17493 16865 17527
rect 16865 17493 16899 17527
rect 16899 17493 16908 17527
rect 16856 17484 16908 17493
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 1768 17280 1820 17332
rect 2412 17323 2464 17332
rect 2412 17289 2421 17323
rect 2421 17289 2455 17323
rect 2455 17289 2464 17323
rect 2412 17280 2464 17289
rect 3056 17280 3108 17332
rect 5540 17280 5592 17332
rect 7380 17280 7432 17332
rect 8668 17323 8720 17332
rect 8668 17289 8677 17323
rect 8677 17289 8711 17323
rect 8711 17289 8720 17323
rect 8668 17280 8720 17289
rect 10876 17323 10928 17332
rect 10876 17289 10885 17323
rect 10885 17289 10919 17323
rect 10919 17289 10928 17323
rect 10876 17280 10928 17289
rect 12532 17280 12584 17332
rect 15752 17280 15804 17332
rect 17408 17323 17460 17332
rect 17408 17289 17417 17323
rect 17417 17289 17451 17323
rect 17451 17289 17460 17323
rect 17408 17280 17460 17289
rect 17500 17280 17552 17332
rect 3148 17212 3200 17264
rect 4620 17255 4672 17264
rect 2044 17187 2096 17196
rect 2044 17153 2053 17187
rect 2053 17153 2087 17187
rect 2087 17153 2096 17187
rect 2044 17144 2096 17153
rect 4620 17221 4629 17255
rect 4629 17221 4663 17255
rect 4663 17221 4672 17255
rect 4620 17212 4672 17221
rect 6184 17212 6236 17264
rect 6644 17212 6696 17264
rect 4896 17144 4948 17196
rect 5448 17144 5500 17196
rect 6092 17144 6144 17196
rect 3608 17119 3660 17128
rect 3608 17085 3617 17119
rect 3617 17085 3651 17119
rect 3651 17085 3660 17119
rect 3608 17076 3660 17085
rect 6000 17076 6052 17128
rect 6552 17076 6604 17128
rect 6920 17076 6972 17128
rect 7840 17076 7892 17128
rect 8760 17119 8812 17128
rect 8760 17085 8769 17119
rect 8769 17085 8803 17119
rect 8803 17085 8812 17119
rect 8760 17076 8812 17085
rect 9588 17076 9640 17128
rect 12440 17076 12492 17128
rect 1676 17008 1728 17060
rect 1860 16983 1912 16992
rect 1860 16949 1869 16983
rect 1869 16949 1903 16983
rect 1903 16949 1912 16983
rect 1860 16940 1912 16949
rect 6368 17008 6420 17060
rect 13176 17076 13228 17128
rect 15016 17119 15068 17128
rect 15016 17085 15025 17119
rect 15025 17085 15059 17119
rect 15059 17085 15068 17119
rect 15016 17076 15068 17085
rect 15568 17076 15620 17128
rect 16764 17076 16816 17128
rect 17684 17119 17736 17128
rect 17684 17085 17693 17119
rect 17693 17085 17727 17119
rect 17727 17085 17736 17119
rect 17684 17076 17736 17085
rect 13084 17008 13136 17060
rect 14740 17008 14792 17060
rect 3516 16983 3568 16992
rect 3516 16949 3525 16983
rect 3525 16949 3559 16983
rect 3559 16949 3568 16983
rect 3516 16940 3568 16949
rect 5080 16983 5132 16992
rect 5080 16949 5089 16983
rect 5089 16949 5123 16983
rect 5123 16949 5132 16983
rect 5080 16940 5132 16949
rect 6460 16940 6512 16992
rect 8300 16983 8352 16992
rect 8300 16949 8309 16983
rect 8309 16949 8343 16983
rect 8343 16949 8352 16983
rect 8300 16940 8352 16949
rect 11520 16940 11572 16992
rect 11704 16983 11756 16992
rect 11704 16949 11713 16983
rect 11713 16949 11747 16983
rect 11747 16949 11756 16983
rect 11704 16940 11756 16949
rect 13544 16940 13596 16992
rect 13912 16983 13964 16992
rect 13912 16949 13921 16983
rect 13921 16949 13955 16983
rect 13955 16949 13964 16983
rect 13912 16940 13964 16949
rect 14280 16940 14332 16992
rect 15568 16940 15620 16992
rect 15936 16940 15988 16992
rect 16672 16940 16724 16992
rect 17868 16940 17920 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 2780 16736 2832 16788
rect 3516 16779 3568 16788
rect 3516 16745 3525 16779
rect 3525 16745 3559 16779
rect 3559 16745 3568 16779
rect 3516 16736 3568 16745
rect 4896 16779 4948 16788
rect 4896 16745 4905 16779
rect 4905 16745 4939 16779
rect 4939 16745 4948 16779
rect 4896 16736 4948 16745
rect 7288 16736 7340 16788
rect 9772 16736 9824 16788
rect 10048 16736 10100 16788
rect 10876 16779 10928 16788
rect 10876 16745 10885 16779
rect 10885 16745 10919 16779
rect 10919 16745 10928 16779
rect 10876 16736 10928 16745
rect 11152 16779 11204 16788
rect 11152 16745 11161 16779
rect 11161 16745 11195 16779
rect 11195 16745 11204 16779
rect 11152 16736 11204 16745
rect 12624 16779 12676 16788
rect 12624 16745 12633 16779
rect 12633 16745 12667 16779
rect 12667 16745 12676 16779
rect 12624 16736 12676 16745
rect 13544 16736 13596 16788
rect 14832 16736 14884 16788
rect 15844 16736 15896 16788
rect 17132 16736 17184 16788
rect 17684 16736 17736 16788
rect 5356 16668 5408 16720
rect 1492 16643 1544 16652
rect 1492 16609 1501 16643
rect 1501 16609 1535 16643
rect 1535 16609 1544 16643
rect 1492 16600 1544 16609
rect 2504 16600 2556 16652
rect 3056 16600 3108 16652
rect 3792 16600 3844 16652
rect 5080 16600 5132 16652
rect 6828 16668 6880 16720
rect 7012 16668 7064 16720
rect 8300 16711 8352 16720
rect 8300 16677 8309 16711
rect 8309 16677 8343 16711
rect 8343 16677 8352 16711
rect 8300 16668 8352 16677
rect 8760 16668 8812 16720
rect 12440 16668 12492 16720
rect 5816 16643 5868 16652
rect 5816 16609 5825 16643
rect 5825 16609 5859 16643
rect 5859 16609 5868 16643
rect 5816 16600 5868 16609
rect 6644 16600 6696 16652
rect 8944 16643 8996 16652
rect 8944 16609 8953 16643
rect 8953 16609 8987 16643
rect 8987 16609 8996 16643
rect 8944 16600 8996 16609
rect 10048 16600 10100 16652
rect 11520 16643 11572 16652
rect 11520 16609 11529 16643
rect 11529 16609 11563 16643
rect 11563 16609 11572 16643
rect 11520 16600 11572 16609
rect 11612 16643 11664 16652
rect 11612 16609 11621 16643
rect 11621 16609 11655 16643
rect 11655 16609 11664 16643
rect 11612 16600 11664 16609
rect 12808 16600 12860 16652
rect 13544 16600 13596 16652
rect 14004 16643 14056 16652
rect 14004 16609 14013 16643
rect 14013 16609 14047 16643
rect 14047 16609 14056 16643
rect 14004 16600 14056 16609
rect 6092 16575 6144 16584
rect 6092 16541 6101 16575
rect 6101 16541 6135 16575
rect 6135 16541 6144 16575
rect 6092 16532 6144 16541
rect 8484 16575 8536 16584
rect 8484 16541 8493 16575
rect 8493 16541 8527 16575
rect 8527 16541 8536 16575
rect 8484 16532 8536 16541
rect 9772 16532 9824 16584
rect 11888 16532 11940 16584
rect 13176 16532 13228 16584
rect 14648 16668 14700 16720
rect 14924 16668 14976 16720
rect 15292 16668 15344 16720
rect 14372 16600 14424 16652
rect 6276 16464 6328 16516
rect 15568 16532 15620 16584
rect 17316 16575 17368 16584
rect 17316 16541 17325 16575
rect 17325 16541 17359 16575
rect 17359 16541 17368 16575
rect 17316 16532 17368 16541
rect 17500 16575 17552 16584
rect 17500 16541 17509 16575
rect 17509 16541 17543 16575
rect 17543 16541 17552 16575
rect 17500 16532 17552 16541
rect 3056 16396 3108 16448
rect 6460 16396 6512 16448
rect 7840 16439 7892 16448
rect 7840 16405 7849 16439
rect 7849 16405 7883 16439
rect 7883 16405 7892 16439
rect 7840 16396 7892 16405
rect 13084 16396 13136 16448
rect 14280 16396 14332 16448
rect 14740 16396 14792 16448
rect 16488 16439 16540 16448
rect 16488 16405 16497 16439
rect 16497 16405 16531 16439
rect 16531 16405 16540 16439
rect 16488 16396 16540 16405
rect 16948 16396 17000 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 4620 16235 4672 16244
rect 4620 16201 4629 16235
rect 4629 16201 4663 16235
rect 4663 16201 4672 16235
rect 4620 16192 4672 16201
rect 7012 16235 7064 16244
rect 7012 16201 7021 16235
rect 7021 16201 7055 16235
rect 7055 16201 7064 16235
rect 7012 16192 7064 16201
rect 7564 16192 7616 16244
rect 9772 16192 9824 16244
rect 10968 16192 11020 16244
rect 11520 16192 11572 16244
rect 13176 16235 13228 16244
rect 13176 16201 13185 16235
rect 13185 16201 13219 16235
rect 13219 16201 13228 16235
rect 13176 16192 13228 16201
rect 13636 16235 13688 16244
rect 13636 16201 13645 16235
rect 13645 16201 13679 16235
rect 13679 16201 13688 16235
rect 13636 16192 13688 16201
rect 4068 16124 4120 16176
rect 11152 16124 11204 16176
rect 1768 16056 1820 16108
rect 4252 16099 4304 16108
rect 4252 16065 4261 16099
rect 4261 16065 4295 16099
rect 4295 16065 4304 16099
rect 4252 16056 4304 16065
rect 6460 16056 6512 16108
rect 7564 16099 7616 16108
rect 7564 16065 7573 16099
rect 7573 16065 7607 16099
rect 7607 16065 7616 16099
rect 7564 16056 7616 16065
rect 9220 16099 9272 16108
rect 9220 16065 9229 16099
rect 9229 16065 9263 16099
rect 9263 16065 9272 16099
rect 9220 16056 9272 16065
rect 10784 16056 10836 16108
rect 11244 16099 11296 16108
rect 11244 16065 11253 16099
rect 11253 16065 11287 16099
rect 11287 16065 11296 16099
rect 11244 16056 11296 16065
rect 12624 16124 12676 16176
rect 2412 16031 2464 16040
rect 2412 15997 2421 16031
rect 2421 15997 2455 16031
rect 2455 15997 2464 16031
rect 2412 15988 2464 15997
rect 3608 15988 3660 16040
rect 4160 15988 4212 16040
rect 16764 16192 16816 16244
rect 17132 16235 17184 16244
rect 17132 16201 17141 16235
rect 17141 16201 17175 16235
rect 17175 16201 17184 16235
rect 17132 16192 17184 16201
rect 13912 16056 13964 16108
rect 14096 16031 14148 16040
rect 14096 15997 14105 16031
rect 14105 15997 14139 16031
rect 14139 15997 14148 16031
rect 14096 15988 14148 15997
rect 2320 15920 2372 15972
rect 2504 15963 2556 15972
rect 2504 15929 2513 15963
rect 2513 15929 2547 15963
rect 2547 15929 2556 15963
rect 2504 15920 2556 15929
rect 4436 15920 4488 15972
rect 4896 15920 4948 15972
rect 2044 15895 2096 15904
rect 2044 15861 2053 15895
rect 2053 15861 2087 15895
rect 2087 15861 2096 15895
rect 2044 15852 2096 15861
rect 3884 15852 3936 15904
rect 4712 15852 4764 15904
rect 11520 15920 11572 15972
rect 13544 15920 13596 15972
rect 16396 15988 16448 16040
rect 15844 15920 15896 15972
rect 5172 15895 5224 15904
rect 5172 15861 5181 15895
rect 5181 15861 5215 15895
rect 5215 15861 5224 15895
rect 5172 15852 5224 15861
rect 5356 15852 5408 15904
rect 6276 15895 6328 15904
rect 6276 15861 6285 15895
rect 6285 15861 6319 15895
rect 6319 15861 6328 15895
rect 6276 15852 6328 15861
rect 6736 15852 6788 15904
rect 6920 15852 6972 15904
rect 9128 15852 9180 15904
rect 9772 15852 9824 15904
rect 10048 15852 10100 15904
rect 12624 15852 12676 15904
rect 14740 15895 14792 15904
rect 14740 15861 14749 15895
rect 14749 15861 14783 15895
rect 14783 15861 14792 15895
rect 14740 15852 14792 15861
rect 15292 15852 15344 15904
rect 17500 15920 17552 15972
rect 17868 15852 17920 15904
rect 17960 15852 18012 15904
rect 18696 15852 18748 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 1768 15691 1820 15700
rect 1768 15657 1777 15691
rect 1777 15657 1811 15691
rect 1811 15657 1820 15691
rect 1768 15648 1820 15657
rect 2412 15648 2464 15700
rect 4160 15648 4212 15700
rect 4436 15691 4488 15700
rect 4436 15657 4445 15691
rect 4445 15657 4479 15691
rect 4479 15657 4488 15691
rect 4436 15648 4488 15657
rect 5448 15648 5500 15700
rect 6000 15648 6052 15700
rect 6920 15648 6972 15700
rect 7748 15691 7800 15700
rect 7748 15657 7757 15691
rect 7757 15657 7791 15691
rect 7791 15657 7800 15691
rect 7748 15648 7800 15657
rect 7840 15648 7892 15700
rect 9680 15691 9732 15700
rect 9680 15657 9689 15691
rect 9689 15657 9723 15691
rect 9723 15657 9732 15691
rect 9680 15648 9732 15657
rect 10784 15691 10836 15700
rect 10784 15657 10793 15691
rect 10793 15657 10827 15691
rect 10827 15657 10836 15691
rect 10784 15648 10836 15657
rect 11152 15691 11204 15700
rect 11152 15657 11161 15691
rect 11161 15657 11195 15691
rect 11195 15657 11204 15691
rect 11152 15648 11204 15657
rect 11612 15648 11664 15700
rect 12440 15691 12492 15700
rect 12440 15657 12449 15691
rect 12449 15657 12483 15691
rect 12483 15657 12492 15691
rect 12440 15648 12492 15657
rect 12624 15648 12676 15700
rect 13176 15648 13228 15700
rect 13452 15691 13504 15700
rect 13452 15657 13461 15691
rect 13461 15657 13495 15691
rect 13495 15657 13504 15691
rect 13452 15648 13504 15657
rect 14096 15691 14148 15700
rect 14096 15657 14105 15691
rect 14105 15657 14139 15691
rect 14139 15657 14148 15691
rect 14096 15648 14148 15657
rect 14832 15648 14884 15700
rect 15568 15691 15620 15700
rect 15568 15657 15577 15691
rect 15577 15657 15611 15691
rect 15611 15657 15620 15691
rect 15568 15648 15620 15657
rect 15844 15691 15896 15700
rect 15844 15657 15853 15691
rect 15853 15657 15887 15691
rect 15887 15657 15896 15691
rect 15844 15648 15896 15657
rect 18512 15691 18564 15700
rect 18512 15657 18521 15691
rect 18521 15657 18555 15691
rect 18555 15657 18564 15691
rect 18512 15648 18564 15657
rect 3148 15580 3200 15632
rect 5356 15580 5408 15632
rect 12808 15623 12860 15632
rect 12808 15589 12817 15623
rect 12817 15589 12851 15623
rect 12851 15589 12860 15623
rect 12808 15580 12860 15589
rect 16304 15580 16356 15632
rect 16948 15623 17000 15632
rect 16948 15589 16957 15623
rect 16957 15589 16991 15623
rect 16991 15589 17000 15623
rect 16948 15580 17000 15589
rect 17316 15580 17368 15632
rect 17960 15580 18012 15632
rect 3240 15512 3292 15564
rect 4528 15555 4580 15564
rect 4528 15521 4537 15555
rect 4537 15521 4571 15555
rect 4571 15521 4580 15555
rect 4528 15512 4580 15521
rect 5448 15512 5500 15564
rect 6460 15512 6512 15564
rect 6920 15512 6972 15564
rect 8208 15512 8260 15564
rect 10140 15512 10192 15564
rect 11428 15512 11480 15564
rect 11704 15512 11756 15564
rect 12716 15512 12768 15564
rect 18052 15512 18104 15564
rect 18236 15512 18288 15564
rect 3056 15487 3108 15496
rect 1952 15376 2004 15428
rect 3056 15453 3065 15487
rect 3065 15453 3099 15487
rect 3099 15453 3108 15487
rect 3056 15444 3108 15453
rect 4436 15444 4488 15496
rect 6000 15487 6052 15496
rect 6000 15453 6009 15487
rect 6009 15453 6043 15487
rect 6043 15453 6052 15487
rect 6000 15444 6052 15453
rect 6184 15444 6236 15496
rect 8116 15376 8168 15428
rect 10784 15444 10836 15496
rect 11152 15444 11204 15496
rect 11980 15487 12032 15496
rect 11980 15453 11989 15487
rect 11989 15453 12023 15487
rect 12023 15453 12032 15487
rect 11980 15444 12032 15453
rect 13728 15444 13780 15496
rect 17224 15444 17276 15496
rect 16488 15419 16540 15428
rect 16488 15385 16497 15419
rect 16497 15385 16531 15419
rect 16531 15385 16540 15419
rect 16488 15376 16540 15385
rect 3976 15308 4028 15360
rect 6828 15308 6880 15360
rect 7564 15351 7616 15360
rect 7564 15317 7573 15351
rect 7573 15317 7607 15351
rect 7607 15317 7616 15351
rect 7564 15308 7616 15317
rect 9220 15308 9272 15360
rect 9588 15308 9640 15360
rect 14372 15351 14424 15360
rect 14372 15317 14381 15351
rect 14381 15317 14415 15351
rect 14415 15317 14424 15351
rect 14372 15308 14424 15317
rect 17868 15351 17920 15360
rect 17868 15317 17877 15351
rect 17877 15317 17911 15351
rect 17911 15317 17920 15351
rect 17868 15308 17920 15317
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 3240 15104 3292 15156
rect 5356 15104 5408 15156
rect 6920 15104 6972 15156
rect 1492 14968 1544 15020
rect 4160 14968 4212 15020
rect 5172 15011 5224 15020
rect 5172 14977 5181 15011
rect 5181 14977 5215 15011
rect 5215 14977 5224 15011
rect 5172 14968 5224 14977
rect 8484 15104 8536 15156
rect 10784 15147 10836 15156
rect 10784 15113 10793 15147
rect 10793 15113 10827 15147
rect 10827 15113 10836 15147
rect 10784 15104 10836 15113
rect 11704 15104 11756 15156
rect 11888 15104 11940 15156
rect 11980 15104 12032 15156
rect 13636 15104 13688 15156
rect 14740 15104 14792 15156
rect 16120 15104 16172 15156
rect 17500 15147 17552 15156
rect 17500 15113 17509 15147
rect 17509 15113 17543 15147
rect 17543 15113 17552 15147
rect 17500 15104 17552 15113
rect 17960 15104 18012 15156
rect 12624 15036 12676 15088
rect 13176 15036 13228 15088
rect 16304 15036 16356 15088
rect 17592 15036 17644 15088
rect 18052 15036 18104 15088
rect 2136 14832 2188 14884
rect 5080 14875 5132 14884
rect 5080 14841 5089 14875
rect 5089 14841 5123 14875
rect 5123 14841 5132 14875
rect 5080 14832 5132 14841
rect 3056 14807 3108 14816
rect 3056 14773 3065 14807
rect 3065 14773 3099 14807
rect 3099 14773 3108 14807
rect 3056 14764 3108 14773
rect 3792 14807 3844 14816
rect 3792 14773 3801 14807
rect 3801 14773 3835 14807
rect 3835 14773 3844 14807
rect 3792 14764 3844 14773
rect 4436 14764 4488 14816
rect 16580 14968 16632 15020
rect 6920 14900 6972 14952
rect 8760 14943 8812 14952
rect 8760 14909 8769 14943
rect 8769 14909 8803 14943
rect 8803 14909 8812 14943
rect 8760 14900 8812 14909
rect 12440 14900 12492 14952
rect 13084 14900 13136 14952
rect 13912 14943 13964 14952
rect 13912 14909 13946 14943
rect 13946 14909 13964 14943
rect 13912 14900 13964 14909
rect 14372 14900 14424 14952
rect 7104 14832 7156 14884
rect 8116 14832 8168 14884
rect 8944 14832 8996 14884
rect 18696 14900 18748 14952
rect 18328 14875 18380 14884
rect 18328 14841 18340 14875
rect 18340 14841 18380 14875
rect 18328 14832 18380 14841
rect 6184 14807 6236 14816
rect 6184 14773 6193 14807
rect 6193 14773 6227 14807
rect 6227 14773 6236 14807
rect 6184 14764 6236 14773
rect 6460 14764 6512 14816
rect 8300 14764 8352 14816
rect 9588 14764 9640 14816
rect 10048 14764 10100 14816
rect 11060 14807 11112 14816
rect 11060 14773 11069 14807
rect 11069 14773 11103 14807
rect 11103 14773 11112 14807
rect 11060 14764 11112 14773
rect 11428 14807 11480 14816
rect 11428 14773 11437 14807
rect 11437 14773 11471 14807
rect 11471 14773 11480 14807
rect 11428 14764 11480 14773
rect 12716 14764 12768 14816
rect 13360 14764 13412 14816
rect 15384 14764 15436 14816
rect 16764 14807 16816 14816
rect 16764 14773 16773 14807
rect 16773 14773 16807 14807
rect 16807 14773 16816 14807
rect 16764 14764 16816 14773
rect 19432 14807 19484 14816
rect 19432 14773 19441 14807
rect 19441 14773 19475 14807
rect 19475 14773 19484 14807
rect 19432 14764 19484 14773
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 1676 14560 1728 14612
rect 2412 14603 2464 14612
rect 2412 14569 2421 14603
rect 2421 14569 2455 14603
rect 2455 14569 2464 14603
rect 2412 14560 2464 14569
rect 3056 14560 3108 14612
rect 5448 14560 5500 14612
rect 6920 14560 6972 14612
rect 11152 14560 11204 14612
rect 12992 14560 13044 14612
rect 14188 14560 14240 14612
rect 18328 14603 18380 14612
rect 18328 14569 18337 14603
rect 18337 14569 18371 14603
rect 18371 14569 18380 14603
rect 18328 14560 18380 14569
rect 3148 14492 3200 14544
rect 3332 14492 3384 14544
rect 5540 14492 5592 14544
rect 7104 14492 7156 14544
rect 7564 14492 7616 14544
rect 8208 14492 8260 14544
rect 9956 14492 10008 14544
rect 12532 14492 12584 14544
rect 14556 14492 14608 14544
rect 15660 14535 15712 14544
rect 15660 14501 15669 14535
rect 15669 14501 15703 14535
rect 15703 14501 15712 14535
rect 15660 14492 15712 14501
rect 2780 14467 2832 14476
rect 2780 14433 2789 14467
rect 2789 14433 2823 14467
rect 2823 14433 2832 14467
rect 2780 14424 2832 14433
rect 4252 14424 4304 14476
rect 6552 14424 6604 14476
rect 4160 14399 4212 14408
rect 4160 14365 4169 14399
rect 4169 14365 4203 14399
rect 4203 14365 4212 14399
rect 4160 14356 4212 14365
rect 2136 14288 2188 14340
rect 3792 14288 3844 14340
rect 1768 14220 1820 14272
rect 11060 14424 11112 14476
rect 12348 14424 12400 14476
rect 15752 14467 15804 14476
rect 15752 14433 15761 14467
rect 15761 14433 15795 14467
rect 15795 14433 15804 14467
rect 15752 14424 15804 14433
rect 17224 14467 17276 14476
rect 17224 14433 17258 14467
rect 17258 14433 17276 14467
rect 17224 14424 17276 14433
rect 11520 14399 11572 14408
rect 11520 14365 11529 14399
rect 11529 14365 11563 14399
rect 11563 14365 11572 14399
rect 11520 14356 11572 14365
rect 11704 14399 11756 14408
rect 11704 14365 11713 14399
rect 11713 14365 11747 14399
rect 11747 14365 11756 14399
rect 11704 14356 11756 14365
rect 14280 14399 14332 14408
rect 14280 14365 14289 14399
rect 14289 14365 14323 14399
rect 14323 14365 14332 14399
rect 14280 14356 14332 14365
rect 14556 14356 14608 14408
rect 15936 14399 15988 14408
rect 15936 14365 15945 14399
rect 15945 14365 15979 14399
rect 15979 14365 15988 14399
rect 15936 14356 15988 14365
rect 7748 14288 7800 14340
rect 8484 14288 8536 14340
rect 9772 14288 9824 14340
rect 13176 14331 13228 14340
rect 13176 14297 13185 14331
rect 13185 14297 13219 14331
rect 13219 14297 13228 14331
rect 13176 14288 13228 14297
rect 8208 14220 8260 14272
rect 8300 14220 8352 14272
rect 9404 14220 9456 14272
rect 12072 14263 12124 14272
rect 12072 14229 12081 14263
rect 12081 14229 12115 14263
rect 12115 14229 12124 14263
rect 12072 14220 12124 14229
rect 12440 14263 12492 14272
rect 12440 14229 12449 14263
rect 12449 14229 12483 14263
rect 12483 14229 12492 14263
rect 12440 14220 12492 14229
rect 15384 14220 15436 14272
rect 16488 14220 16540 14272
rect 18696 14220 18748 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 1400 14059 1452 14068
rect 1400 14025 1409 14059
rect 1409 14025 1443 14059
rect 1443 14025 1452 14059
rect 1400 14016 1452 14025
rect 3148 14016 3200 14068
rect 4344 14016 4396 14068
rect 2780 13991 2832 14000
rect 2780 13957 2789 13991
rect 2789 13957 2823 13991
rect 2823 13957 2832 13991
rect 5172 14016 5224 14068
rect 6092 14016 6144 14068
rect 7748 14016 7800 14068
rect 8944 14059 8996 14068
rect 8944 14025 8953 14059
rect 8953 14025 8987 14059
rect 8987 14025 8996 14059
rect 8944 14016 8996 14025
rect 9772 14059 9824 14068
rect 9772 14025 9781 14059
rect 9781 14025 9815 14059
rect 9815 14025 9824 14059
rect 9772 14016 9824 14025
rect 11060 14016 11112 14068
rect 11704 14016 11756 14068
rect 13912 14016 13964 14068
rect 14188 14016 14240 14068
rect 14372 14059 14424 14068
rect 14372 14025 14381 14059
rect 14381 14025 14415 14059
rect 14415 14025 14424 14059
rect 14372 14016 14424 14025
rect 15752 14016 15804 14068
rect 16764 14016 16816 14068
rect 17960 14016 18012 14068
rect 25504 14059 25556 14068
rect 25504 14025 25513 14059
rect 25513 14025 25547 14059
rect 25547 14025 25556 14059
rect 25504 14016 25556 14025
rect 2780 13948 2832 13957
rect 2136 13880 2188 13932
rect 6552 13948 6604 14000
rect 15660 13948 15712 14000
rect 2964 13855 3016 13864
rect 2964 13821 2973 13855
rect 2973 13821 3007 13855
rect 3007 13821 3016 13855
rect 2964 13812 3016 13821
rect 3240 13855 3292 13864
rect 3240 13821 3249 13855
rect 3249 13821 3283 13855
rect 3283 13821 3292 13855
rect 3240 13812 3292 13821
rect 6092 13880 6144 13932
rect 11980 13880 12032 13932
rect 5080 13812 5132 13864
rect 7104 13855 7156 13864
rect 7104 13821 7113 13855
rect 7113 13821 7147 13855
rect 7147 13821 7156 13855
rect 7104 13812 7156 13821
rect 7840 13855 7892 13864
rect 1768 13719 1820 13728
rect 1768 13685 1777 13719
rect 1777 13685 1811 13719
rect 1811 13685 1820 13719
rect 1768 13676 1820 13685
rect 2320 13676 2372 13728
rect 3516 13676 3568 13728
rect 7380 13744 7432 13796
rect 7840 13821 7874 13855
rect 7874 13821 7892 13855
rect 7840 13812 7892 13821
rect 8760 13812 8812 13864
rect 9220 13812 9272 13864
rect 10692 13855 10744 13864
rect 10692 13821 10701 13855
rect 10701 13821 10735 13855
rect 10735 13821 10744 13855
rect 11244 13855 11296 13864
rect 10692 13812 10744 13821
rect 11244 13821 11253 13855
rect 11253 13821 11287 13855
rect 11287 13821 11296 13855
rect 11244 13812 11296 13821
rect 12440 13855 12492 13864
rect 12440 13821 12449 13855
rect 12449 13821 12483 13855
rect 12483 13821 12492 13855
rect 12440 13812 12492 13821
rect 15476 13880 15528 13932
rect 15936 13880 15988 13932
rect 16764 13923 16816 13932
rect 16764 13889 16773 13923
rect 16773 13889 16807 13923
rect 16807 13889 16816 13923
rect 16764 13880 16816 13889
rect 13728 13812 13780 13864
rect 17224 13812 17276 13864
rect 11152 13787 11204 13796
rect 11152 13753 11161 13787
rect 11161 13753 11195 13787
rect 11195 13753 11204 13787
rect 11152 13744 11204 13753
rect 14188 13744 14240 13796
rect 16028 13744 16080 13796
rect 18696 13855 18748 13864
rect 18696 13821 18705 13855
rect 18705 13821 18739 13855
rect 18739 13821 18748 13855
rect 18696 13812 18748 13821
rect 24124 13855 24176 13864
rect 24124 13821 24133 13855
rect 24133 13821 24167 13855
rect 24167 13821 24176 13855
rect 24124 13812 24176 13821
rect 24400 13855 24452 13864
rect 24400 13821 24434 13855
rect 24434 13821 24452 13855
rect 24400 13812 24452 13821
rect 18512 13744 18564 13796
rect 4252 13719 4304 13728
rect 4252 13685 4261 13719
rect 4261 13685 4295 13719
rect 4295 13685 4304 13719
rect 4252 13676 4304 13685
rect 10968 13676 11020 13728
rect 11796 13676 11848 13728
rect 14004 13676 14056 13728
rect 17224 13676 17276 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 2412 13515 2464 13524
rect 2412 13481 2421 13515
rect 2421 13481 2455 13515
rect 2455 13481 2464 13515
rect 2412 13472 2464 13481
rect 3792 13472 3844 13524
rect 5540 13515 5592 13524
rect 5540 13481 5549 13515
rect 5549 13481 5583 13515
rect 5583 13481 5592 13515
rect 5540 13472 5592 13481
rect 8024 13472 8076 13524
rect 8300 13472 8352 13524
rect 9220 13515 9272 13524
rect 9220 13481 9229 13515
rect 9229 13481 9263 13515
rect 9263 13481 9272 13515
rect 9220 13472 9272 13481
rect 11520 13472 11572 13524
rect 12072 13515 12124 13524
rect 12072 13481 12081 13515
rect 12081 13481 12115 13515
rect 12115 13481 12124 13515
rect 12072 13472 12124 13481
rect 13268 13472 13320 13524
rect 14280 13515 14332 13524
rect 14280 13481 14289 13515
rect 14289 13481 14323 13515
rect 14323 13481 14332 13515
rect 14280 13472 14332 13481
rect 15476 13472 15528 13524
rect 16672 13515 16724 13524
rect 16672 13481 16681 13515
rect 16681 13481 16715 13515
rect 16715 13481 16724 13515
rect 16672 13472 16724 13481
rect 24124 13515 24176 13524
rect 24124 13481 24133 13515
rect 24133 13481 24167 13515
rect 24167 13481 24176 13515
rect 24124 13472 24176 13481
rect 3976 13404 4028 13456
rect 5356 13404 5408 13456
rect 2044 13379 2096 13388
rect 2044 13345 2053 13379
rect 2053 13345 2087 13379
rect 2087 13345 2096 13379
rect 2044 13336 2096 13345
rect 2964 13311 3016 13320
rect 2964 13277 2973 13311
rect 2973 13277 3007 13311
rect 3007 13277 3016 13311
rect 2964 13268 3016 13277
rect 4252 13336 4304 13388
rect 4528 13379 4580 13388
rect 4528 13345 4537 13379
rect 4537 13345 4571 13379
rect 4571 13345 4580 13379
rect 5632 13379 5684 13388
rect 4528 13336 4580 13345
rect 5632 13345 5641 13379
rect 5641 13345 5675 13379
rect 5675 13345 5684 13379
rect 5632 13336 5684 13345
rect 6184 13336 6236 13388
rect 7104 13336 7156 13388
rect 12164 13404 12216 13456
rect 12440 13404 12492 13456
rect 9956 13379 10008 13388
rect 9956 13345 9990 13379
rect 9990 13345 10008 13379
rect 9956 13336 10008 13345
rect 12808 13379 12860 13388
rect 12808 13345 12817 13379
rect 12817 13345 12851 13379
rect 12851 13345 12860 13379
rect 12808 13336 12860 13345
rect 16488 13404 16540 13456
rect 15568 13379 15620 13388
rect 15568 13345 15602 13379
rect 15602 13345 15620 13379
rect 15568 13336 15620 13345
rect 17500 13336 17552 13388
rect 4620 13311 4672 13320
rect 4620 13277 4629 13311
rect 4629 13277 4663 13311
rect 4663 13277 4672 13311
rect 4620 13268 4672 13277
rect 7564 13311 7616 13320
rect 7564 13277 7573 13311
rect 7573 13277 7607 13311
rect 7607 13277 7616 13311
rect 7564 13268 7616 13277
rect 7656 13311 7708 13320
rect 7656 13277 7665 13311
rect 7665 13277 7699 13311
rect 7699 13277 7708 13311
rect 18236 13311 18288 13320
rect 7656 13268 7708 13277
rect 18236 13277 18245 13311
rect 18245 13277 18279 13311
rect 18279 13277 18288 13311
rect 18236 13268 18288 13277
rect 18328 13311 18380 13320
rect 18328 13277 18337 13311
rect 18337 13277 18371 13311
rect 18371 13277 18380 13311
rect 18328 13268 18380 13277
rect 5816 13243 5868 13252
rect 5816 13209 5825 13243
rect 5825 13209 5859 13243
rect 5859 13209 5868 13243
rect 5816 13200 5868 13209
rect 2320 13132 2372 13184
rect 6552 13175 6604 13184
rect 6552 13141 6561 13175
rect 6561 13141 6595 13175
rect 6595 13141 6604 13175
rect 6552 13132 6604 13141
rect 7104 13132 7156 13184
rect 8116 13175 8168 13184
rect 8116 13141 8125 13175
rect 8125 13141 8159 13175
rect 8159 13141 8168 13175
rect 8116 13132 8168 13141
rect 11060 13175 11112 13184
rect 11060 13141 11069 13175
rect 11069 13141 11103 13175
rect 11103 13141 11112 13175
rect 11060 13132 11112 13141
rect 12440 13175 12492 13184
rect 12440 13141 12449 13175
rect 12449 13141 12483 13175
rect 12483 13141 12492 13175
rect 12440 13132 12492 13141
rect 15292 13132 15344 13184
rect 15660 13132 15712 13184
rect 17224 13175 17276 13184
rect 17224 13141 17233 13175
rect 17233 13141 17267 13175
rect 17267 13141 17276 13175
rect 17224 13132 17276 13141
rect 18788 13175 18840 13184
rect 18788 13141 18797 13175
rect 18797 13141 18831 13175
rect 18831 13141 18840 13175
rect 18788 13132 18840 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 1400 12971 1452 12980
rect 1400 12937 1409 12971
rect 1409 12937 1443 12971
rect 1443 12937 1452 12971
rect 1400 12928 1452 12937
rect 2596 12928 2648 12980
rect 2964 12928 3016 12980
rect 4528 12928 4580 12980
rect 6184 12971 6236 12980
rect 6184 12937 6193 12971
rect 6193 12937 6227 12971
rect 6227 12937 6236 12971
rect 6184 12928 6236 12937
rect 7564 12928 7616 12980
rect 7656 12928 7708 12980
rect 9956 12928 10008 12980
rect 12808 12928 12860 12980
rect 13636 12928 13688 12980
rect 13820 12971 13872 12980
rect 13820 12937 13829 12971
rect 13829 12937 13863 12971
rect 13863 12937 13872 12971
rect 13820 12928 13872 12937
rect 17500 12971 17552 12980
rect 17500 12937 17509 12971
rect 17509 12937 17543 12971
rect 17543 12937 17552 12971
rect 17500 12928 17552 12937
rect 17960 12928 18012 12980
rect 12440 12860 12492 12912
rect 2044 12656 2096 12708
rect 6460 12792 6512 12844
rect 7656 12792 7708 12844
rect 8116 12835 8168 12844
rect 8116 12801 8125 12835
rect 8125 12801 8159 12835
rect 8159 12801 8168 12835
rect 8116 12792 8168 12801
rect 11060 12792 11112 12844
rect 3056 12724 3108 12776
rect 4160 12724 4212 12776
rect 5448 12724 5500 12776
rect 10876 12724 10928 12776
rect 12164 12724 12216 12776
rect 18604 12835 18656 12844
rect 18604 12801 18613 12835
rect 18613 12801 18647 12835
rect 18647 12801 18656 12835
rect 18604 12792 18656 12801
rect 8024 12699 8076 12708
rect 8024 12665 8033 12699
rect 8033 12665 8067 12699
rect 8067 12665 8076 12699
rect 8024 12656 8076 12665
rect 10968 12656 11020 12708
rect 15752 12724 15804 12776
rect 17224 12724 17276 12776
rect 18788 12724 18840 12776
rect 14648 12656 14700 12708
rect 16764 12656 16816 12708
rect 18236 12656 18288 12708
rect 3516 12588 3568 12640
rect 4344 12631 4396 12640
rect 4344 12597 4353 12631
rect 4353 12597 4387 12631
rect 4387 12597 4396 12631
rect 4344 12588 4396 12597
rect 4620 12588 4672 12640
rect 7012 12631 7064 12640
rect 7012 12597 7021 12631
rect 7021 12597 7055 12631
rect 7055 12597 7064 12631
rect 7012 12588 7064 12597
rect 11060 12588 11112 12640
rect 11888 12631 11940 12640
rect 11888 12597 11897 12631
rect 11897 12597 11931 12631
rect 11931 12597 11940 12631
rect 11888 12588 11940 12597
rect 13268 12588 13320 12640
rect 15016 12588 15068 12640
rect 15200 12588 15252 12640
rect 15568 12631 15620 12640
rect 15568 12597 15577 12631
rect 15577 12597 15611 12631
rect 15611 12597 15620 12631
rect 15568 12588 15620 12597
rect 16856 12588 16908 12640
rect 17868 12588 17920 12640
rect 18328 12588 18380 12640
rect 18420 12588 18472 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 2872 12427 2924 12436
rect 2872 12393 2881 12427
rect 2881 12393 2915 12427
rect 2915 12393 2924 12427
rect 2872 12384 2924 12393
rect 3976 12384 4028 12436
rect 5448 12427 5500 12436
rect 5448 12393 5457 12427
rect 5457 12393 5491 12427
rect 5491 12393 5500 12427
rect 6092 12427 6144 12436
rect 5448 12384 5500 12393
rect 6092 12393 6101 12427
rect 6101 12393 6135 12427
rect 6135 12393 6144 12427
rect 6092 12384 6144 12393
rect 6552 12384 6604 12436
rect 7104 12384 7156 12436
rect 9680 12427 9732 12436
rect 9680 12393 9689 12427
rect 9689 12393 9723 12427
rect 9723 12393 9732 12427
rect 9680 12384 9732 12393
rect 11152 12427 11204 12436
rect 11152 12393 11161 12427
rect 11161 12393 11195 12427
rect 11195 12393 11204 12427
rect 11152 12384 11204 12393
rect 11520 12384 11572 12436
rect 12900 12427 12952 12436
rect 12900 12393 12909 12427
rect 12909 12393 12943 12427
rect 12943 12393 12952 12427
rect 12900 12384 12952 12393
rect 13544 12384 13596 12436
rect 14004 12384 14056 12436
rect 14648 12427 14700 12436
rect 2044 12316 2096 12368
rect 3056 12316 3108 12368
rect 3332 12316 3384 12368
rect 8852 12316 8904 12368
rect 1768 12291 1820 12300
rect 1768 12257 1802 12291
rect 1802 12257 1820 12291
rect 1768 12248 1820 12257
rect 4252 12248 4304 12300
rect 4436 12291 4488 12300
rect 4436 12257 4445 12291
rect 4445 12257 4479 12291
rect 4479 12257 4488 12291
rect 4436 12248 4488 12257
rect 7012 12248 7064 12300
rect 7380 12291 7432 12300
rect 7380 12257 7389 12291
rect 7389 12257 7423 12291
rect 7423 12257 7432 12291
rect 7380 12248 7432 12257
rect 10048 12291 10100 12300
rect 10048 12257 10057 12291
rect 10057 12257 10091 12291
rect 10091 12257 10100 12291
rect 10048 12248 10100 12257
rect 12072 12248 12124 12300
rect 14004 12291 14056 12300
rect 14004 12257 14013 12291
rect 14013 12257 14047 12291
rect 14047 12257 14056 12291
rect 14004 12248 14056 12257
rect 14648 12393 14657 12427
rect 14657 12393 14691 12427
rect 14691 12393 14700 12427
rect 14648 12384 14700 12393
rect 15016 12427 15068 12436
rect 15016 12393 15025 12427
rect 15025 12393 15059 12427
rect 15059 12393 15068 12427
rect 15016 12384 15068 12393
rect 15752 12427 15804 12436
rect 15752 12393 15761 12427
rect 15761 12393 15795 12427
rect 15795 12393 15804 12427
rect 15752 12384 15804 12393
rect 18604 12427 18656 12436
rect 18604 12393 18613 12427
rect 18613 12393 18647 12427
rect 18647 12393 18656 12427
rect 18604 12384 18656 12393
rect 18512 12316 18564 12368
rect 15752 12248 15804 12300
rect 16580 12291 16632 12300
rect 16580 12257 16589 12291
rect 16589 12257 16623 12291
rect 16623 12257 16632 12291
rect 16580 12248 16632 12257
rect 16856 12291 16908 12300
rect 16856 12257 16890 12291
rect 16890 12257 16908 12291
rect 16856 12248 16908 12257
rect 4528 12223 4580 12232
rect 4528 12189 4537 12223
rect 4537 12189 4571 12223
rect 4571 12189 4580 12223
rect 4528 12180 4580 12189
rect 3792 12112 3844 12164
rect 4344 12112 4396 12164
rect 4896 12180 4948 12232
rect 7196 12180 7248 12232
rect 6276 12112 6328 12164
rect 8024 12180 8076 12232
rect 9680 12180 9732 12232
rect 10784 12180 10836 12232
rect 11060 12180 11112 12232
rect 11244 12180 11296 12232
rect 11980 12223 12032 12232
rect 11980 12189 11989 12223
rect 11989 12189 12023 12223
rect 12023 12189 12032 12223
rect 11980 12180 12032 12189
rect 14280 12223 14332 12232
rect 14280 12189 14289 12223
rect 14289 12189 14323 12223
rect 14323 12189 14332 12223
rect 14280 12180 14332 12189
rect 14372 12180 14424 12232
rect 14740 12180 14792 12232
rect 3516 12087 3568 12096
rect 3516 12053 3525 12087
rect 3525 12053 3559 12087
rect 3559 12053 3568 12087
rect 3516 12044 3568 12053
rect 5080 12044 5132 12096
rect 6552 12044 6604 12096
rect 7840 12044 7892 12096
rect 8116 12044 8168 12096
rect 8392 12087 8444 12096
rect 8392 12053 8401 12087
rect 8401 12053 8435 12087
rect 8435 12053 8444 12087
rect 8392 12044 8444 12053
rect 10876 12087 10928 12096
rect 10876 12053 10885 12087
rect 10885 12053 10919 12087
rect 10919 12053 10928 12087
rect 10876 12044 10928 12053
rect 13176 12044 13228 12096
rect 14648 12044 14700 12096
rect 14832 12044 14884 12096
rect 16304 12044 16356 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 3516 11840 3568 11892
rect 4436 11840 4488 11892
rect 6276 11883 6328 11892
rect 6276 11849 6285 11883
rect 6285 11849 6319 11883
rect 6319 11849 6328 11883
rect 6276 11840 6328 11849
rect 7380 11840 7432 11892
rect 8116 11840 8168 11892
rect 8576 11840 8628 11892
rect 9680 11883 9732 11892
rect 9680 11849 9689 11883
rect 9689 11849 9723 11883
rect 9723 11849 9732 11883
rect 9680 11840 9732 11849
rect 11980 11840 12032 11892
rect 14280 11840 14332 11892
rect 14648 11883 14700 11892
rect 14648 11849 14657 11883
rect 14657 11849 14691 11883
rect 14691 11849 14700 11883
rect 14648 11840 14700 11849
rect 14832 11840 14884 11892
rect 16120 11883 16172 11892
rect 16120 11849 16129 11883
rect 16129 11849 16163 11883
rect 16163 11849 16172 11883
rect 16120 11840 16172 11849
rect 18512 11883 18564 11892
rect 18512 11849 18521 11883
rect 18521 11849 18555 11883
rect 18555 11849 18564 11883
rect 18512 11840 18564 11849
rect 4988 11772 5040 11824
rect 7196 11772 7248 11824
rect 15292 11772 15344 11824
rect 4344 11704 4396 11756
rect 4620 11704 4672 11756
rect 5080 11747 5132 11756
rect 5080 11713 5089 11747
rect 5089 11713 5123 11747
rect 5123 11713 5132 11747
rect 5080 11704 5132 11713
rect 9496 11704 9548 11756
rect 13268 11747 13320 11756
rect 13268 11713 13284 11747
rect 13284 11713 13318 11747
rect 13318 11713 13320 11747
rect 13268 11704 13320 11713
rect 16856 11704 16908 11756
rect 2044 11679 2096 11688
rect 2044 11645 2053 11679
rect 2053 11645 2087 11679
rect 2087 11645 2096 11679
rect 2044 11636 2096 11645
rect 4896 11679 4948 11688
rect 4896 11645 4905 11679
rect 4905 11645 4939 11679
rect 4939 11645 4948 11679
rect 4896 11636 4948 11645
rect 7380 11636 7432 11688
rect 10048 11636 10100 11688
rect 12072 11636 12124 11688
rect 2412 11568 2464 11620
rect 4620 11568 4672 11620
rect 7840 11568 7892 11620
rect 9864 11568 9916 11620
rect 1400 11500 1452 11552
rect 7288 11500 7340 11552
rect 9312 11500 9364 11552
rect 10692 11500 10744 11552
rect 12348 11568 12400 11620
rect 13544 11611 13596 11620
rect 13544 11577 13578 11611
rect 13578 11577 13596 11611
rect 13544 11568 13596 11577
rect 15936 11611 15988 11620
rect 15936 11577 15945 11611
rect 15945 11577 15979 11611
rect 15979 11577 15988 11611
rect 15936 11568 15988 11577
rect 16396 11568 16448 11620
rect 17960 11568 18012 11620
rect 11888 11500 11940 11552
rect 13636 11500 13688 11552
rect 13912 11500 13964 11552
rect 16304 11500 16356 11552
rect 18052 11543 18104 11552
rect 18052 11509 18061 11543
rect 18061 11509 18095 11543
rect 18095 11509 18104 11543
rect 18052 11500 18104 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 1768 11296 1820 11348
rect 3792 11339 3844 11348
rect 3792 11305 3801 11339
rect 3801 11305 3835 11339
rect 3835 11305 3844 11339
rect 3792 11296 3844 11305
rect 4528 11296 4580 11348
rect 6092 11339 6144 11348
rect 6092 11305 6101 11339
rect 6101 11305 6135 11339
rect 6135 11305 6144 11339
rect 6092 11296 6144 11305
rect 7840 11339 7892 11348
rect 7840 11305 7849 11339
rect 7849 11305 7883 11339
rect 7883 11305 7892 11339
rect 9496 11339 9548 11348
rect 7840 11296 7892 11305
rect 9496 11305 9505 11339
rect 9505 11305 9539 11339
rect 9539 11305 9548 11339
rect 9496 11296 9548 11305
rect 11244 11339 11296 11348
rect 11244 11305 11253 11339
rect 11253 11305 11287 11339
rect 11287 11305 11296 11339
rect 11244 11296 11296 11305
rect 12716 11339 12768 11348
rect 12716 11305 12725 11339
rect 12725 11305 12759 11339
rect 12759 11305 12768 11339
rect 12716 11296 12768 11305
rect 13176 11339 13228 11348
rect 13176 11305 13185 11339
rect 13185 11305 13219 11339
rect 13219 11305 13228 11339
rect 13176 11296 13228 11305
rect 14004 11296 14056 11348
rect 15752 11296 15804 11348
rect 16396 11339 16448 11348
rect 16396 11305 16405 11339
rect 16405 11305 16439 11339
rect 16439 11305 16448 11339
rect 16396 11296 16448 11305
rect 16672 11296 16724 11348
rect 18052 11296 18104 11348
rect 3516 11228 3568 11280
rect 6644 11228 6696 11280
rect 7380 11228 7432 11280
rect 9128 11228 9180 11280
rect 9864 11228 9916 11280
rect 10692 11228 10744 11280
rect 10876 11228 10928 11280
rect 12532 11228 12584 11280
rect 13360 11228 13412 11280
rect 14372 11271 14424 11280
rect 1492 11160 1544 11212
rect 1860 11160 1912 11212
rect 3240 11160 3292 11212
rect 4804 11160 4856 11212
rect 5448 11160 5500 11212
rect 6552 11160 6604 11212
rect 8392 11160 8444 11212
rect 10048 11203 10100 11212
rect 10048 11169 10057 11203
rect 10057 11169 10091 11203
rect 10091 11169 10100 11203
rect 10048 11160 10100 11169
rect 11612 11160 11664 11212
rect 14004 11160 14056 11212
rect 14372 11237 14381 11271
rect 14381 11237 14415 11271
rect 14415 11237 14424 11271
rect 14372 11228 14424 11237
rect 15568 11228 15620 11280
rect 17132 11160 17184 11212
rect 17408 11228 17460 11280
rect 17684 11160 17736 11212
rect 2136 11024 2188 11076
rect 2780 11024 2832 11076
rect 3884 11024 3936 11076
rect 5080 11092 5132 11144
rect 10324 11135 10376 11144
rect 10324 11101 10333 11135
rect 10333 11101 10367 11135
rect 10367 11101 10376 11135
rect 10324 11092 10376 11101
rect 12164 11135 12216 11144
rect 12164 11101 12173 11135
rect 12173 11101 12207 11135
rect 12207 11101 12216 11135
rect 12164 11092 12216 11101
rect 12348 11135 12400 11144
rect 12348 11101 12357 11135
rect 12357 11101 12391 11135
rect 12391 11101 12400 11135
rect 12348 11092 12400 11101
rect 13728 11135 13780 11144
rect 4896 11024 4948 11076
rect 5172 11024 5224 11076
rect 8208 11024 8260 11076
rect 5540 10956 5592 11008
rect 6092 10956 6144 11008
rect 8392 10999 8444 11008
rect 8392 10965 8401 10999
rect 8401 10965 8435 10999
rect 8435 10965 8444 10999
rect 8392 10956 8444 10965
rect 13728 11101 13737 11135
rect 13737 11101 13771 11135
rect 13771 11101 13780 11135
rect 13728 11092 13780 11101
rect 13176 11024 13228 11076
rect 15292 11092 15344 11144
rect 16304 11092 16356 11144
rect 18052 11135 18104 11144
rect 15568 11024 15620 11076
rect 18052 11101 18061 11135
rect 18061 11101 18095 11135
rect 18095 11101 18104 11135
rect 18052 11092 18104 11101
rect 18604 11135 18656 11144
rect 18604 11101 18613 11135
rect 18613 11101 18647 11135
rect 18647 11101 18656 11135
rect 18604 11092 18656 11101
rect 17408 11067 17460 11076
rect 14648 10999 14700 11008
rect 14648 10965 14657 10999
rect 14657 10965 14691 10999
rect 14691 10965 14700 10999
rect 14648 10956 14700 10965
rect 15844 10999 15896 11008
rect 15844 10965 15853 10999
rect 15853 10965 15887 10999
rect 15887 10965 15896 10999
rect 17408 11033 17417 11067
rect 17417 11033 17451 11067
rect 17451 11033 17460 11067
rect 17408 11024 17460 11033
rect 15844 10956 15896 10965
rect 18512 10956 18564 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 2688 10795 2740 10804
rect 2688 10761 2697 10795
rect 2697 10761 2731 10795
rect 2731 10761 2740 10795
rect 2688 10752 2740 10761
rect 5172 10795 5224 10804
rect 5172 10761 5181 10795
rect 5181 10761 5215 10795
rect 5215 10761 5224 10795
rect 5172 10752 5224 10761
rect 5448 10752 5500 10804
rect 7564 10752 7616 10804
rect 10324 10752 10376 10804
rect 10692 10752 10744 10804
rect 11612 10752 11664 10804
rect 11980 10752 12032 10804
rect 14004 10795 14056 10804
rect 14004 10761 14013 10795
rect 14013 10761 14047 10795
rect 14047 10761 14056 10795
rect 14004 10752 14056 10761
rect 14648 10752 14700 10804
rect 16396 10752 16448 10804
rect 17684 10795 17736 10804
rect 17684 10761 17693 10795
rect 17693 10761 17727 10795
rect 17727 10761 17736 10795
rect 17684 10752 17736 10761
rect 5816 10727 5868 10736
rect 5816 10693 5825 10727
rect 5825 10693 5859 10727
rect 5859 10693 5868 10727
rect 5816 10684 5868 10693
rect 13912 10727 13964 10736
rect 13912 10693 13921 10727
rect 13921 10693 13955 10727
rect 13955 10693 13964 10727
rect 13912 10684 13964 10693
rect 2228 10659 2280 10668
rect 2228 10625 2237 10659
rect 2237 10625 2271 10659
rect 2271 10625 2280 10659
rect 2228 10616 2280 10625
rect 8576 10659 8628 10668
rect 8576 10625 8585 10659
rect 8585 10625 8619 10659
rect 8619 10625 8628 10659
rect 8576 10616 8628 10625
rect 2044 10548 2096 10600
rect 2780 10548 2832 10600
rect 5540 10548 5592 10600
rect 9312 10548 9364 10600
rect 12716 10616 12768 10668
rect 12992 10659 13044 10668
rect 12992 10625 13001 10659
rect 13001 10625 13035 10659
rect 13035 10625 13044 10659
rect 13544 10659 13596 10668
rect 12992 10616 13044 10625
rect 13544 10625 13553 10659
rect 13553 10625 13587 10659
rect 13587 10625 13596 10659
rect 14556 10659 14608 10668
rect 13544 10616 13596 10625
rect 14556 10625 14565 10659
rect 14565 10625 14599 10659
rect 14599 10625 14608 10659
rect 14556 10616 14608 10625
rect 16764 10659 16816 10668
rect 16764 10625 16773 10659
rect 16773 10625 16807 10659
rect 16807 10625 16816 10659
rect 16764 10616 16816 10625
rect 16948 10659 17000 10668
rect 16948 10625 16957 10659
rect 16957 10625 16991 10659
rect 16991 10625 17000 10659
rect 16948 10616 17000 10625
rect 18604 10659 18656 10668
rect 18604 10625 18613 10659
rect 18613 10625 18647 10659
rect 18647 10625 18656 10659
rect 18604 10616 18656 10625
rect 9956 10591 10008 10600
rect 9956 10557 9979 10591
rect 9979 10557 10008 10591
rect 2872 10480 2924 10532
rect 3424 10523 3476 10532
rect 3424 10489 3436 10523
rect 3436 10489 3476 10523
rect 6828 10523 6880 10532
rect 3424 10480 3476 10489
rect 6828 10489 6837 10523
rect 6837 10489 6871 10523
rect 6871 10489 6880 10523
rect 6828 10480 6880 10489
rect 9956 10548 10008 10557
rect 14096 10548 14148 10600
rect 14740 10548 14792 10600
rect 16672 10591 16724 10600
rect 16672 10557 16681 10591
rect 16681 10557 16715 10591
rect 16715 10557 16724 10591
rect 16672 10548 16724 10557
rect 18052 10548 18104 10600
rect 10140 10480 10192 10532
rect 11980 10480 12032 10532
rect 13912 10480 13964 10532
rect 1584 10455 1636 10464
rect 1584 10421 1593 10455
rect 1593 10421 1627 10455
rect 1627 10421 1636 10455
rect 1584 10412 1636 10421
rect 1860 10412 1912 10464
rect 2044 10455 2096 10464
rect 2044 10421 2053 10455
rect 2053 10421 2087 10455
rect 2087 10421 2096 10455
rect 2044 10412 2096 10421
rect 3240 10412 3292 10464
rect 4436 10412 4488 10464
rect 6644 10412 6696 10464
rect 7104 10412 7156 10464
rect 8944 10412 8996 10464
rect 12440 10455 12492 10464
rect 12440 10421 12449 10455
rect 12449 10421 12483 10455
rect 12483 10421 12492 10455
rect 12440 10412 12492 10421
rect 12716 10412 12768 10464
rect 15476 10480 15528 10532
rect 18420 10523 18472 10532
rect 18420 10489 18429 10523
rect 18429 10489 18463 10523
rect 18463 10489 18472 10523
rect 18420 10480 18472 10489
rect 14740 10412 14792 10464
rect 15292 10455 15344 10464
rect 15292 10421 15301 10455
rect 15301 10421 15335 10455
rect 15335 10421 15344 10455
rect 15292 10412 15344 10421
rect 16304 10455 16356 10464
rect 16304 10421 16313 10455
rect 16313 10421 16347 10455
rect 16347 10421 16356 10455
rect 16304 10412 16356 10421
rect 17960 10412 18012 10464
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 3424 10251 3476 10260
rect 3424 10217 3433 10251
rect 3433 10217 3467 10251
rect 3467 10217 3476 10251
rect 3424 10208 3476 10217
rect 3516 10208 3568 10260
rect 5632 10208 5684 10260
rect 8208 10208 8260 10260
rect 9864 10251 9916 10260
rect 9864 10217 9873 10251
rect 9873 10217 9907 10251
rect 9907 10217 9916 10251
rect 9864 10208 9916 10217
rect 10048 10208 10100 10260
rect 12440 10208 12492 10260
rect 13084 10208 13136 10260
rect 13728 10208 13780 10260
rect 14096 10251 14148 10260
rect 14096 10217 14105 10251
rect 14105 10217 14139 10251
rect 14139 10217 14148 10251
rect 14096 10208 14148 10217
rect 15292 10208 15344 10260
rect 15752 10208 15804 10260
rect 17960 10208 18012 10260
rect 2596 10140 2648 10192
rect 3332 10140 3384 10192
rect 6092 10140 6144 10192
rect 8576 10140 8628 10192
rect 9956 10140 10008 10192
rect 10692 10140 10744 10192
rect 17132 10140 17184 10192
rect 18052 10183 18104 10192
rect 18052 10149 18061 10183
rect 18061 10149 18095 10183
rect 18095 10149 18104 10183
rect 18052 10140 18104 10149
rect 18512 10140 18564 10192
rect 19340 10140 19392 10192
rect 3700 10072 3752 10124
rect 5448 10072 5500 10124
rect 10140 10072 10192 10124
rect 11060 10072 11112 10124
rect 13360 10115 13412 10124
rect 13360 10081 13369 10115
rect 13369 10081 13403 10115
rect 13403 10081 13412 10115
rect 13360 10072 13412 10081
rect 4528 10047 4580 10056
rect 2228 9936 2280 9988
rect 2688 9936 2740 9988
rect 4528 10013 4537 10047
rect 4537 10013 4571 10047
rect 4571 10013 4580 10047
rect 4528 10004 4580 10013
rect 4712 10047 4764 10056
rect 4712 10013 4721 10047
rect 4721 10013 4755 10047
rect 4755 10013 4764 10047
rect 4712 10004 4764 10013
rect 5172 10004 5224 10056
rect 13728 10004 13780 10056
rect 3056 9936 3108 9988
rect 4436 9936 4488 9988
rect 7104 9979 7156 9988
rect 7104 9945 7113 9979
rect 7113 9945 7147 9979
rect 7147 9945 7156 9979
rect 7104 9936 7156 9945
rect 12900 9979 12952 9988
rect 12900 9945 12909 9979
rect 12909 9945 12943 9979
rect 12943 9945 12952 9979
rect 12900 9936 12952 9945
rect 1952 9868 2004 9920
rect 3148 9868 3200 9920
rect 4160 9868 4212 9920
rect 8392 9868 8444 9920
rect 9404 9868 9456 9920
rect 11428 9868 11480 9920
rect 12164 9868 12216 9920
rect 12440 9911 12492 9920
rect 12440 9877 12449 9911
rect 12449 9877 12483 9911
rect 12483 9877 12492 9911
rect 12992 9911 13044 9920
rect 12440 9868 12492 9877
rect 12992 9877 13001 9911
rect 13001 9877 13035 9911
rect 13035 9877 13044 9911
rect 12992 9868 13044 9877
rect 15476 9868 15528 9920
rect 15844 10072 15896 10124
rect 16948 10072 17000 10124
rect 15936 10047 15988 10056
rect 15936 10013 15945 10047
rect 15945 10013 15979 10047
rect 15979 10013 15988 10047
rect 15936 10004 15988 10013
rect 18972 10047 19024 10056
rect 18972 10013 18981 10047
rect 18981 10013 19015 10047
rect 19015 10013 19024 10047
rect 18972 10004 19024 10013
rect 18144 9936 18196 9988
rect 16580 9868 16632 9920
rect 19432 9911 19484 9920
rect 19432 9877 19441 9911
rect 19441 9877 19475 9911
rect 19475 9877 19484 9911
rect 19432 9868 19484 9877
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 2596 9664 2648 9716
rect 4252 9664 4304 9716
rect 4712 9707 4764 9716
rect 4712 9673 4721 9707
rect 4721 9673 4755 9707
rect 4755 9673 4764 9707
rect 4712 9664 4764 9673
rect 4804 9664 4856 9716
rect 6092 9707 6144 9716
rect 6092 9673 6101 9707
rect 6101 9673 6135 9707
rect 6135 9673 6144 9707
rect 6092 9664 6144 9673
rect 7196 9596 7248 9648
rect 7748 9596 7800 9648
rect 9128 9639 9180 9648
rect 9128 9605 9137 9639
rect 9137 9605 9171 9639
rect 9171 9605 9180 9639
rect 9128 9596 9180 9605
rect 15384 9664 15436 9716
rect 15936 9664 15988 9716
rect 2044 9528 2096 9580
rect 2780 9571 2832 9580
rect 2780 9537 2789 9571
rect 2789 9537 2823 9571
rect 2823 9537 2832 9571
rect 2780 9528 2832 9537
rect 5080 9571 5132 9580
rect 5080 9537 5089 9571
rect 5089 9537 5123 9571
rect 5123 9537 5132 9571
rect 5080 9528 5132 9537
rect 5540 9571 5592 9580
rect 5540 9537 5549 9571
rect 5549 9537 5583 9571
rect 5583 9537 5592 9571
rect 5540 9528 5592 9537
rect 8116 9571 8168 9580
rect 8116 9537 8125 9571
rect 8125 9537 8159 9571
rect 8159 9537 8168 9571
rect 8116 9528 8168 9537
rect 9220 9528 9272 9580
rect 10784 9596 10836 9648
rect 11152 9596 11204 9648
rect 15568 9639 15620 9648
rect 15568 9605 15577 9639
rect 15577 9605 15611 9639
rect 15611 9605 15620 9639
rect 15568 9596 15620 9605
rect 9956 9528 10008 9580
rect 14280 9528 14332 9580
rect 14556 9528 14608 9580
rect 17040 9596 17092 9648
rect 17868 9596 17920 9648
rect 19340 9596 19392 9648
rect 16580 9571 16632 9580
rect 16580 9537 16589 9571
rect 16589 9537 16623 9571
rect 16623 9537 16632 9571
rect 16580 9528 16632 9537
rect 1400 9503 1452 9512
rect 1400 9469 1409 9503
rect 1409 9469 1443 9503
rect 1443 9469 1452 9503
rect 1400 9460 1452 9469
rect 2504 9460 2556 9512
rect 3056 9503 3108 9512
rect 3056 9469 3090 9503
rect 3090 9469 3108 9503
rect 3056 9460 3108 9469
rect 3608 9460 3660 9512
rect 8208 9460 8260 9512
rect 10140 9460 10192 9512
rect 10600 9503 10652 9512
rect 10600 9469 10609 9503
rect 10609 9469 10643 9503
rect 10643 9469 10652 9503
rect 10600 9460 10652 9469
rect 10692 9460 10744 9512
rect 12532 9460 12584 9512
rect 13268 9503 13320 9512
rect 13268 9469 13277 9503
rect 13277 9469 13311 9503
rect 13311 9469 13320 9503
rect 13268 9460 13320 9469
rect 16304 9460 16356 9512
rect 17040 9460 17092 9512
rect 5080 9392 5132 9444
rect 9956 9392 10008 9444
rect 10048 9392 10100 9444
rect 4160 9367 4212 9376
rect 4160 9333 4169 9367
rect 4169 9333 4203 9367
rect 4203 9333 4212 9367
rect 4160 9324 4212 9333
rect 9496 9367 9548 9376
rect 9496 9333 9505 9367
rect 9505 9333 9539 9367
rect 9539 9333 9548 9367
rect 9496 9324 9548 9333
rect 10784 9392 10836 9444
rect 10968 9392 11020 9444
rect 13360 9392 13412 9444
rect 11244 9324 11296 9376
rect 12808 9367 12860 9376
rect 12808 9333 12817 9367
rect 12817 9333 12851 9367
rect 12851 9333 12860 9367
rect 12808 9324 12860 9333
rect 12900 9324 12952 9376
rect 14280 9392 14332 9444
rect 19340 9392 19392 9444
rect 13728 9324 13780 9376
rect 15476 9324 15528 9376
rect 16028 9367 16080 9376
rect 16028 9333 16037 9367
rect 16037 9333 16071 9367
rect 16071 9333 16080 9367
rect 16028 9324 16080 9333
rect 17224 9324 17276 9376
rect 19432 9367 19484 9376
rect 19432 9333 19441 9367
rect 19441 9333 19475 9367
rect 19475 9333 19484 9367
rect 19432 9324 19484 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 2780 9163 2832 9172
rect 2780 9129 2789 9163
rect 2789 9129 2823 9163
rect 2823 9129 2832 9163
rect 2780 9120 2832 9129
rect 5080 9120 5132 9172
rect 8484 9163 8536 9172
rect 8484 9129 8493 9163
rect 8493 9129 8527 9163
rect 8527 9129 8536 9163
rect 8484 9120 8536 9129
rect 9220 9163 9272 9172
rect 9220 9129 9229 9163
rect 9229 9129 9263 9163
rect 9263 9129 9272 9163
rect 9220 9120 9272 9129
rect 9404 9120 9456 9172
rect 10968 9120 11020 9172
rect 13084 9163 13136 9172
rect 13084 9129 13093 9163
rect 13093 9129 13127 9163
rect 13127 9129 13136 9163
rect 13084 9120 13136 9129
rect 13360 9120 13412 9172
rect 16304 9120 16356 9172
rect 2228 9052 2280 9104
rect 4620 9052 4672 9104
rect 11336 9052 11388 9104
rect 15292 9052 15344 9104
rect 17224 9120 17276 9172
rect 17960 9163 18012 9172
rect 17960 9129 17969 9163
rect 17969 9129 18003 9163
rect 18003 9129 18012 9163
rect 17960 9120 18012 9129
rect 18972 9120 19024 9172
rect 16856 9095 16908 9104
rect 16856 9061 16890 9095
rect 16890 9061 16908 9095
rect 16856 9052 16908 9061
rect 17040 9052 17092 9104
rect 2044 8984 2096 9036
rect 4804 8984 4856 9036
rect 6644 8984 6696 9036
rect 8208 8984 8260 9036
rect 13268 8984 13320 9036
rect 19432 9027 19484 9036
rect 19432 8993 19441 9027
rect 19441 8993 19475 9027
rect 19475 8993 19484 9027
rect 19432 8984 19484 8993
rect 3424 8891 3476 8900
rect 3424 8857 3433 8891
rect 3433 8857 3467 8891
rect 3467 8857 3476 8891
rect 3424 8848 3476 8857
rect 4436 8848 4488 8900
rect 5540 8916 5592 8968
rect 5172 8848 5224 8900
rect 3516 8780 3568 8832
rect 5540 8823 5592 8832
rect 5540 8789 5549 8823
rect 5549 8789 5583 8823
rect 5583 8789 5592 8823
rect 5540 8780 5592 8789
rect 6552 8916 6604 8968
rect 6828 8916 6880 8968
rect 9864 8916 9916 8968
rect 11060 8916 11112 8968
rect 13544 8916 13596 8968
rect 14280 8959 14332 8968
rect 14280 8925 14289 8959
rect 14289 8925 14323 8959
rect 14323 8925 14332 8959
rect 14280 8916 14332 8925
rect 19340 8916 19392 8968
rect 12900 8848 12952 8900
rect 6276 8780 6328 8832
rect 6552 8823 6604 8832
rect 6552 8789 6561 8823
rect 6561 8789 6595 8823
rect 6595 8789 6604 8823
rect 6552 8780 6604 8789
rect 6920 8823 6972 8832
rect 6920 8789 6929 8823
rect 6929 8789 6963 8823
rect 6963 8789 6972 8823
rect 6920 8780 6972 8789
rect 10784 8823 10836 8832
rect 10784 8789 10793 8823
rect 10793 8789 10827 8823
rect 10827 8789 10836 8823
rect 10784 8780 10836 8789
rect 12440 8780 12492 8832
rect 12808 8780 12860 8832
rect 13728 8780 13780 8832
rect 18604 8848 18656 8900
rect 20076 8891 20128 8900
rect 20076 8857 20085 8891
rect 20085 8857 20119 8891
rect 20119 8857 20128 8891
rect 20076 8848 20128 8857
rect 15384 8780 15436 8832
rect 15568 8780 15620 8832
rect 16580 8780 16632 8832
rect 18788 8780 18840 8832
rect 19064 8823 19116 8832
rect 19064 8789 19073 8823
rect 19073 8789 19107 8823
rect 19107 8789 19116 8823
rect 19064 8780 19116 8789
rect 19524 8780 19576 8832
rect 20444 8823 20496 8832
rect 20444 8789 20453 8823
rect 20453 8789 20487 8823
rect 20487 8789 20496 8823
rect 20444 8780 20496 8789
rect 21180 8823 21232 8832
rect 21180 8789 21189 8823
rect 21189 8789 21223 8823
rect 21223 8789 21232 8823
rect 21180 8780 21232 8789
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 1860 8576 1912 8628
rect 4068 8576 4120 8628
rect 9864 8619 9916 8628
rect 9864 8585 9873 8619
rect 9873 8585 9907 8619
rect 9907 8585 9916 8619
rect 9864 8576 9916 8585
rect 9956 8619 10008 8628
rect 9956 8585 9965 8619
rect 9965 8585 9999 8619
rect 9999 8585 10008 8619
rect 9956 8576 10008 8585
rect 11336 8576 11388 8628
rect 11428 8576 11480 8628
rect 12900 8576 12952 8628
rect 13268 8619 13320 8628
rect 13268 8585 13277 8619
rect 13277 8585 13311 8619
rect 13311 8585 13320 8619
rect 13268 8576 13320 8585
rect 13544 8619 13596 8628
rect 13544 8585 13553 8619
rect 13553 8585 13587 8619
rect 13587 8585 13596 8619
rect 13544 8576 13596 8585
rect 2964 8508 3016 8560
rect 3424 8508 3476 8560
rect 3884 8508 3936 8560
rect 6000 8551 6052 8560
rect 6000 8517 6009 8551
rect 6009 8517 6043 8551
rect 6043 8517 6052 8551
rect 6000 8508 6052 8517
rect 6828 8508 6880 8560
rect 8208 8551 8260 8560
rect 8208 8517 8217 8551
rect 8217 8517 8251 8551
rect 8251 8517 8260 8551
rect 8208 8508 8260 8517
rect 8852 8551 8904 8560
rect 8852 8517 8861 8551
rect 8861 8517 8895 8551
rect 8895 8517 8904 8551
rect 8852 8508 8904 8517
rect 1952 8483 2004 8492
rect 1952 8449 1961 8483
rect 1961 8449 1995 8483
rect 1995 8449 2004 8483
rect 1952 8440 2004 8449
rect 2228 8440 2280 8492
rect 3516 8483 3568 8492
rect 3516 8449 3525 8483
rect 3525 8449 3559 8483
rect 3559 8449 3568 8483
rect 3516 8440 3568 8449
rect 3608 8440 3660 8492
rect 4160 8440 4212 8492
rect 5172 8483 5224 8492
rect 5172 8449 5181 8483
rect 5181 8449 5215 8483
rect 5215 8449 5224 8483
rect 5172 8440 5224 8449
rect 6644 8415 6696 8424
rect 2412 8304 2464 8356
rect 4804 8304 4856 8356
rect 3884 8236 3936 8288
rect 4712 8236 4764 8288
rect 4988 8279 5040 8288
rect 4988 8245 4997 8279
rect 4997 8245 5031 8279
rect 5031 8245 5040 8279
rect 4988 8236 5040 8245
rect 6644 8381 6653 8415
rect 6653 8381 6687 8415
rect 6687 8381 6696 8415
rect 6644 8372 6696 8381
rect 10692 8440 10744 8492
rect 8576 8372 8628 8424
rect 9864 8372 9916 8424
rect 14096 8576 14148 8628
rect 16028 8576 16080 8628
rect 16856 8576 16908 8628
rect 20720 8576 20772 8628
rect 13360 8440 13412 8492
rect 17960 8508 18012 8560
rect 19340 8508 19392 8560
rect 19616 8551 19668 8560
rect 19616 8517 19625 8551
rect 19625 8517 19659 8551
rect 19659 8517 19668 8551
rect 19616 8508 19668 8517
rect 20076 8508 20128 8560
rect 20996 8551 21048 8560
rect 13544 8372 13596 8424
rect 18604 8483 18656 8492
rect 6368 8236 6420 8288
rect 6644 8236 6696 8288
rect 6920 8304 6972 8356
rect 9128 8304 9180 8356
rect 10140 8304 10192 8356
rect 16028 8372 16080 8424
rect 16672 8347 16724 8356
rect 8576 8236 8628 8288
rect 9404 8236 9456 8288
rect 10692 8236 10744 8288
rect 11060 8236 11112 8288
rect 11244 8236 11296 8288
rect 12532 8236 12584 8288
rect 13544 8236 13596 8288
rect 13728 8236 13780 8288
rect 14648 8236 14700 8288
rect 16212 8279 16264 8288
rect 16212 8245 16221 8279
rect 16221 8245 16255 8279
rect 16255 8245 16264 8279
rect 16212 8236 16264 8245
rect 16672 8313 16681 8347
rect 16681 8313 16715 8347
rect 16715 8313 16724 8347
rect 16672 8304 16724 8313
rect 18604 8449 18613 8483
rect 18613 8449 18647 8483
rect 18647 8449 18656 8483
rect 18604 8440 18656 8449
rect 19432 8483 19484 8492
rect 19432 8449 19441 8483
rect 19441 8449 19475 8483
rect 19475 8449 19484 8483
rect 19432 8440 19484 8449
rect 20996 8517 21005 8551
rect 21005 8517 21039 8551
rect 21039 8517 21048 8551
rect 20996 8508 21048 8517
rect 19064 8372 19116 8424
rect 18788 8304 18840 8356
rect 19340 8304 19392 8356
rect 20444 8372 20496 8424
rect 21180 8440 21232 8492
rect 18052 8279 18104 8288
rect 18052 8245 18061 8279
rect 18061 8245 18095 8279
rect 18095 8245 18104 8279
rect 18052 8236 18104 8245
rect 18696 8236 18748 8288
rect 19524 8236 19576 8288
rect 21640 8279 21692 8288
rect 21640 8245 21649 8279
rect 21649 8245 21683 8279
rect 21683 8245 21692 8279
rect 21640 8236 21692 8245
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 2228 8032 2280 8084
rect 2412 8075 2464 8084
rect 2412 8041 2421 8075
rect 2421 8041 2455 8075
rect 2455 8041 2464 8075
rect 2412 8032 2464 8041
rect 3608 8032 3660 8084
rect 3884 8075 3936 8084
rect 3884 8041 3893 8075
rect 3893 8041 3927 8075
rect 3927 8041 3936 8075
rect 3884 8032 3936 8041
rect 4620 8075 4672 8084
rect 4620 8041 4629 8075
rect 4629 8041 4663 8075
rect 4663 8041 4672 8075
rect 4620 8032 4672 8041
rect 8208 8032 8260 8084
rect 8852 8075 8904 8084
rect 8852 8041 8861 8075
rect 8861 8041 8895 8075
rect 8895 8041 8904 8075
rect 8852 8032 8904 8041
rect 10140 8075 10192 8084
rect 10140 8041 10149 8075
rect 10149 8041 10183 8075
rect 10183 8041 10192 8075
rect 10140 8032 10192 8041
rect 12348 8032 12400 8084
rect 14280 8032 14332 8084
rect 15108 8075 15160 8084
rect 15108 8041 15117 8075
rect 15117 8041 15151 8075
rect 15151 8041 15160 8075
rect 15108 8032 15160 8041
rect 19064 8075 19116 8084
rect 2872 8007 2924 8016
rect 2872 7973 2881 8007
rect 2881 7973 2915 8007
rect 2915 7973 2924 8007
rect 2872 7964 2924 7973
rect 2780 7939 2832 7948
rect 2780 7905 2789 7939
rect 2789 7905 2823 7939
rect 2823 7905 2832 7939
rect 6828 7964 6880 8016
rect 13820 7964 13872 8016
rect 2780 7896 2832 7905
rect 5540 7939 5592 7948
rect 5540 7905 5574 7939
rect 5574 7905 5592 7939
rect 5540 7896 5592 7905
rect 8116 7939 8168 7948
rect 8116 7905 8125 7939
rect 8125 7905 8159 7939
rect 8159 7905 8168 7939
rect 8116 7896 8168 7905
rect 9680 7939 9732 7948
rect 9680 7905 9689 7939
rect 9689 7905 9723 7939
rect 9723 7905 9732 7939
rect 9680 7896 9732 7905
rect 11244 7896 11296 7948
rect 12348 7896 12400 7948
rect 12440 7896 12492 7948
rect 14740 7896 14792 7948
rect 15752 7896 15804 7948
rect 17040 7964 17092 8016
rect 16764 7896 16816 7948
rect 19064 8041 19073 8075
rect 19073 8041 19107 8075
rect 19107 8041 19116 8075
rect 19064 8032 19116 8041
rect 19248 8032 19300 8084
rect 19984 8032 20036 8084
rect 18880 7964 18932 8016
rect 21640 7896 21692 7948
rect 2964 7871 3016 7880
rect 2964 7837 2973 7871
rect 2973 7837 3007 7871
rect 3007 7837 3016 7871
rect 2964 7828 3016 7837
rect 7840 7828 7892 7880
rect 8668 7828 8720 7880
rect 1308 7760 1360 7812
rect 4712 7760 4764 7812
rect 7012 7760 7064 7812
rect 9312 7803 9364 7812
rect 9312 7769 9321 7803
rect 9321 7769 9355 7803
rect 9355 7769 9364 7803
rect 9312 7760 9364 7769
rect 2320 7735 2372 7744
rect 2320 7701 2329 7735
rect 2329 7701 2363 7735
rect 2363 7701 2372 7735
rect 2320 7692 2372 7701
rect 2688 7692 2740 7744
rect 6644 7735 6696 7744
rect 6644 7701 6653 7735
rect 6653 7701 6687 7735
rect 6687 7701 6696 7735
rect 6644 7692 6696 7701
rect 7564 7735 7616 7744
rect 7564 7701 7573 7735
rect 7573 7701 7607 7735
rect 7607 7701 7616 7735
rect 7564 7692 7616 7701
rect 10692 7692 10744 7744
rect 12072 7692 12124 7744
rect 13360 7828 13412 7880
rect 14280 7871 14332 7880
rect 13636 7803 13688 7812
rect 13636 7769 13645 7803
rect 13645 7769 13679 7803
rect 13679 7769 13688 7803
rect 13636 7760 13688 7769
rect 14280 7837 14289 7871
rect 14289 7837 14323 7871
rect 14323 7837 14332 7871
rect 14280 7828 14332 7837
rect 15384 7828 15436 7880
rect 13268 7692 13320 7744
rect 16396 7760 16448 7812
rect 19524 7760 19576 7812
rect 15292 7692 15344 7744
rect 16028 7692 16080 7744
rect 16672 7692 16724 7744
rect 18144 7692 18196 7744
rect 18696 7735 18748 7744
rect 18696 7701 18705 7735
rect 18705 7701 18739 7735
rect 18739 7701 18748 7735
rect 18696 7692 18748 7701
rect 20076 7692 20128 7744
rect 20536 7735 20588 7744
rect 20536 7701 20545 7735
rect 20545 7701 20579 7735
rect 20579 7701 20588 7735
rect 20536 7692 20588 7701
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 1676 7531 1728 7540
rect 1676 7497 1685 7531
rect 1685 7497 1719 7531
rect 1719 7497 1728 7531
rect 1676 7488 1728 7497
rect 2964 7488 3016 7540
rect 6460 7488 6512 7540
rect 6736 7488 6788 7540
rect 7840 7531 7892 7540
rect 7840 7497 7849 7531
rect 7849 7497 7883 7531
rect 7883 7497 7892 7531
rect 7840 7488 7892 7497
rect 8668 7531 8720 7540
rect 8668 7497 8677 7531
rect 8677 7497 8711 7531
rect 8711 7497 8720 7531
rect 8668 7488 8720 7497
rect 12348 7488 12400 7540
rect 13176 7488 13228 7540
rect 13820 7488 13872 7540
rect 16672 7488 16724 7540
rect 18880 7488 18932 7540
rect 19616 7531 19668 7540
rect 19616 7497 19625 7531
rect 19625 7497 19659 7531
rect 19659 7497 19668 7531
rect 19616 7488 19668 7497
rect 20720 7488 20772 7540
rect 1584 7352 1636 7404
rect 2044 7352 2096 7404
rect 2320 7284 2372 7336
rect 2964 7284 3016 7336
rect 3976 7420 4028 7472
rect 5172 7463 5224 7472
rect 5172 7429 5181 7463
rect 5181 7429 5215 7463
rect 5215 7429 5224 7463
rect 5172 7420 5224 7429
rect 6092 7352 6144 7404
rect 7380 7395 7432 7404
rect 7380 7361 7389 7395
rect 7389 7361 7423 7395
rect 7423 7361 7432 7395
rect 7380 7352 7432 7361
rect 8668 7352 8720 7404
rect 11152 7420 11204 7472
rect 12808 7352 12860 7404
rect 13636 7395 13688 7404
rect 13636 7361 13645 7395
rect 13645 7361 13679 7395
rect 13679 7361 13688 7395
rect 13636 7352 13688 7361
rect 3424 7284 3476 7336
rect 4344 7284 4396 7336
rect 6736 7284 6788 7336
rect 9588 7284 9640 7336
rect 13728 7284 13780 7336
rect 18420 7352 18472 7404
rect 19524 7352 19576 7404
rect 20996 7395 21048 7404
rect 20996 7361 21005 7395
rect 21005 7361 21039 7395
rect 21039 7361 21048 7395
rect 20996 7352 21048 7361
rect 14648 7327 14700 7336
rect 14648 7293 14657 7327
rect 14657 7293 14691 7327
rect 14691 7293 14700 7327
rect 14648 7284 14700 7293
rect 17040 7284 17092 7336
rect 17408 7327 17460 7336
rect 17408 7293 17417 7327
rect 17417 7293 17451 7327
rect 17451 7293 17460 7327
rect 17408 7284 17460 7293
rect 1124 7148 1176 7200
rect 2872 7148 2924 7200
rect 3700 7148 3752 7200
rect 6000 7216 6052 7268
rect 6460 7216 6512 7268
rect 9312 7216 9364 7268
rect 6828 7191 6880 7200
rect 6828 7157 6837 7191
rect 6837 7157 6871 7191
rect 6871 7157 6880 7191
rect 6828 7148 6880 7157
rect 8208 7191 8260 7200
rect 8208 7157 8217 7191
rect 8217 7157 8251 7191
rect 8251 7157 8260 7191
rect 8208 7148 8260 7157
rect 9496 7148 9548 7200
rect 10140 7216 10192 7268
rect 10692 7216 10744 7268
rect 14096 7216 14148 7268
rect 16580 7216 16632 7268
rect 20168 7216 20220 7268
rect 21180 7216 21232 7268
rect 9864 7148 9916 7200
rect 10968 7148 11020 7200
rect 11980 7148 12032 7200
rect 13176 7191 13228 7200
rect 13176 7157 13185 7191
rect 13185 7157 13219 7191
rect 13219 7157 13228 7191
rect 13176 7148 13228 7157
rect 13544 7191 13596 7200
rect 13544 7157 13553 7191
rect 13553 7157 13587 7191
rect 13587 7157 13596 7191
rect 13544 7148 13596 7157
rect 15384 7148 15436 7200
rect 16764 7148 16816 7200
rect 17040 7148 17092 7200
rect 18052 7191 18104 7200
rect 18052 7157 18061 7191
rect 18061 7157 18095 7191
rect 18095 7157 18104 7191
rect 18052 7148 18104 7157
rect 18512 7191 18564 7200
rect 18512 7157 18521 7191
rect 18521 7157 18555 7191
rect 18555 7157 18564 7191
rect 18512 7148 18564 7157
rect 20076 7191 20128 7200
rect 20076 7157 20085 7191
rect 20085 7157 20119 7191
rect 20119 7157 20128 7191
rect 20076 7148 20128 7157
rect 21548 7191 21600 7200
rect 21548 7157 21557 7191
rect 21557 7157 21591 7191
rect 21591 7157 21600 7191
rect 21548 7148 21600 7157
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 1676 6944 1728 6996
rect 2780 6987 2832 6996
rect 2780 6953 2789 6987
rect 2789 6953 2823 6987
rect 2823 6953 2832 6987
rect 2780 6944 2832 6953
rect 7380 6944 7432 6996
rect 8668 6987 8720 6996
rect 8668 6953 8677 6987
rect 8677 6953 8711 6987
rect 8711 6953 8720 6987
rect 8668 6944 8720 6953
rect 9588 6944 9640 6996
rect 11060 6944 11112 6996
rect 11980 6987 12032 6996
rect 11980 6953 11989 6987
rect 11989 6953 12023 6987
rect 12023 6953 12032 6987
rect 11980 6944 12032 6953
rect 13544 6944 13596 6996
rect 1492 6876 1544 6928
rect 4712 6876 4764 6928
rect 8300 6876 8352 6928
rect 4988 6851 5040 6860
rect 4988 6817 4997 6851
rect 4997 6817 5031 6851
rect 5031 6817 5040 6851
rect 4988 6808 5040 6817
rect 6092 6808 6144 6860
rect 8024 6851 8076 6860
rect 8024 6817 8033 6851
rect 8033 6817 8067 6851
rect 8067 6817 8076 6851
rect 8024 6808 8076 6817
rect 10324 6808 10376 6860
rect 12072 6808 12124 6860
rect 12992 6808 13044 6860
rect 13268 6851 13320 6860
rect 13268 6817 13277 6851
rect 13277 6817 13311 6851
rect 13311 6817 13320 6851
rect 13268 6808 13320 6817
rect 1768 6672 1820 6724
rect 2504 6740 2556 6792
rect 5080 6783 5132 6792
rect 5080 6749 5089 6783
rect 5089 6749 5123 6783
rect 5123 6749 5132 6783
rect 5080 6740 5132 6749
rect 7656 6740 7708 6792
rect 6552 6672 6604 6724
rect 9404 6672 9456 6724
rect 12532 6740 12584 6792
rect 13636 6740 13688 6792
rect 14280 6944 14332 6996
rect 15752 6987 15804 6996
rect 15752 6953 15761 6987
rect 15761 6953 15795 6987
rect 15795 6953 15804 6987
rect 15752 6944 15804 6953
rect 18420 6944 18472 6996
rect 19524 6944 19576 6996
rect 16120 6851 16172 6860
rect 16120 6817 16129 6851
rect 16129 6817 16163 6851
rect 16163 6817 16172 6851
rect 16120 6808 16172 6817
rect 16948 6808 17000 6860
rect 18512 6876 18564 6928
rect 19984 6876 20036 6928
rect 18144 6851 18196 6860
rect 18144 6817 18178 6851
rect 18178 6817 18196 6851
rect 18144 6808 18196 6817
rect 16212 6740 16264 6792
rect 11152 6672 11204 6724
rect 15936 6672 15988 6724
rect 16488 6672 16540 6724
rect 1860 6604 1912 6656
rect 2596 6604 2648 6656
rect 3516 6647 3568 6656
rect 3516 6613 3525 6647
rect 3525 6613 3559 6647
rect 3559 6613 3568 6647
rect 3516 6604 3568 6613
rect 3884 6647 3936 6656
rect 3884 6613 3893 6647
rect 3893 6613 3927 6647
rect 3927 6613 3936 6647
rect 3884 6604 3936 6613
rect 4620 6647 4672 6656
rect 4620 6613 4629 6647
rect 4629 6613 4663 6647
rect 4663 6613 4672 6647
rect 4620 6604 4672 6613
rect 6276 6604 6328 6656
rect 7380 6647 7432 6656
rect 7380 6613 7389 6647
rect 7389 6613 7423 6647
rect 7423 6613 7432 6647
rect 7380 6604 7432 6613
rect 14832 6647 14884 6656
rect 14832 6613 14841 6647
rect 14841 6613 14875 6647
rect 14875 6613 14884 6647
rect 14832 6604 14884 6613
rect 16120 6604 16172 6656
rect 16856 6783 16908 6792
rect 16856 6749 16865 6783
rect 16865 6749 16899 6783
rect 16899 6749 16908 6783
rect 17316 6783 17368 6792
rect 16856 6740 16908 6749
rect 17316 6749 17325 6783
rect 17325 6749 17359 6783
rect 17359 6749 17368 6783
rect 17316 6740 17368 6749
rect 21180 6783 21232 6792
rect 17040 6672 17092 6724
rect 21180 6749 21189 6783
rect 21189 6749 21223 6783
rect 21223 6749 21232 6783
rect 21180 6740 21232 6749
rect 20536 6647 20588 6656
rect 20536 6613 20545 6647
rect 20545 6613 20579 6647
rect 20579 6613 20588 6647
rect 20536 6604 20588 6613
rect 21548 6647 21600 6656
rect 21548 6613 21557 6647
rect 21557 6613 21591 6647
rect 21591 6613 21600 6647
rect 21548 6604 21600 6613
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 2688 6400 2740 6452
rect 4160 6400 4212 6452
rect 4988 6443 5040 6452
rect 4988 6409 4997 6443
rect 4997 6409 5031 6443
rect 5031 6409 5040 6443
rect 4988 6400 5040 6409
rect 8024 6400 8076 6452
rect 8300 6443 8352 6452
rect 8300 6409 8309 6443
rect 8309 6409 8343 6443
rect 8343 6409 8352 6443
rect 8300 6400 8352 6409
rect 2872 6332 2924 6384
rect 6828 6375 6880 6384
rect 1584 6307 1636 6316
rect 1584 6273 1593 6307
rect 1593 6273 1627 6307
rect 1627 6273 1636 6307
rect 1584 6264 1636 6273
rect 4620 6307 4672 6316
rect 4620 6273 4629 6307
rect 4629 6273 4663 6307
rect 4663 6273 4672 6307
rect 4620 6264 4672 6273
rect 5540 6264 5592 6316
rect 6276 6264 6328 6316
rect 6828 6341 6837 6375
rect 6837 6341 6871 6375
rect 6871 6341 6880 6375
rect 6828 6332 6880 6341
rect 6092 6196 6144 6248
rect 6368 6196 6420 6248
rect 7656 6264 7708 6316
rect 8576 6400 8628 6452
rect 9404 6400 9456 6452
rect 10324 6443 10376 6452
rect 10324 6409 10333 6443
rect 10333 6409 10367 6443
rect 10367 6409 10376 6443
rect 10324 6400 10376 6409
rect 11060 6443 11112 6452
rect 11060 6409 11069 6443
rect 11069 6409 11103 6443
rect 11103 6409 11112 6443
rect 11060 6400 11112 6409
rect 13636 6400 13688 6452
rect 14096 6400 14148 6452
rect 16212 6443 16264 6452
rect 16212 6409 16221 6443
rect 16221 6409 16255 6443
rect 16255 6409 16264 6443
rect 16212 6400 16264 6409
rect 16948 6400 17000 6452
rect 10692 6307 10744 6316
rect 10692 6273 10701 6307
rect 10701 6273 10735 6307
rect 10735 6273 10744 6307
rect 10692 6264 10744 6273
rect 13176 6264 13228 6316
rect 13728 6307 13780 6316
rect 13728 6273 13737 6307
rect 13737 6273 13771 6307
rect 13771 6273 13780 6307
rect 13728 6264 13780 6273
rect 14740 6375 14792 6384
rect 14740 6341 14749 6375
rect 14749 6341 14783 6375
rect 14783 6341 14792 6375
rect 14740 6332 14792 6341
rect 8668 6239 8720 6248
rect 8668 6205 8702 6239
rect 8702 6205 8720 6239
rect 8668 6196 8720 6205
rect 12992 6196 13044 6248
rect 14832 6264 14884 6316
rect 15384 6307 15436 6316
rect 15384 6273 15393 6307
rect 15393 6273 15427 6307
rect 15427 6273 15436 6307
rect 15384 6264 15436 6273
rect 16580 6264 16632 6316
rect 16856 6264 16908 6316
rect 18144 6400 18196 6452
rect 18420 6443 18472 6452
rect 18420 6409 18429 6443
rect 18429 6409 18463 6443
rect 18463 6409 18472 6443
rect 18420 6400 18472 6409
rect 20444 6443 20496 6452
rect 20444 6409 20453 6443
rect 20453 6409 20487 6443
rect 20487 6409 20496 6443
rect 20444 6400 20496 6409
rect 20812 6375 20864 6384
rect 20812 6341 20821 6375
rect 20821 6341 20855 6375
rect 20855 6341 20864 6375
rect 20812 6332 20864 6341
rect 20996 6375 21048 6384
rect 20996 6341 21005 6375
rect 21005 6341 21039 6375
rect 21039 6341 21048 6375
rect 20996 6332 21048 6341
rect 16212 6196 16264 6248
rect 17040 6196 17092 6248
rect 18512 6239 18564 6248
rect 18512 6205 18521 6239
rect 18521 6205 18555 6239
rect 18555 6205 18564 6239
rect 18512 6196 18564 6205
rect 21640 6307 21692 6316
rect 21640 6273 21649 6307
rect 21649 6273 21683 6307
rect 21683 6273 21692 6307
rect 21640 6264 21692 6273
rect 22008 6196 22060 6248
rect 1952 6128 2004 6180
rect 2872 6128 2924 6180
rect 5172 6128 5224 6180
rect 16856 6171 16908 6180
rect 3608 6103 3660 6112
rect 3608 6069 3617 6103
rect 3617 6069 3651 6103
rect 3651 6069 3660 6103
rect 3608 6060 3660 6069
rect 4068 6103 4120 6112
rect 4068 6069 4077 6103
rect 4077 6069 4111 6103
rect 4111 6069 4120 6103
rect 4068 6060 4120 6069
rect 5080 6103 5132 6112
rect 5080 6069 5089 6103
rect 5089 6069 5123 6103
rect 5123 6069 5132 6103
rect 5080 6060 5132 6069
rect 6828 6060 6880 6112
rect 6920 6060 6972 6112
rect 10140 6060 10192 6112
rect 12532 6060 12584 6112
rect 13084 6060 13136 6112
rect 16856 6137 16865 6171
rect 16865 6137 16899 6171
rect 16899 6137 16908 6171
rect 16856 6128 16908 6137
rect 15292 6103 15344 6112
rect 15292 6069 15301 6103
rect 15301 6069 15335 6103
rect 15335 6069 15344 6103
rect 15292 6060 15344 6069
rect 16764 6103 16816 6112
rect 16764 6069 16773 6103
rect 16773 6069 16807 6103
rect 16807 6069 16816 6103
rect 16764 6060 16816 6069
rect 19340 6060 19392 6112
rect 22100 6103 22152 6112
rect 22100 6069 22109 6103
rect 22109 6069 22143 6103
rect 22143 6069 22152 6103
rect 22100 6060 22152 6069
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 2872 5899 2924 5908
rect 2872 5865 2881 5899
rect 2881 5865 2915 5899
rect 2915 5865 2924 5899
rect 2872 5856 2924 5865
rect 3516 5856 3568 5908
rect 5908 5856 5960 5908
rect 6552 5856 6604 5908
rect 6920 5899 6972 5908
rect 6920 5865 6929 5899
rect 6929 5865 6963 5899
rect 6963 5865 6972 5899
rect 6920 5856 6972 5865
rect 7656 5856 7708 5908
rect 8024 5899 8076 5908
rect 8024 5865 8033 5899
rect 8033 5865 8067 5899
rect 8067 5865 8076 5899
rect 8024 5856 8076 5865
rect 9680 5856 9732 5908
rect 11060 5856 11112 5908
rect 11520 5899 11572 5908
rect 1768 5831 1820 5840
rect 1768 5797 1802 5831
rect 1802 5797 1820 5831
rect 1768 5788 1820 5797
rect 1860 5788 1912 5840
rect 10048 5831 10100 5840
rect 10048 5797 10057 5831
rect 10057 5797 10091 5831
rect 10091 5797 10100 5831
rect 10048 5788 10100 5797
rect 10692 5831 10744 5840
rect 10692 5797 10701 5831
rect 10701 5797 10735 5831
rect 10735 5797 10744 5831
rect 10692 5788 10744 5797
rect 11520 5865 11529 5899
rect 11529 5865 11563 5899
rect 11563 5865 11572 5899
rect 11520 5856 11572 5865
rect 12992 5899 13044 5908
rect 12992 5865 13001 5899
rect 13001 5865 13035 5899
rect 13035 5865 13044 5899
rect 12992 5856 13044 5865
rect 13268 5856 13320 5908
rect 13452 5856 13504 5908
rect 13728 5856 13780 5908
rect 15384 5856 15436 5908
rect 15936 5899 15988 5908
rect 15936 5865 15945 5899
rect 15945 5865 15979 5899
rect 15979 5865 15988 5899
rect 16580 5899 16632 5908
rect 15936 5856 15988 5865
rect 16580 5865 16589 5899
rect 16589 5865 16623 5899
rect 16623 5865 16632 5899
rect 16580 5856 16632 5865
rect 16856 5899 16908 5908
rect 16856 5865 16865 5899
rect 16865 5865 16899 5899
rect 16899 5865 16908 5899
rect 16856 5856 16908 5865
rect 18512 5856 18564 5908
rect 20536 5856 20588 5908
rect 12440 5788 12492 5840
rect 17224 5788 17276 5840
rect 1584 5720 1636 5772
rect 2688 5720 2740 5772
rect 3884 5720 3936 5772
rect 5448 5720 5500 5772
rect 6092 5763 6144 5772
rect 6092 5729 6101 5763
rect 6101 5729 6135 5763
rect 6135 5729 6144 5763
rect 6092 5720 6144 5729
rect 8392 5763 8444 5772
rect 8392 5729 8401 5763
rect 8401 5729 8435 5763
rect 8435 5729 8444 5763
rect 8392 5720 8444 5729
rect 11888 5763 11940 5772
rect 4160 5652 4212 5704
rect 6276 5695 6328 5704
rect 6276 5661 6285 5695
rect 6285 5661 6319 5695
rect 6319 5661 6328 5695
rect 6276 5652 6328 5661
rect 8300 5652 8352 5704
rect 11888 5729 11897 5763
rect 11897 5729 11931 5763
rect 11931 5729 11940 5763
rect 11888 5720 11940 5729
rect 13728 5720 13780 5772
rect 14556 5720 14608 5772
rect 15292 5720 15344 5772
rect 15844 5720 15896 5772
rect 19524 5763 19576 5772
rect 19524 5729 19533 5763
rect 19533 5729 19567 5763
rect 19567 5729 19576 5763
rect 19524 5720 19576 5729
rect 10232 5695 10284 5704
rect 4068 5627 4120 5636
rect 4068 5593 4077 5627
rect 4077 5593 4111 5627
rect 4111 5593 4120 5627
rect 4068 5584 4120 5593
rect 10232 5661 10241 5695
rect 10241 5661 10275 5695
rect 10275 5661 10284 5695
rect 10232 5652 10284 5661
rect 11980 5695 12032 5704
rect 11980 5661 11989 5695
rect 11989 5661 12023 5695
rect 12023 5661 12032 5695
rect 11980 5652 12032 5661
rect 12072 5695 12124 5704
rect 12072 5661 12081 5695
rect 12081 5661 12115 5695
rect 12115 5661 12124 5695
rect 12072 5652 12124 5661
rect 12808 5652 12860 5704
rect 9036 5627 9088 5636
rect 9036 5593 9045 5627
rect 9045 5593 9079 5627
rect 9079 5593 9088 5627
rect 9036 5584 9088 5593
rect 11152 5584 11204 5636
rect 13268 5584 13320 5636
rect 15568 5652 15620 5704
rect 16120 5695 16172 5704
rect 16120 5661 16129 5695
rect 16129 5661 16163 5695
rect 16163 5661 16172 5695
rect 16120 5652 16172 5661
rect 16580 5652 16632 5704
rect 17040 5695 17092 5704
rect 17040 5661 17049 5695
rect 17049 5661 17083 5695
rect 17083 5661 17092 5695
rect 17040 5652 17092 5661
rect 13728 5584 13780 5636
rect 2964 5516 3016 5568
rect 5356 5516 5408 5568
rect 7840 5559 7892 5568
rect 7840 5525 7849 5559
rect 7849 5525 7883 5559
rect 7883 5525 7892 5559
rect 7840 5516 7892 5525
rect 10140 5516 10192 5568
rect 13636 5516 13688 5568
rect 14648 5516 14700 5568
rect 16028 5516 16080 5568
rect 18328 5516 18380 5568
rect 18512 5516 18564 5568
rect 19432 5516 19484 5568
rect 20720 5516 20772 5568
rect 21640 5516 21692 5568
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 2596 5312 2648 5364
rect 2964 5355 3016 5364
rect 2964 5321 2973 5355
rect 2973 5321 3007 5355
rect 3007 5321 3016 5355
rect 2964 5312 3016 5321
rect 4160 5355 4212 5364
rect 4160 5321 4169 5355
rect 4169 5321 4203 5355
rect 4203 5321 4212 5355
rect 4160 5312 4212 5321
rect 5448 5312 5500 5364
rect 7288 5312 7340 5364
rect 9956 5312 10008 5364
rect 10968 5312 11020 5364
rect 11152 5355 11204 5364
rect 11152 5321 11161 5355
rect 11161 5321 11195 5355
rect 11195 5321 11204 5355
rect 11152 5312 11204 5321
rect 11888 5312 11940 5364
rect 13452 5355 13504 5364
rect 13452 5321 13461 5355
rect 13461 5321 13495 5355
rect 13495 5321 13504 5355
rect 13452 5312 13504 5321
rect 13912 5355 13964 5364
rect 13912 5321 13921 5355
rect 13921 5321 13955 5355
rect 13955 5321 13964 5355
rect 13912 5312 13964 5321
rect 15384 5312 15436 5364
rect 16120 5312 16172 5364
rect 18052 5355 18104 5364
rect 18052 5321 18061 5355
rect 18061 5321 18095 5355
rect 18095 5321 18104 5355
rect 18052 5312 18104 5321
rect 20076 5312 20128 5364
rect 20536 5312 20588 5364
rect 1768 5244 1820 5296
rect 1952 5219 2004 5228
rect 1952 5185 1961 5219
rect 1961 5185 1995 5219
rect 1995 5185 2004 5219
rect 1952 5176 2004 5185
rect 13820 5244 13872 5296
rect 15476 5244 15528 5296
rect 2228 5176 2280 5228
rect 3608 5219 3660 5228
rect 3608 5185 3617 5219
rect 3617 5185 3651 5219
rect 3651 5185 3660 5219
rect 3608 5176 3660 5185
rect 5632 5176 5684 5228
rect 6368 5176 6420 5228
rect 1860 5151 1912 5160
rect 1860 5117 1869 5151
rect 1869 5117 1903 5151
rect 1903 5117 1912 5151
rect 1860 5108 1912 5117
rect 6552 5108 6604 5160
rect 7196 5151 7248 5160
rect 7196 5117 7205 5151
rect 7205 5117 7239 5151
rect 7239 5117 7248 5151
rect 7196 5108 7248 5117
rect 1676 5040 1728 5092
rect 2504 5040 2556 5092
rect 8576 5219 8628 5228
rect 8576 5185 8585 5219
rect 8585 5185 8619 5219
rect 8619 5185 8628 5219
rect 8576 5176 8628 5185
rect 12900 5219 12952 5228
rect 12900 5185 12909 5219
rect 12909 5185 12943 5219
rect 12943 5185 12952 5219
rect 12900 5176 12952 5185
rect 13268 5176 13320 5228
rect 16764 5219 16816 5228
rect 16764 5185 16773 5219
rect 16773 5185 16807 5219
rect 16807 5185 16816 5219
rect 16764 5176 16816 5185
rect 18328 5176 18380 5228
rect 18972 5176 19024 5228
rect 20720 5176 20772 5228
rect 11152 5108 11204 5160
rect 12440 5108 12492 5160
rect 16304 5108 16356 5160
rect 19248 5108 19300 5160
rect 21180 5151 21232 5160
rect 21180 5117 21189 5151
rect 21189 5117 21223 5151
rect 21223 5117 21232 5151
rect 21180 5108 21232 5117
rect 8668 5040 8720 5092
rect 10232 5040 10284 5092
rect 11336 5040 11388 5092
rect 11980 5040 12032 5092
rect 14556 5040 14608 5092
rect 15384 5083 15436 5092
rect 15384 5049 15393 5083
rect 15393 5049 15427 5083
rect 15427 5049 15436 5083
rect 15384 5040 15436 5049
rect 21456 5083 21508 5092
rect 21456 5049 21465 5083
rect 21465 5049 21499 5083
rect 21499 5049 21508 5083
rect 21456 5040 21508 5049
rect 2596 4972 2648 5024
rect 3884 4972 3936 5024
rect 5356 4972 5408 5024
rect 6000 4972 6052 5024
rect 6368 4972 6420 5024
rect 6828 5015 6880 5024
rect 6828 4981 6837 5015
rect 6837 4981 6871 5015
rect 6871 4981 6880 5015
rect 6828 4972 6880 4981
rect 7288 5015 7340 5024
rect 7288 4981 7297 5015
rect 7297 4981 7331 5015
rect 7331 4981 7340 5015
rect 7288 4972 7340 4981
rect 7932 4972 7984 5024
rect 8208 4972 8260 5024
rect 8392 5015 8444 5024
rect 8392 4981 8401 5015
rect 8401 4981 8435 5015
rect 8435 4981 8444 5015
rect 8392 4972 8444 4981
rect 9956 5015 10008 5024
rect 9956 4981 9965 5015
rect 9965 4981 9999 5015
rect 9999 4981 10008 5015
rect 9956 4972 10008 4981
rect 11612 4972 11664 5024
rect 12440 5015 12492 5024
rect 12440 4981 12449 5015
rect 12449 4981 12483 5015
rect 12483 4981 12492 5015
rect 12440 4972 12492 4981
rect 14924 4972 14976 5024
rect 16396 4972 16448 5024
rect 16856 4972 16908 5024
rect 17224 5015 17276 5024
rect 17224 4981 17233 5015
rect 17233 4981 17267 5015
rect 17267 4981 17276 5015
rect 17224 4972 17276 4981
rect 18512 5015 18564 5024
rect 18512 4981 18521 5015
rect 18521 4981 18555 5015
rect 18555 4981 18564 5015
rect 19064 5015 19116 5024
rect 18512 4972 18564 4981
rect 19064 4981 19073 5015
rect 19073 4981 19107 5015
rect 19107 4981 19116 5015
rect 19064 4972 19116 4981
rect 19340 4972 19392 5024
rect 21364 4972 21416 5024
rect 22100 4972 22152 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 1676 4811 1728 4820
rect 1676 4777 1685 4811
rect 1685 4777 1719 4811
rect 1719 4777 1728 4811
rect 1676 4768 1728 4777
rect 2964 4768 3016 4820
rect 3608 4768 3660 4820
rect 4068 4768 4120 4820
rect 5632 4811 5684 4820
rect 5632 4777 5641 4811
rect 5641 4777 5675 4811
rect 5675 4777 5684 4811
rect 5632 4768 5684 4777
rect 6276 4811 6328 4820
rect 6276 4777 6285 4811
rect 6285 4777 6319 4811
rect 6319 4777 6328 4811
rect 6276 4768 6328 4777
rect 6828 4768 6880 4820
rect 7288 4768 7340 4820
rect 8668 4811 8720 4820
rect 8668 4777 8677 4811
rect 8677 4777 8711 4811
rect 8711 4777 8720 4811
rect 8668 4768 8720 4777
rect 9496 4811 9548 4820
rect 9496 4777 9505 4811
rect 9505 4777 9539 4811
rect 9539 4777 9548 4811
rect 9496 4768 9548 4777
rect 9772 4768 9824 4820
rect 10048 4811 10100 4820
rect 10048 4777 10057 4811
rect 10057 4777 10091 4811
rect 10091 4777 10100 4811
rect 10048 4768 10100 4777
rect 10968 4768 11020 4820
rect 12900 4768 12952 4820
rect 13636 4811 13688 4820
rect 13636 4777 13645 4811
rect 13645 4777 13679 4811
rect 13679 4777 13688 4811
rect 13636 4768 13688 4777
rect 17224 4768 17276 4820
rect 18328 4811 18380 4820
rect 18328 4777 18337 4811
rect 18337 4777 18371 4811
rect 18371 4777 18380 4811
rect 18328 4768 18380 4777
rect 18604 4811 18656 4820
rect 18604 4777 18613 4811
rect 18613 4777 18647 4811
rect 18647 4777 18656 4811
rect 18604 4768 18656 4777
rect 18788 4811 18840 4820
rect 18788 4777 18797 4811
rect 18797 4777 18831 4811
rect 18831 4777 18840 4811
rect 18788 4768 18840 4777
rect 20536 4811 20588 4820
rect 20536 4777 20545 4811
rect 20545 4777 20579 4811
rect 20579 4777 20588 4811
rect 20536 4768 20588 4777
rect 21364 4768 21416 4820
rect 3884 4700 3936 4752
rect 4436 4700 4488 4752
rect 9956 4700 10008 4752
rect 2136 4632 2188 4684
rect 4068 4632 4120 4684
rect 4988 4632 5040 4684
rect 7196 4632 7248 4684
rect 7932 4675 7984 4684
rect 7932 4641 7941 4675
rect 7941 4641 7975 4675
rect 7975 4641 7984 4675
rect 7932 4632 7984 4641
rect 8208 4632 8260 4684
rect 14464 4700 14516 4752
rect 14924 4743 14976 4752
rect 14924 4709 14933 4743
rect 14933 4709 14967 4743
rect 14967 4709 14976 4743
rect 14924 4700 14976 4709
rect 16304 4700 16356 4752
rect 12348 4632 12400 4684
rect 13452 4632 13504 4684
rect 16212 4632 16264 4684
rect 19156 4675 19208 4684
rect 19156 4641 19165 4675
rect 19165 4641 19199 4675
rect 19199 4641 19208 4675
rect 19156 4632 19208 4641
rect 21456 4632 21508 4684
rect 22376 4675 22428 4684
rect 22376 4641 22385 4675
rect 22385 4641 22419 4675
rect 22419 4641 22428 4675
rect 22376 4632 22428 4641
rect 1952 4564 2004 4616
rect 2780 4564 2832 4616
rect 8116 4607 8168 4616
rect 8116 4573 8125 4607
rect 8125 4573 8159 4607
rect 8159 4573 8168 4607
rect 8116 4564 8168 4573
rect 10232 4607 10284 4616
rect 10232 4573 10241 4607
rect 10241 4573 10275 4607
rect 10275 4573 10284 4607
rect 10232 4564 10284 4573
rect 2688 4496 2740 4548
rect 9772 4496 9824 4548
rect 11980 4496 12032 4548
rect 13268 4564 13320 4616
rect 19248 4607 19300 4616
rect 15292 4496 15344 4548
rect 19248 4573 19257 4607
rect 19257 4573 19291 4607
rect 19291 4573 19300 4607
rect 19248 4564 19300 4573
rect 9680 4471 9732 4480
rect 9680 4437 9689 4471
rect 9689 4437 9723 4471
rect 9723 4437 9732 4471
rect 9680 4428 9732 4437
rect 10692 4471 10744 4480
rect 10692 4437 10701 4471
rect 10701 4437 10735 4471
rect 10735 4437 10744 4471
rect 10692 4428 10744 4437
rect 11152 4428 11204 4480
rect 12072 4428 12124 4480
rect 13176 4471 13228 4480
rect 13176 4437 13185 4471
rect 13185 4437 13219 4471
rect 13219 4437 13228 4471
rect 13176 4428 13228 4437
rect 14096 4428 14148 4480
rect 15844 4471 15896 4480
rect 15844 4437 15853 4471
rect 15853 4437 15887 4471
rect 15887 4437 15896 4471
rect 15844 4428 15896 4437
rect 16212 4471 16264 4480
rect 16212 4437 16221 4471
rect 16221 4437 16255 4471
rect 16255 4437 16264 4471
rect 16212 4428 16264 4437
rect 18972 4496 19024 4548
rect 23480 4564 23532 4616
rect 16580 4428 16632 4480
rect 20260 4471 20312 4480
rect 20260 4437 20269 4471
rect 20269 4437 20303 4471
rect 20303 4437 20312 4471
rect 20260 4428 20312 4437
rect 20628 4428 20680 4480
rect 23112 4428 23164 4480
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 2228 4088 2280 4140
rect 2780 4088 2832 4140
rect 4160 4088 4212 4140
rect 5264 4088 5316 4140
rect 6368 4224 6420 4276
rect 10048 4224 10100 4276
rect 7288 4131 7340 4140
rect 7288 4097 7297 4131
rect 7297 4097 7331 4131
rect 7331 4097 7340 4131
rect 7288 4088 7340 4097
rect 2320 4020 2372 4072
rect 3056 4020 3108 4072
rect 3424 4020 3476 4072
rect 8576 4088 8628 4140
rect 2136 3952 2188 4004
rect 2964 3952 3016 4004
rect 3792 3995 3844 4004
rect 3792 3961 3801 3995
rect 3801 3961 3835 3995
rect 3835 3961 3844 3995
rect 3792 3952 3844 3961
rect 5540 3995 5592 4004
rect 5540 3961 5549 3995
rect 5549 3961 5583 3995
rect 5583 3961 5592 3995
rect 5540 3952 5592 3961
rect 8116 4020 8168 4072
rect 11244 4063 11296 4072
rect 11244 4029 11253 4063
rect 11253 4029 11287 4063
rect 11287 4029 11296 4063
rect 13452 4267 13504 4276
rect 13452 4233 13461 4267
rect 13461 4233 13495 4267
rect 13495 4233 13504 4267
rect 13452 4224 13504 4233
rect 16396 4267 16448 4276
rect 16396 4233 16405 4267
rect 16405 4233 16439 4267
rect 16439 4233 16448 4267
rect 16396 4224 16448 4233
rect 19156 4267 19208 4276
rect 19156 4233 19165 4267
rect 19165 4233 19199 4267
rect 19199 4233 19208 4267
rect 19156 4224 19208 4233
rect 21456 4224 21508 4276
rect 22376 4267 22428 4276
rect 22376 4233 22385 4267
rect 22385 4233 22419 4267
rect 22419 4233 22428 4267
rect 22376 4224 22428 4233
rect 15844 4156 15896 4208
rect 15936 4088 15988 4140
rect 17224 4156 17276 4208
rect 18604 4156 18656 4208
rect 17132 4088 17184 4140
rect 17868 4131 17920 4140
rect 17868 4097 17877 4131
rect 17877 4097 17911 4131
rect 17911 4097 17920 4131
rect 17868 4088 17920 4097
rect 18420 4088 18472 4140
rect 11244 4020 11296 4029
rect 13452 4020 13504 4072
rect 13912 4020 13964 4072
rect 14372 4020 14424 4072
rect 15752 4020 15804 4072
rect 19984 4020 20036 4072
rect 20352 4020 20404 4072
rect 21824 4063 21876 4072
rect 21824 4029 21833 4063
rect 21833 4029 21867 4063
rect 21867 4029 21876 4063
rect 21824 4020 21876 4029
rect 23480 4020 23532 4072
rect 9496 3952 9548 4004
rect 10232 3952 10284 4004
rect 11060 3952 11112 4004
rect 11888 3952 11940 4004
rect 13268 3952 13320 4004
rect 14096 3995 14148 4004
rect 14096 3961 14108 3995
rect 14108 3961 14148 3995
rect 14096 3952 14148 3961
rect 16764 3995 16816 4004
rect 16764 3961 16773 3995
rect 16773 3961 16807 3995
rect 16807 3961 16816 3995
rect 16764 3952 16816 3961
rect 20260 3952 20312 4004
rect 1952 3884 2004 3936
rect 2320 3927 2372 3936
rect 2320 3893 2329 3927
rect 2329 3893 2363 3927
rect 2363 3893 2372 3927
rect 3424 3927 3476 3936
rect 2320 3884 2372 3893
rect 3424 3893 3433 3927
rect 3433 3893 3467 3927
rect 3467 3893 3476 3927
rect 3424 3884 3476 3893
rect 3884 3927 3936 3936
rect 3884 3893 3893 3927
rect 3893 3893 3927 3927
rect 3927 3893 3936 3927
rect 3884 3884 3936 3893
rect 5172 3927 5224 3936
rect 5172 3893 5181 3927
rect 5181 3893 5215 3927
rect 5215 3893 5224 3927
rect 5172 3884 5224 3893
rect 6644 3927 6696 3936
rect 6644 3893 6653 3927
rect 6653 3893 6687 3927
rect 6687 3893 6696 3927
rect 6644 3884 6696 3893
rect 6828 3927 6880 3936
rect 6828 3893 6837 3927
rect 6837 3893 6871 3927
rect 6871 3893 6880 3927
rect 6828 3884 6880 3893
rect 7196 3927 7248 3936
rect 7196 3893 7205 3927
rect 7205 3893 7239 3927
rect 7239 3893 7248 3927
rect 7196 3884 7248 3893
rect 8300 3927 8352 3936
rect 8300 3893 8309 3927
rect 8309 3893 8343 3927
rect 8343 3893 8352 3927
rect 8300 3884 8352 3893
rect 10048 3884 10100 3936
rect 11428 3927 11480 3936
rect 11428 3893 11437 3927
rect 11437 3893 11471 3927
rect 11471 3893 11480 3927
rect 11428 3884 11480 3893
rect 13636 3884 13688 3936
rect 13728 3884 13780 3936
rect 15200 3927 15252 3936
rect 15200 3893 15209 3927
rect 15209 3893 15243 3927
rect 15243 3893 15252 3927
rect 15200 3884 15252 3893
rect 17960 3884 18012 3936
rect 19248 3884 19300 3936
rect 19524 3927 19576 3936
rect 19524 3893 19533 3927
rect 19533 3893 19567 3927
rect 19567 3893 19576 3927
rect 19524 3884 19576 3893
rect 20076 3884 20128 3936
rect 22008 3927 22060 3936
rect 22008 3893 22017 3927
rect 22017 3893 22051 3927
rect 22051 3893 22060 3927
rect 22008 3884 22060 3893
rect 25320 3884 25372 3936
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 1952 3723 2004 3732
rect 1952 3689 1961 3723
rect 1961 3689 1995 3723
rect 1995 3689 2004 3723
rect 1952 3680 2004 3689
rect 2228 3723 2280 3732
rect 2228 3689 2237 3723
rect 2237 3689 2271 3723
rect 2271 3689 2280 3723
rect 2228 3680 2280 3689
rect 2412 3723 2464 3732
rect 2412 3689 2421 3723
rect 2421 3689 2455 3723
rect 2455 3689 2464 3723
rect 2412 3680 2464 3689
rect 3424 3680 3476 3732
rect 5172 3680 5224 3732
rect 7196 3680 7248 3732
rect 7932 3680 7984 3732
rect 8300 3680 8352 3732
rect 11244 3723 11296 3732
rect 11244 3689 11253 3723
rect 11253 3689 11287 3723
rect 11287 3689 11296 3723
rect 11244 3680 11296 3689
rect 12532 3680 12584 3732
rect 13176 3680 13228 3732
rect 13820 3680 13872 3732
rect 18328 3680 18380 3732
rect 18972 3680 19024 3732
rect 20168 3680 20220 3732
rect 20352 3723 20404 3732
rect 20352 3689 20361 3723
rect 20361 3689 20395 3723
rect 20395 3689 20404 3723
rect 20352 3680 20404 3689
rect 20720 3723 20772 3732
rect 20720 3689 20729 3723
rect 20729 3689 20763 3723
rect 20763 3689 20772 3723
rect 20720 3680 20772 3689
rect 21364 3680 21416 3732
rect 3148 3612 3200 3664
rect 4160 3612 4212 3664
rect 6368 3612 6420 3664
rect 4068 3587 4120 3596
rect 4068 3553 4077 3587
rect 4077 3553 4111 3587
rect 4111 3553 4120 3587
rect 4068 3544 4120 3553
rect 6736 3587 6788 3596
rect 6736 3553 6745 3587
rect 6745 3553 6779 3587
rect 6779 3553 6788 3587
rect 6736 3544 6788 3553
rect 7104 3544 7156 3596
rect 6092 3519 6144 3528
rect 2504 3408 2556 3460
rect 2872 3340 2924 3392
rect 3056 3340 3108 3392
rect 6092 3485 6101 3519
rect 6101 3485 6135 3519
rect 6135 3485 6144 3519
rect 6092 3476 6144 3485
rect 6828 3476 6880 3528
rect 10140 3612 10192 3664
rect 10876 3655 10928 3664
rect 10876 3621 10885 3655
rect 10885 3621 10919 3655
rect 10919 3621 10928 3655
rect 10876 3612 10928 3621
rect 15200 3612 15252 3664
rect 15936 3612 15988 3664
rect 8392 3587 8444 3596
rect 8392 3553 8401 3587
rect 8401 3553 8435 3587
rect 8435 3553 8444 3587
rect 8392 3544 8444 3553
rect 8760 3544 8812 3596
rect 10048 3544 10100 3596
rect 9680 3476 9732 3528
rect 11520 3544 11572 3596
rect 12440 3544 12492 3596
rect 13636 3544 13688 3596
rect 15292 3587 15344 3596
rect 15292 3553 15301 3587
rect 15301 3553 15335 3587
rect 15335 3553 15344 3587
rect 15292 3544 15344 3553
rect 19156 3587 19208 3596
rect 11796 3519 11848 3528
rect 6460 3408 6512 3460
rect 7104 3408 7156 3460
rect 11796 3485 11805 3519
rect 11805 3485 11839 3519
rect 11839 3485 11848 3519
rect 11796 3476 11848 3485
rect 12716 3476 12768 3528
rect 11060 3408 11112 3460
rect 12348 3408 12400 3460
rect 12900 3408 12952 3460
rect 13728 3408 13780 3460
rect 16304 3476 16356 3528
rect 19156 3553 19165 3587
rect 19165 3553 19199 3587
rect 19199 3553 19208 3587
rect 19156 3544 19208 3553
rect 19340 3587 19392 3596
rect 19340 3553 19349 3587
rect 19349 3553 19383 3587
rect 19383 3553 19392 3587
rect 19340 3544 19392 3553
rect 20904 3587 20956 3596
rect 20904 3553 20913 3587
rect 20913 3553 20947 3587
rect 20947 3553 20956 3587
rect 20904 3544 20956 3553
rect 16580 3408 16632 3460
rect 18604 3476 18656 3528
rect 4436 3340 4488 3392
rect 9496 3383 9548 3392
rect 9496 3349 9505 3383
rect 9505 3349 9539 3383
rect 9539 3349 9548 3383
rect 9496 3340 9548 3349
rect 12440 3340 12492 3392
rect 12716 3340 12768 3392
rect 13268 3383 13320 3392
rect 13268 3349 13277 3383
rect 13277 3349 13311 3383
rect 13311 3349 13320 3383
rect 13268 3340 13320 3349
rect 14556 3383 14608 3392
rect 14556 3349 14565 3383
rect 14565 3349 14599 3383
rect 14599 3349 14608 3383
rect 14556 3340 14608 3349
rect 14832 3340 14884 3392
rect 15476 3340 15528 3392
rect 16212 3340 16264 3392
rect 17592 3383 17644 3392
rect 17592 3349 17601 3383
rect 17601 3349 17635 3383
rect 17635 3349 17644 3383
rect 22100 3408 22152 3460
rect 19524 3383 19576 3392
rect 17592 3340 17644 3349
rect 19524 3349 19533 3383
rect 19533 3349 19567 3383
rect 19567 3349 19576 3383
rect 19524 3340 19576 3349
rect 20812 3340 20864 3392
rect 21824 3383 21876 3392
rect 21824 3349 21833 3383
rect 21833 3349 21867 3383
rect 21867 3349 21876 3383
rect 21824 3340 21876 3349
rect 22192 3383 22244 3392
rect 22192 3349 22201 3383
rect 22201 3349 22235 3383
rect 22235 3349 22244 3383
rect 22192 3340 22244 3349
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 2504 3179 2556 3188
rect 2504 3145 2513 3179
rect 2513 3145 2547 3179
rect 2547 3145 2556 3179
rect 2504 3136 2556 3145
rect 3884 3136 3936 3188
rect 6736 3136 6788 3188
rect 8392 3136 8444 3188
rect 9312 3179 9364 3188
rect 9312 3145 9321 3179
rect 9321 3145 9355 3179
rect 9355 3145 9364 3179
rect 9312 3136 9364 3145
rect 9496 3136 9548 3188
rect 11796 3136 11848 3188
rect 15936 3179 15988 3188
rect 15936 3145 15945 3179
rect 15945 3145 15979 3179
rect 15979 3145 15988 3179
rect 15936 3136 15988 3145
rect 16304 3179 16356 3188
rect 16304 3145 16313 3179
rect 16313 3145 16347 3179
rect 16347 3145 16356 3179
rect 16304 3136 16356 3145
rect 18328 3136 18380 3188
rect 19064 3179 19116 3188
rect 19064 3145 19073 3179
rect 19073 3145 19107 3179
rect 19107 3145 19116 3179
rect 19064 3136 19116 3145
rect 19340 3136 19392 3188
rect 1492 3068 1544 3120
rect 4160 3068 4212 3120
rect 5632 3111 5684 3120
rect 5632 3077 5641 3111
rect 5641 3077 5675 3111
rect 5675 3077 5684 3111
rect 5632 3068 5684 3077
rect 6368 3068 6420 3120
rect 5540 3000 5592 3052
rect 11520 3068 11572 3120
rect 9772 3043 9824 3052
rect 2412 2932 2464 2984
rect 4068 2932 4120 2984
rect 6828 2975 6880 2984
rect 6828 2941 6837 2975
rect 6837 2941 6871 2975
rect 6871 2941 6880 2975
rect 6828 2932 6880 2941
rect 9772 3009 9781 3043
rect 9781 3009 9815 3043
rect 9815 3009 9824 3043
rect 9772 3000 9824 3009
rect 9864 3000 9916 3052
rect 11152 3043 11204 3052
rect 11152 3009 11161 3043
rect 11161 3009 11195 3043
rect 11195 3009 11204 3043
rect 11152 3000 11204 3009
rect 15476 3043 15528 3052
rect 15476 3009 15485 3043
rect 15485 3009 15519 3043
rect 15519 3009 15528 3043
rect 15476 3000 15528 3009
rect 10692 2932 10744 2984
rect 10876 2975 10928 2984
rect 10876 2941 10885 2975
rect 10885 2941 10919 2975
rect 10919 2941 10928 2975
rect 10876 2932 10928 2941
rect 13452 2932 13504 2984
rect 13728 2932 13780 2984
rect 14556 2932 14608 2984
rect 16764 3043 16816 3052
rect 16764 3009 16773 3043
rect 16773 3009 16807 3043
rect 16807 3009 16816 3043
rect 16764 3000 16816 3009
rect 18604 3043 18656 3052
rect 18604 3009 18613 3043
rect 18613 3009 18647 3043
rect 18647 3009 18656 3043
rect 18604 3000 18656 3009
rect 20904 3136 20956 3188
rect 21732 3136 21784 3188
rect 22100 3136 22152 3188
rect 21364 3068 21416 3120
rect 3056 2864 3108 2916
rect 8208 2839 8260 2848
rect 8208 2805 8217 2839
rect 8217 2805 8251 2839
rect 8251 2805 8260 2839
rect 8208 2796 8260 2805
rect 8760 2839 8812 2848
rect 8760 2805 8769 2839
rect 8769 2805 8803 2839
rect 8803 2805 8812 2839
rect 8760 2796 8812 2805
rect 11612 2839 11664 2848
rect 11612 2805 11621 2839
rect 11621 2805 11655 2839
rect 11655 2805 11664 2839
rect 11612 2796 11664 2805
rect 12348 2864 12400 2916
rect 13176 2864 13228 2916
rect 14832 2864 14884 2916
rect 12440 2796 12492 2848
rect 13268 2796 13320 2848
rect 15108 2796 15160 2848
rect 19248 2932 19300 2984
rect 19340 2932 19392 2984
rect 20720 2932 20772 2984
rect 21732 2932 21784 2984
rect 17868 2907 17920 2916
rect 17868 2873 17877 2907
rect 17877 2873 17911 2907
rect 17911 2873 17920 2907
rect 17868 2864 17920 2873
rect 16580 2796 16632 2848
rect 18052 2839 18104 2848
rect 18052 2805 18061 2839
rect 18061 2805 18095 2839
rect 18095 2805 18104 2839
rect 18052 2796 18104 2805
rect 22468 2864 22520 2916
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 1676 2592 1728 2644
rect 2872 2635 2924 2644
rect 2872 2601 2881 2635
rect 2881 2601 2915 2635
rect 2915 2601 2924 2635
rect 2872 2592 2924 2601
rect 2964 2592 3016 2644
rect 3976 2592 4028 2644
rect 4712 2635 4764 2644
rect 4712 2601 4721 2635
rect 4721 2601 4755 2635
rect 4755 2601 4764 2635
rect 4712 2592 4764 2601
rect 6644 2592 6696 2644
rect 8208 2592 8260 2644
rect 9956 2592 10008 2644
rect 10968 2592 11020 2644
rect 11060 2592 11112 2644
rect 13176 2635 13228 2644
rect 13176 2601 13185 2635
rect 13185 2601 13219 2635
rect 13219 2601 13228 2635
rect 13176 2592 13228 2601
rect 13820 2592 13872 2644
rect 15200 2635 15252 2644
rect 15200 2601 15209 2635
rect 15209 2601 15243 2635
rect 15243 2601 15252 2635
rect 16580 2635 16632 2644
rect 15200 2592 15252 2601
rect 11244 2524 11296 2576
rect 3608 2456 3660 2508
rect 5172 2499 5224 2508
rect 5172 2465 5181 2499
rect 5181 2465 5215 2499
rect 5215 2465 5224 2499
rect 5172 2456 5224 2465
rect 6092 2456 6144 2508
rect 6828 2456 6880 2508
rect 8576 2456 8628 2508
rect 3056 2431 3108 2440
rect 3056 2397 3065 2431
rect 3065 2397 3099 2431
rect 3099 2397 3108 2431
rect 3056 2388 3108 2397
rect 6368 2431 6420 2440
rect 6368 2397 6377 2431
rect 6377 2397 6411 2431
rect 6411 2397 6420 2431
rect 6368 2388 6420 2397
rect 12072 2456 12124 2508
rect 13544 2499 13596 2508
rect 13544 2465 13553 2499
rect 13553 2465 13587 2499
rect 13587 2465 13596 2499
rect 13544 2456 13596 2465
rect 15844 2499 15896 2508
rect 5264 2363 5316 2372
rect 5264 2329 5273 2363
rect 5273 2329 5307 2363
rect 5307 2329 5316 2363
rect 5264 2320 5316 2329
rect 13728 2431 13780 2440
rect 13728 2397 13737 2431
rect 13737 2397 13771 2431
rect 13771 2397 13780 2431
rect 13728 2388 13780 2397
rect 9864 2320 9916 2372
rect 11244 2363 11296 2372
rect 11244 2329 11253 2363
rect 11253 2329 11287 2363
rect 11287 2329 11296 2363
rect 11244 2320 11296 2329
rect 12348 2320 12400 2372
rect 15844 2465 15853 2499
rect 15853 2465 15887 2499
rect 15887 2465 15896 2499
rect 15844 2456 15896 2465
rect 16580 2601 16589 2635
rect 16589 2601 16623 2635
rect 16623 2601 16632 2635
rect 16580 2592 16632 2601
rect 18144 2635 18196 2644
rect 18144 2601 18153 2635
rect 18153 2601 18187 2635
rect 18187 2601 18196 2635
rect 18144 2592 18196 2601
rect 22008 2592 22060 2644
rect 22100 2635 22152 2644
rect 22100 2601 22109 2635
rect 22109 2601 22143 2635
rect 22143 2601 22152 2635
rect 22100 2592 22152 2601
rect 16120 2524 16172 2576
rect 18052 2524 18104 2576
rect 19892 2499 19944 2508
rect 14648 2320 14700 2372
rect 17040 2388 17092 2440
rect 19892 2465 19901 2499
rect 19901 2465 19935 2499
rect 19935 2465 19944 2499
rect 19892 2456 19944 2465
rect 21180 2499 21232 2508
rect 21180 2465 21189 2499
rect 21189 2465 21223 2499
rect 21223 2465 21232 2499
rect 21180 2456 21232 2465
rect 22284 2499 22336 2508
rect 22284 2465 22293 2499
rect 22293 2465 22327 2499
rect 22327 2465 22336 2499
rect 22284 2456 22336 2465
rect 24032 2499 24084 2508
rect 24032 2465 24041 2499
rect 24041 2465 24075 2499
rect 24075 2465 24084 2499
rect 24032 2456 24084 2465
rect 16488 2320 16540 2372
rect 17316 2363 17368 2372
rect 17316 2329 17325 2363
rect 17325 2329 17359 2363
rect 17359 2329 17368 2363
rect 17316 2320 17368 2329
rect 18604 2320 18656 2372
rect 21916 2320 21968 2372
rect 23664 2320 23716 2372
rect 18328 2295 18380 2304
rect 18328 2261 18337 2295
rect 18337 2261 18371 2295
rect 18371 2261 18380 2295
rect 18328 2252 18380 2261
rect 20720 2252 20772 2304
rect 23480 2252 23532 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 6000 552 6052 604
rect 6184 552 6236 604
<< metal2 >>
rect 294 27520 350 28000
rect 846 27520 902 28000
rect 1398 27520 1454 28000
rect 1950 27520 2006 28000
rect 2502 27520 2558 28000
rect 3146 27520 3202 28000
rect 3514 27704 3570 27713
rect 3514 27639 3570 27648
rect 308 21049 336 27520
rect 294 21040 350 21049
rect 294 20975 350 20984
rect 860 17746 888 27520
rect 1412 19394 1440 27520
rect 1964 26874 1992 27520
rect 2516 26874 2544 27520
rect 1872 26846 1992 26874
rect 2332 26846 2544 26874
rect 1584 25356 1636 25362
rect 1584 25298 1636 25304
rect 1596 24750 1624 25298
rect 1584 24744 1636 24750
rect 1584 24686 1636 24692
rect 1766 24712 1822 24721
rect 1766 24647 1768 24656
rect 1820 24647 1822 24656
rect 1768 24618 1820 24624
rect 1766 24304 1822 24313
rect 1676 24268 1728 24274
rect 1766 24239 1822 24248
rect 1676 24210 1728 24216
rect 1688 23322 1716 24210
rect 1780 23730 1808 24239
rect 1768 23724 1820 23730
rect 1768 23666 1820 23672
rect 1676 23316 1728 23322
rect 1676 23258 1728 23264
rect 1584 22092 1636 22098
rect 1584 22034 1636 22040
rect 1596 22001 1624 22034
rect 1582 21992 1638 22001
rect 1582 21927 1638 21936
rect 1596 21146 1624 21927
rect 1768 21344 1820 21350
rect 1768 21286 1820 21292
rect 1584 21140 1636 21146
rect 1584 21082 1636 21088
rect 1674 20904 1730 20913
rect 1674 20839 1730 20848
rect 1688 20602 1716 20839
rect 1676 20596 1728 20602
rect 1676 20538 1728 20544
rect 1688 20398 1716 20538
rect 1780 20505 1808 21286
rect 1766 20496 1822 20505
rect 1766 20431 1822 20440
rect 1676 20392 1728 20398
rect 1676 20334 1728 20340
rect 1412 19366 1624 19394
rect 1400 19304 1452 19310
rect 1400 19246 1452 19252
rect 1490 19272 1546 19281
rect 1412 18970 1440 19246
rect 1490 19207 1546 19216
rect 1504 19174 1532 19207
rect 1492 19168 1544 19174
rect 1492 19110 1544 19116
rect 1400 18964 1452 18970
rect 1400 18906 1452 18912
rect 1400 18760 1452 18766
rect 1400 18702 1452 18708
rect 848 17740 900 17746
rect 848 17682 900 17688
rect 1412 14074 1440 18702
rect 1492 18216 1544 18222
rect 1492 18158 1544 18164
rect 1504 16658 1532 18158
rect 1492 16652 1544 16658
rect 1492 16594 1544 16600
rect 1504 15026 1532 16594
rect 1596 16425 1624 19366
rect 1768 18828 1820 18834
rect 1768 18770 1820 18776
rect 1676 17536 1728 17542
rect 1676 17478 1728 17484
rect 1688 17066 1716 17478
rect 1780 17338 1808 18770
rect 1872 18086 1900 26846
rect 2044 25424 2096 25430
rect 2044 25366 2096 25372
rect 1950 24576 2006 24585
rect 1950 24511 2006 24520
rect 1964 24342 1992 24511
rect 1952 24336 2004 24342
rect 1952 24278 2004 24284
rect 2056 22642 2084 25366
rect 2136 25152 2188 25158
rect 2136 25094 2188 25100
rect 2148 24818 2176 25094
rect 2136 24812 2188 24818
rect 2136 24754 2188 24760
rect 2044 22636 2096 22642
rect 2044 22578 2096 22584
rect 2042 21584 2098 21593
rect 2042 21519 2098 21528
rect 1952 21004 2004 21010
rect 1952 20946 2004 20952
rect 1964 20602 1992 20946
rect 1952 20596 2004 20602
rect 1952 20538 2004 20544
rect 2056 20466 2084 21519
rect 2148 21457 2176 24754
rect 2228 24268 2280 24274
rect 2228 24210 2280 24216
rect 2240 21554 2268 24210
rect 2228 21548 2280 21554
rect 2228 21490 2280 21496
rect 2134 21448 2190 21457
rect 2134 21383 2190 21392
rect 2044 20460 2096 20466
rect 2044 20402 2096 20408
rect 2228 19848 2280 19854
rect 2226 19816 2228 19825
rect 2280 19816 2282 19825
rect 2226 19751 2282 19760
rect 1952 19712 2004 19718
rect 1952 19654 2004 19660
rect 1964 19174 1992 19654
rect 1952 19168 2004 19174
rect 1952 19110 2004 19116
rect 1860 18080 1912 18086
rect 1860 18022 1912 18028
rect 1860 17672 1912 17678
rect 1860 17614 1912 17620
rect 1768 17332 1820 17338
rect 1768 17274 1820 17280
rect 1676 17060 1728 17066
rect 1676 17002 1728 17008
rect 1582 16416 1638 16425
rect 1582 16351 1638 16360
rect 1492 15020 1544 15026
rect 1492 14962 1544 14968
rect 1688 14618 1716 17002
rect 1872 16998 1900 17614
rect 1860 16992 1912 16998
rect 1860 16934 1912 16940
rect 1768 16108 1820 16114
rect 1768 16050 1820 16056
rect 1780 15706 1808 16050
rect 1768 15700 1820 15706
rect 1768 15642 1820 15648
rect 1676 14612 1728 14618
rect 1676 14554 1728 14560
rect 1768 14272 1820 14278
rect 1768 14214 1820 14220
rect 1400 14068 1452 14074
rect 1400 14010 1452 14016
rect 1780 13734 1808 14214
rect 1768 13728 1820 13734
rect 1768 13670 1820 13676
rect 1398 13288 1454 13297
rect 1398 13223 1454 13232
rect 1412 12986 1440 13223
rect 1582 13152 1638 13161
rect 1582 13087 1638 13096
rect 1400 12980 1452 12986
rect 1400 12922 1452 12928
rect 1596 12356 1624 13087
rect 1780 12900 1808 13670
rect 1872 13161 1900 16934
rect 1964 15434 1992 19110
rect 2044 17604 2096 17610
rect 2044 17546 2096 17552
rect 2056 17202 2084 17546
rect 2044 17196 2096 17202
rect 2096 17156 2176 17184
rect 2044 17138 2096 17144
rect 2044 15904 2096 15910
rect 2044 15846 2096 15852
rect 2056 15609 2084 15846
rect 2042 15600 2098 15609
rect 2042 15535 2098 15544
rect 1952 15428 2004 15434
rect 1952 15370 2004 15376
rect 2148 14890 2176 17156
rect 2332 15978 2360 26846
rect 3056 25492 3108 25498
rect 3056 25434 3108 25440
rect 2596 25356 2648 25362
rect 2596 25298 2648 25304
rect 2504 24676 2556 24682
rect 2504 24618 2556 24624
rect 2410 23896 2466 23905
rect 2410 23831 2412 23840
rect 2464 23831 2466 23840
rect 2412 23802 2464 23808
rect 2412 23180 2464 23186
rect 2412 23122 2464 23128
rect 2424 22778 2452 23122
rect 2412 22772 2464 22778
rect 2412 22714 2464 22720
rect 2516 22658 2544 24618
rect 2608 24614 2636 25298
rect 2872 25288 2924 25294
rect 2872 25230 2924 25236
rect 2688 24744 2740 24750
rect 2688 24686 2740 24692
rect 2596 24608 2648 24614
rect 2596 24550 2648 24556
rect 2424 22630 2544 22658
rect 2424 22098 2452 22630
rect 2412 22092 2464 22098
rect 2412 22034 2464 22040
rect 2608 21078 2636 24550
rect 2700 23769 2728 24686
rect 2884 24410 2912 25230
rect 2964 24744 3016 24750
rect 2964 24686 3016 24692
rect 2872 24404 2924 24410
rect 2872 24346 2924 24352
rect 2686 23760 2742 23769
rect 2686 23695 2742 23704
rect 2688 23520 2740 23526
rect 2688 23462 2740 23468
rect 2700 22778 2728 23462
rect 2872 23112 2924 23118
rect 2872 23054 2924 23060
rect 2780 23044 2832 23050
rect 2780 22986 2832 22992
rect 2688 22772 2740 22778
rect 2688 22714 2740 22720
rect 2700 22574 2728 22714
rect 2792 22574 2820 22986
rect 2884 22710 2912 23054
rect 2872 22704 2924 22710
rect 2872 22646 2924 22652
rect 2688 22568 2740 22574
rect 2688 22510 2740 22516
rect 2780 22568 2832 22574
rect 2780 22510 2832 22516
rect 2792 22420 2820 22510
rect 2872 22500 2924 22506
rect 2872 22442 2924 22448
rect 2700 22392 2820 22420
rect 2700 22098 2728 22392
rect 2688 22092 2740 22098
rect 2688 22034 2740 22040
rect 2780 22092 2832 22098
rect 2780 22034 2832 22040
rect 2792 21690 2820 22034
rect 2780 21684 2832 21690
rect 2780 21626 2832 21632
rect 2792 21298 2820 21626
rect 2700 21270 2820 21298
rect 2596 21072 2648 21078
rect 2596 21014 2648 21020
rect 2504 20596 2556 20602
rect 2504 20538 2556 20544
rect 2516 20369 2544 20538
rect 2502 20360 2558 20369
rect 2700 20346 2728 21270
rect 2884 20777 2912 22442
rect 2870 20768 2926 20777
rect 2870 20703 2926 20712
rect 2502 20295 2558 20304
rect 2608 20318 2728 20346
rect 2608 19990 2636 20318
rect 2872 20256 2924 20262
rect 2686 20224 2742 20233
rect 2872 20198 2924 20204
rect 2686 20159 2742 20168
rect 2596 19984 2648 19990
rect 2596 19926 2648 19932
rect 2700 19922 2728 20159
rect 2688 19916 2740 19922
rect 2688 19858 2740 19864
rect 2780 19916 2832 19922
rect 2780 19858 2832 19864
rect 2596 19712 2648 19718
rect 2596 19654 2648 19660
rect 2504 19304 2556 19310
rect 2608 19292 2636 19654
rect 2556 19264 2636 19292
rect 2504 19246 2556 19252
rect 2688 19168 2740 19174
rect 2688 19110 2740 19116
rect 2504 18624 2556 18630
rect 2504 18566 2556 18572
rect 2412 17740 2464 17746
rect 2412 17682 2464 17688
rect 2424 17338 2452 17682
rect 2412 17332 2464 17338
rect 2412 17274 2464 17280
rect 2516 16658 2544 18566
rect 2700 18154 2728 19110
rect 2792 18970 2820 19858
rect 2780 18964 2832 18970
rect 2780 18906 2832 18912
rect 2688 18148 2740 18154
rect 2740 18108 2820 18136
rect 2688 18090 2740 18096
rect 2594 18048 2650 18057
rect 2594 17983 2650 17992
rect 2504 16652 2556 16658
rect 2504 16594 2556 16600
rect 2502 16144 2558 16153
rect 2502 16079 2558 16088
rect 2412 16040 2464 16046
rect 2412 15982 2464 15988
rect 2320 15972 2372 15978
rect 2320 15914 2372 15920
rect 2424 15706 2452 15982
rect 2516 15978 2544 16079
rect 2504 15972 2556 15978
rect 2504 15914 2556 15920
rect 2412 15700 2464 15706
rect 2412 15642 2464 15648
rect 2410 15192 2466 15201
rect 2410 15127 2466 15136
rect 2136 14884 2188 14890
rect 2136 14826 2188 14832
rect 2148 14346 2176 14826
rect 2424 14618 2452 15127
rect 2412 14612 2464 14618
rect 2412 14554 2464 14560
rect 2136 14340 2188 14346
rect 2136 14282 2188 14288
rect 2148 13938 2176 14282
rect 2502 13968 2558 13977
rect 2136 13932 2188 13938
rect 2502 13903 2558 13912
rect 2136 13874 2188 13880
rect 2320 13728 2372 13734
rect 2320 13670 2372 13676
rect 2410 13696 2466 13705
rect 2042 13424 2098 13433
rect 2042 13359 2044 13368
rect 2096 13359 2098 13368
rect 2044 13330 2096 13336
rect 1858 13152 1914 13161
rect 1858 13087 1914 13096
rect 1780 12872 1900 12900
rect 1596 12328 1716 12356
rect 1400 11552 1452 11558
rect 1400 11494 1452 11500
rect 1412 9602 1440 11494
rect 1492 11212 1544 11218
rect 1492 11154 1544 11160
rect 1320 9574 1440 9602
rect 1320 9330 1348 9574
rect 1400 9512 1452 9518
rect 1398 9480 1400 9489
rect 1452 9480 1454 9489
rect 1398 9415 1454 9424
rect 1320 9302 1440 9330
rect 1308 7812 1360 7818
rect 1308 7754 1360 7760
rect 1124 7200 1176 7206
rect 1124 7142 1176 7148
rect 1136 4457 1164 7142
rect 1122 4448 1178 4457
rect 1122 4383 1178 4392
rect 846 2136 902 2145
rect 846 2071 902 2080
rect 294 1728 350 1737
rect 294 1663 350 1672
rect 308 480 336 1663
rect 860 480 888 2071
rect 1320 921 1348 7754
rect 1412 3482 1440 9302
rect 1504 9081 1532 11154
rect 1584 10464 1636 10470
rect 1584 10406 1636 10412
rect 1596 9625 1624 10406
rect 1582 9616 1638 9625
rect 1582 9551 1638 9560
rect 1490 9072 1546 9081
rect 1490 9007 1546 9016
rect 1504 6934 1532 9007
rect 1688 7546 1716 12328
rect 1768 12300 1820 12306
rect 1768 12242 1820 12248
rect 1780 11354 1808 12242
rect 1768 11348 1820 11354
rect 1768 11290 1820 11296
rect 1872 11218 1900 12872
rect 2056 12714 2084 13330
rect 2332 13190 2360 13670
rect 2410 13631 2466 13640
rect 2424 13530 2452 13631
rect 2412 13524 2464 13530
rect 2412 13466 2464 13472
rect 2320 13184 2372 13190
rect 2320 13126 2372 13132
rect 2044 12708 2096 12714
rect 2044 12650 2096 12656
rect 2044 12368 2096 12374
rect 2044 12310 2096 12316
rect 2056 11694 2084 12310
rect 2044 11688 2096 11694
rect 2044 11630 2096 11636
rect 1860 11212 1912 11218
rect 1860 11154 1912 11160
rect 2056 10606 2084 11630
rect 2136 11076 2188 11082
rect 2136 11018 2188 11024
rect 2044 10600 2096 10606
rect 2044 10542 2096 10548
rect 1860 10464 1912 10470
rect 2044 10464 2096 10470
rect 1860 10406 1912 10412
rect 2042 10432 2044 10441
rect 2096 10432 2098 10441
rect 1872 10305 1900 10406
rect 2042 10367 2098 10376
rect 1858 10296 1914 10305
rect 1858 10231 1914 10240
rect 1872 8634 1900 10231
rect 1952 9920 2004 9926
rect 1952 9862 2004 9868
rect 1964 8673 1992 9862
rect 2044 9580 2096 9586
rect 2044 9522 2096 9528
rect 2056 9042 2084 9522
rect 2044 9036 2096 9042
rect 2044 8978 2096 8984
rect 1950 8664 2006 8673
rect 1860 8628 1912 8634
rect 1950 8599 2006 8608
rect 1860 8570 1912 8576
rect 1964 8498 1992 8599
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 1676 7540 1728 7546
rect 1676 7482 1728 7488
rect 1584 7404 1636 7410
rect 1584 7346 1636 7352
rect 1492 6928 1544 6934
rect 1492 6870 1544 6876
rect 1596 6322 1624 7346
rect 1688 7002 1716 7482
rect 1766 7440 1822 7449
rect 2056 7410 2084 8978
rect 1766 7375 1822 7384
rect 2044 7404 2096 7410
rect 1676 6996 1728 7002
rect 1676 6938 1728 6944
rect 1780 6882 1808 7375
rect 2044 7346 2096 7352
rect 1688 6854 1808 6882
rect 1584 6316 1636 6322
rect 1584 6258 1636 6264
rect 1596 5778 1624 6258
rect 1584 5772 1636 5778
rect 1584 5714 1636 5720
rect 1688 5250 1716 6854
rect 1768 6724 1820 6730
rect 1768 6666 1820 6672
rect 1780 5846 1808 6666
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 1872 5846 1900 6598
rect 1952 6180 2004 6186
rect 1952 6122 2004 6128
rect 1768 5840 1820 5846
rect 1768 5782 1820 5788
rect 1860 5840 1912 5846
rect 1860 5782 1912 5788
rect 1780 5302 1808 5782
rect 1504 5222 1716 5250
rect 1768 5296 1820 5302
rect 1768 5238 1820 5244
rect 1504 4706 1532 5222
rect 1872 5166 1900 5782
rect 1964 5234 1992 6122
rect 1952 5228 2004 5234
rect 1952 5170 2004 5176
rect 1860 5160 1912 5166
rect 1860 5102 1912 5108
rect 1676 5092 1728 5098
rect 1676 5034 1728 5040
rect 1688 4826 1716 5034
rect 1858 4992 1914 5001
rect 1858 4927 1914 4936
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1504 4678 1716 4706
rect 1412 3454 1532 3482
rect 1398 3360 1454 3369
rect 1398 3295 1454 3304
rect 1306 912 1362 921
rect 1306 847 1362 856
rect 1412 480 1440 3295
rect 1504 3126 1532 3454
rect 1492 3120 1544 3126
rect 1492 3062 1544 3068
rect 1688 2650 1716 4678
rect 1676 2644 1728 2650
rect 1676 2586 1728 2592
rect 1872 626 1900 4927
rect 1964 4622 1992 5170
rect 2148 4808 2176 11018
rect 2228 10668 2280 10674
rect 2228 10610 2280 10616
rect 2240 9994 2268 10610
rect 2228 9988 2280 9994
rect 2228 9930 2280 9936
rect 2228 9104 2280 9110
rect 2228 9046 2280 9052
rect 2240 8498 2268 9046
rect 2228 8492 2280 8498
rect 2228 8434 2280 8440
rect 2240 8090 2268 8434
rect 2228 8084 2280 8090
rect 2228 8026 2280 8032
rect 2332 7834 2360 13126
rect 2412 11620 2464 11626
rect 2412 11562 2464 11568
rect 2424 9330 2452 11562
rect 2516 9518 2544 13903
rect 2608 12986 2636 17983
rect 2792 16794 2820 18108
rect 2780 16788 2832 16794
rect 2780 16730 2832 16736
rect 2700 16510 2820 16538
rect 2700 16425 2728 16510
rect 2686 16416 2742 16425
rect 2686 16351 2742 16360
rect 2792 15881 2820 16510
rect 2778 15872 2834 15881
rect 2778 15807 2834 15816
rect 2686 15464 2742 15473
rect 2686 15399 2742 15408
rect 2596 12980 2648 12986
rect 2596 12922 2648 12928
rect 2700 12753 2728 15399
rect 2792 14482 2820 15807
rect 2780 14476 2832 14482
rect 2780 14418 2832 14424
rect 2792 14006 2820 14418
rect 2780 14000 2832 14006
rect 2884 13977 2912 20198
rect 2976 19990 3004 24686
rect 3068 22506 3096 25434
rect 3160 24698 3188 27520
rect 3528 27266 3556 27639
rect 3698 27520 3754 28000
rect 4250 27520 4306 28000
rect 4802 27520 4858 28000
rect 5354 27520 5410 28000
rect 5998 27520 6054 28000
rect 6550 27520 6606 28000
rect 7102 27520 7158 28000
rect 7654 27520 7710 28000
rect 8206 27520 8262 28000
rect 8850 27520 8906 28000
rect 9402 27520 9458 28000
rect 9954 27520 10010 28000
rect 10506 27520 10562 28000
rect 11058 27520 11114 28000
rect 11702 27520 11758 28000
rect 12254 27520 12310 28000
rect 12806 27520 12862 28000
rect 13358 27520 13414 28000
rect 13910 27520 13966 28000
rect 14554 27520 14610 28000
rect 15106 27520 15162 28000
rect 15658 27520 15714 28000
rect 16210 27520 16266 28000
rect 16762 27520 16818 28000
rect 17406 27520 17462 28000
rect 17958 27520 18014 28000
rect 18510 27520 18566 28000
rect 19062 27520 19118 28000
rect 19614 27520 19670 28000
rect 20258 27520 20314 28000
rect 20810 27520 20866 28000
rect 21362 27520 21418 28000
rect 21914 27520 21970 28000
rect 22466 27520 22522 28000
rect 23110 27520 23166 28000
rect 23662 27520 23718 28000
rect 24214 27520 24270 28000
rect 24766 27520 24822 28000
rect 25318 27520 25374 28000
rect 25962 27520 26018 28000
rect 26514 27520 26570 28000
rect 27066 27520 27122 28000
rect 27618 27520 27674 28000
rect 3516 27260 3568 27266
rect 3516 27202 3568 27208
rect 3514 27160 3570 27169
rect 3514 27095 3570 27104
rect 3528 26314 3556 27095
rect 3516 26308 3568 26314
rect 3516 26250 3568 26256
rect 3330 25392 3386 25401
rect 3330 25327 3386 25336
rect 3344 24954 3372 25327
rect 3516 25152 3568 25158
rect 3516 25094 3568 25100
rect 3332 24948 3384 24954
rect 3332 24890 3384 24896
rect 3160 24670 3372 24698
rect 3240 24608 3292 24614
rect 3240 24550 3292 24556
rect 3148 24404 3200 24410
rect 3148 24346 3200 24352
rect 3056 22500 3108 22506
rect 3056 22442 3108 22448
rect 3056 21888 3108 21894
rect 3160 21865 3188 24346
rect 3056 21830 3108 21836
rect 3146 21856 3202 21865
rect 2964 19984 3016 19990
rect 2964 19926 3016 19932
rect 3068 19553 3096 21830
rect 3146 21791 3202 21800
rect 3252 21321 3280 24550
rect 3344 24290 3372 24670
rect 3344 24262 3464 24290
rect 3332 24200 3384 24206
rect 3332 24142 3384 24148
rect 3344 23866 3372 24142
rect 3332 23860 3384 23866
rect 3332 23802 3384 23808
rect 3344 23118 3372 23802
rect 3332 23112 3384 23118
rect 3332 23054 3384 23060
rect 3332 22432 3384 22438
rect 3332 22374 3384 22380
rect 3344 22166 3372 22374
rect 3332 22160 3384 22166
rect 3436 22148 3464 24262
rect 3528 24177 3556 25094
rect 3514 24168 3570 24177
rect 3514 24103 3570 24112
rect 3516 22976 3568 22982
rect 3516 22918 3568 22924
rect 3528 22438 3556 22918
rect 3606 22672 3662 22681
rect 3606 22607 3608 22616
rect 3660 22607 3662 22616
rect 3608 22578 3660 22584
rect 3516 22432 3568 22438
rect 3516 22374 3568 22380
rect 3332 22102 3384 22108
rect 3427 22120 3464 22148
rect 3344 21554 3372 22102
rect 3427 22080 3455 22120
rect 3427 22052 3464 22080
rect 3436 22012 3464 22052
rect 3436 21984 3556 22012
rect 3332 21548 3384 21554
rect 3332 21490 3384 21496
rect 3424 21344 3476 21350
rect 3238 21312 3294 21321
rect 3424 21286 3476 21292
rect 3238 21247 3294 21256
rect 3330 21040 3386 21049
rect 3330 20975 3386 20984
rect 3240 20256 3292 20262
rect 3240 20198 3292 20204
rect 3054 19544 3110 19553
rect 3054 19479 3110 19488
rect 3148 19304 3200 19310
rect 3148 19246 3200 19252
rect 3056 19168 3108 19174
rect 3056 19110 3108 19116
rect 3068 18086 3096 19110
rect 3160 18222 3188 19246
rect 3252 19009 3280 20198
rect 3238 19000 3294 19009
rect 3238 18935 3294 18944
rect 3148 18216 3200 18222
rect 3148 18158 3200 18164
rect 2964 18080 3016 18086
rect 2964 18022 3016 18028
rect 3056 18080 3108 18086
rect 3056 18022 3108 18028
rect 2976 17882 3004 18022
rect 2964 17876 3016 17882
rect 2964 17818 3016 17824
rect 2964 17740 3016 17746
rect 2964 17682 3016 17688
rect 2976 17649 3004 17682
rect 3068 17678 3096 18022
rect 3148 17876 3200 17882
rect 3148 17818 3200 17824
rect 3056 17672 3108 17678
rect 2962 17640 3018 17649
rect 3056 17614 3108 17620
rect 2962 17575 3018 17584
rect 3068 17338 3096 17614
rect 3056 17332 3108 17338
rect 3056 17274 3108 17280
rect 3160 17270 3188 17818
rect 3148 17264 3200 17270
rect 2962 17232 3018 17241
rect 3148 17206 3200 17212
rect 2962 17167 3018 17176
rect 2976 14498 3004 17167
rect 3056 16652 3108 16658
rect 3056 16594 3108 16600
rect 3068 16454 3096 16594
rect 3056 16448 3108 16454
rect 3056 16390 3108 16396
rect 3068 15502 3096 16390
rect 3160 15638 3188 17206
rect 3148 15632 3200 15638
rect 3148 15574 3200 15580
rect 3240 15564 3292 15570
rect 3240 15506 3292 15512
rect 3056 15496 3108 15502
rect 3056 15438 3108 15444
rect 3068 14822 3096 15438
rect 3252 15162 3280 15506
rect 3240 15156 3292 15162
rect 3240 15098 3292 15104
rect 3056 14816 3108 14822
rect 3056 14758 3108 14764
rect 3068 14618 3096 14758
rect 3056 14612 3108 14618
rect 3056 14554 3108 14560
rect 3344 14550 3372 20975
rect 3148 14544 3200 14550
rect 2976 14470 3096 14498
rect 3148 14486 3200 14492
rect 3332 14544 3384 14550
rect 3332 14486 3384 14492
rect 2780 13942 2832 13948
rect 2870 13968 2926 13977
rect 2870 13903 2926 13912
rect 2964 13864 3016 13870
rect 2964 13806 3016 13812
rect 2976 13705 3004 13806
rect 2962 13696 3018 13705
rect 2962 13631 3018 13640
rect 2964 13320 3016 13326
rect 2964 13262 3016 13268
rect 2976 12986 3004 13262
rect 2964 12980 3016 12986
rect 2884 12940 2964 12968
rect 2686 12744 2742 12753
rect 2686 12679 2742 12688
rect 2884 12442 2912 12940
rect 2964 12922 3016 12928
rect 3068 12866 3096 14470
rect 3160 14074 3188 14486
rect 3148 14068 3200 14074
rect 3148 14010 3200 14016
rect 3240 13864 3292 13870
rect 3238 13832 3240 13841
rect 3292 13832 3294 13841
rect 3238 13767 3294 13776
rect 3436 13716 3464 21286
rect 3528 17377 3556 21984
rect 3712 19990 3740 27520
rect 4066 26616 4122 26625
rect 4066 26551 4068 26560
rect 4120 26551 4122 26560
rect 4068 26522 4120 26528
rect 4066 25936 4122 25945
rect 4066 25871 4122 25880
rect 4080 25498 4108 25871
rect 4068 25492 4120 25498
rect 4068 25434 4120 25440
rect 4068 25220 4120 25226
rect 4068 25162 4120 25168
rect 4080 24857 4108 25162
rect 4066 24848 4122 24857
rect 4066 24783 4122 24792
rect 4068 24608 4120 24614
rect 4068 24550 4120 24556
rect 3976 24064 4028 24070
rect 3976 24006 4028 24012
rect 3884 23112 3936 23118
rect 3884 23054 3936 23060
rect 3896 21894 3924 23054
rect 3988 22545 4016 24006
rect 4080 23633 4108 24550
rect 4066 23624 4122 23633
rect 4066 23559 4122 23568
rect 4068 23520 4120 23526
rect 4120 23480 4200 23508
rect 4068 23462 4120 23468
rect 4172 22642 4200 23480
rect 4160 22636 4212 22642
rect 4160 22578 4212 22584
rect 3974 22536 4030 22545
rect 3974 22471 4030 22480
rect 4068 22432 4120 22438
rect 4120 22392 4200 22420
rect 4068 22374 4120 22380
rect 3884 21888 3936 21894
rect 3884 21830 3936 21836
rect 3896 21010 3924 21830
rect 4172 21690 4200 22392
rect 4160 21684 4212 21690
rect 4160 21626 4212 21632
rect 3884 21004 3936 21010
rect 3884 20946 3936 20952
rect 3896 20058 3924 20946
rect 3884 20052 3936 20058
rect 3884 19994 3936 20000
rect 3700 19984 3752 19990
rect 3700 19926 3752 19932
rect 3608 17536 3660 17542
rect 3608 17478 3660 17484
rect 3514 17368 3570 17377
rect 3514 17303 3570 17312
rect 3528 16998 3556 17303
rect 3620 17134 3648 17478
rect 3608 17128 3660 17134
rect 3608 17070 3660 17076
rect 3516 16992 3568 16998
rect 3516 16934 3568 16940
rect 3528 16794 3556 16934
rect 3516 16788 3568 16794
rect 3712 16776 3740 19926
rect 3896 19310 3924 19994
rect 3884 19304 3936 19310
rect 3884 19246 3936 19252
rect 4264 19145 4292 27520
rect 4436 25356 4488 25362
rect 4436 25298 4488 25304
rect 4448 24614 4476 25298
rect 4436 24608 4488 24614
rect 4436 24550 4488 24556
rect 4344 23520 4396 23526
rect 4344 23462 4396 23468
rect 4356 23186 4384 23462
rect 4344 23180 4396 23186
rect 4344 23122 4396 23128
rect 4344 21548 4396 21554
rect 4344 21490 4396 21496
rect 4356 21146 4384 21490
rect 4344 21140 4396 21146
rect 4344 21082 4396 21088
rect 4344 20324 4396 20330
rect 4344 20266 4396 20272
rect 4356 20058 4384 20266
rect 4344 20052 4396 20058
rect 4344 19994 4396 20000
rect 4344 19848 4396 19854
rect 4344 19790 4396 19796
rect 4250 19136 4306 19145
rect 4250 19071 4306 19080
rect 4264 18902 4292 19071
rect 4252 18896 4304 18902
rect 4252 18838 4304 18844
rect 4160 18828 4212 18834
rect 4160 18770 4212 18776
rect 4172 18426 4200 18770
rect 4264 18426 4292 18838
rect 4160 18420 4212 18426
rect 4160 18362 4212 18368
rect 4252 18420 4304 18426
rect 4252 18362 4304 18368
rect 3516 16730 3568 16736
rect 3620 16748 3740 16776
rect 3620 16046 3648 16748
rect 3698 16688 3754 16697
rect 3698 16623 3754 16632
rect 3792 16652 3844 16658
rect 3608 16040 3660 16046
rect 3608 15982 3660 15988
rect 2976 12838 3096 12866
rect 3252 13688 3464 13716
rect 3516 13728 3568 13734
rect 2872 12436 2924 12442
rect 2872 12378 2924 12384
rect 2780 11076 2832 11082
rect 2780 11018 2832 11024
rect 2792 10826 2820 11018
rect 2700 10810 2820 10826
rect 2688 10804 2820 10810
rect 2740 10798 2820 10804
rect 2688 10746 2740 10752
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 2596 10192 2648 10198
rect 2596 10134 2648 10140
rect 2608 9722 2636 10134
rect 2688 9988 2740 9994
rect 2688 9930 2740 9936
rect 2596 9716 2648 9722
rect 2596 9658 2648 9664
rect 2504 9512 2556 9518
rect 2504 9454 2556 9460
rect 2424 9302 2544 9330
rect 2410 8392 2466 8401
rect 2410 8327 2412 8336
rect 2464 8327 2466 8336
rect 2412 8298 2464 8304
rect 2424 8090 2452 8298
rect 2412 8084 2464 8090
rect 2412 8026 2464 8032
rect 2240 7806 2360 7834
rect 2240 5386 2268 7806
rect 2320 7744 2372 7750
rect 2320 7686 2372 7692
rect 2332 7342 2360 7686
rect 2516 7562 2544 9302
rect 2700 9194 2728 9930
rect 2792 9586 2820 10542
rect 2884 10538 2912 12378
rect 2976 10713 3004 12838
rect 3056 12776 3108 12782
rect 3056 12718 3108 12724
rect 3068 12374 3096 12718
rect 3056 12368 3108 12374
rect 3056 12310 3108 12316
rect 3252 11336 3280 13688
rect 3516 13670 3568 13676
rect 3422 13424 3478 13433
rect 3422 13359 3478 13368
rect 3436 12481 3464 13359
rect 3528 13161 3556 13670
rect 3606 13560 3662 13569
rect 3606 13495 3662 13504
rect 3514 13152 3570 13161
rect 3514 13087 3570 13096
rect 3516 12640 3568 12646
rect 3516 12582 3568 12588
rect 3422 12472 3478 12481
rect 3422 12407 3478 12416
rect 3332 12368 3384 12374
rect 3332 12310 3384 12316
rect 3160 11308 3280 11336
rect 2962 10704 3018 10713
rect 2962 10639 3018 10648
rect 2872 10532 2924 10538
rect 2872 10474 2924 10480
rect 3160 10112 3188 11308
rect 3240 11212 3292 11218
rect 3240 11154 3292 11160
rect 3252 10470 3280 11154
rect 3240 10464 3292 10470
rect 3240 10406 3292 10412
rect 2884 10084 3188 10112
rect 2780 9580 2832 9586
rect 2780 9522 2832 9528
rect 2700 9178 2820 9194
rect 2700 9172 2832 9178
rect 2700 9166 2780 9172
rect 2700 7750 2728 9166
rect 2780 9114 2832 9120
rect 2884 8022 2912 10084
rect 3056 9988 3108 9994
rect 3056 9930 3108 9936
rect 3068 9518 3096 9930
rect 3148 9920 3200 9926
rect 3148 9862 3200 9868
rect 3056 9512 3108 9518
rect 3056 9454 3108 9460
rect 3054 9072 3110 9081
rect 3054 9007 3110 9016
rect 2964 8560 3016 8566
rect 2964 8502 3016 8508
rect 2872 8016 2924 8022
rect 2872 7958 2924 7964
rect 2780 7948 2832 7954
rect 2780 7890 2832 7896
rect 2688 7744 2740 7750
rect 2688 7686 2740 7692
rect 2516 7534 2728 7562
rect 2320 7336 2372 7342
rect 2320 7278 2372 7284
rect 2504 6792 2556 6798
rect 2504 6734 2556 6740
rect 2410 5808 2466 5817
rect 2410 5743 2466 5752
rect 2240 5358 2360 5386
rect 2228 5228 2280 5234
rect 2228 5170 2280 5176
rect 2056 4780 2176 4808
rect 1952 4616 2004 4622
rect 1952 4558 2004 4564
rect 1950 4176 2006 4185
rect 1950 4111 2006 4120
rect 1964 3942 1992 4111
rect 2056 4049 2084 4780
rect 2136 4684 2188 4690
rect 2136 4626 2188 4632
rect 2042 4040 2098 4049
rect 2148 4010 2176 4626
rect 2240 4146 2268 5170
rect 2332 5137 2360 5358
rect 2318 5128 2374 5137
rect 2318 5063 2374 5072
rect 2332 4185 2360 5063
rect 2318 4176 2374 4185
rect 2228 4140 2280 4146
rect 2318 4111 2374 4120
rect 2228 4082 2280 4088
rect 2042 3975 2098 3984
rect 2136 4004 2188 4010
rect 2136 3946 2188 3952
rect 1952 3936 2004 3942
rect 1952 3878 2004 3884
rect 1964 3738 1992 3878
rect 2240 3738 2268 4082
rect 2320 4072 2372 4078
rect 2320 4014 2372 4020
rect 2332 3942 2360 4014
rect 2320 3936 2372 3942
rect 2320 3878 2372 3884
rect 1952 3732 2004 3738
rect 1952 3674 2004 3680
rect 2228 3732 2280 3738
rect 2228 3674 2280 3680
rect 2332 2961 2360 3878
rect 2424 3738 2452 5743
rect 2516 5098 2544 6734
rect 2596 6656 2648 6662
rect 2596 6598 2648 6604
rect 2608 5370 2636 6598
rect 2700 6458 2728 7534
rect 2792 7002 2820 7890
rect 2884 7206 2912 7958
rect 2976 7886 3004 8502
rect 2964 7880 3016 7886
rect 2964 7822 3016 7828
rect 2976 7546 3004 7822
rect 2964 7540 3016 7546
rect 2964 7482 3016 7488
rect 2964 7336 3016 7342
rect 2964 7278 3016 7284
rect 2872 7200 2924 7206
rect 2872 7142 2924 7148
rect 2780 6996 2832 7002
rect 2780 6938 2832 6944
rect 2688 6452 2740 6458
rect 2688 6394 2740 6400
rect 2884 6390 2912 7142
rect 2872 6384 2924 6390
rect 2872 6326 2924 6332
rect 2872 6180 2924 6186
rect 2872 6122 2924 6128
rect 2884 5914 2912 6122
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 2596 5364 2648 5370
rect 2596 5306 2648 5312
rect 2504 5092 2556 5098
rect 2504 5034 2556 5040
rect 2596 5024 2648 5030
rect 2596 4966 2648 4972
rect 2412 3732 2464 3738
rect 2412 3674 2464 3680
rect 2424 2990 2452 3674
rect 2504 3460 2556 3466
rect 2504 3402 2556 3408
rect 2516 3194 2544 3402
rect 2608 3369 2636 4966
rect 2700 4554 2728 5714
rect 2976 5658 3004 7278
rect 2884 5630 3004 5658
rect 2780 4616 2832 4622
rect 2780 4558 2832 4564
rect 2688 4548 2740 4554
rect 2688 4490 2740 4496
rect 2792 4146 2820 4558
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 2884 3398 2912 5630
rect 2964 5568 3016 5574
rect 3068 5545 3096 9007
rect 2964 5510 3016 5516
rect 3054 5536 3110 5545
rect 2976 5370 3004 5510
rect 3054 5471 3110 5480
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 2976 4826 3004 5306
rect 2964 4820 3016 4826
rect 2964 4762 3016 4768
rect 3056 4072 3108 4078
rect 3056 4014 3108 4020
rect 2964 4004 3016 4010
rect 2964 3946 3016 3952
rect 2872 3392 2924 3398
rect 2594 3360 2650 3369
rect 2872 3334 2924 3340
rect 2594 3295 2650 3304
rect 2504 3188 2556 3194
rect 2504 3130 2556 3136
rect 2870 3088 2926 3097
rect 2870 3023 2926 3032
rect 2412 2984 2464 2990
rect 2318 2952 2374 2961
rect 2412 2926 2464 2932
rect 2318 2887 2374 2896
rect 2502 2816 2558 2825
rect 2502 2751 2558 2760
rect 1872 598 1992 626
rect 1964 480 1992 598
rect 2516 480 2544 2751
rect 2884 2650 2912 3023
rect 2976 2650 3004 3946
rect 3068 3777 3096 4014
rect 3054 3768 3110 3777
rect 3054 3703 3110 3712
rect 3160 3670 3188 9862
rect 3148 3664 3200 3670
rect 3148 3606 3200 3612
rect 3056 3392 3108 3398
rect 3056 3334 3108 3340
rect 3068 2922 3096 3334
rect 3160 3097 3188 3606
rect 3146 3088 3202 3097
rect 3146 3023 3202 3032
rect 3056 2916 3108 2922
rect 3056 2858 3108 2864
rect 2872 2644 2924 2650
rect 2872 2586 2924 2592
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 3068 2446 3096 2858
rect 3252 2553 3280 10406
rect 3344 10198 3372 12310
rect 3528 12102 3556 12582
rect 3516 12096 3568 12102
rect 3516 12038 3568 12044
rect 3528 11898 3556 12038
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 3528 11286 3556 11834
rect 3516 11280 3568 11286
rect 3516 11222 3568 11228
rect 3424 10532 3476 10538
rect 3424 10474 3476 10480
rect 3436 10266 3464 10474
rect 3528 10266 3556 11222
rect 3424 10260 3476 10266
rect 3424 10202 3476 10208
rect 3516 10260 3568 10266
rect 3516 10202 3568 10208
rect 3332 10192 3384 10198
rect 3332 10134 3384 10140
rect 3344 8072 3372 10134
rect 3620 9518 3648 13495
rect 3712 13433 3740 16623
rect 3792 16594 3844 16600
rect 3804 15473 3832 16594
rect 4158 16552 4214 16561
rect 4158 16487 4214 16496
rect 4068 16176 4120 16182
rect 4068 16118 4120 16124
rect 3884 15904 3936 15910
rect 3884 15846 3936 15852
rect 3896 15745 3924 15846
rect 3882 15736 3938 15745
rect 3882 15671 3938 15680
rect 3790 15464 3846 15473
rect 3790 15399 3846 15408
rect 3976 15360 4028 15366
rect 3976 15302 4028 15308
rect 3988 15065 4016 15302
rect 3974 15056 4030 15065
rect 4080 15042 4108 16118
rect 4172 16046 4200 16487
rect 4252 16108 4304 16114
rect 4252 16050 4304 16056
rect 4160 16040 4212 16046
rect 4160 15982 4212 15988
rect 4172 15706 4200 15982
rect 4160 15700 4212 15706
rect 4160 15642 4212 15648
rect 4080 15026 4200 15042
rect 4080 15020 4212 15026
rect 4080 15014 4160 15020
rect 3974 14991 4030 15000
rect 4160 14962 4212 14968
rect 3882 14920 3938 14929
rect 3882 14855 3938 14864
rect 3792 14816 3844 14822
rect 3792 14758 3844 14764
rect 3804 14346 3832 14758
rect 3792 14340 3844 14346
rect 3792 14282 3844 14288
rect 3804 13530 3832 14282
rect 3792 13524 3844 13530
rect 3792 13466 3844 13472
rect 3698 13424 3754 13433
rect 3698 13359 3754 13368
rect 3896 12889 3924 14855
rect 4264 14482 4292 16050
rect 4356 15858 4384 19790
rect 4448 15978 4476 24550
rect 4528 22432 4580 22438
rect 4528 22374 4580 22380
rect 4540 21894 4568 22374
rect 4816 22148 4844 27520
rect 5368 27470 5396 27520
rect 5264 27464 5316 27470
rect 5264 27406 5316 27412
rect 5356 27464 5408 27470
rect 5356 27406 5408 27412
rect 5172 24608 5224 24614
rect 5172 24550 5224 24556
rect 4896 24404 4948 24410
rect 4896 24346 4948 24352
rect 4724 22120 4844 22148
rect 4724 22012 4752 22120
rect 4632 21984 4752 22012
rect 4528 21888 4580 21894
rect 4528 21830 4580 21836
rect 4540 21321 4568 21830
rect 4526 21312 4582 21321
rect 4526 21247 4582 21256
rect 4540 19854 4568 21247
rect 4528 19848 4580 19854
rect 4528 19790 4580 19796
rect 4528 19168 4580 19174
rect 4528 19110 4580 19116
rect 4540 18698 4568 19110
rect 4528 18692 4580 18698
rect 4528 18634 4580 18640
rect 4632 18057 4660 21984
rect 4804 20256 4856 20262
rect 4802 20224 4804 20233
rect 4856 20224 4858 20233
rect 4802 20159 4858 20168
rect 4712 19916 4764 19922
rect 4712 19858 4764 19864
rect 4724 18970 4752 19858
rect 4804 19780 4856 19786
rect 4908 19768 4936 24346
rect 5184 23905 5212 24550
rect 5170 23896 5226 23905
rect 5170 23831 5226 23840
rect 4986 23352 5042 23361
rect 4986 23287 5042 23296
rect 5000 22574 5028 23287
rect 4988 22568 5040 22574
rect 4988 22510 5040 22516
rect 5276 22148 5304 27406
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 5540 24608 5592 24614
rect 5540 24550 5592 24556
rect 5448 22976 5500 22982
rect 5448 22918 5500 22924
rect 5460 22166 5488 22918
rect 5184 22120 5304 22148
rect 5448 22160 5500 22166
rect 5184 21486 5212 22120
rect 5448 22102 5500 22108
rect 5460 21690 5488 22102
rect 5448 21684 5500 21690
rect 5448 21626 5500 21632
rect 5552 21554 5580 24550
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 5816 23520 5868 23526
rect 5816 23462 5868 23468
rect 5828 23225 5856 23462
rect 5814 23216 5870 23225
rect 5814 23151 5870 23160
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5540 21548 5592 21554
rect 5540 21490 5592 21496
rect 5172 21480 5224 21486
rect 5172 21422 5224 21428
rect 5632 21344 5684 21350
rect 5632 21286 5684 21292
rect 5080 21072 5132 21078
rect 5080 21014 5132 21020
rect 5170 21040 5226 21049
rect 5092 20534 5120 21014
rect 5644 21010 5672 21286
rect 5170 20975 5226 20984
rect 5632 21004 5684 21010
rect 5080 20528 5132 20534
rect 5080 20470 5132 20476
rect 5092 19786 5120 20470
rect 4856 19740 4936 19768
rect 5080 19780 5132 19786
rect 4804 19722 4856 19728
rect 5080 19722 5132 19728
rect 4816 19174 4844 19722
rect 4804 19168 4856 19174
rect 4804 19110 4856 19116
rect 4712 18964 4764 18970
rect 4712 18906 4764 18912
rect 4712 18760 4764 18766
rect 4712 18702 4764 18708
rect 4618 18048 4674 18057
rect 4618 17983 4674 17992
rect 4620 17808 4672 17814
rect 4724 17796 4752 18702
rect 4672 17768 4752 17796
rect 4620 17750 4672 17756
rect 4632 17542 4660 17750
rect 4620 17536 4672 17542
rect 4620 17478 4672 17484
rect 4632 17270 4660 17478
rect 4620 17264 4672 17270
rect 4620 17206 4672 17212
rect 4632 16250 4660 17206
rect 4620 16244 4672 16250
rect 4620 16186 4672 16192
rect 4436 15972 4488 15978
rect 4436 15914 4488 15920
rect 4712 15904 4764 15910
rect 4710 15872 4712 15881
rect 4764 15872 4766 15881
rect 4356 15830 4660 15858
rect 4342 15736 4398 15745
rect 4342 15671 4398 15680
rect 4436 15700 4488 15706
rect 4252 14476 4304 14482
rect 4252 14418 4304 14424
rect 4160 14408 4212 14414
rect 4160 14350 4212 14356
rect 3976 13456 4028 13462
rect 3976 13398 4028 13404
rect 3882 12880 3938 12889
rect 3882 12815 3938 12824
rect 3988 12442 4016 13398
rect 4172 12782 4200 14350
rect 4356 14074 4384 15671
rect 4436 15642 4488 15648
rect 4448 15609 4476 15642
rect 4434 15600 4490 15609
rect 4434 15535 4490 15544
rect 4528 15564 4580 15570
rect 4528 15506 4580 15512
rect 4436 15496 4488 15502
rect 4436 15438 4488 15444
rect 4448 14822 4476 15438
rect 4540 15201 4568 15506
rect 4526 15192 4582 15201
rect 4526 15127 4582 15136
rect 4436 14816 4488 14822
rect 4436 14758 4488 14764
rect 4344 14068 4396 14074
rect 4344 14010 4396 14016
rect 4252 13728 4304 13734
rect 4252 13670 4304 13676
rect 4264 13394 4292 13670
rect 4632 13512 4660 15830
rect 4710 15807 4766 15816
rect 4448 13484 4660 13512
rect 4252 13388 4304 13394
rect 4252 13330 4304 13336
rect 4160 12776 4212 12782
rect 4160 12718 4212 12724
rect 3976 12436 4028 12442
rect 3976 12378 4028 12384
rect 4264 12306 4292 13330
rect 4344 12640 4396 12646
rect 4344 12582 4396 12588
rect 4252 12300 4304 12306
rect 4252 12242 4304 12248
rect 4356 12170 4384 12582
rect 4448 12458 4476 13484
rect 4528 13388 4580 13394
rect 4528 13330 4580 13336
rect 4540 13297 4568 13330
rect 4620 13320 4672 13326
rect 4526 13288 4582 13297
rect 4620 13262 4672 13268
rect 4526 13223 4582 13232
rect 4540 12986 4568 13223
rect 4528 12980 4580 12986
rect 4528 12922 4580 12928
rect 4632 12646 4660 13262
rect 4620 12640 4672 12646
rect 4620 12582 4672 12588
rect 4448 12430 4568 12458
rect 4540 12322 4568 12430
rect 4436 12300 4488 12306
rect 4540 12294 4660 12322
rect 4436 12242 4488 12248
rect 3792 12164 3844 12170
rect 3792 12106 3844 12112
rect 4344 12164 4396 12170
rect 4344 12106 4396 12112
rect 3804 11354 3832 12106
rect 4448 11898 4476 12242
rect 4528 12232 4580 12238
rect 4528 12174 4580 12180
rect 4436 11892 4488 11898
rect 4436 11834 4488 11840
rect 4344 11756 4396 11762
rect 4344 11698 4396 11704
rect 3792 11348 3844 11354
rect 3792 11290 3844 11296
rect 3974 11248 4030 11257
rect 3974 11183 4030 11192
rect 3884 11076 3936 11082
rect 3884 11018 3936 11024
rect 3790 10976 3846 10985
rect 3790 10911 3846 10920
rect 3700 10124 3752 10130
rect 3700 10066 3752 10072
rect 3608 9512 3660 9518
rect 3608 9454 3660 9460
rect 3424 8900 3476 8906
rect 3424 8842 3476 8848
rect 3436 8566 3464 8842
rect 3516 8832 3568 8838
rect 3516 8774 3568 8780
rect 3424 8560 3476 8566
rect 3424 8502 3476 8508
rect 3528 8498 3556 8774
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3608 8492 3660 8498
rect 3608 8434 3660 8440
rect 3620 8090 3648 8434
rect 3608 8084 3660 8090
rect 3344 8044 3464 8072
rect 3330 7984 3386 7993
rect 3330 7919 3386 7928
rect 3344 5658 3372 7919
rect 3436 7342 3464 8044
rect 3608 8026 3660 8032
rect 3424 7336 3476 7342
rect 3424 7278 3476 7284
rect 3712 7206 3740 10066
rect 3804 7857 3832 10911
rect 3896 9874 3924 11018
rect 3988 10169 4016 11183
rect 4066 10432 4122 10441
rect 4066 10367 4122 10376
rect 3974 10160 4030 10169
rect 3974 10095 4030 10104
rect 4080 9908 4108 10367
rect 4160 9920 4212 9926
rect 4080 9880 4160 9908
rect 3896 9846 4016 9874
rect 3884 8560 3936 8566
rect 3884 8502 3936 8508
rect 3896 8294 3924 8502
rect 3884 8288 3936 8294
rect 3884 8230 3936 8236
rect 3896 8090 3924 8230
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 3988 7857 4016 9846
rect 4080 8634 4108 9880
rect 4160 9862 4212 9868
rect 4252 9716 4304 9722
rect 4252 9658 4304 9664
rect 4160 9376 4212 9382
rect 4160 9318 4212 9324
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 4172 8498 4200 9318
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 3790 7848 3846 7857
rect 3790 7783 3846 7792
rect 3974 7848 4030 7857
rect 3974 7783 4030 7792
rect 3988 7478 4016 7783
rect 3976 7472 4028 7478
rect 3976 7414 4028 7420
rect 3700 7200 3752 7206
rect 3700 7142 3752 7148
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3528 5914 3556 6598
rect 3608 6112 3660 6118
rect 3608 6054 3660 6060
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 3344 5630 3464 5658
rect 3330 4992 3386 5001
rect 3330 4927 3386 4936
rect 3238 2544 3294 2553
rect 3238 2479 3294 2488
rect 3056 2440 3108 2446
rect 3056 2382 3108 2388
rect 3344 762 3372 4927
rect 3436 4078 3464 5630
rect 3620 5273 3648 6054
rect 3606 5264 3662 5273
rect 3606 5199 3608 5208
rect 3660 5199 3662 5208
rect 3608 5170 3660 5176
rect 3620 4826 3648 5170
rect 3608 4820 3660 4826
rect 3608 4762 3660 4768
rect 3424 4072 3476 4078
rect 3424 4014 3476 4020
rect 3424 3936 3476 3942
rect 3422 3904 3424 3913
rect 3476 3904 3478 3913
rect 3422 3839 3478 3848
rect 3436 3738 3464 3839
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 3712 3233 3740 7142
rect 3974 6896 4030 6905
rect 3974 6831 4030 6840
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3896 5778 3924 6598
rect 3884 5772 3936 5778
rect 3884 5714 3936 5720
rect 3884 5024 3936 5030
rect 3884 4966 3936 4972
rect 3896 4758 3924 4966
rect 3884 4752 3936 4758
rect 3884 4694 3936 4700
rect 3896 4593 3924 4694
rect 3882 4584 3938 4593
rect 3882 4519 3938 4528
rect 3882 4040 3938 4049
rect 3792 4004 3844 4010
rect 3882 3975 3938 3984
rect 3792 3946 3844 3952
rect 3804 3777 3832 3946
rect 3896 3942 3924 3975
rect 3884 3936 3936 3942
rect 3884 3878 3936 3884
rect 3790 3768 3846 3777
rect 3790 3703 3846 3712
rect 3698 3224 3754 3233
rect 3896 3194 3924 3878
rect 3698 3159 3754 3168
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 3698 2952 3754 2961
rect 3698 2887 3754 2896
rect 3608 2508 3660 2514
rect 3608 2450 3660 2456
rect 3620 2417 3648 2450
rect 3606 2408 3662 2417
rect 3606 2343 3662 2352
rect 3160 734 3372 762
rect 3160 480 3188 734
rect 3712 480 3740 2887
rect 3988 2650 4016 6831
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 4080 5953 4108 6054
rect 4066 5944 4122 5953
rect 4066 5879 4122 5888
rect 4172 5710 4200 6394
rect 4160 5704 4212 5710
rect 4066 5672 4122 5681
rect 4160 5646 4212 5652
rect 4066 5607 4068 5616
rect 4120 5607 4122 5616
rect 4068 5578 4120 5584
rect 4172 5370 4200 5646
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 4264 4842 4292 9658
rect 4356 7993 4384 11698
rect 4540 11354 4568 12174
rect 4632 11762 4660 12294
rect 4620 11756 4672 11762
rect 4620 11698 4672 11704
rect 4632 11626 4660 11698
rect 4620 11620 4672 11626
rect 4620 11562 4672 11568
rect 4528 11348 4580 11354
rect 4528 11290 4580 11296
rect 4816 11218 4844 19110
rect 5092 18902 5120 19722
rect 5080 18896 5132 18902
rect 5080 18838 5132 18844
rect 5080 18624 5132 18630
rect 5080 18566 5132 18572
rect 4896 17196 4948 17202
rect 4896 17138 4948 17144
rect 4908 16794 4936 17138
rect 5092 16998 5120 18566
rect 5184 18426 5212 20975
rect 5632 20946 5684 20952
rect 5540 20800 5592 20806
rect 5460 20748 5540 20754
rect 5460 20742 5592 20748
rect 5460 20726 5580 20742
rect 5460 20466 5488 20726
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5448 20460 5500 20466
rect 5448 20402 5500 20408
rect 5908 20392 5960 20398
rect 5908 20334 5960 20340
rect 5920 20058 5948 20334
rect 5908 20052 5960 20058
rect 5908 19994 5960 20000
rect 5264 19712 5316 19718
rect 5264 19654 5316 19660
rect 5172 18420 5224 18426
rect 5172 18362 5224 18368
rect 5276 18086 5304 19654
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5540 19304 5592 19310
rect 5460 19264 5540 19292
rect 5356 19168 5408 19174
rect 5356 19110 5408 19116
rect 5368 18970 5396 19110
rect 5356 18964 5408 18970
rect 5356 18906 5408 18912
rect 5356 18624 5408 18630
rect 5460 18612 5488 19264
rect 5540 19246 5592 19252
rect 5540 19168 5592 19174
rect 5540 19110 5592 19116
rect 5408 18584 5488 18612
rect 5356 18566 5408 18572
rect 5264 18080 5316 18086
rect 5264 18022 5316 18028
rect 5080 16992 5132 16998
rect 5080 16934 5132 16940
rect 4896 16788 4948 16794
rect 4896 16730 4948 16736
rect 5092 16658 5120 16934
rect 5368 16726 5396 18566
rect 5446 18456 5502 18465
rect 5552 18442 5580 19110
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5502 18414 5580 18442
rect 5446 18391 5502 18400
rect 5448 18352 5500 18358
rect 5448 18294 5500 18300
rect 5460 17746 5488 18294
rect 5540 18216 5592 18222
rect 5540 18158 5592 18164
rect 5448 17740 5500 17746
rect 5448 17682 5500 17688
rect 5552 17610 5580 18158
rect 5540 17604 5592 17610
rect 5540 17546 5592 17552
rect 5448 17536 5500 17542
rect 5448 17478 5500 17484
rect 5460 17202 5488 17478
rect 5552 17338 5580 17546
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5540 17332 5592 17338
rect 5540 17274 5592 17280
rect 5448 17196 5500 17202
rect 5448 17138 5500 17144
rect 6012 17134 6040 27520
rect 6276 24812 6328 24818
rect 6276 24754 6328 24760
rect 6288 24614 6316 24754
rect 6276 24608 6328 24614
rect 6276 24550 6328 24556
rect 6288 24274 6316 24550
rect 6276 24268 6328 24274
rect 6276 24210 6328 24216
rect 6288 23866 6316 24210
rect 6276 23860 6328 23866
rect 6276 23802 6328 23808
rect 6182 23624 6238 23633
rect 6182 23559 6238 23568
rect 6092 23520 6144 23526
rect 6092 23462 6144 23468
rect 6104 21593 6132 23462
rect 6090 21584 6146 21593
rect 6090 21519 6146 21528
rect 6196 21049 6224 23559
rect 6564 23361 6592 27520
rect 7012 27260 7064 27266
rect 7012 27202 7064 27208
rect 6920 25356 6972 25362
rect 6920 25298 6972 25304
rect 6932 24886 6960 25298
rect 7024 25226 7052 27202
rect 7012 25220 7064 25226
rect 7012 25162 7064 25168
rect 6920 24880 6972 24886
rect 6920 24822 6972 24828
rect 6932 24721 6960 24822
rect 6918 24712 6974 24721
rect 6918 24647 6974 24656
rect 6828 24608 6880 24614
rect 6828 24550 6880 24556
rect 6644 24064 6696 24070
rect 6644 24006 6696 24012
rect 6550 23352 6606 23361
rect 6550 23287 6606 23296
rect 6552 23180 6604 23186
rect 6552 23122 6604 23128
rect 6458 23080 6514 23089
rect 6458 23015 6514 23024
rect 6274 22672 6330 22681
rect 6274 22607 6330 22616
rect 6288 21962 6316 22607
rect 6276 21956 6328 21962
rect 6276 21898 6328 21904
rect 6274 21584 6330 21593
rect 6274 21519 6330 21528
rect 6288 21418 6316 21519
rect 6276 21412 6328 21418
rect 6276 21354 6328 21360
rect 6182 21040 6238 21049
rect 6182 20975 6238 20984
rect 6276 21004 6328 21010
rect 6276 20946 6328 20952
rect 6288 20262 6316 20946
rect 6276 20256 6328 20262
rect 6276 20198 6328 20204
rect 6184 18896 6236 18902
rect 6184 18838 6236 18844
rect 6196 18086 6224 18838
rect 6288 18834 6316 20198
rect 6472 18970 6500 23015
rect 6564 21350 6592 23122
rect 6656 22778 6684 24006
rect 6734 23352 6790 23361
rect 6734 23287 6790 23296
rect 6644 22772 6696 22778
rect 6644 22714 6696 22720
rect 6644 22024 6696 22030
rect 6644 21966 6696 21972
rect 6656 21690 6684 21966
rect 6644 21684 6696 21690
rect 6644 21626 6696 21632
rect 6552 21344 6604 21350
rect 6552 21286 6604 21292
rect 6552 20392 6604 20398
rect 6552 20334 6604 20340
rect 6564 20233 6592 20334
rect 6550 20224 6606 20233
rect 6550 20159 6606 20168
rect 6644 19916 6696 19922
rect 6644 19858 6696 19864
rect 6552 19848 6604 19854
rect 6552 19790 6604 19796
rect 6460 18964 6512 18970
rect 6460 18906 6512 18912
rect 6276 18828 6328 18834
rect 6276 18770 6328 18776
rect 6288 18358 6316 18770
rect 6276 18352 6328 18358
rect 6276 18294 6328 18300
rect 6288 18222 6316 18294
rect 6276 18216 6328 18222
rect 6276 18158 6328 18164
rect 6184 18080 6236 18086
rect 6184 18022 6236 18028
rect 6196 17542 6224 18022
rect 6472 17626 6500 18906
rect 6564 18737 6592 19790
rect 6656 19553 6684 19858
rect 6642 19544 6698 19553
rect 6642 19479 6644 19488
rect 6696 19479 6698 19488
rect 6644 19450 6696 19456
rect 6550 18728 6606 18737
rect 6550 18663 6606 18672
rect 6288 17598 6500 17626
rect 6184 17536 6236 17542
rect 6184 17478 6236 17484
rect 6196 17270 6224 17478
rect 6184 17264 6236 17270
rect 6184 17206 6236 17212
rect 6092 17196 6144 17202
rect 6092 17138 6144 17144
rect 6000 17128 6052 17134
rect 6000 17070 6052 17076
rect 5814 16824 5870 16833
rect 5814 16759 5870 16768
rect 5356 16720 5408 16726
rect 5356 16662 5408 16668
rect 5828 16658 5856 16759
rect 5080 16652 5132 16658
rect 5080 16594 5132 16600
rect 5816 16652 5868 16658
rect 5868 16612 6040 16640
rect 5816 16594 5868 16600
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5170 16008 5226 16017
rect 4896 15972 4948 15978
rect 5170 15943 5226 15952
rect 4896 15914 4948 15920
rect 4908 12458 4936 15914
rect 5184 15910 5212 15943
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 5356 15904 5408 15910
rect 5356 15846 5408 15852
rect 5368 15638 5396 15846
rect 6012 15706 6040 16612
rect 6104 16590 6132 17138
rect 6288 17116 6316 17598
rect 6368 17536 6420 17542
rect 6368 17478 6420 17484
rect 6644 17536 6696 17542
rect 6644 17478 6696 17484
rect 6196 17088 6316 17116
rect 6092 16584 6144 16590
rect 6092 16526 6144 16532
rect 6196 15722 6224 17088
rect 6380 17066 6408 17478
rect 6656 17270 6684 17478
rect 6644 17264 6696 17270
rect 6644 17206 6696 17212
rect 6552 17128 6604 17134
rect 6552 17070 6604 17076
rect 6368 17060 6420 17066
rect 6368 17002 6420 17008
rect 6460 16992 6512 16998
rect 6380 16940 6460 16946
rect 6380 16934 6512 16940
rect 6380 16918 6500 16934
rect 6276 16516 6328 16522
rect 6276 16458 6328 16464
rect 6288 15910 6316 16458
rect 6276 15904 6328 15910
rect 6276 15846 6328 15852
rect 5448 15700 5500 15706
rect 6000 15700 6052 15706
rect 5500 15660 5580 15688
rect 5448 15642 5500 15648
rect 5356 15632 5408 15638
rect 5356 15574 5408 15580
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 5356 15156 5408 15162
rect 5356 15098 5408 15104
rect 5172 15020 5224 15026
rect 5172 14962 5224 14968
rect 5078 14920 5134 14929
rect 5078 14855 5080 14864
rect 5132 14855 5134 14864
rect 5080 14826 5132 14832
rect 5184 14074 5212 14962
rect 5262 14240 5318 14249
rect 5262 14175 5318 14184
rect 5172 14068 5224 14074
rect 5172 14010 5224 14016
rect 5080 13864 5132 13870
rect 5080 13806 5132 13812
rect 4908 12430 5028 12458
rect 4896 12232 4948 12238
rect 4896 12174 4948 12180
rect 4908 11694 4936 12174
rect 5000 11830 5028 12430
rect 5092 12102 5120 13806
rect 5170 12200 5226 12209
rect 5170 12135 5226 12144
rect 5080 12096 5132 12102
rect 5080 12038 5132 12044
rect 4988 11824 5040 11830
rect 4988 11766 5040 11772
rect 4896 11688 4948 11694
rect 4896 11630 4948 11636
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 4896 11076 4948 11082
rect 4896 11018 4948 11024
rect 4436 10464 4488 10470
rect 4436 10406 4488 10412
rect 4448 9994 4476 10406
rect 4528 10056 4580 10062
rect 4528 9998 4580 10004
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4436 9988 4488 9994
rect 4436 9930 4488 9936
rect 4448 8906 4476 9930
rect 4540 9602 4568 9998
rect 4724 9722 4752 9998
rect 4712 9716 4764 9722
rect 4712 9658 4764 9664
rect 4804 9716 4856 9722
rect 4804 9658 4856 9664
rect 4816 9602 4844 9658
rect 4540 9574 4844 9602
rect 4436 8900 4488 8906
rect 4436 8842 4488 8848
rect 4342 7984 4398 7993
rect 4342 7919 4398 7928
rect 4540 7449 4568 9574
rect 4620 9104 4672 9110
rect 4620 9046 4672 9052
rect 4632 8265 4660 9046
rect 4804 9036 4856 9042
rect 4804 8978 4856 8984
rect 4816 8362 4844 8978
rect 4804 8356 4856 8362
rect 4804 8298 4856 8304
rect 4712 8288 4764 8294
rect 4618 8256 4674 8265
rect 4712 8230 4764 8236
rect 4618 8191 4674 8200
rect 4632 8090 4660 8191
rect 4620 8084 4672 8090
rect 4620 8026 4672 8032
rect 4724 7818 4752 8230
rect 4712 7812 4764 7818
rect 4712 7754 4764 7760
rect 4526 7440 4582 7449
rect 4526 7375 4582 7384
rect 4344 7336 4396 7342
rect 4344 7278 4396 7284
rect 4080 4826 4292 4842
rect 4068 4820 4292 4826
rect 4120 4814 4292 4820
rect 4068 4762 4120 4768
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 4080 3602 4108 4626
rect 4172 4146 4200 4814
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 4172 3670 4200 4082
rect 4160 3664 4212 3670
rect 4160 3606 4212 3612
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 4080 2990 4108 3538
rect 4172 3126 4200 3606
rect 4160 3120 4212 3126
rect 4160 3062 4212 3068
rect 4068 2984 4120 2990
rect 4068 2926 4120 2932
rect 3976 2644 4028 2650
rect 3976 2586 4028 2592
rect 4356 2009 4384 7278
rect 4724 6934 4752 7754
rect 4712 6928 4764 6934
rect 4712 6870 4764 6876
rect 4620 6656 4672 6662
rect 4620 6598 4672 6604
rect 4632 6322 4660 6598
rect 4620 6316 4672 6322
rect 4620 6258 4672 6264
rect 4436 4752 4488 4758
rect 4436 4694 4488 4700
rect 4526 4720 4582 4729
rect 4448 3398 4476 4694
rect 4526 4655 4582 4664
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 4342 2000 4398 2009
rect 4342 1935 4398 1944
rect 4540 626 4568 4655
rect 4710 3360 4766 3369
rect 4710 3295 4766 3304
rect 4724 2650 4752 3295
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 4264 598 4568 626
rect 4264 480 4292 598
rect 4816 480 4844 8298
rect 4908 1465 4936 11018
rect 5000 8294 5028 11766
rect 5092 11762 5120 12038
rect 5080 11756 5132 11762
rect 5080 11698 5132 11704
rect 5092 11150 5120 11698
rect 5080 11144 5132 11150
rect 5080 11086 5132 11092
rect 5184 11082 5212 12135
rect 5172 11076 5224 11082
rect 5172 11018 5224 11024
rect 5184 10810 5212 11018
rect 5172 10804 5224 10810
rect 5172 10746 5224 10752
rect 5172 10056 5224 10062
rect 5172 9998 5224 10004
rect 5078 9616 5134 9625
rect 5078 9551 5080 9560
rect 5132 9551 5134 9560
rect 5080 9522 5132 9528
rect 5080 9444 5132 9450
rect 5184 9432 5212 9998
rect 5132 9404 5212 9432
rect 5080 9386 5132 9392
rect 5092 9178 5120 9386
rect 5080 9172 5132 9178
rect 5080 9114 5132 9120
rect 4988 8288 5040 8294
rect 4988 8230 5040 8236
rect 4988 6860 5040 6866
rect 4988 6802 5040 6808
rect 5000 6458 5028 6802
rect 5092 6798 5120 9114
rect 5172 8900 5224 8906
rect 5172 8842 5224 8848
rect 5184 8498 5212 8842
rect 5172 8492 5224 8498
rect 5172 8434 5224 8440
rect 5172 7472 5224 7478
rect 5170 7440 5172 7449
rect 5224 7440 5226 7449
rect 5170 7375 5226 7384
rect 5080 6792 5132 6798
rect 5080 6734 5132 6740
rect 4988 6452 5040 6458
rect 4988 6394 5040 6400
rect 5092 6202 5120 6734
rect 5000 6174 5120 6202
rect 5184 6186 5212 7375
rect 5172 6180 5224 6186
rect 5000 4690 5028 6174
rect 5172 6122 5224 6128
rect 5080 6112 5132 6118
rect 5080 6054 5132 6060
rect 5092 5817 5120 6054
rect 5078 5808 5134 5817
rect 5078 5743 5134 5752
rect 4988 4684 5040 4690
rect 4988 4626 5040 4632
rect 5276 4146 5304 14175
rect 5368 13462 5396 15098
rect 5460 14618 5488 15506
rect 5448 14612 5500 14618
rect 5448 14554 5500 14560
rect 5552 14550 5580 15660
rect 6196 15694 6316 15722
rect 6000 15642 6052 15648
rect 6000 15496 6052 15502
rect 5998 15464 6000 15473
rect 6184 15496 6236 15502
rect 6052 15464 6054 15473
rect 6184 15438 6236 15444
rect 5998 15399 6054 15408
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5998 15192 6054 15201
rect 5998 15127 6054 15136
rect 5540 14544 5592 14550
rect 5540 14486 5592 14492
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5630 13832 5686 13841
rect 5630 13767 5686 13776
rect 5538 13696 5594 13705
rect 5538 13631 5594 13640
rect 5552 13530 5580 13631
rect 5540 13524 5592 13530
rect 5540 13466 5592 13472
rect 5356 13456 5408 13462
rect 5356 13398 5408 13404
rect 5644 13394 5672 13767
rect 5814 13424 5870 13433
rect 5632 13388 5684 13394
rect 5814 13359 5870 13368
rect 5632 13330 5684 13336
rect 5828 13258 5856 13359
rect 5816 13252 5868 13258
rect 5816 13194 5868 13200
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 5460 12442 5488 12718
rect 5448 12436 5500 12442
rect 5448 12378 5500 12384
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 5460 10810 5488 11154
rect 5540 11008 5592 11014
rect 5540 10950 5592 10956
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5552 10606 5580 10950
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5816 10736 5868 10742
rect 5814 10704 5816 10713
rect 5868 10704 5870 10713
rect 5814 10639 5870 10648
rect 5540 10600 5592 10606
rect 5540 10542 5592 10548
rect 5448 10124 5500 10130
rect 5448 10066 5500 10072
rect 5460 9466 5488 10066
rect 5552 9586 5580 10542
rect 5630 10296 5686 10305
rect 5630 10231 5632 10240
rect 5684 10231 5686 10240
rect 5632 10202 5684 10208
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 5460 9438 5580 9466
rect 5552 8974 5580 9438
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 5552 8401 5580 8774
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 6012 8650 6040 15127
rect 6090 15056 6146 15065
rect 6090 14991 6146 15000
rect 6104 14074 6132 14991
rect 6196 14822 6224 15438
rect 6184 14816 6236 14822
rect 6184 14758 6236 14764
rect 6196 14385 6224 14758
rect 6182 14376 6238 14385
rect 6182 14311 6238 14320
rect 6092 14068 6144 14074
rect 6092 14010 6144 14016
rect 6092 13932 6144 13938
rect 6092 13874 6144 13880
rect 6104 12866 6132 13874
rect 6184 13388 6236 13394
rect 6184 13330 6236 13336
rect 6196 12986 6224 13330
rect 6184 12980 6236 12986
rect 6184 12922 6236 12928
rect 6104 12838 6224 12866
rect 6092 12436 6144 12442
rect 6092 12378 6144 12384
rect 6104 11354 6132 12378
rect 6092 11348 6144 11354
rect 6092 11290 6144 11296
rect 6104 11014 6132 11290
rect 6092 11008 6144 11014
rect 6092 10950 6144 10956
rect 6104 10198 6132 10229
rect 6092 10192 6144 10198
rect 6090 10160 6092 10169
rect 6144 10160 6146 10169
rect 6090 10095 6146 10104
rect 6104 9722 6132 10095
rect 6092 9716 6144 9722
rect 6092 9658 6144 9664
rect 6012 8622 6132 8650
rect 6000 8560 6052 8566
rect 5998 8528 6000 8537
rect 6052 8528 6054 8537
rect 5998 8463 6054 8472
rect 5538 8392 5594 8401
rect 6104 8378 6132 8622
rect 5538 8327 5594 8336
rect 6012 8350 6132 8378
rect 5540 7948 5592 7954
rect 5540 7890 5592 7896
rect 5552 6322 5580 7890
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 6012 7274 6040 8350
rect 6092 7404 6144 7410
rect 6092 7346 6144 7352
rect 6000 7268 6052 7274
rect 6000 7210 6052 7216
rect 6104 6866 6132 7346
rect 6092 6860 6144 6866
rect 6092 6802 6144 6808
rect 5998 6760 6054 6769
rect 5998 6695 6054 6704
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 6012 5930 6040 6695
rect 6104 6254 6132 6802
rect 6092 6248 6144 6254
rect 6092 6190 6144 6196
rect 5920 5914 6040 5930
rect 5908 5908 6040 5914
rect 5960 5902 6040 5908
rect 5908 5850 5960 5856
rect 6090 5808 6146 5817
rect 5448 5772 5500 5778
rect 6090 5743 6092 5752
rect 5448 5714 5500 5720
rect 6144 5743 6146 5752
rect 6092 5714 6144 5720
rect 5356 5568 5408 5574
rect 5356 5510 5408 5516
rect 5368 5030 5396 5510
rect 5460 5370 5488 5714
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5448 5364 5500 5370
rect 5448 5306 5500 5312
rect 5632 5228 5684 5234
rect 5632 5170 5684 5176
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 5644 4826 5672 5170
rect 6000 5024 6052 5030
rect 6000 4966 6052 4972
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 6012 4457 6040 4966
rect 5998 4448 6054 4457
rect 5622 4380 5918 4400
rect 5998 4383 6054 4392
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 5540 4004 5592 4010
rect 5540 3946 5592 3952
rect 5172 3936 5224 3942
rect 5172 3878 5224 3884
rect 5184 3738 5212 3878
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 5552 3058 5580 3946
rect 6090 3768 6146 3777
rect 6090 3703 6146 3712
rect 6104 3534 6132 3703
rect 6092 3528 6144 3534
rect 6092 3470 6144 3476
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5632 3120 5684 3126
rect 5630 3088 5632 3097
rect 5684 3088 5686 3097
rect 5540 3052 5592 3058
rect 5630 3023 5686 3032
rect 5540 2994 5592 3000
rect 5262 2544 5318 2553
rect 5172 2508 5224 2514
rect 5262 2479 5318 2488
rect 6092 2508 6144 2514
rect 5172 2450 5224 2456
rect 5184 2145 5212 2450
rect 5276 2378 5304 2479
rect 6092 2450 6144 2456
rect 5354 2408 5410 2417
rect 5264 2372 5316 2378
rect 5354 2343 5410 2352
rect 5264 2314 5316 2320
rect 5170 2136 5226 2145
rect 5170 2071 5226 2080
rect 4894 1456 4950 1465
rect 4894 1391 4950 1400
rect 5368 480 5396 2343
rect 6104 2281 6132 2450
rect 6090 2272 6146 2281
rect 5622 2204 5918 2224
rect 6090 2207 6146 2216
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 6196 610 6224 12838
rect 6288 12628 6316 15694
rect 6380 12730 6408 16918
rect 6458 16688 6514 16697
rect 6458 16623 6514 16632
rect 6472 16454 6500 16623
rect 6460 16448 6512 16454
rect 6460 16390 6512 16396
rect 6472 16114 6500 16390
rect 6460 16108 6512 16114
rect 6460 16050 6512 16056
rect 6564 15586 6592 17070
rect 6656 16658 6684 17206
rect 6644 16652 6696 16658
rect 6644 16594 6696 16600
rect 6748 15994 6776 23287
rect 6840 22778 6868 24550
rect 7012 24064 7064 24070
rect 6918 24032 6974 24041
rect 7012 24006 7064 24012
rect 6918 23967 6974 23976
rect 6932 23089 6960 23967
rect 7024 23730 7052 24006
rect 7012 23724 7064 23730
rect 7012 23666 7064 23672
rect 7024 23322 7052 23666
rect 7012 23316 7064 23322
rect 7012 23258 7064 23264
rect 6918 23080 6974 23089
rect 6918 23015 6974 23024
rect 6828 22772 6880 22778
rect 7116 22760 7144 27520
rect 7196 26308 7248 26314
rect 7196 26250 7248 26256
rect 7208 25498 7236 26250
rect 7196 25492 7248 25498
rect 7196 25434 7248 25440
rect 7668 23712 7696 27520
rect 8116 26580 8168 26586
rect 8116 26522 8168 26528
rect 7748 25356 7800 25362
rect 7748 25298 7800 25304
rect 7760 24449 7788 25298
rect 8128 24954 8156 26522
rect 8116 24948 8168 24954
rect 8116 24890 8168 24896
rect 8220 24834 8248 27520
rect 7944 24806 8248 24834
rect 7840 24744 7892 24750
rect 7840 24686 7892 24692
rect 7746 24440 7802 24449
rect 7746 24375 7802 24384
rect 7852 24313 7880 24686
rect 7838 24304 7894 24313
rect 7838 24239 7894 24248
rect 7484 23684 7696 23712
rect 7116 22732 7236 22760
rect 6828 22714 6880 22720
rect 7104 22432 7156 22438
rect 7104 22374 7156 22380
rect 7116 21894 7144 22374
rect 7104 21888 7156 21894
rect 7104 21830 7156 21836
rect 7116 20942 7144 21830
rect 7104 20936 7156 20942
rect 7104 20878 7156 20884
rect 6920 20800 6972 20806
rect 6920 20742 6972 20748
rect 6932 20398 6960 20742
rect 6920 20392 6972 20398
rect 6920 20334 6972 20340
rect 7010 20360 7066 20369
rect 7010 20295 7066 20304
rect 6828 20052 6880 20058
rect 6828 19994 6880 20000
rect 6840 19310 6868 19994
rect 7024 19786 7052 20295
rect 7012 19780 7064 19786
rect 7012 19722 7064 19728
rect 6828 19304 6880 19310
rect 6880 19264 6960 19292
rect 6828 19246 6880 19252
rect 6828 19168 6880 19174
rect 6828 19110 6880 19116
rect 6840 18465 6868 19110
rect 6826 18456 6882 18465
rect 6826 18391 6882 18400
rect 6932 18306 6960 19264
rect 7012 19168 7064 19174
rect 7010 19136 7012 19145
rect 7064 19136 7066 19145
rect 7010 19071 7066 19080
rect 7012 18624 7064 18630
rect 7012 18566 7064 18572
rect 6840 18278 6960 18306
rect 7024 18290 7052 18566
rect 7012 18284 7064 18290
rect 6840 17762 6868 18278
rect 7012 18226 7064 18232
rect 6920 18148 6972 18154
rect 6920 18090 6972 18096
rect 6932 17882 6960 18090
rect 7012 18080 7064 18086
rect 7012 18022 7064 18028
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 6840 17734 6960 17762
rect 6932 17134 6960 17734
rect 6920 17128 6972 17134
rect 6920 17070 6972 17076
rect 6932 16946 6960 17070
rect 6840 16918 6960 16946
rect 6840 16726 6868 16918
rect 7024 16810 7052 18022
rect 6932 16782 7052 16810
rect 6828 16720 6880 16726
rect 6828 16662 6880 16668
rect 6656 15966 6776 15994
rect 6656 15745 6684 15966
rect 6932 15910 6960 16782
rect 7012 16720 7064 16726
rect 7012 16662 7064 16668
rect 7024 16250 7052 16662
rect 7012 16244 7064 16250
rect 7012 16186 7064 16192
rect 6736 15904 6788 15910
rect 6736 15846 6788 15852
rect 6920 15904 6972 15910
rect 6920 15846 6972 15852
rect 6642 15736 6698 15745
rect 6642 15671 6698 15680
rect 6460 15564 6512 15570
rect 6564 15558 6684 15586
rect 6460 15506 6512 15512
rect 6472 14822 6500 15506
rect 6550 15056 6606 15065
rect 6550 14991 6606 15000
rect 6460 14816 6512 14822
rect 6460 14758 6512 14764
rect 6472 12850 6500 14758
rect 6564 14482 6592 14991
rect 6552 14476 6604 14482
rect 6552 14418 6604 14424
rect 6564 14006 6592 14418
rect 6552 14000 6604 14006
rect 6552 13942 6604 13948
rect 6656 13705 6684 15558
rect 6642 13696 6698 13705
rect 6642 13631 6698 13640
rect 6552 13184 6604 13190
rect 6552 13126 6604 13132
rect 6460 12844 6512 12850
rect 6460 12786 6512 12792
rect 6380 12702 6500 12730
rect 6288 12600 6408 12628
rect 6276 12164 6328 12170
rect 6276 12106 6328 12112
rect 6288 11898 6316 12106
rect 6276 11892 6328 11898
rect 6276 11834 6328 11840
rect 6276 8832 6328 8838
rect 6274 8800 6276 8809
rect 6328 8800 6330 8809
rect 6274 8735 6330 8744
rect 6380 8294 6408 12600
rect 6368 8288 6420 8294
rect 6368 8230 6420 8236
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6380 6610 6408 8230
rect 6472 8129 6500 12702
rect 6564 12442 6592 13126
rect 6748 12617 6776 15846
rect 6932 15706 6960 15846
rect 6920 15700 6972 15706
rect 6920 15642 6972 15648
rect 6920 15564 6972 15570
rect 6920 15506 6972 15512
rect 6828 15360 6880 15366
rect 6828 15302 6880 15308
rect 6840 15042 6868 15302
rect 6932 15162 6960 15506
rect 7116 15201 7144 20878
rect 7102 15192 7158 15201
rect 6920 15156 6972 15162
rect 7102 15127 7158 15136
rect 6920 15098 6972 15104
rect 6840 15014 6960 15042
rect 6932 14958 6960 15014
rect 6920 14952 6972 14958
rect 6920 14894 6972 14900
rect 6932 14618 6960 14894
rect 7104 14884 7156 14890
rect 7104 14826 7156 14832
rect 6920 14612 6972 14618
rect 6920 14554 6972 14560
rect 7116 14550 7144 14826
rect 7104 14544 7156 14550
rect 7104 14486 7156 14492
rect 7116 13870 7144 14486
rect 7104 13864 7156 13870
rect 7102 13832 7104 13841
rect 7156 13832 7158 13841
rect 7102 13767 7158 13776
rect 6826 13696 6882 13705
rect 7208 13682 7236 22732
rect 7380 22160 7432 22166
rect 7380 22102 7432 22108
rect 7392 21690 7420 22102
rect 7380 21684 7432 21690
rect 7380 21626 7432 21632
rect 7380 20800 7432 20806
rect 7380 20742 7432 20748
rect 7392 20058 7420 20742
rect 7380 20052 7432 20058
rect 7380 19994 7432 20000
rect 7288 19984 7340 19990
rect 7288 19926 7340 19932
rect 7300 19378 7328 19926
rect 7380 19712 7432 19718
rect 7380 19654 7432 19660
rect 7288 19372 7340 19378
rect 7288 19314 7340 19320
rect 7300 18086 7328 19314
rect 7392 19174 7420 19654
rect 7380 19168 7432 19174
rect 7380 19110 7432 19116
rect 7288 18080 7340 18086
rect 7288 18022 7340 18028
rect 7288 17740 7340 17746
rect 7288 17682 7340 17688
rect 7300 16794 7328 17682
rect 7380 17672 7432 17678
rect 7380 17614 7432 17620
rect 7392 17338 7420 17614
rect 7380 17332 7432 17338
rect 7380 17274 7432 17280
rect 7288 16788 7340 16794
rect 7288 16730 7340 16736
rect 7286 15600 7342 15609
rect 7286 15535 7342 15544
rect 6826 13631 6882 13640
rect 6932 13654 7236 13682
rect 6734 12608 6790 12617
rect 6734 12543 6790 12552
rect 6552 12436 6604 12442
rect 6552 12378 6604 12384
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 6564 11218 6592 12038
rect 6644 11280 6696 11286
rect 6644 11222 6696 11228
rect 6552 11212 6604 11218
rect 6552 11154 6604 11160
rect 6564 8974 6592 11154
rect 6656 10470 6684 11222
rect 6644 10464 6696 10470
rect 6644 10406 6696 10412
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6552 8832 6604 8838
rect 6552 8774 6604 8780
rect 6458 8120 6514 8129
rect 6458 8055 6514 8064
rect 6472 7546 6500 8055
rect 6460 7540 6512 7546
rect 6460 7482 6512 7488
rect 6472 7274 6500 7482
rect 6460 7268 6512 7274
rect 6460 7210 6512 7216
rect 6564 6730 6592 8774
rect 6656 8430 6684 8978
rect 6644 8424 6696 8430
rect 6642 8392 6644 8401
rect 6696 8392 6698 8401
rect 6642 8327 6698 8336
rect 6644 8288 6696 8294
rect 6644 8230 6696 8236
rect 6656 7750 6684 8230
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 6656 7585 6684 7686
rect 6642 7576 6698 7585
rect 6748 7546 6776 12543
rect 6840 12481 6868 13631
rect 6826 12472 6882 12481
rect 6826 12407 6882 12416
rect 6826 10568 6882 10577
rect 6826 10503 6828 10512
rect 6880 10503 6882 10512
rect 6828 10474 6880 10480
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 6932 8922 6960 13654
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 7116 13190 7144 13330
rect 7104 13184 7156 13190
rect 7104 13126 7156 13132
rect 7012 12640 7064 12646
rect 7012 12582 7064 12588
rect 7024 12306 7052 12582
rect 7116 12442 7144 13126
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 7208 11830 7236 12174
rect 7196 11824 7248 11830
rect 7196 11766 7248 11772
rect 7300 11558 7328 15535
rect 7380 13796 7432 13802
rect 7380 13738 7432 13744
rect 7392 13161 7420 13738
rect 7378 13152 7434 13161
rect 7378 13087 7434 13096
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 7392 11898 7420 12242
rect 7380 11892 7432 11898
rect 7380 11834 7432 11840
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 7288 11552 7340 11558
rect 7288 11494 7340 11500
rect 7392 11286 7420 11630
rect 7380 11280 7432 11286
rect 7010 11248 7066 11257
rect 7380 11222 7432 11228
rect 7010 11183 7066 11192
rect 7024 9024 7052 11183
rect 7194 10704 7250 10713
rect 7194 10639 7250 10648
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 7116 10033 7144 10406
rect 7102 10024 7158 10033
rect 7102 9959 7104 9968
rect 7156 9959 7158 9968
rect 7104 9930 7156 9936
rect 7208 9654 7236 10639
rect 7196 9648 7248 9654
rect 7196 9590 7248 9596
rect 7208 9489 7236 9590
rect 7194 9480 7250 9489
rect 7194 9415 7250 9424
rect 7024 8996 7236 9024
rect 6840 8566 6868 8910
rect 6932 8894 7144 8922
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 6840 8022 6868 8502
rect 6932 8362 6960 8774
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 7116 8265 7144 8894
rect 7102 8256 7158 8265
rect 7102 8191 7158 8200
rect 6828 8016 6880 8022
rect 6828 7958 6880 7964
rect 7012 7812 7064 7818
rect 7012 7754 7064 7760
rect 6642 7511 6698 7520
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6748 7342 6776 7482
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 6826 7304 6882 7313
rect 6826 7239 6882 7248
rect 6840 7206 6868 7239
rect 6828 7200 6880 7206
rect 6828 7142 6880 7148
rect 6552 6724 6604 6730
rect 6552 6666 6604 6672
rect 6288 6322 6316 6598
rect 6380 6582 6500 6610
rect 6276 6316 6328 6322
rect 6276 6258 6328 6264
rect 6288 5710 6316 6258
rect 6368 6248 6420 6254
rect 6368 6190 6420 6196
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 6288 4826 6316 5646
rect 6380 5234 6408 6190
rect 6368 5228 6420 5234
rect 6368 5170 6420 5176
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6276 4820 6328 4826
rect 6276 4762 6328 4768
rect 6380 4282 6408 4966
rect 6368 4276 6420 4282
rect 6368 4218 6420 4224
rect 6380 3670 6408 4218
rect 6368 3664 6420 3670
rect 6368 3606 6420 3612
rect 6380 3126 6408 3606
rect 6472 3466 6500 6582
rect 6564 5914 6592 6666
rect 6828 6384 6880 6390
rect 6826 6352 6828 6361
rect 6880 6352 6882 6361
rect 6826 6287 6882 6296
rect 6840 6118 6868 6287
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6920 6112 6972 6118
rect 6920 6054 6972 6060
rect 6932 5953 6960 6054
rect 6918 5944 6974 5953
rect 6552 5908 6604 5914
rect 6918 5879 6920 5888
rect 6552 5850 6604 5856
rect 6972 5879 6974 5888
rect 6920 5850 6972 5856
rect 6552 5160 6604 5166
rect 6552 5102 6604 5108
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 6368 3120 6420 3126
rect 6368 3062 6420 3068
rect 6368 2440 6420 2446
rect 6366 2408 6368 2417
rect 6420 2408 6422 2417
rect 6366 2343 6422 2352
rect 6000 604 6052 610
rect 6000 546 6052 552
rect 6184 604 6236 610
rect 6184 546 6236 552
rect 6012 480 6040 546
rect 6564 480 6592 5102
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6840 4826 6868 4966
rect 6828 4820 6880 4826
rect 6828 4762 6880 4768
rect 6826 4040 6882 4049
rect 6826 3975 6882 3984
rect 6840 3942 6868 3975
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 6656 2650 6684 3878
rect 7024 3618 7052 7754
rect 7102 7712 7158 7721
rect 7102 7647 7158 7656
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 6840 3590 7052 3618
rect 7116 3602 7144 7647
rect 7208 5166 7236 8996
rect 7380 7404 7432 7410
rect 7380 7346 7432 7352
rect 7392 7002 7420 7346
rect 7380 6996 7432 7002
rect 7300 6956 7380 6984
rect 7300 6497 7328 6956
rect 7380 6938 7432 6944
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7286 6488 7342 6497
rect 7286 6423 7342 6432
rect 7286 6080 7342 6089
rect 7286 6015 7342 6024
rect 7300 5370 7328 6015
rect 7288 5364 7340 5370
rect 7288 5306 7340 5312
rect 7196 5160 7248 5166
rect 7196 5102 7248 5108
rect 7208 4690 7236 5102
rect 7300 5030 7328 5306
rect 7288 5024 7340 5030
rect 7288 4966 7340 4972
rect 7288 4820 7340 4826
rect 7288 4762 7340 4768
rect 7196 4684 7248 4690
rect 7196 4626 7248 4632
rect 7300 4146 7328 4762
rect 7288 4140 7340 4146
rect 7288 4082 7340 4088
rect 7196 3936 7248 3942
rect 7392 3913 7420 6598
rect 7196 3878 7248 3884
rect 7378 3904 7434 3913
rect 7208 3738 7236 3878
rect 7378 3839 7434 3848
rect 7196 3732 7248 3738
rect 7196 3674 7248 3680
rect 7104 3596 7156 3602
rect 6748 3505 6776 3538
rect 6840 3534 6868 3590
rect 7104 3538 7156 3544
rect 6828 3528 6880 3534
rect 6734 3496 6790 3505
rect 6828 3470 6880 3476
rect 6734 3431 6790 3440
rect 7104 3460 7156 3466
rect 6748 3194 6776 3431
rect 7104 3402 7156 3408
rect 6736 3188 6788 3194
rect 6736 3130 6788 3136
rect 6828 2984 6880 2990
rect 6828 2926 6880 2932
rect 6644 2644 6696 2650
rect 6644 2586 6696 2592
rect 6840 2514 6868 2926
rect 6828 2508 6880 2514
rect 6828 2450 6880 2456
rect 7116 480 7144 3402
rect 7484 3097 7512 23684
rect 7564 23588 7616 23594
rect 7564 23530 7616 23536
rect 7576 23322 7604 23530
rect 7564 23316 7616 23322
rect 7564 23258 7616 23264
rect 7576 22642 7604 23258
rect 7656 23180 7708 23186
rect 7656 23122 7708 23128
rect 7564 22636 7616 22642
rect 7564 22578 7616 22584
rect 7668 22574 7696 23122
rect 7656 22568 7708 22574
rect 7656 22510 7708 22516
rect 7668 22098 7696 22510
rect 7656 22092 7708 22098
rect 7656 22034 7708 22040
rect 7656 21888 7708 21894
rect 7656 21830 7708 21836
rect 7668 21457 7696 21830
rect 7654 21448 7710 21457
rect 7654 21383 7710 21392
rect 7840 20936 7892 20942
rect 7840 20878 7892 20884
rect 7852 20534 7880 20878
rect 7840 20528 7892 20534
rect 7840 20470 7892 20476
rect 7748 20324 7800 20330
rect 7748 20266 7800 20272
rect 7760 19854 7788 20266
rect 7748 19848 7800 19854
rect 7748 19790 7800 19796
rect 7564 19168 7616 19174
rect 7564 19110 7616 19116
rect 7576 16250 7604 19110
rect 7760 18970 7788 19790
rect 7748 18964 7800 18970
rect 7748 18906 7800 18912
rect 7654 18184 7710 18193
rect 7654 18119 7710 18128
rect 7840 18148 7892 18154
rect 7564 16244 7616 16250
rect 7564 16186 7616 16192
rect 7564 16108 7616 16114
rect 7564 16050 7616 16056
rect 7576 15366 7604 16050
rect 7564 15360 7616 15366
rect 7564 15302 7616 15308
rect 7576 14550 7604 15302
rect 7564 14544 7616 14550
rect 7564 14486 7616 14492
rect 7668 13410 7696 18119
rect 7840 18090 7892 18096
rect 7746 18048 7802 18057
rect 7746 17983 7802 17992
rect 7760 15706 7788 17983
rect 7852 17542 7880 18090
rect 7840 17536 7892 17542
rect 7840 17478 7892 17484
rect 7838 17232 7894 17241
rect 7838 17167 7894 17176
rect 7852 17134 7880 17167
rect 7840 17128 7892 17134
rect 7840 17070 7892 17076
rect 7840 16448 7892 16454
rect 7840 16390 7892 16396
rect 7852 15706 7880 16390
rect 7748 15700 7800 15706
rect 7748 15642 7800 15648
rect 7840 15700 7892 15706
rect 7840 15642 7892 15648
rect 7748 14340 7800 14346
rect 7748 14282 7800 14288
rect 7760 14074 7788 14282
rect 7748 14068 7800 14074
rect 7748 14010 7800 14016
rect 7760 13954 7788 14010
rect 7760 13926 7880 13954
rect 7852 13870 7880 13926
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 7668 13382 7788 13410
rect 7564 13320 7616 13326
rect 7564 13262 7616 13268
rect 7656 13320 7708 13326
rect 7656 13262 7708 13268
rect 7576 12986 7604 13262
rect 7668 12986 7696 13262
rect 7564 12980 7616 12986
rect 7564 12922 7616 12928
rect 7656 12980 7708 12986
rect 7656 12922 7708 12928
rect 7576 10810 7604 12922
rect 7668 12850 7696 12922
rect 7656 12844 7708 12850
rect 7656 12786 7708 12792
rect 7564 10804 7616 10810
rect 7564 10746 7616 10752
rect 7760 9654 7788 13382
rect 7840 12096 7892 12102
rect 7840 12038 7892 12044
rect 7852 11626 7880 12038
rect 7840 11620 7892 11626
rect 7840 11562 7892 11568
rect 7852 11354 7880 11562
rect 7840 11348 7892 11354
rect 7840 11290 7892 11296
rect 7748 9648 7800 9654
rect 7748 9590 7800 9596
rect 7944 8072 7972 24806
rect 8864 24698 8892 27520
rect 9416 27470 9444 27520
rect 8944 27464 8996 27470
rect 8944 27406 8996 27412
rect 9404 27464 9456 27470
rect 9404 27406 9456 27412
rect 8772 24670 8892 24698
rect 8668 24200 8720 24206
rect 8666 24168 8668 24177
rect 8720 24168 8722 24177
rect 8666 24103 8722 24112
rect 8116 24064 8168 24070
rect 8116 24006 8168 24012
rect 8024 22160 8076 22166
rect 8022 22128 8024 22137
rect 8076 22128 8078 22137
rect 8022 22063 8078 22072
rect 8128 22030 8156 24006
rect 8576 22772 8628 22778
rect 8680 22760 8708 24103
rect 8628 22732 8708 22760
rect 8576 22714 8628 22720
rect 8680 22574 8708 22732
rect 8668 22568 8720 22574
rect 8482 22536 8538 22545
rect 8668 22510 8720 22516
rect 8482 22471 8538 22480
rect 8392 22092 8444 22098
rect 8392 22034 8444 22040
rect 8116 22024 8168 22030
rect 8116 21966 8168 21972
rect 8024 21956 8076 21962
rect 8024 21898 8076 21904
rect 8036 21418 8064 21898
rect 8024 21412 8076 21418
rect 8024 21354 8076 21360
rect 8036 20942 8064 21354
rect 8404 21146 8432 22034
rect 8392 21140 8444 21146
rect 8392 21082 8444 21088
rect 8208 21004 8260 21010
rect 8208 20946 8260 20952
rect 8024 20936 8076 20942
rect 8024 20878 8076 20884
rect 8036 20262 8064 20878
rect 8220 20602 8248 20946
rect 8208 20596 8260 20602
rect 8208 20538 8260 20544
rect 8024 20256 8076 20262
rect 8024 20198 8076 20204
rect 8390 20088 8446 20097
rect 8390 20023 8446 20032
rect 8300 19916 8352 19922
rect 8300 19858 8352 19864
rect 8022 19816 8078 19825
rect 8022 19751 8078 19760
rect 8036 13530 8064 19751
rect 8208 19372 8260 19378
rect 8208 19314 8260 19320
rect 8220 19009 8248 19314
rect 8312 19174 8340 19858
rect 8300 19168 8352 19174
rect 8300 19110 8352 19116
rect 8206 19000 8262 19009
rect 8312 18970 8340 19110
rect 8206 18935 8208 18944
rect 8260 18935 8262 18944
rect 8300 18964 8352 18970
rect 8208 18906 8260 18912
rect 8300 18906 8352 18912
rect 8220 18426 8248 18906
rect 8404 18698 8432 20023
rect 8392 18692 8444 18698
rect 8392 18634 8444 18640
rect 8208 18420 8260 18426
rect 8208 18362 8260 18368
rect 8496 18193 8524 22471
rect 8772 22438 8800 24670
rect 8852 24608 8904 24614
rect 8852 24550 8904 24556
rect 8864 24449 8892 24550
rect 8850 24440 8906 24449
rect 8850 24375 8906 24384
rect 8956 23304 8984 27406
rect 9496 25424 9548 25430
rect 9496 25366 9548 25372
rect 9508 24750 9536 25366
rect 9968 24834 9996 27520
rect 10520 25786 10548 27520
rect 10520 25758 10824 25786
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 9876 24806 9996 24834
rect 9496 24744 9548 24750
rect 9496 24686 9548 24692
rect 9312 24404 9364 24410
rect 9312 24346 9364 24352
rect 9036 24268 9088 24274
rect 9036 24210 9088 24216
rect 9048 23905 9076 24210
rect 9034 23896 9090 23905
rect 9324 23866 9352 24346
rect 9678 24304 9734 24313
rect 9678 24239 9734 24248
rect 9034 23831 9036 23840
rect 9088 23831 9090 23840
rect 9312 23860 9364 23866
rect 9036 23802 9088 23808
rect 9312 23802 9364 23808
rect 9494 23760 9550 23769
rect 9494 23695 9550 23704
rect 8864 23276 8984 23304
rect 8760 22432 8812 22438
rect 8760 22374 8812 22380
rect 8576 20256 8628 20262
rect 8576 20198 8628 20204
rect 8588 19718 8616 20198
rect 8864 19825 8892 23276
rect 8942 23216 8998 23225
rect 8942 23151 8998 23160
rect 8850 19816 8906 19825
rect 8850 19751 8906 19760
rect 8576 19712 8628 19718
rect 8576 19654 8628 19660
rect 8588 19378 8616 19654
rect 8576 19372 8628 19378
rect 8576 19314 8628 19320
rect 8760 19304 8812 19310
rect 8760 19246 8812 19252
rect 8576 18828 8628 18834
rect 8576 18770 8628 18776
rect 8482 18184 8538 18193
rect 8482 18119 8538 18128
rect 8588 18086 8616 18770
rect 8668 18420 8720 18426
rect 8668 18362 8720 18368
rect 8576 18080 8628 18086
rect 8576 18022 8628 18028
rect 8484 17672 8536 17678
rect 8484 17614 8536 17620
rect 8392 17536 8444 17542
rect 8392 17478 8444 17484
rect 8300 16992 8352 16998
rect 8300 16934 8352 16940
rect 8312 16726 8340 16934
rect 8300 16720 8352 16726
rect 8300 16662 8352 16668
rect 8208 15564 8260 15570
rect 8208 15506 8260 15512
rect 8116 15428 8168 15434
rect 8116 15370 8168 15376
rect 8128 14890 8156 15370
rect 8116 14884 8168 14890
rect 8116 14826 8168 14832
rect 8220 14550 8248 15506
rect 8300 14816 8352 14822
rect 8300 14758 8352 14764
rect 8208 14544 8260 14550
rect 8208 14486 8260 14492
rect 8312 14278 8340 14758
rect 8208 14272 8260 14278
rect 8208 14214 8260 14220
rect 8300 14272 8352 14278
rect 8300 14214 8352 14220
rect 8220 14090 8248 14214
rect 8404 14090 8432 17478
rect 8496 16833 8524 17614
rect 8680 17338 8708 18362
rect 8772 18329 8800 19246
rect 8852 19168 8904 19174
rect 8852 19110 8904 19116
rect 8864 18873 8892 19110
rect 8850 18864 8906 18873
rect 8850 18799 8906 18808
rect 8850 18592 8906 18601
rect 8850 18527 8906 18536
rect 8758 18320 8814 18329
rect 8758 18255 8814 18264
rect 8760 17604 8812 17610
rect 8760 17546 8812 17552
rect 8668 17332 8720 17338
rect 8668 17274 8720 17280
rect 8482 16824 8538 16833
rect 8482 16759 8538 16768
rect 8680 16697 8708 17274
rect 8772 17134 8800 17546
rect 8760 17128 8812 17134
rect 8760 17070 8812 17076
rect 8772 16726 8800 17070
rect 8760 16720 8812 16726
rect 8666 16688 8722 16697
rect 8760 16662 8812 16668
rect 8666 16623 8722 16632
rect 8484 16584 8536 16590
rect 8484 16526 8536 16532
rect 8496 15162 8524 16526
rect 8484 15156 8536 15162
rect 8484 15098 8536 15104
rect 8496 14346 8524 15098
rect 8772 14958 8800 16662
rect 8760 14952 8812 14958
rect 8760 14894 8812 14900
rect 8484 14340 8536 14346
rect 8484 14282 8536 14288
rect 8220 14062 8432 14090
rect 8312 13530 8340 14062
rect 8772 13870 8800 14894
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 8024 13524 8076 13530
rect 8024 13466 8076 13472
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 8206 13288 8262 13297
rect 8206 13223 8262 13232
rect 8116 13184 8168 13190
rect 8116 13126 8168 13132
rect 8128 12850 8156 13126
rect 8116 12844 8168 12850
rect 8116 12786 8168 12792
rect 8024 12708 8076 12714
rect 8024 12650 8076 12656
rect 8036 12238 8064 12650
rect 8024 12232 8076 12238
rect 8024 12174 8076 12180
rect 8036 11914 8064 12174
rect 8128 12102 8156 12786
rect 8116 12096 8168 12102
rect 8116 12038 8168 12044
rect 8036 11898 8156 11914
rect 8036 11892 8168 11898
rect 8036 11886 8116 11892
rect 8116 11834 8168 11840
rect 8220 11234 8248 13223
rect 8864 12374 8892 18527
rect 8956 18057 8984 23151
rect 9036 23112 9088 23118
rect 9036 23054 9088 23060
rect 9048 22506 9076 23054
rect 9036 22500 9088 22506
rect 9036 22442 9088 22448
rect 9048 21894 9076 22442
rect 9128 22024 9180 22030
rect 9128 21966 9180 21972
rect 9036 21888 9088 21894
rect 9036 21830 9088 21836
rect 9048 21486 9076 21830
rect 9036 21480 9088 21486
rect 9036 21422 9088 21428
rect 9048 20806 9076 21422
rect 9140 21418 9168 21966
rect 9128 21412 9180 21418
rect 9128 21354 9180 21360
rect 9140 21185 9168 21354
rect 9312 21344 9364 21350
rect 9364 21304 9444 21332
rect 9312 21286 9364 21292
rect 9126 21176 9182 21185
rect 9126 21111 9182 21120
rect 9416 20806 9444 21304
rect 9036 20800 9088 20806
rect 9036 20742 9088 20748
rect 9404 20800 9456 20806
rect 9404 20742 9456 20748
rect 9048 20398 9076 20742
rect 9036 20392 9088 20398
rect 9036 20334 9088 20340
rect 9048 19718 9076 20334
rect 9416 20330 9444 20742
rect 9508 20641 9536 23695
rect 9692 23361 9720 24239
rect 9678 23352 9734 23361
rect 9678 23287 9734 23296
rect 9588 22432 9640 22438
rect 9588 22374 9640 22380
rect 9600 22098 9628 22374
rect 9588 22092 9640 22098
rect 9588 22034 9640 22040
rect 9772 21480 9824 21486
rect 9772 21422 9824 21428
rect 9680 21412 9732 21418
rect 9680 21354 9732 21360
rect 9494 20632 9550 20641
rect 9494 20567 9550 20576
rect 9404 20324 9456 20330
rect 9404 20266 9456 20272
rect 9126 20224 9182 20233
rect 9126 20159 9182 20168
rect 9140 19922 9168 20159
rect 9128 19916 9180 19922
rect 9128 19858 9180 19864
rect 9036 19712 9088 19718
rect 9036 19654 9088 19660
rect 8942 18048 8998 18057
rect 8942 17983 8998 17992
rect 9048 17610 9076 19654
rect 9140 19394 9168 19858
rect 9494 19544 9550 19553
rect 9494 19479 9550 19488
rect 9218 19408 9274 19417
rect 9140 19366 9218 19394
rect 9218 19343 9274 19352
rect 9232 18970 9260 19343
rect 9220 18964 9272 18970
rect 9220 18906 9272 18912
rect 9036 17604 9088 17610
rect 9036 17546 9088 17552
rect 9508 16946 9536 19479
rect 9692 18290 9720 21354
rect 9784 21350 9812 21422
rect 9772 21344 9824 21350
rect 9770 21312 9772 21321
rect 9824 21312 9826 21321
rect 9770 21247 9826 21256
rect 9772 20256 9824 20262
rect 9772 20198 9824 20204
rect 9680 18284 9732 18290
rect 9680 18226 9732 18232
rect 9784 17882 9812 20198
rect 9772 17876 9824 17882
rect 9772 17818 9824 17824
rect 9770 17776 9826 17785
rect 9770 17711 9826 17720
rect 9680 17536 9732 17542
rect 9680 17478 9732 17484
rect 9588 17128 9640 17134
rect 9586 17096 9588 17105
rect 9640 17096 9642 17105
rect 9586 17031 9642 17040
rect 9508 16918 9628 16946
rect 8942 16688 8998 16697
rect 8942 16623 8944 16632
rect 8996 16623 8998 16632
rect 8944 16594 8996 16600
rect 9220 16108 9272 16114
rect 9220 16050 9272 16056
rect 9128 15904 9180 15910
rect 9128 15846 9180 15852
rect 8944 14884 8996 14890
rect 8944 14826 8996 14832
rect 8956 14074 8984 14826
rect 8944 14068 8996 14074
rect 8944 14010 8996 14016
rect 8852 12368 8904 12374
rect 8852 12310 8904 12316
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 7760 8044 7972 8072
rect 8036 11206 8248 11234
rect 8404 11218 8432 12038
rect 8576 11892 8628 11898
rect 8576 11834 8628 11840
rect 8392 11212 8444 11218
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7576 7449 7604 7686
rect 7562 7440 7618 7449
rect 7562 7375 7618 7384
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 7668 6322 7696 6734
rect 7656 6316 7708 6322
rect 7656 6258 7708 6264
rect 7668 5914 7696 6258
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 7760 4457 7788 8044
rect 7838 7984 7894 7993
rect 7838 7919 7894 7928
rect 7852 7886 7880 7919
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 7852 7546 7880 7822
rect 7840 7540 7892 7546
rect 7840 7482 7892 7488
rect 8036 6866 8064 11206
rect 8392 11154 8444 11160
rect 8208 11076 8260 11082
rect 8208 11018 8260 11024
rect 8220 10266 8248 11018
rect 8392 11008 8444 11014
rect 8392 10950 8444 10956
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 8116 9580 8168 9586
rect 8116 9522 8168 9528
rect 8128 9489 8156 9522
rect 8220 9518 8248 10202
rect 8404 9926 8432 10950
rect 8588 10674 8616 11834
rect 9140 11286 9168 15846
rect 9232 15366 9260 16050
rect 9600 15586 9628 16918
rect 9692 15706 9720 17478
rect 9784 16794 9812 17711
rect 9772 16788 9824 16794
rect 9772 16730 9824 16736
rect 9772 16584 9824 16590
rect 9772 16526 9824 16532
rect 9784 16250 9812 16526
rect 9772 16244 9824 16250
rect 9772 16186 9824 16192
rect 9772 15904 9824 15910
rect 9772 15846 9824 15852
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 9784 15609 9812 15846
rect 9770 15600 9826 15609
rect 9600 15558 9720 15586
rect 9220 15360 9272 15366
rect 9220 15302 9272 15308
rect 9588 15360 9640 15366
rect 9588 15302 9640 15308
rect 9600 14822 9628 15302
rect 9588 14816 9640 14822
rect 9588 14758 9640 14764
rect 9404 14272 9456 14278
rect 9404 14214 9456 14220
rect 9220 13864 9272 13870
rect 9220 13806 9272 13812
rect 9232 13530 9260 13806
rect 9220 13524 9272 13530
rect 9220 13466 9272 13472
rect 9416 13002 9444 14214
rect 9692 13954 9720 15558
rect 9770 15535 9826 15544
rect 9772 14340 9824 14346
rect 9772 14282 9824 14288
rect 9784 14074 9812 14282
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9692 13926 9812 13954
rect 9416 12974 9720 13002
rect 9692 12442 9720 12974
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9692 11898 9720 12174
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9496 11756 9548 11762
rect 9496 11698 9548 11704
rect 9312 11552 9364 11558
rect 9312 11494 9364 11500
rect 9128 11280 9180 11286
rect 9128 11222 9180 11228
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 8588 10198 8616 10610
rect 9324 10606 9352 11494
rect 9508 11354 9536 11698
rect 9496 11348 9548 11354
rect 9692 11336 9720 11834
rect 9496 11290 9548 11296
rect 9600 11308 9720 11336
rect 9312 10600 9364 10606
rect 9312 10542 9364 10548
rect 8944 10464 8996 10470
rect 8944 10406 8996 10412
rect 8576 10192 8628 10198
rect 8482 10160 8538 10169
rect 8576 10134 8628 10140
rect 8482 10095 8538 10104
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8208 9512 8260 9518
rect 8114 9480 8170 9489
rect 8208 9454 8260 9460
rect 8114 9415 8170 9424
rect 8496 9178 8524 10095
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 8208 9036 8260 9042
rect 8208 8978 8260 8984
rect 8220 8566 8248 8978
rect 8208 8560 8260 8566
rect 8206 8528 8208 8537
rect 8852 8560 8904 8566
rect 8260 8528 8262 8537
rect 8852 8502 8904 8508
rect 8206 8463 8262 8472
rect 8220 8090 8248 8463
rect 8576 8424 8628 8430
rect 8864 8401 8892 8502
rect 8576 8366 8628 8372
rect 8850 8392 8906 8401
rect 8588 8294 8616 8366
rect 8850 8327 8906 8336
rect 8576 8288 8628 8294
rect 8576 8230 8628 8236
rect 8864 8090 8892 8327
rect 8208 8084 8260 8090
rect 8208 8026 8260 8032
rect 8852 8084 8904 8090
rect 8852 8026 8904 8032
rect 8116 7948 8168 7954
rect 8168 7908 8248 7936
rect 8116 7890 8168 7896
rect 8220 7206 8248 7908
rect 8668 7880 8720 7886
rect 8666 7848 8668 7857
rect 8720 7848 8722 7857
rect 8666 7783 8722 7792
rect 8680 7585 8708 7783
rect 8666 7576 8722 7585
rect 8666 7511 8668 7520
rect 8720 7511 8722 7520
rect 8668 7482 8720 7488
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 8208 7200 8260 7206
rect 8208 7142 8260 7148
rect 8220 6905 8248 7142
rect 8680 7002 8708 7346
rect 8668 6996 8720 7002
rect 8668 6938 8720 6944
rect 8300 6928 8352 6934
rect 8206 6896 8262 6905
rect 8024 6860 8076 6866
rect 8300 6870 8352 6876
rect 8206 6831 8262 6840
rect 8024 6802 8076 6808
rect 8036 6458 8064 6802
rect 8312 6458 8340 6870
rect 8024 6452 8076 6458
rect 8300 6452 8352 6458
rect 8076 6412 8156 6440
rect 8024 6394 8076 6400
rect 8022 6216 8078 6225
rect 8022 6151 8078 6160
rect 8036 5914 8064 6151
rect 8024 5908 8076 5914
rect 8024 5850 8076 5856
rect 8128 5794 8156 6412
rect 8300 6394 8352 6400
rect 8576 6452 8628 6458
rect 8576 6394 8628 6400
rect 8036 5766 8156 5794
rect 8392 5772 8444 5778
rect 7840 5568 7892 5574
rect 7840 5510 7892 5516
rect 7746 4448 7802 4457
rect 7746 4383 7802 4392
rect 7470 3088 7526 3097
rect 7470 3023 7526 3032
rect 7852 2417 7880 5510
rect 7932 5024 7984 5030
rect 7930 4992 7932 5001
rect 7984 4992 7986 5001
rect 7930 4927 7986 4936
rect 7932 4684 7984 4690
rect 7932 4626 7984 4632
rect 7944 3738 7972 4626
rect 7932 3732 7984 3738
rect 7932 3674 7984 3680
rect 7838 2408 7894 2417
rect 7838 2343 7894 2352
rect 7654 1864 7710 1873
rect 7654 1799 7710 1808
rect 7668 480 7696 1799
rect 8036 1306 8064 5766
rect 8392 5714 8444 5720
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8208 5024 8260 5030
rect 8312 5012 8340 5646
rect 8404 5030 8432 5714
rect 8588 5234 8616 6394
rect 8680 6254 8708 6938
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 8576 5228 8628 5234
rect 8576 5170 8628 5176
rect 8260 4984 8340 5012
rect 8392 5024 8444 5030
rect 8208 4966 8260 4972
rect 8392 4966 8444 4972
rect 8208 4684 8260 4690
rect 8208 4626 8260 4632
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 8128 4078 8156 4558
rect 8116 4072 8168 4078
rect 8116 4014 8168 4020
rect 8220 3924 8248 4626
rect 8300 3936 8352 3942
rect 8220 3896 8300 3924
rect 8300 3878 8352 3884
rect 8312 3738 8340 3878
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 8404 3602 8432 4966
rect 8588 4146 8616 5170
rect 8668 5092 8720 5098
rect 8668 5034 8720 5040
rect 8680 4826 8708 5034
rect 8668 4820 8720 4826
rect 8668 4762 8720 4768
rect 8850 4176 8906 4185
rect 8576 4140 8628 4146
rect 8850 4111 8906 4120
rect 8576 4082 8628 4088
rect 8392 3596 8444 3602
rect 8392 3538 8444 3544
rect 8404 3194 8432 3538
rect 8392 3188 8444 3194
rect 8392 3130 8444 3136
rect 8404 2961 8432 3130
rect 8390 2952 8446 2961
rect 8390 2887 8446 2896
rect 8208 2848 8260 2854
rect 8208 2790 8260 2796
rect 8220 2650 8248 2790
rect 8208 2644 8260 2650
rect 8208 2586 8260 2592
rect 8588 2514 8616 4082
rect 8760 3596 8812 3602
rect 8760 3538 8812 3544
rect 8772 3233 8800 3538
rect 8758 3224 8814 3233
rect 8758 3159 8814 3168
rect 8772 2854 8800 3159
rect 8760 2848 8812 2854
rect 8758 2816 8760 2825
rect 8812 2816 8814 2825
rect 8758 2751 8814 2760
rect 8576 2508 8628 2514
rect 8576 2450 8628 2456
rect 8036 1278 8248 1306
rect 8220 480 8248 1278
rect 8864 480 8892 4111
rect 8956 2961 8984 10406
rect 9600 10146 9628 11308
rect 9600 10118 9720 10146
rect 9404 9920 9456 9926
rect 9404 9862 9456 9868
rect 9128 9648 9180 9654
rect 9128 9590 9180 9596
rect 9140 8362 9168 9590
rect 9220 9580 9272 9586
rect 9220 9522 9272 9528
rect 9232 9353 9260 9522
rect 9218 9344 9274 9353
rect 9218 9279 9274 9288
rect 9232 9178 9260 9279
rect 9416 9178 9444 9862
rect 9496 9376 9548 9382
rect 9496 9318 9548 9324
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 9404 9172 9456 9178
rect 9404 9114 9456 9120
rect 9508 8945 9536 9318
rect 9494 8936 9550 8945
rect 9494 8871 9550 8880
rect 9128 8356 9180 8362
rect 9128 8298 9180 8304
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 9310 7848 9366 7857
rect 9310 7783 9312 7792
rect 9364 7783 9366 7792
rect 9312 7754 9364 7760
rect 9324 7274 9352 7754
rect 9312 7268 9364 7274
rect 9312 7210 9364 7216
rect 9416 6730 9444 8230
rect 9692 8072 9720 10118
rect 9600 8044 9720 8072
rect 9600 7834 9628 8044
rect 9678 7984 9734 7993
rect 9678 7919 9680 7928
rect 9732 7919 9734 7928
rect 9680 7890 9732 7896
rect 9600 7806 9720 7834
rect 9588 7336 9640 7342
rect 9588 7278 9640 7284
rect 9496 7200 9548 7206
rect 9496 7142 9548 7148
rect 9404 6724 9456 6730
rect 9404 6666 9456 6672
rect 9416 6458 9444 6666
rect 9404 6452 9456 6458
rect 9404 6394 9456 6400
rect 9508 5930 9536 7142
rect 9600 7041 9628 7278
rect 9586 7032 9642 7041
rect 9586 6967 9588 6976
rect 9640 6967 9642 6976
rect 9588 6938 9640 6944
rect 9600 6907 9628 6938
rect 9692 6089 9720 7806
rect 9678 6080 9734 6089
rect 9678 6015 9734 6024
rect 9508 5914 9720 5930
rect 9508 5908 9732 5914
rect 9508 5902 9680 5908
rect 9034 5672 9090 5681
rect 9034 5607 9036 5616
rect 9088 5607 9090 5616
rect 9036 5578 9088 5584
rect 9508 4826 9536 5902
rect 9680 5850 9732 5856
rect 9784 4826 9812 13926
rect 9876 11626 9904 24806
rect 9956 24744 10008 24750
rect 9956 24686 10008 24692
rect 9968 24138 9996 24686
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10324 24268 10376 24274
rect 10324 24210 10376 24216
rect 10140 24200 10192 24206
rect 10140 24142 10192 24148
rect 9956 24132 10008 24138
rect 9956 24074 10008 24080
rect 9956 23656 10008 23662
rect 9956 23598 10008 23604
rect 9968 23118 9996 23598
rect 10152 23594 10180 24142
rect 10336 23594 10364 24210
rect 10140 23588 10192 23594
rect 10140 23530 10192 23536
rect 10324 23588 10376 23594
rect 10324 23530 10376 23536
rect 10152 23322 10180 23530
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10140 23316 10192 23322
rect 10140 23258 10192 23264
rect 10508 23248 10560 23254
rect 10508 23190 10560 23196
rect 9956 23112 10008 23118
rect 9956 23054 10008 23060
rect 10232 23112 10284 23118
rect 10232 23054 10284 23060
rect 10244 22506 10272 23054
rect 10520 22778 10548 23190
rect 10508 22772 10560 22778
rect 10508 22714 10560 22720
rect 10232 22500 10284 22506
rect 10232 22442 10284 22448
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10048 22092 10100 22098
rect 10048 22034 10100 22040
rect 9956 21344 10008 21350
rect 9956 21286 10008 21292
rect 9968 20058 9996 21286
rect 10060 21078 10088 22034
rect 10232 22024 10284 22030
rect 10232 21966 10284 21972
rect 10416 22024 10468 22030
rect 10416 21966 10468 21972
rect 10244 21865 10272 21966
rect 10230 21856 10286 21865
rect 10230 21791 10286 21800
rect 10428 21690 10456 21966
rect 10692 21888 10744 21894
rect 10692 21830 10744 21836
rect 10140 21684 10192 21690
rect 10140 21626 10192 21632
rect 10416 21684 10468 21690
rect 10416 21626 10468 21632
rect 10048 21072 10100 21078
rect 10048 21014 10100 21020
rect 10046 20496 10102 20505
rect 10046 20431 10102 20440
rect 9956 20052 10008 20058
rect 9956 19994 10008 20000
rect 9968 18970 9996 19994
rect 10060 19786 10088 20431
rect 10048 19780 10100 19786
rect 10048 19722 10100 19728
rect 10152 19009 10180 21626
rect 10704 21554 10732 21830
rect 10692 21548 10744 21554
rect 10692 21490 10744 21496
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10704 21010 10732 21490
rect 10692 21004 10744 21010
rect 10692 20946 10744 20952
rect 10704 20262 10732 20946
rect 10692 20256 10744 20262
rect 10692 20198 10744 20204
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10600 19984 10652 19990
rect 10600 19926 10652 19932
rect 10232 19848 10284 19854
rect 10232 19790 10284 19796
rect 10324 19848 10376 19854
rect 10324 19790 10376 19796
rect 10244 19446 10272 19790
rect 10336 19514 10364 19790
rect 10324 19508 10376 19514
rect 10324 19450 10376 19456
rect 10232 19440 10284 19446
rect 10232 19382 10284 19388
rect 10244 19310 10272 19382
rect 10232 19304 10284 19310
rect 10232 19246 10284 19252
rect 10612 19156 10640 19926
rect 10704 19378 10732 20198
rect 10692 19372 10744 19378
rect 10692 19314 10744 19320
rect 10612 19128 10732 19156
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10138 19000 10194 19009
rect 9956 18964 10008 18970
rect 9956 18906 10008 18912
rect 10048 18964 10100 18970
rect 10289 18992 10585 19012
rect 10138 18935 10194 18944
rect 10048 18906 10100 18912
rect 9954 18456 10010 18465
rect 10060 18426 10088 18906
rect 10140 18828 10192 18834
rect 10140 18770 10192 18776
rect 9954 18391 10010 18400
rect 10048 18420 10100 18426
rect 9968 18170 9996 18391
rect 10048 18362 10100 18368
rect 9968 18142 10088 18170
rect 9956 18080 10008 18086
rect 9956 18022 10008 18028
rect 9968 14550 9996 18022
rect 10060 16794 10088 18142
rect 10152 17542 10180 18770
rect 10600 18760 10652 18766
rect 10600 18702 10652 18708
rect 10612 18290 10640 18702
rect 10704 18358 10732 19128
rect 10692 18352 10744 18358
rect 10692 18294 10744 18300
rect 10600 18284 10652 18290
rect 10600 18226 10652 18232
rect 10612 18154 10640 18226
rect 10796 18170 10824 25758
rect 11072 23905 11100 27520
rect 11242 24168 11298 24177
rect 11242 24103 11298 24112
rect 11058 23896 11114 23905
rect 11256 23866 11284 24103
rect 11716 23905 11744 27520
rect 12268 24834 12296 27520
rect 12820 27418 12848 27520
rect 12728 27390 12848 27418
rect 12624 25288 12676 25294
rect 12624 25230 12676 25236
rect 11992 24806 12296 24834
rect 12636 24818 12664 25230
rect 12624 24812 12676 24818
rect 11702 23896 11758 23905
rect 11058 23831 11114 23840
rect 11244 23860 11296 23866
rect 11702 23831 11758 23840
rect 11244 23802 11296 23808
rect 10968 23520 11020 23526
rect 10968 23462 11020 23468
rect 10980 22234 11008 23462
rect 11242 22672 11298 22681
rect 11242 22607 11298 22616
rect 11060 22432 11112 22438
rect 11060 22374 11112 22380
rect 10968 22228 11020 22234
rect 10968 22170 11020 22176
rect 11072 22137 11100 22374
rect 11256 22137 11284 22607
rect 11058 22128 11114 22137
rect 11058 22063 11114 22072
rect 11242 22128 11298 22137
rect 11242 22063 11298 22072
rect 10968 21956 11020 21962
rect 10968 21898 11020 21904
rect 10876 21072 10928 21078
rect 10876 21014 10928 21020
rect 10888 19990 10916 21014
rect 10876 19984 10928 19990
rect 10876 19926 10928 19932
rect 10876 19712 10928 19718
rect 10876 19654 10928 19660
rect 10888 19553 10916 19654
rect 10874 19544 10930 19553
rect 10874 19479 10930 19488
rect 10980 18902 11008 21898
rect 11888 21548 11940 21554
rect 11888 21490 11940 21496
rect 11900 21350 11928 21490
rect 11888 21344 11940 21350
rect 11888 21286 11940 21292
rect 11612 20800 11664 20806
rect 11612 20742 11664 20748
rect 11336 20392 11388 20398
rect 11336 20334 11388 20340
rect 11348 19718 11376 20334
rect 11624 19922 11652 20742
rect 11900 20602 11928 21286
rect 11888 20596 11940 20602
rect 11888 20538 11940 20544
rect 11794 20360 11850 20369
rect 11794 20295 11850 20304
rect 11612 19916 11664 19922
rect 11612 19858 11664 19864
rect 11336 19712 11388 19718
rect 11336 19654 11388 19660
rect 11242 19544 11298 19553
rect 11242 19479 11298 19488
rect 11256 19310 11284 19479
rect 11244 19304 11296 19310
rect 11150 19272 11206 19281
rect 11244 19246 11296 19252
rect 11348 19242 11376 19654
rect 11624 19514 11652 19858
rect 11612 19508 11664 19514
rect 11612 19450 11664 19456
rect 11150 19207 11152 19216
rect 11204 19207 11206 19216
rect 11336 19236 11388 19242
rect 11152 19178 11204 19184
rect 11336 19178 11388 19184
rect 11242 19000 11298 19009
rect 11242 18935 11298 18944
rect 10968 18896 11020 18902
rect 10968 18838 11020 18844
rect 10876 18624 10928 18630
rect 10876 18566 10928 18572
rect 11152 18624 11204 18630
rect 11256 18601 11284 18935
rect 11152 18566 11204 18572
rect 11242 18592 11298 18601
rect 10600 18148 10652 18154
rect 10600 18090 10652 18096
rect 10704 18142 10824 18170
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10140 17536 10192 17542
rect 10140 17478 10192 17484
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10048 16788 10100 16794
rect 10100 16748 10180 16776
rect 10048 16730 10100 16736
rect 10048 16652 10100 16658
rect 10048 16594 10100 16600
rect 10060 15910 10088 16594
rect 10048 15904 10100 15910
rect 10048 15846 10100 15852
rect 10152 15570 10180 16748
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10704 15586 10732 18142
rect 10784 18080 10836 18086
rect 10784 18022 10836 18028
rect 10796 17785 10824 18022
rect 10888 17921 10916 18566
rect 11164 18222 11192 18566
rect 11242 18527 11298 18536
rect 11244 18352 11296 18358
rect 11244 18294 11296 18300
rect 11152 18216 11204 18222
rect 11152 18158 11204 18164
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 10874 17912 10930 17921
rect 10874 17847 10930 17856
rect 10968 17876 11020 17882
rect 11072 17864 11100 18022
rect 11020 17836 11100 17864
rect 10968 17818 11020 17824
rect 10876 17808 10928 17814
rect 10782 17776 10838 17785
rect 10876 17750 10928 17756
rect 10782 17711 10838 17720
rect 10888 17338 10916 17750
rect 10876 17332 10928 17338
rect 10796 17292 10876 17320
rect 10796 16114 10824 17292
rect 10876 17274 10928 17280
rect 10874 16824 10930 16833
rect 10874 16759 10876 16768
rect 10928 16759 10930 16768
rect 10876 16730 10928 16736
rect 10980 16250 11008 17818
rect 11164 16794 11192 18158
rect 11256 17649 11284 18294
rect 11348 17746 11376 19178
rect 11704 18828 11756 18834
rect 11704 18770 11756 18776
rect 11336 17740 11388 17746
rect 11336 17682 11388 17688
rect 11242 17640 11298 17649
rect 11242 17575 11298 17584
rect 11716 16998 11744 18770
rect 11520 16992 11572 16998
rect 11520 16934 11572 16940
rect 11704 16992 11756 16998
rect 11704 16934 11756 16940
rect 11242 16824 11298 16833
rect 11152 16788 11204 16794
rect 11242 16759 11298 16768
rect 11152 16730 11204 16736
rect 10968 16244 11020 16250
rect 10968 16186 11020 16192
rect 11152 16176 11204 16182
rect 11152 16118 11204 16124
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 10782 15736 10838 15745
rect 11164 15706 11192 16118
rect 11256 16114 11284 16759
rect 11532 16658 11560 16934
rect 11520 16652 11572 16658
rect 11520 16594 11572 16600
rect 11612 16652 11664 16658
rect 11612 16594 11664 16600
rect 11532 16250 11560 16594
rect 11520 16244 11572 16250
rect 11520 16186 11572 16192
rect 11244 16108 11296 16114
rect 11244 16050 11296 16056
rect 11520 15972 11572 15978
rect 11520 15914 11572 15920
rect 10782 15671 10784 15680
rect 10836 15671 10838 15680
rect 11152 15700 11204 15706
rect 10784 15642 10836 15648
rect 11152 15642 11204 15648
rect 10140 15564 10192 15570
rect 10704 15558 10916 15586
rect 10140 15506 10192 15512
rect 10784 15496 10836 15502
rect 10784 15438 10836 15444
rect 10796 15162 10824 15438
rect 10784 15156 10836 15162
rect 10784 15098 10836 15104
rect 10048 14816 10100 14822
rect 10048 14758 10100 14764
rect 9956 14544 10008 14550
rect 9956 14486 10008 14492
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 9968 12986 9996 13330
rect 9956 12980 10008 12986
rect 9956 12922 10008 12928
rect 10060 12424 10088 14758
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10692 13864 10744 13870
rect 10692 13806 10744 13812
rect 10782 13832 10838 13841
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 9968 12396 10088 12424
rect 10138 12472 10194 12481
rect 10289 12464 10585 12484
rect 10138 12407 10194 12416
rect 9864 11620 9916 11626
rect 9864 11562 9916 11568
rect 9864 11280 9916 11286
rect 9864 11222 9916 11228
rect 9876 10266 9904 11222
rect 9968 10606 9996 12396
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 10060 11694 10088 12242
rect 10048 11688 10100 11694
rect 10048 11630 10100 11636
rect 10060 11393 10088 11630
rect 10046 11384 10102 11393
rect 10046 11319 10102 11328
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 9956 10600 10008 10606
rect 9956 10542 10008 10548
rect 9864 10260 9916 10266
rect 9864 10202 9916 10208
rect 9968 10198 9996 10542
rect 10060 10266 10088 11154
rect 10152 11121 10180 12407
rect 10704 12209 10732 13806
rect 10782 13767 10838 13776
rect 10796 12238 10824 13767
rect 10888 12782 10916 15558
rect 11164 15502 11192 15642
rect 11428 15564 11480 15570
rect 11428 15506 11480 15512
rect 11152 15496 11204 15502
rect 11152 15438 11204 15444
rect 11242 15328 11298 15337
rect 11242 15263 11298 15272
rect 11060 14816 11112 14822
rect 11060 14758 11112 14764
rect 11072 14482 11100 14758
rect 11152 14612 11204 14618
rect 11152 14554 11204 14560
rect 11060 14476 11112 14482
rect 11060 14418 11112 14424
rect 11072 14074 11100 14418
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 11164 13802 11192 14554
rect 11256 13870 11284 15263
rect 11440 14822 11468 15506
rect 11532 14906 11560 15914
rect 11624 15706 11652 16594
rect 11716 16017 11744 16934
rect 11702 16008 11758 16017
rect 11702 15943 11758 15952
rect 11612 15700 11664 15706
rect 11612 15642 11664 15648
rect 11702 15600 11758 15609
rect 11702 15535 11704 15544
rect 11756 15535 11758 15544
rect 11704 15506 11756 15512
rect 11716 15162 11744 15506
rect 11704 15156 11756 15162
rect 11704 15098 11756 15104
rect 11610 14920 11666 14929
rect 11532 14878 11610 14906
rect 11610 14855 11666 14864
rect 11428 14816 11480 14822
rect 11334 14784 11390 14793
rect 11428 14758 11480 14764
rect 11334 14719 11390 14728
rect 11244 13864 11296 13870
rect 11244 13806 11296 13812
rect 11152 13796 11204 13802
rect 11152 13738 11204 13744
rect 10968 13728 11020 13734
rect 10968 13670 11020 13676
rect 10876 12776 10928 12782
rect 10876 12718 10928 12724
rect 10784 12232 10836 12238
rect 10690 12200 10746 12209
rect 10784 12174 10836 12180
rect 10690 12135 10746 12144
rect 10888 12102 10916 12718
rect 10980 12714 11008 13670
rect 11348 13297 11376 14719
rect 11334 13288 11390 13297
rect 11334 13223 11390 13232
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 11072 12850 11100 13126
rect 11060 12844 11112 12850
rect 11060 12786 11112 12792
rect 11072 12730 11100 12786
rect 10968 12708 11020 12714
rect 11072 12702 11192 12730
rect 10968 12650 11020 12656
rect 10876 12096 10928 12102
rect 10796 12044 10876 12050
rect 10796 12038 10928 12044
rect 10796 12022 10916 12038
rect 10692 11552 10744 11558
rect 10692 11494 10744 11500
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10704 11286 10732 11494
rect 10692 11280 10744 11286
rect 10692 11222 10744 11228
rect 10324 11144 10376 11150
rect 10138 11112 10194 11121
rect 10324 11086 10376 11092
rect 10138 11047 10194 11056
rect 10336 10810 10364 11086
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 10140 10532 10192 10538
rect 10140 10474 10192 10480
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 9956 10192 10008 10198
rect 9956 10134 10008 10140
rect 9968 9586 9996 10134
rect 9956 9580 10008 9586
rect 9956 9522 10008 9528
rect 10060 9450 10088 10202
rect 10152 10130 10180 10474
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10704 10198 10732 10746
rect 10692 10192 10744 10198
rect 10692 10134 10744 10140
rect 10140 10124 10192 10130
rect 10140 10066 10192 10072
rect 10598 9616 10654 9625
rect 10598 9551 10654 9560
rect 10612 9518 10640 9551
rect 10704 9518 10732 10134
rect 10796 9654 10824 12022
rect 10888 11973 10916 12022
rect 10876 11280 10928 11286
rect 10876 11222 10928 11228
rect 10784 9648 10836 9654
rect 10784 9590 10836 9596
rect 10140 9512 10192 9518
rect 10140 9454 10192 9460
rect 10600 9512 10652 9518
rect 10600 9454 10652 9460
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 9956 9444 10008 9450
rect 9956 9386 10008 9392
rect 10048 9444 10100 9450
rect 10048 9386 10100 9392
rect 9864 8968 9916 8974
rect 9864 8910 9916 8916
rect 9876 8634 9904 8910
rect 9968 8634 9996 9386
rect 10152 9081 10180 9454
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10138 9072 10194 9081
rect 10138 9007 10194 9016
rect 10046 8800 10102 8809
rect 10046 8735 10102 8744
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 9956 8628 10008 8634
rect 9956 8570 10008 8576
rect 9876 8430 9904 8570
rect 9864 8424 9916 8430
rect 9864 8366 9916 8372
rect 9954 8256 10010 8265
rect 9954 8191 10010 8200
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9496 4820 9548 4826
rect 9496 4762 9548 4768
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9876 4729 9904 7142
rect 9968 5370 9996 8191
rect 10060 5846 10088 8735
rect 10704 8498 10732 9454
rect 10784 9444 10836 9450
rect 10784 9386 10836 9392
rect 10796 8838 10824 9386
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10692 8492 10744 8498
rect 10692 8434 10744 8440
rect 10140 8356 10192 8362
rect 10140 8298 10192 8304
rect 10152 8090 10180 8298
rect 10692 8288 10744 8294
rect 10690 8256 10692 8265
rect 10744 8256 10746 8265
rect 10289 8188 10585 8208
rect 10690 8191 10746 8200
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10140 8084 10192 8090
rect 10140 8026 10192 8032
rect 10692 7744 10744 7750
rect 10692 7686 10744 7692
rect 10704 7274 10732 7686
rect 10140 7268 10192 7274
rect 10140 7210 10192 7216
rect 10692 7268 10744 7274
rect 10692 7210 10744 7216
rect 10152 7177 10180 7210
rect 10138 7168 10194 7177
rect 10138 7103 10194 7112
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 10336 6458 10364 6802
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 10690 6352 10746 6361
rect 10690 6287 10692 6296
rect 10744 6287 10746 6296
rect 10692 6258 10744 6264
rect 10140 6112 10192 6118
rect 10140 6054 10192 6060
rect 10048 5840 10100 5846
rect 10048 5782 10100 5788
rect 10152 5794 10180 6054
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10692 5840 10744 5846
rect 10690 5808 10692 5817
rect 10744 5808 10746 5817
rect 10152 5766 10272 5794
rect 10244 5710 10272 5766
rect 10690 5743 10746 5752
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 10140 5568 10192 5574
rect 10140 5510 10192 5516
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 9956 5024 10008 5030
rect 9956 4966 10008 4972
rect 9968 4758 9996 4966
rect 10048 4820 10100 4826
rect 10048 4762 10100 4768
rect 9956 4752 10008 4758
rect 9862 4720 9918 4729
rect 9956 4694 10008 4700
rect 9862 4655 9918 4664
rect 9772 4548 9824 4554
rect 9772 4490 9824 4496
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9496 4004 9548 4010
rect 9496 3946 9548 3952
rect 9402 3632 9458 3641
rect 9402 3567 9458 3576
rect 9310 3496 9366 3505
rect 9310 3431 9366 3440
rect 9324 3194 9352 3431
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 8942 2952 8998 2961
rect 8942 2887 8998 2896
rect 9416 480 9444 3567
rect 9508 3398 9536 3946
rect 9692 3534 9720 4422
rect 9680 3528 9732 3534
rect 9680 3470 9732 3476
rect 9496 3392 9548 3398
rect 9496 3334 9548 3340
rect 9508 3194 9536 3334
rect 9496 3188 9548 3194
rect 9496 3130 9548 3136
rect 9784 3058 9812 4490
rect 10060 4282 10088 4762
rect 10048 4276 10100 4282
rect 10048 4218 10100 4224
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 10060 3602 10088 3878
rect 10152 3670 10180 5510
rect 10244 5098 10272 5646
rect 10232 5092 10284 5098
rect 10232 5034 10284 5040
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 10244 4010 10272 4558
rect 10692 4480 10744 4486
rect 10692 4422 10744 4428
rect 10704 4049 10732 4422
rect 10690 4040 10746 4049
rect 10232 4004 10284 4010
rect 10690 3975 10746 3984
rect 10232 3946 10284 3952
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10140 3664 10192 3670
rect 10140 3606 10192 3612
rect 10048 3596 10100 3602
rect 10048 3538 10100 3544
rect 9772 3052 9824 3058
rect 9772 2994 9824 3000
rect 9864 3052 9916 3058
rect 9864 2994 9916 3000
rect 9876 2378 9904 2994
rect 10704 2990 10732 3975
rect 10692 2984 10744 2990
rect 10692 2926 10744 2932
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 9956 2644 10008 2650
rect 9956 2586 10008 2592
rect 9864 2372 9916 2378
rect 9864 2314 9916 2320
rect 9968 480 9996 2586
rect 10796 762 10824 8774
rect 10888 3754 10916 11222
rect 10980 9450 11008 12650
rect 11060 12640 11112 12646
rect 11060 12582 11112 12588
rect 11072 12238 11100 12582
rect 11164 12442 11192 12702
rect 11152 12436 11204 12442
rect 11152 12378 11204 12384
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 11244 12232 11296 12238
rect 11244 12174 11296 12180
rect 11256 11354 11284 12174
rect 11440 11801 11468 14758
rect 11520 14408 11572 14414
rect 11520 14350 11572 14356
rect 11532 13530 11560 14350
rect 11624 13954 11652 14855
rect 11704 14408 11756 14414
rect 11704 14350 11756 14356
rect 11716 14074 11744 14350
rect 11704 14068 11756 14074
rect 11704 14010 11756 14016
rect 11624 13926 11744 13954
rect 11520 13524 11572 13530
rect 11520 13466 11572 13472
rect 11532 12442 11560 13466
rect 11520 12436 11572 12442
rect 11520 12378 11572 12384
rect 11426 11792 11482 11801
rect 11426 11727 11482 11736
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 11612 11212 11664 11218
rect 11612 11154 11664 11160
rect 11624 10849 11652 11154
rect 11610 10840 11666 10849
rect 11610 10775 11612 10784
rect 11664 10775 11666 10784
rect 11612 10746 11664 10752
rect 11060 10124 11112 10130
rect 11060 10066 11112 10072
rect 10968 9444 11020 9450
rect 10968 9386 11020 9392
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 10980 7834 11008 9114
rect 11072 8974 11100 10066
rect 11428 9920 11480 9926
rect 11348 9880 11428 9908
rect 11152 9648 11204 9654
rect 11152 9590 11204 9596
rect 11242 9616 11298 9625
rect 11164 9194 11192 9590
rect 11242 9551 11298 9560
rect 11256 9382 11284 9551
rect 11348 9489 11376 9880
rect 11428 9862 11480 9868
rect 11334 9480 11390 9489
rect 11334 9415 11390 9424
rect 11244 9376 11296 9382
rect 11242 9344 11244 9353
rect 11296 9344 11298 9353
rect 11242 9279 11298 9288
rect 11164 9166 11284 9194
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 11150 8936 11206 8945
rect 11072 8294 11100 8910
rect 11150 8871 11206 8880
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 10980 7806 11100 7834
rect 10968 7200 11020 7206
rect 10968 7142 11020 7148
rect 10980 5930 11008 7142
rect 11072 7002 11100 7806
rect 11164 7478 11192 8871
rect 11256 8514 11284 9166
rect 11348 9110 11376 9415
rect 11336 9104 11388 9110
rect 11336 9046 11388 9052
rect 11348 8634 11376 9046
rect 11336 8628 11388 8634
rect 11336 8570 11388 8576
rect 11428 8628 11480 8634
rect 11428 8570 11480 8576
rect 11256 8486 11376 8514
rect 11244 8288 11296 8294
rect 11244 8230 11296 8236
rect 11256 7954 11284 8230
rect 11244 7948 11296 7954
rect 11244 7890 11296 7896
rect 11152 7472 11204 7478
rect 11152 7414 11204 7420
rect 11060 6996 11112 7002
rect 11060 6938 11112 6944
rect 11072 6458 11100 6938
rect 11164 6730 11192 7414
rect 11152 6724 11204 6730
rect 11152 6666 11204 6672
rect 11150 6488 11206 6497
rect 11060 6452 11112 6458
rect 11150 6423 11206 6432
rect 11060 6394 11112 6400
rect 10980 5914 11100 5930
rect 10980 5908 11112 5914
rect 10980 5902 11060 5908
rect 11060 5850 11112 5856
rect 11164 5642 11192 6423
rect 11242 5672 11298 5681
rect 11152 5636 11204 5642
rect 11242 5607 11298 5616
rect 11152 5578 11204 5584
rect 11164 5370 11192 5578
rect 10968 5364 11020 5370
rect 10968 5306 11020 5312
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 10980 4826 11008 5306
rect 11152 5160 11204 5166
rect 11152 5102 11204 5108
rect 10968 4820 11020 4826
rect 10968 4762 11020 4768
rect 10980 4706 11008 4762
rect 10980 4678 11100 4706
rect 11072 4010 11100 4678
rect 11164 4486 11192 5102
rect 11152 4480 11204 4486
rect 11152 4422 11204 4428
rect 11060 4004 11112 4010
rect 11060 3946 11112 3952
rect 10888 3726 11008 3754
rect 10876 3664 10928 3670
rect 10876 3606 10928 3612
rect 10888 2990 10916 3606
rect 10876 2984 10928 2990
rect 10876 2926 10928 2932
rect 10980 2650 11008 3726
rect 11060 3460 11112 3466
rect 11060 3402 11112 3408
rect 11072 2650 11100 3402
rect 11164 3058 11192 4422
rect 11256 4078 11284 5607
rect 11348 5545 11376 8486
rect 11440 8265 11468 8570
rect 11426 8256 11482 8265
rect 11426 8191 11482 8200
rect 11518 6080 11574 6089
rect 11518 6015 11574 6024
rect 11532 5914 11560 6015
rect 11520 5908 11572 5914
rect 11520 5850 11572 5856
rect 11334 5536 11390 5545
rect 11334 5471 11390 5480
rect 11336 5092 11388 5098
rect 11336 5034 11388 5040
rect 11348 4593 11376 5034
rect 11612 5024 11664 5030
rect 11612 4966 11664 4972
rect 11334 4584 11390 4593
rect 11334 4519 11390 4528
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 11244 3732 11296 3738
rect 11244 3674 11296 3680
rect 11152 3052 11204 3058
rect 11152 2994 11204 3000
rect 11150 2952 11206 2961
rect 11150 2887 11206 2896
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 11164 1034 11192 2887
rect 11256 2582 11284 3674
rect 11244 2576 11296 2582
rect 11244 2518 11296 2524
rect 11242 2408 11298 2417
rect 11242 2343 11244 2352
rect 11296 2343 11298 2352
rect 11244 2314 11296 2320
rect 11348 2281 11376 4519
rect 11428 3936 11480 3942
rect 11428 3878 11480 3884
rect 11440 2961 11468 3878
rect 11520 3596 11572 3602
rect 11520 3538 11572 3544
rect 11532 3369 11560 3538
rect 11518 3360 11574 3369
rect 11518 3295 11574 3304
rect 11532 3126 11560 3295
rect 11520 3120 11572 3126
rect 11624 3097 11652 4966
rect 11520 3062 11572 3068
rect 11610 3088 11666 3097
rect 11610 3023 11666 3032
rect 11426 2952 11482 2961
rect 11426 2887 11482 2896
rect 11612 2848 11664 2854
rect 11612 2790 11664 2796
rect 11334 2272 11390 2281
rect 11334 2207 11390 2216
rect 11624 1737 11652 2790
rect 11610 1728 11666 1737
rect 11610 1663 11666 1672
rect 10520 734 10824 762
rect 11072 1006 11192 1034
rect 10520 480 10548 734
rect 11072 480 11100 1006
rect 11716 480 11744 13926
rect 11808 13734 11836 20295
rect 11992 19689 12020 24806
rect 12624 24754 12676 24760
rect 12070 24712 12126 24721
rect 12070 24647 12126 24656
rect 12084 24410 12112 24647
rect 12072 24404 12124 24410
rect 12072 24346 12124 24352
rect 12084 23866 12112 24346
rect 12256 24268 12308 24274
rect 12256 24210 12308 24216
rect 12072 23860 12124 23866
rect 12072 23802 12124 23808
rect 12072 23656 12124 23662
rect 12072 23598 12124 23604
rect 11978 19680 12034 19689
rect 11978 19615 12034 19624
rect 11888 18420 11940 18426
rect 11888 18362 11940 18368
rect 11900 17814 11928 18362
rect 11888 17808 11940 17814
rect 11888 17750 11940 17756
rect 12084 17762 12112 23598
rect 12268 23526 12296 24210
rect 12348 24200 12400 24206
rect 12348 24142 12400 24148
rect 12256 23520 12308 23526
rect 12256 23462 12308 23468
rect 12164 21616 12216 21622
rect 12162 21584 12164 21593
rect 12216 21584 12218 21593
rect 12162 21519 12218 21528
rect 12176 21418 12204 21519
rect 12164 21412 12216 21418
rect 12164 21354 12216 21360
rect 12268 19009 12296 23462
rect 12360 23322 12388 24142
rect 12624 23792 12676 23798
rect 12622 23760 12624 23769
rect 12676 23760 12678 23769
rect 12622 23695 12678 23704
rect 12348 23316 12400 23322
rect 12348 23258 12400 23264
rect 12532 23112 12584 23118
rect 12532 23054 12584 23060
rect 12544 22438 12572 23054
rect 12532 22432 12584 22438
rect 12532 22374 12584 22380
rect 12728 22114 12756 27390
rect 13372 24721 13400 27520
rect 13358 24712 13414 24721
rect 13358 24647 13414 24656
rect 13084 24608 13136 24614
rect 13084 24550 13136 24556
rect 13636 24608 13688 24614
rect 13636 24550 13688 24556
rect 13096 24410 13124 24550
rect 13084 24404 13136 24410
rect 13084 24346 13136 24352
rect 13360 24268 13412 24274
rect 13360 24210 13412 24216
rect 12992 24132 13044 24138
rect 12992 24074 13044 24080
rect 13004 23186 13032 24074
rect 13372 23526 13400 24210
rect 13544 24200 13596 24206
rect 13544 24142 13596 24148
rect 13360 23520 13412 23526
rect 13452 23520 13504 23526
rect 13360 23462 13412 23468
rect 13450 23488 13452 23497
rect 13504 23488 13506 23497
rect 12992 23180 13044 23186
rect 12992 23122 13044 23128
rect 13004 22778 13032 23122
rect 12992 22772 13044 22778
rect 12992 22714 13044 22720
rect 13268 22568 13320 22574
rect 13268 22510 13320 22516
rect 12636 22086 12756 22114
rect 12440 21344 12492 21350
rect 12440 21286 12492 21292
rect 12452 21146 12480 21286
rect 12440 21140 12492 21146
rect 12440 21082 12492 21088
rect 12452 21010 12572 21026
rect 12452 21004 12584 21010
rect 12452 20998 12532 21004
rect 12452 20754 12480 20998
rect 12532 20946 12584 20952
rect 12530 20904 12586 20913
rect 12530 20839 12532 20848
rect 12584 20839 12586 20848
rect 12532 20810 12584 20816
rect 12360 20726 12480 20754
rect 12360 20602 12388 20726
rect 12348 20596 12400 20602
rect 12348 20538 12400 20544
rect 12440 19304 12492 19310
rect 12440 19246 12492 19252
rect 12254 19000 12310 19009
rect 12254 18935 12310 18944
rect 12164 18760 12216 18766
rect 12164 18702 12216 18708
rect 12176 18426 12204 18702
rect 12452 18630 12480 19246
rect 12636 18902 12664 22086
rect 13280 21894 13308 22510
rect 13372 22234 13400 23462
rect 13450 23423 13506 23432
rect 13556 23254 13584 24142
rect 13648 23662 13676 24550
rect 13728 24200 13780 24206
rect 13728 24142 13780 24148
rect 13740 23866 13768 24142
rect 13820 24064 13872 24070
rect 13820 24006 13872 24012
rect 13924 24018 13952 27520
rect 14568 27418 14596 27520
rect 14568 27390 14688 27418
rect 13832 23882 13860 24006
rect 13924 23990 14320 24018
rect 13728 23860 13780 23866
rect 13832 23854 13952 23882
rect 13728 23802 13780 23808
rect 13636 23656 13688 23662
rect 13636 23598 13688 23604
rect 13544 23248 13596 23254
rect 13544 23190 13596 23196
rect 13556 22778 13584 23190
rect 13544 22772 13596 22778
rect 13544 22714 13596 22720
rect 13360 22228 13412 22234
rect 13360 22170 13412 22176
rect 13452 22092 13504 22098
rect 13452 22034 13504 22040
rect 12808 21888 12860 21894
rect 12808 21830 12860 21836
rect 13268 21888 13320 21894
rect 13268 21830 13320 21836
rect 12820 21350 12848 21830
rect 12808 21344 12860 21350
rect 12808 21286 12860 21292
rect 12820 20505 12848 21286
rect 12992 20936 13044 20942
rect 12992 20878 13044 20884
rect 12806 20496 12862 20505
rect 12806 20431 12862 20440
rect 12716 20324 12768 20330
rect 12716 20266 12768 20272
rect 12728 20058 12756 20266
rect 12716 20052 12768 20058
rect 12716 19994 12768 20000
rect 12898 19816 12954 19825
rect 12898 19751 12954 19760
rect 12806 19408 12862 19417
rect 12806 19343 12862 19352
rect 12624 18896 12676 18902
rect 12622 18864 12624 18873
rect 12676 18864 12678 18873
rect 12622 18799 12678 18808
rect 12440 18624 12492 18630
rect 12440 18566 12492 18572
rect 12164 18420 12216 18426
rect 12164 18362 12216 18368
rect 12164 18284 12216 18290
rect 12164 18226 12216 18232
rect 12176 17882 12204 18226
rect 12452 18222 12480 18566
rect 12440 18216 12492 18222
rect 12440 18158 12492 18164
rect 12164 17876 12216 17882
rect 12164 17818 12216 17824
rect 12452 17814 12480 18158
rect 12714 17912 12770 17921
rect 12714 17847 12716 17856
rect 12768 17847 12770 17856
rect 12716 17818 12768 17824
rect 12440 17808 12492 17814
rect 11900 16590 11928 17750
rect 12084 17734 12296 17762
rect 12440 17750 12492 17756
rect 12622 17776 12678 17785
rect 12268 17241 12296 17734
rect 12346 17640 12402 17649
rect 12346 17575 12402 17584
rect 12254 17232 12310 17241
rect 12254 17167 12310 17176
rect 11978 17096 12034 17105
rect 11978 17031 12034 17040
rect 11888 16584 11940 16590
rect 11888 16526 11940 16532
rect 11992 15502 12020 17031
rect 11980 15496 12032 15502
rect 11980 15438 12032 15444
rect 11992 15162 12020 15438
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 11980 15156 12032 15162
rect 11980 15098 12032 15104
rect 11796 13728 11848 13734
rect 11796 13670 11848 13676
rect 11900 13546 11928 15098
rect 12072 14272 12124 14278
rect 12072 14214 12124 14220
rect 11980 13932 12032 13938
rect 11980 13874 12032 13880
rect 11808 13518 11928 13546
rect 11808 8673 11836 13518
rect 11888 12640 11940 12646
rect 11888 12582 11940 12588
rect 11900 12481 11928 12582
rect 11886 12472 11942 12481
rect 11886 12407 11942 12416
rect 11992 12238 12020 13874
rect 12084 13530 12112 14214
rect 12072 13524 12124 13530
rect 12072 13466 12124 13472
rect 12164 13456 12216 13462
rect 12164 13398 12216 13404
rect 12176 12782 12204 13398
rect 12164 12776 12216 12782
rect 12164 12718 12216 12724
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 11980 12232 12032 12238
rect 11980 12174 12032 12180
rect 11992 11898 12020 12174
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 11978 11792 12034 11801
rect 11978 11727 12034 11736
rect 11888 11552 11940 11558
rect 11888 11494 11940 11500
rect 11900 11121 11928 11494
rect 11886 11112 11942 11121
rect 11886 11047 11942 11056
rect 11992 10810 12020 11727
rect 12084 11694 12112 12242
rect 12072 11688 12124 11694
rect 12072 11630 12124 11636
rect 11980 10804 12032 10810
rect 11980 10746 12032 10752
rect 11992 10538 12020 10746
rect 11980 10532 12032 10538
rect 11980 10474 12032 10480
rect 11794 8664 11850 8673
rect 11794 8599 11850 8608
rect 12084 8242 12112 11630
rect 12164 11144 12216 11150
rect 12164 11086 12216 11092
rect 12176 9926 12204 11086
rect 12164 9920 12216 9926
rect 12164 9862 12216 9868
rect 12084 8214 12204 8242
rect 12072 7744 12124 7750
rect 12072 7686 12124 7692
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 11992 7002 12020 7142
rect 11980 6996 12032 7002
rect 11980 6938 12032 6944
rect 12084 6866 12112 7686
rect 12072 6860 12124 6866
rect 12072 6802 12124 6808
rect 12070 6216 12126 6225
rect 12070 6151 12126 6160
rect 11888 5772 11940 5778
rect 11888 5714 11940 5720
rect 11900 5370 11928 5714
rect 12084 5710 12112 6151
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 12072 5704 12124 5710
rect 12072 5646 12124 5652
rect 11888 5364 11940 5370
rect 11888 5306 11940 5312
rect 11900 5001 11928 5306
rect 11992 5098 12020 5646
rect 11980 5092 12032 5098
rect 11980 5034 12032 5040
rect 11886 4992 11942 5001
rect 11886 4927 11942 4936
rect 11980 4548 12032 4554
rect 11980 4490 12032 4496
rect 11888 4004 11940 4010
rect 11888 3946 11940 3952
rect 11796 3528 11848 3534
rect 11796 3470 11848 3476
rect 11808 3194 11836 3470
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 11900 1601 11928 3946
rect 11992 2553 12020 4490
rect 12072 4480 12124 4486
rect 12072 4422 12124 4428
rect 11978 2544 12034 2553
rect 12084 2514 12112 4422
rect 12176 3913 12204 8214
rect 12162 3904 12218 3913
rect 12162 3839 12218 3848
rect 11978 2479 12034 2488
rect 12072 2508 12124 2514
rect 12072 2450 12124 2456
rect 11886 1592 11942 1601
rect 11886 1527 11942 1536
rect 12268 480 12296 17167
rect 12360 14482 12388 17575
rect 12452 17134 12480 17750
rect 12622 17711 12624 17720
rect 12676 17711 12678 17720
rect 12624 17682 12676 17688
rect 12532 17332 12584 17338
rect 12532 17274 12584 17280
rect 12440 17128 12492 17134
rect 12440 17070 12492 17076
rect 12440 16720 12492 16726
rect 12440 16662 12492 16668
rect 12452 15706 12480 16662
rect 12544 16561 12572 17274
rect 12636 16794 12664 17682
rect 12624 16788 12676 16794
rect 12624 16730 12676 16736
rect 12820 16658 12848 19343
rect 12808 16652 12860 16658
rect 12808 16594 12860 16600
rect 12530 16552 12586 16561
rect 12530 16487 12586 16496
rect 12624 16176 12676 16182
rect 12622 16144 12624 16153
rect 12676 16144 12678 16153
rect 12622 16079 12678 16088
rect 12624 15904 12676 15910
rect 12624 15846 12676 15852
rect 12636 15706 12664 15846
rect 12440 15700 12492 15706
rect 12440 15642 12492 15648
rect 12624 15700 12676 15706
rect 12624 15642 12676 15648
rect 12820 15638 12848 16594
rect 12808 15632 12860 15638
rect 12808 15574 12860 15580
rect 12716 15564 12768 15570
rect 12716 15506 12768 15512
rect 12624 15088 12676 15094
rect 12624 15030 12676 15036
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 12348 14476 12400 14482
rect 12348 14418 12400 14424
rect 12452 14278 12480 14894
rect 12532 14544 12584 14550
rect 12532 14486 12584 14492
rect 12440 14272 12492 14278
rect 12440 14214 12492 14220
rect 12452 13870 12480 14214
rect 12440 13864 12492 13870
rect 12440 13806 12492 13812
rect 12452 13462 12480 13806
rect 12440 13456 12492 13462
rect 12440 13398 12492 13404
rect 12440 13184 12492 13190
rect 12440 13126 12492 13132
rect 12452 12918 12480 13126
rect 12440 12912 12492 12918
rect 12440 12854 12492 12860
rect 12348 11620 12400 11626
rect 12348 11562 12400 11568
rect 12360 11150 12388 11562
rect 12544 11286 12572 14486
rect 12532 11280 12584 11286
rect 12532 11222 12584 11228
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12452 10266 12480 10406
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 12440 9920 12492 9926
rect 12360 9880 12440 9908
rect 12360 8090 12388 9880
rect 12440 9862 12492 9868
rect 12532 9512 12584 9518
rect 12532 9454 12584 9460
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12348 8084 12400 8090
rect 12348 8026 12400 8032
rect 12452 7954 12480 8774
rect 12544 8294 12572 9454
rect 12532 8288 12584 8294
rect 12532 8230 12584 8236
rect 12348 7948 12400 7954
rect 12348 7890 12400 7896
rect 12440 7948 12492 7954
rect 12440 7890 12492 7896
rect 12360 7546 12388 7890
rect 12348 7540 12400 7546
rect 12348 7482 12400 7488
rect 12360 7313 12388 7482
rect 12346 7304 12402 7313
rect 12346 7239 12402 7248
rect 12532 6792 12584 6798
rect 12532 6734 12584 6740
rect 12544 6118 12572 6734
rect 12532 6112 12584 6118
rect 12532 6054 12584 6060
rect 12440 5840 12492 5846
rect 12440 5782 12492 5788
rect 12452 5166 12480 5782
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 12348 4684 12400 4690
rect 12348 4626 12400 4632
rect 12360 3466 12388 4626
rect 12452 3602 12480 4966
rect 12544 3738 12572 6054
rect 12532 3732 12584 3738
rect 12532 3674 12584 3680
rect 12440 3596 12492 3602
rect 12440 3538 12492 3544
rect 12348 3460 12400 3466
rect 12348 3402 12400 3408
rect 12440 3392 12492 3398
rect 12440 3334 12492 3340
rect 12452 3210 12480 3334
rect 12360 3182 12480 3210
rect 12360 2922 12388 3182
rect 12544 3074 12572 3674
rect 12636 3210 12664 15030
rect 12728 14822 12756 15506
rect 12716 14816 12768 14822
rect 12716 14758 12768 14764
rect 12728 11354 12756 14758
rect 12912 14498 12940 19751
rect 13004 19514 13032 20878
rect 13174 19952 13230 19961
rect 13174 19887 13230 19896
rect 12992 19508 13044 19514
rect 12992 19450 13044 19456
rect 12990 19272 13046 19281
rect 12990 19207 13046 19216
rect 13004 18873 13032 19207
rect 12990 18864 13046 18873
rect 12990 18799 13046 18808
rect 13188 18329 13216 19887
rect 13174 18320 13230 18329
rect 13174 18255 13230 18264
rect 13176 17672 13228 17678
rect 13176 17614 13228 17620
rect 13188 17134 13216 17614
rect 13176 17128 13228 17134
rect 13176 17070 13228 17076
rect 13084 17060 13136 17066
rect 13084 17002 13136 17008
rect 12990 16688 13046 16697
rect 12990 16623 13046 16632
rect 13004 14618 13032 16623
rect 13096 16454 13124 17002
rect 13176 16584 13228 16590
rect 13176 16526 13228 16532
rect 13084 16448 13136 16454
rect 13084 16390 13136 16396
rect 13096 14958 13124 16390
rect 13188 16250 13216 16526
rect 13176 16244 13228 16250
rect 13176 16186 13228 16192
rect 13176 15700 13228 15706
rect 13176 15642 13228 15648
rect 13188 15094 13216 15642
rect 13280 15337 13308 21830
rect 13464 21350 13492 22034
rect 13648 21554 13676 23598
rect 13924 23594 13952 23854
rect 13912 23588 13964 23594
rect 13912 23530 13964 23536
rect 13726 23488 13782 23497
rect 13726 23423 13782 23432
rect 13740 22642 13768 23423
rect 13924 22681 13952 23530
rect 13910 22672 13966 22681
rect 13728 22636 13780 22642
rect 13910 22607 13912 22616
rect 13728 22578 13780 22584
rect 13964 22607 13966 22616
rect 13912 22578 13964 22584
rect 13924 22522 13952 22578
rect 13740 22494 13952 22522
rect 13740 22234 13768 22494
rect 14188 22432 14240 22438
rect 14188 22374 14240 22380
rect 13728 22228 13780 22234
rect 13728 22170 13780 22176
rect 14002 21856 14058 21865
rect 14002 21791 14058 21800
rect 13636 21548 13688 21554
rect 13636 21490 13688 21496
rect 13912 21548 13964 21554
rect 13912 21490 13964 21496
rect 13452 21344 13504 21350
rect 13452 21286 13504 21292
rect 13360 20800 13412 20806
rect 13360 20742 13412 20748
rect 13372 20398 13400 20742
rect 13360 20392 13412 20398
rect 13360 20334 13412 20340
rect 13358 19408 13414 19417
rect 13358 19343 13414 19352
rect 13266 15328 13322 15337
rect 13266 15263 13322 15272
rect 13176 15088 13228 15094
rect 13176 15030 13228 15036
rect 13372 15042 13400 19343
rect 13464 19145 13492 21286
rect 13544 20052 13596 20058
rect 13544 19994 13596 20000
rect 13556 19378 13584 19994
rect 13544 19372 13596 19378
rect 13544 19314 13596 19320
rect 13648 19310 13676 21490
rect 13820 21344 13872 21350
rect 13820 21286 13872 21292
rect 13832 21010 13860 21286
rect 13924 21146 13952 21490
rect 13912 21140 13964 21146
rect 13912 21082 13964 21088
rect 13820 21004 13872 21010
rect 13820 20946 13872 20952
rect 13832 20602 13860 20946
rect 13820 20596 13872 20602
rect 13820 20538 13872 20544
rect 13820 19916 13872 19922
rect 13820 19858 13872 19864
rect 13636 19304 13688 19310
rect 13542 19272 13598 19281
rect 13636 19246 13688 19252
rect 13728 19304 13780 19310
rect 13728 19246 13780 19252
rect 13542 19207 13598 19216
rect 13556 19174 13584 19207
rect 13544 19168 13596 19174
rect 13450 19136 13506 19145
rect 13544 19110 13596 19116
rect 13636 19168 13688 19174
rect 13636 19110 13688 19116
rect 13450 19071 13506 19080
rect 13556 18630 13584 19110
rect 13648 18970 13676 19110
rect 13636 18964 13688 18970
rect 13636 18906 13688 18912
rect 13544 18624 13596 18630
rect 13544 18566 13596 18572
rect 13450 18320 13506 18329
rect 13450 18255 13506 18264
rect 13464 15706 13492 18255
rect 13740 17610 13768 19246
rect 13832 19174 13860 19858
rect 13912 19236 13964 19242
rect 13912 19178 13964 19184
rect 13820 19168 13872 19174
rect 13924 19145 13952 19178
rect 13820 19110 13872 19116
rect 13910 19136 13966 19145
rect 13910 19071 13966 19080
rect 14016 18986 14044 21791
rect 14094 20632 14150 20641
rect 14094 20567 14150 20576
rect 14108 19990 14136 20567
rect 14096 19984 14148 19990
rect 14096 19926 14148 19932
rect 14016 18958 14136 18986
rect 14004 18828 14056 18834
rect 14004 18770 14056 18776
rect 13912 18624 13964 18630
rect 13912 18566 13964 18572
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 13832 17678 13860 18022
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 13728 17604 13780 17610
rect 13728 17546 13780 17552
rect 13924 17490 13952 18566
rect 14016 18426 14044 18770
rect 14004 18420 14056 18426
rect 14004 18362 14056 18368
rect 14004 17740 14056 17746
rect 14004 17682 14056 17688
rect 13832 17462 13952 17490
rect 13544 16992 13596 16998
rect 13544 16934 13596 16940
rect 13556 16794 13584 16934
rect 13544 16788 13596 16794
rect 13544 16730 13596 16736
rect 13726 16688 13782 16697
rect 13544 16652 13596 16658
rect 13726 16623 13782 16632
rect 13544 16594 13596 16600
rect 13556 15978 13584 16594
rect 13634 16552 13690 16561
rect 13634 16487 13690 16496
rect 13648 16250 13676 16487
rect 13636 16244 13688 16250
rect 13636 16186 13688 16192
rect 13544 15972 13596 15978
rect 13544 15914 13596 15920
rect 13452 15700 13504 15706
rect 13452 15642 13504 15648
rect 13740 15502 13768 16623
rect 13728 15496 13780 15502
rect 13728 15438 13780 15444
rect 13636 15156 13688 15162
rect 13740 15144 13768 15438
rect 13688 15116 13768 15144
rect 13636 15098 13688 15104
rect 13372 15014 13584 15042
rect 13084 14952 13136 14958
rect 13084 14894 13136 14900
rect 13360 14816 13412 14822
rect 13360 14758 13412 14764
rect 12992 14612 13044 14618
rect 12992 14554 13044 14560
rect 12912 14470 13124 14498
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 12820 12986 12848 13330
rect 12898 13288 12954 13297
rect 12898 13223 12954 13232
rect 12808 12980 12860 12986
rect 12808 12922 12860 12928
rect 12912 12481 12940 13223
rect 12898 12472 12954 12481
rect 12898 12407 12900 12416
rect 12952 12407 12954 12416
rect 12900 12378 12952 12384
rect 12716 11348 12768 11354
rect 12716 11290 12768 11296
rect 12728 10985 12756 11290
rect 12714 10976 12770 10985
rect 13096 10962 13124 14470
rect 13176 14340 13228 14346
rect 13176 14282 13228 14288
rect 13188 13841 13216 14282
rect 13174 13832 13230 13841
rect 13174 13767 13230 13776
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 13280 12646 13308 13466
rect 13372 13161 13400 14758
rect 13358 13152 13414 13161
rect 13358 13087 13414 13096
rect 13268 12640 13320 12646
rect 13268 12582 13320 12588
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 13188 11354 13216 12038
rect 13280 11762 13308 12582
rect 13268 11756 13320 11762
rect 13268 11698 13320 11704
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 13188 11082 13216 11290
rect 13176 11076 13228 11082
rect 13176 11018 13228 11024
rect 13096 10934 13216 10962
rect 12714 10911 12770 10920
rect 12728 10674 12756 10911
rect 12716 10668 12768 10674
rect 12716 10610 12768 10616
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12728 3777 12756 10406
rect 13004 10010 13032 10610
rect 13084 10260 13136 10266
rect 13084 10202 13136 10208
rect 12912 9994 13032 10010
rect 12900 9988 13032 9994
rect 12952 9982 13032 9988
rect 12900 9930 12952 9936
rect 12912 9382 12940 9930
rect 12992 9920 13044 9926
rect 12992 9862 13044 9868
rect 12808 9376 12860 9382
rect 12808 9318 12860 9324
rect 12900 9376 12952 9382
rect 12900 9318 12952 9324
rect 12820 8838 12848 9318
rect 12900 8900 12952 8906
rect 12900 8842 12952 8848
rect 12808 8832 12860 8838
rect 12808 8774 12860 8780
rect 12912 8634 12940 8842
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 12808 7404 12860 7410
rect 12808 7346 12860 7352
rect 12820 5710 12848 7346
rect 13004 6866 13032 9862
rect 13096 9178 13124 10202
rect 13084 9172 13136 9178
rect 13084 9114 13136 9120
rect 13188 7732 13216 10934
rect 13280 9518 13308 11698
rect 13372 11286 13400 13087
rect 13556 12442 13584 15014
rect 13832 13954 13860 17462
rect 13912 16992 13964 16998
rect 13912 16934 13964 16940
rect 13924 16114 13952 16934
rect 14016 16658 14044 17682
rect 14004 16652 14056 16658
rect 14004 16594 14056 16600
rect 13912 16108 13964 16114
rect 13912 16050 13964 16056
rect 14108 16046 14136 18958
rect 14096 16040 14148 16046
rect 14096 15982 14148 15988
rect 14108 15706 14136 15982
rect 14096 15700 14148 15706
rect 14096 15642 14148 15648
rect 13912 14952 13964 14958
rect 13912 14894 13964 14900
rect 13924 14074 13952 14894
rect 14200 14618 14228 22374
rect 14292 19825 14320 23990
rect 14370 23896 14426 23905
rect 14370 23831 14426 23840
rect 14278 19816 14334 19825
rect 14278 19751 14334 19760
rect 14280 19236 14332 19242
rect 14280 19178 14332 19184
rect 14292 18766 14320 19178
rect 14384 18970 14412 23831
rect 14464 22772 14516 22778
rect 14464 22714 14516 22720
rect 14372 18964 14424 18970
rect 14372 18906 14424 18912
rect 14372 18828 14424 18834
rect 14372 18770 14424 18776
rect 14280 18760 14332 18766
rect 14280 18702 14332 18708
rect 14292 18358 14320 18702
rect 14280 18352 14332 18358
rect 14280 18294 14332 18300
rect 14384 17542 14412 18770
rect 14372 17536 14424 17542
rect 14372 17478 14424 17484
rect 14280 16992 14332 16998
rect 14280 16934 14332 16940
rect 14292 16454 14320 16934
rect 14384 16658 14412 17478
rect 14372 16652 14424 16658
rect 14372 16594 14424 16600
rect 14280 16448 14332 16454
rect 14280 16390 14332 16396
rect 14188 14612 14240 14618
rect 14188 14554 14240 14560
rect 14200 14074 14228 14554
rect 14292 14498 14320 16390
rect 14372 15360 14424 15366
rect 14372 15302 14424 15308
rect 14384 14958 14412 15302
rect 14372 14952 14424 14958
rect 14372 14894 14424 14900
rect 14476 14521 14504 22714
rect 14556 20936 14608 20942
rect 14556 20878 14608 20884
rect 14568 20602 14596 20878
rect 14556 20596 14608 20602
rect 14556 20538 14608 20544
rect 14568 20398 14596 20538
rect 14556 20392 14608 20398
rect 14556 20334 14608 20340
rect 14660 19281 14688 27390
rect 15120 25242 15148 27520
rect 15672 25514 15700 27520
rect 14752 25214 15148 25242
rect 15580 25486 15700 25514
rect 14752 23322 14780 25214
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 15384 24676 15436 24682
rect 15384 24618 15436 24624
rect 15292 24268 15344 24274
rect 15292 24210 15344 24216
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 15200 23520 15252 23526
rect 14844 23468 15200 23474
rect 15304 23508 15332 24210
rect 15396 23730 15424 24618
rect 15384 23724 15436 23730
rect 15384 23666 15436 23672
rect 15252 23480 15332 23508
rect 15580 23497 15608 25486
rect 15660 25356 15712 25362
rect 15660 25298 15712 25304
rect 15672 24614 15700 25298
rect 16120 24744 16172 24750
rect 16120 24686 16172 24692
rect 15660 24608 15712 24614
rect 15660 24550 15712 24556
rect 15566 23488 15622 23497
rect 14844 23462 15252 23468
rect 14844 23446 15240 23462
rect 14740 23316 14792 23322
rect 14740 23258 14792 23264
rect 14752 22778 14780 23258
rect 14740 22772 14792 22778
rect 14740 22714 14792 22720
rect 14844 22098 14872 23446
rect 15566 23423 15622 23432
rect 15568 23180 15620 23186
rect 15568 23122 15620 23128
rect 15292 22976 15344 22982
rect 15292 22918 15344 22924
rect 15476 22976 15528 22982
rect 15476 22918 15528 22924
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 14832 22092 14884 22098
rect 14832 22034 14884 22040
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 14830 21448 14886 21457
rect 14830 21383 14886 21392
rect 14738 20904 14794 20913
rect 14738 20839 14794 20848
rect 14646 19272 14702 19281
rect 14646 19207 14702 19216
rect 14752 19122 14780 20839
rect 14568 19094 14780 19122
rect 14568 14550 14596 19094
rect 14738 19000 14794 19009
rect 14648 18964 14700 18970
rect 14738 18935 14794 18944
rect 14648 18906 14700 18912
rect 14660 16726 14688 18906
rect 14752 18358 14780 18935
rect 14740 18352 14792 18358
rect 14740 18294 14792 18300
rect 14844 17746 14872 21383
rect 15304 21146 15332 22918
rect 15488 22642 15516 22918
rect 15476 22636 15528 22642
rect 15476 22578 15528 22584
rect 15488 22234 15516 22578
rect 15580 22438 15608 23122
rect 15568 22432 15620 22438
rect 15568 22374 15620 22380
rect 15476 22228 15528 22234
rect 15476 22170 15528 22176
rect 15382 21992 15438 22001
rect 15382 21927 15438 21936
rect 15292 21140 15344 21146
rect 15292 21082 15344 21088
rect 15292 21004 15344 21010
rect 15292 20946 15344 20952
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 15304 20534 15332 20946
rect 15396 20874 15424 21927
rect 15488 21418 15516 22170
rect 15476 21412 15528 21418
rect 15476 21354 15528 21360
rect 15384 20868 15436 20874
rect 15384 20810 15436 20816
rect 15292 20528 15344 20534
rect 15292 20470 15344 20476
rect 15304 20058 15332 20470
rect 15384 20256 15436 20262
rect 15384 20198 15436 20204
rect 15292 20052 15344 20058
rect 15292 19994 15344 20000
rect 15292 19916 15344 19922
rect 15292 19858 15344 19864
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15304 19378 15332 19858
rect 15292 19372 15344 19378
rect 15292 19314 15344 19320
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 15108 18148 15160 18154
rect 15108 18090 15160 18096
rect 15120 17882 15148 18090
rect 15108 17876 15160 17882
rect 15108 17818 15160 17824
rect 14832 17740 14884 17746
rect 14832 17682 14884 17688
rect 14832 17604 14884 17610
rect 14832 17546 14884 17552
rect 14740 17060 14792 17066
rect 14740 17002 14792 17008
rect 14648 16720 14700 16726
rect 14648 16662 14700 16668
rect 14556 14544 14608 14550
rect 14462 14512 14518 14521
rect 14292 14470 14412 14498
rect 14280 14408 14332 14414
rect 14278 14376 14280 14385
rect 14332 14376 14334 14385
rect 14278 14311 14334 14320
rect 14384 14226 14412 14470
rect 14556 14486 14608 14492
rect 14462 14447 14518 14456
rect 14556 14408 14608 14414
rect 14556 14350 14608 14356
rect 14292 14198 14412 14226
rect 13912 14068 13964 14074
rect 13912 14010 13964 14016
rect 14188 14068 14240 14074
rect 14188 14010 14240 14016
rect 13832 13926 13952 13954
rect 13728 13864 13780 13870
rect 13780 13812 13860 13818
rect 13728 13806 13860 13812
rect 13740 13790 13860 13806
rect 13634 13016 13690 13025
rect 13832 12986 13860 13790
rect 13634 12951 13636 12960
rect 13688 12951 13690 12960
rect 13820 12980 13872 12986
rect 13636 12922 13688 12928
rect 13820 12922 13872 12928
rect 13818 12880 13874 12889
rect 13818 12815 13874 12824
rect 13544 12436 13596 12442
rect 13544 12378 13596 12384
rect 13544 11620 13596 11626
rect 13544 11562 13596 11568
rect 13360 11280 13412 11286
rect 13360 11222 13412 11228
rect 13450 10840 13506 10849
rect 13450 10775 13506 10784
rect 13360 10124 13412 10130
rect 13360 10066 13412 10072
rect 13268 9512 13320 9518
rect 13268 9454 13320 9460
rect 13372 9450 13400 10066
rect 13360 9444 13412 9450
rect 13360 9386 13412 9392
rect 13372 9178 13400 9386
rect 13360 9172 13412 9178
rect 13360 9114 13412 9120
rect 13268 9036 13320 9042
rect 13268 8978 13320 8984
rect 13280 8634 13308 8978
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 13360 8492 13412 8498
rect 13360 8434 13412 8440
rect 13372 7886 13400 8434
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 13268 7744 13320 7750
rect 13188 7704 13268 7732
rect 13188 7546 13216 7704
rect 13268 7686 13320 7692
rect 13176 7540 13228 7546
rect 13176 7482 13228 7488
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 12992 6860 13044 6866
rect 12992 6802 13044 6808
rect 12898 6352 12954 6361
rect 12898 6287 12954 6296
rect 12808 5704 12860 5710
rect 12808 5646 12860 5652
rect 12714 3768 12770 3777
rect 12714 3703 12770 3712
rect 12820 3618 12848 5646
rect 12912 5234 12940 6287
rect 13004 6254 13032 6802
rect 13188 6322 13216 7142
rect 13268 6860 13320 6866
rect 13268 6802 13320 6808
rect 13176 6316 13228 6322
rect 13176 6258 13228 6264
rect 12992 6248 13044 6254
rect 12992 6190 13044 6196
rect 13084 6112 13136 6118
rect 13084 6054 13136 6060
rect 12992 5908 13044 5914
rect 12992 5850 13044 5856
rect 12900 5228 12952 5234
rect 12900 5170 12952 5176
rect 12912 4826 12940 5170
rect 12900 4820 12952 4826
rect 12900 4762 12952 4768
rect 12728 3590 12848 3618
rect 12728 3534 12756 3590
rect 12716 3528 12768 3534
rect 12714 3496 12716 3505
rect 12768 3496 12770 3505
rect 12714 3431 12770 3440
rect 12900 3460 12952 3466
rect 12728 3398 12756 3431
rect 12900 3402 12952 3408
rect 12716 3392 12768 3398
rect 12716 3334 12768 3340
rect 12636 3182 12848 3210
rect 12452 3046 12572 3074
rect 12348 2916 12400 2922
rect 12348 2858 12400 2864
rect 12360 2378 12388 2858
rect 12452 2854 12480 3046
rect 12440 2848 12492 2854
rect 12438 2816 12440 2825
rect 12492 2816 12494 2825
rect 12438 2751 12494 2760
rect 12348 2372 12400 2378
rect 12348 2314 12400 2320
rect 12820 480 12848 3182
rect 12912 2009 12940 3402
rect 13004 3233 13032 5850
rect 12990 3224 13046 3233
rect 12990 3159 13046 3168
rect 13004 2553 13032 3159
rect 13096 2689 13124 6054
rect 13280 5914 13308 6802
rect 13464 5914 13492 10775
rect 13556 10674 13584 11562
rect 13636 11552 13688 11558
rect 13832 11506 13860 12815
rect 13924 11558 13952 13926
rect 14188 13796 14240 13802
rect 14188 13738 14240 13744
rect 14004 13728 14056 13734
rect 14004 13670 14056 13676
rect 14016 12442 14044 13670
rect 14004 12436 14056 12442
rect 14004 12378 14056 12384
rect 14004 12300 14056 12306
rect 14004 12242 14056 12248
rect 13636 11494 13688 11500
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 13648 10146 13676 11494
rect 13740 11478 13860 11506
rect 13912 11552 13964 11558
rect 13912 11494 13964 11500
rect 13740 11234 13768 11478
rect 14016 11354 14044 12242
rect 14004 11348 14056 11354
rect 14004 11290 14056 11296
rect 13740 11206 13952 11234
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13740 10266 13768 11086
rect 13924 10742 13952 11206
rect 14004 11212 14056 11218
rect 14004 11154 14056 11160
rect 14016 10810 14044 11154
rect 14004 10804 14056 10810
rect 14004 10746 14056 10752
rect 13912 10736 13964 10742
rect 13912 10678 13964 10684
rect 13924 10538 13952 10678
rect 14096 10600 14148 10606
rect 14096 10542 14148 10548
rect 13912 10532 13964 10538
rect 13912 10474 13964 10480
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 13648 10118 13860 10146
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 13740 9382 13768 9998
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13556 8673 13584 8910
rect 13740 8838 13768 9318
rect 13728 8832 13780 8838
rect 13728 8774 13780 8780
rect 13542 8664 13598 8673
rect 13542 8599 13544 8608
rect 13596 8599 13598 8608
rect 13544 8570 13596 8576
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 13556 8294 13584 8366
rect 13740 8294 13768 8774
rect 13544 8288 13596 8294
rect 13544 8230 13596 8236
rect 13728 8288 13780 8294
rect 13728 8230 13780 8236
rect 13556 7290 13584 8230
rect 13636 7812 13688 7818
rect 13636 7754 13688 7760
rect 13648 7410 13676 7754
rect 13636 7404 13688 7410
rect 13636 7346 13688 7352
rect 13740 7342 13768 8230
rect 13832 8022 13860 10118
rect 13820 8016 13872 8022
rect 13820 7958 13872 7964
rect 13832 7546 13860 7958
rect 13820 7540 13872 7546
rect 13820 7482 13872 7488
rect 13728 7336 13780 7342
rect 13556 7262 13676 7290
rect 13728 7278 13780 7284
rect 13544 7200 13596 7206
rect 13544 7142 13596 7148
rect 13556 7002 13584 7142
rect 13544 6996 13596 7002
rect 13544 6938 13596 6944
rect 13648 6882 13676 7262
rect 13556 6854 13676 6882
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 13452 5908 13504 5914
rect 13452 5850 13504 5856
rect 13268 5636 13320 5642
rect 13268 5578 13320 5584
rect 13280 5234 13308 5578
rect 13464 5370 13492 5850
rect 13452 5364 13504 5370
rect 13452 5306 13504 5312
rect 13268 5228 13320 5234
rect 13268 5170 13320 5176
rect 13280 4622 13308 5170
rect 13452 4684 13504 4690
rect 13452 4626 13504 4632
rect 13268 4616 13320 4622
rect 13268 4558 13320 4564
rect 13176 4480 13228 4486
rect 13176 4422 13228 4428
rect 13188 3738 13216 4422
rect 13280 4010 13308 4558
rect 13464 4282 13492 4626
rect 13452 4276 13504 4282
rect 13452 4218 13504 4224
rect 13452 4072 13504 4078
rect 13556 4060 13584 6854
rect 13636 6792 13688 6798
rect 13636 6734 13688 6740
rect 13648 6458 13676 6734
rect 13636 6452 13688 6458
rect 13636 6394 13688 6400
rect 13728 6316 13780 6322
rect 13728 6258 13780 6264
rect 13740 5914 13768 6258
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 13728 5772 13780 5778
rect 13924 5760 13952 10474
rect 14108 10266 14136 10542
rect 14096 10260 14148 10266
rect 14096 10202 14148 10208
rect 14094 9752 14150 9761
rect 14094 9687 14150 9696
rect 14108 8634 14136 9687
rect 14096 8628 14148 8634
rect 14096 8570 14148 8576
rect 14108 8129 14136 8570
rect 14094 8120 14150 8129
rect 14094 8055 14150 8064
rect 14096 7268 14148 7274
rect 14096 7210 14148 7216
rect 14108 6458 14136 7210
rect 14096 6452 14148 6458
rect 14096 6394 14148 6400
rect 13780 5732 13952 5760
rect 13728 5714 13780 5720
rect 13728 5636 13780 5642
rect 13728 5578 13780 5584
rect 13636 5568 13688 5574
rect 13636 5510 13688 5516
rect 13648 4826 13676 5510
rect 13740 5386 13768 5578
rect 13740 5358 13860 5386
rect 13924 5370 13952 5732
rect 13832 5302 13860 5358
rect 13912 5364 13964 5370
rect 13912 5306 13964 5312
rect 13820 5296 13872 5302
rect 13820 5238 13872 5244
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 14096 4480 14148 4486
rect 14096 4422 14148 4428
rect 13504 4032 13584 4060
rect 13912 4072 13964 4078
rect 13452 4014 13504 4020
rect 13912 4014 13964 4020
rect 13268 4004 13320 4010
rect 13268 3946 13320 3952
rect 13176 3732 13228 3738
rect 13176 3674 13228 3680
rect 13280 3398 13308 3946
rect 13358 3904 13414 3913
rect 13358 3839 13414 3848
rect 13268 3392 13320 3398
rect 13268 3334 13320 3340
rect 13176 2916 13228 2922
rect 13176 2858 13228 2864
rect 13082 2680 13138 2689
rect 13188 2650 13216 2858
rect 13280 2854 13308 3334
rect 13268 2848 13320 2854
rect 13268 2790 13320 2796
rect 13082 2615 13138 2624
rect 13176 2644 13228 2650
rect 13176 2586 13228 2592
rect 12990 2544 13046 2553
rect 12990 2479 13046 2488
rect 12898 2000 12954 2009
rect 12898 1935 12954 1944
rect 13372 480 13400 3839
rect 13464 2990 13492 4014
rect 13636 3936 13688 3942
rect 13636 3878 13688 3884
rect 13728 3936 13780 3942
rect 13728 3878 13780 3884
rect 13648 3777 13676 3878
rect 13634 3768 13690 3777
rect 13634 3703 13690 3712
rect 13634 3632 13690 3641
rect 13634 3567 13636 3576
rect 13688 3567 13690 3576
rect 13636 3538 13688 3544
rect 13740 3466 13768 3878
rect 13820 3732 13872 3738
rect 13820 3674 13872 3680
rect 13728 3460 13780 3466
rect 13728 3402 13780 3408
rect 13740 2990 13768 3402
rect 13452 2984 13504 2990
rect 13452 2926 13504 2932
rect 13728 2984 13780 2990
rect 13728 2926 13780 2932
rect 13544 2508 13596 2514
rect 13544 2450 13596 2456
rect 13556 2417 13584 2450
rect 13740 2446 13768 2926
rect 13832 2650 13860 3674
rect 13820 2644 13872 2650
rect 13820 2586 13872 2592
rect 13728 2440 13780 2446
rect 13542 2408 13598 2417
rect 13728 2382 13780 2388
rect 13542 2343 13598 2352
rect 13924 480 13952 4014
rect 14108 4010 14136 4422
rect 14200 4060 14228 13738
rect 14292 13530 14320 14198
rect 14372 14068 14424 14074
rect 14372 14010 14424 14016
rect 14280 13524 14332 13530
rect 14280 13466 14332 13472
rect 14292 12345 14320 13466
rect 14384 12424 14412 14010
rect 14384 12396 14504 12424
rect 14278 12336 14334 12345
rect 14278 12271 14334 12280
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 14372 12232 14424 12238
rect 14372 12174 14424 12180
rect 14292 11898 14320 12174
rect 14280 11892 14332 11898
rect 14280 11834 14332 11840
rect 14384 11286 14412 12174
rect 14372 11280 14424 11286
rect 14372 11222 14424 11228
rect 14370 11112 14426 11121
rect 14370 11047 14426 11056
rect 14278 10976 14334 10985
rect 14278 10911 14334 10920
rect 14292 9586 14320 10911
rect 14280 9580 14332 9586
rect 14280 9522 14332 9528
rect 14278 9480 14334 9489
rect 14278 9415 14280 9424
rect 14332 9415 14334 9424
rect 14280 9386 14332 9392
rect 14292 8974 14320 9386
rect 14280 8968 14332 8974
rect 14280 8910 14332 8916
rect 14292 8090 14320 8910
rect 14280 8084 14332 8090
rect 14280 8026 14332 8032
rect 14292 7886 14320 8026
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14292 7002 14320 7822
rect 14280 6996 14332 7002
rect 14280 6938 14332 6944
rect 14384 4078 14412 11047
rect 14476 5658 14504 12396
rect 14568 10674 14596 14350
rect 14660 12866 14688 16662
rect 14752 16454 14780 17002
rect 14844 16946 14872 17546
rect 15292 17536 15344 17542
rect 15292 17478 15344 17484
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15016 17128 15068 17134
rect 15014 17096 15016 17105
rect 15068 17096 15070 17105
rect 15014 17031 15070 17040
rect 14844 16918 14964 16946
rect 14832 16788 14884 16794
rect 14832 16730 14884 16736
rect 14740 16448 14792 16454
rect 14740 16390 14792 16396
rect 14752 15910 14780 16390
rect 14740 15904 14792 15910
rect 14740 15846 14792 15852
rect 14752 15162 14780 15846
rect 14844 15706 14872 16730
rect 14936 16726 14964 16918
rect 15304 16833 15332 17478
rect 15290 16824 15346 16833
rect 15290 16759 15346 16768
rect 14924 16720 14976 16726
rect 14922 16688 14924 16697
rect 15292 16720 15344 16726
rect 14976 16688 14978 16697
rect 15292 16662 15344 16668
rect 14922 16623 14978 16632
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15304 15910 15332 16662
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 14832 15700 14884 15706
rect 14832 15642 14884 15648
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14740 15156 14792 15162
rect 14740 15098 14792 15104
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15304 13190 15332 15846
rect 15396 14822 15424 20198
rect 15476 19304 15528 19310
rect 15476 19246 15528 19252
rect 15488 19174 15516 19246
rect 15476 19168 15528 19174
rect 15672 19145 15700 24550
rect 16132 23186 16160 24686
rect 16224 24410 16252 27520
rect 16776 24834 16804 27520
rect 16500 24806 16804 24834
rect 16500 24682 16528 24806
rect 16488 24676 16540 24682
rect 16488 24618 16540 24624
rect 16396 24608 16448 24614
rect 16396 24550 16448 24556
rect 16408 24426 16436 24550
rect 16212 24404 16264 24410
rect 16408 24398 16528 24426
rect 16212 24346 16264 24352
rect 16394 24304 16450 24313
rect 16394 24239 16396 24248
rect 16448 24239 16450 24248
rect 16396 24210 16448 24216
rect 16408 23866 16436 24210
rect 16500 24041 16528 24398
rect 16486 24032 16542 24041
rect 16486 23967 16542 23976
rect 16396 23860 16448 23866
rect 16396 23802 16448 23808
rect 17132 23520 17184 23526
rect 17132 23462 17184 23468
rect 17144 23254 17172 23462
rect 17132 23248 17184 23254
rect 17132 23190 17184 23196
rect 16120 23180 16172 23186
rect 16120 23122 16172 23128
rect 16764 23180 16816 23186
rect 16764 23122 16816 23128
rect 15936 23112 15988 23118
rect 15936 23054 15988 23060
rect 15752 22500 15804 22506
rect 15752 22442 15804 22448
rect 15764 21894 15792 22442
rect 15948 22098 15976 23054
rect 16776 22506 16804 23122
rect 16856 22704 16908 22710
rect 16854 22672 16856 22681
rect 16908 22672 16910 22681
rect 16854 22607 16910 22616
rect 16120 22500 16172 22506
rect 16120 22442 16172 22448
rect 16764 22500 16816 22506
rect 16764 22442 16816 22448
rect 15936 22092 15988 22098
rect 15936 22034 15988 22040
rect 15752 21888 15804 21894
rect 15752 21830 15804 21836
rect 15764 21298 15792 21830
rect 15948 21350 15976 22034
rect 15936 21344 15988 21350
rect 15764 21270 15884 21298
rect 15936 21286 15988 21292
rect 15856 20942 15884 21270
rect 15844 20936 15896 20942
rect 15844 20878 15896 20884
rect 15856 20602 15884 20878
rect 15844 20596 15896 20602
rect 15844 20538 15896 20544
rect 15948 20466 15976 21286
rect 16028 21140 16080 21146
rect 16028 21082 16080 21088
rect 15936 20460 15988 20466
rect 15936 20402 15988 20408
rect 16040 20058 16068 21082
rect 16028 20052 16080 20058
rect 16028 19994 16080 20000
rect 15476 19110 15528 19116
rect 15658 19136 15714 19145
rect 15488 18630 15516 19110
rect 15658 19071 15714 19080
rect 15672 18952 15700 19071
rect 15672 18924 16068 18952
rect 15936 18828 15988 18834
rect 15936 18770 15988 18776
rect 15476 18624 15528 18630
rect 15476 18566 15528 18572
rect 15948 18290 15976 18770
rect 15936 18284 15988 18290
rect 15936 18226 15988 18232
rect 15474 18184 15530 18193
rect 15474 18119 15530 18128
rect 15384 14816 15436 14822
rect 15384 14758 15436 14764
rect 15384 14272 15436 14278
rect 15384 14214 15436 14220
rect 15396 13297 15424 14214
rect 15488 13938 15516 18119
rect 15948 18086 15976 18226
rect 15936 18080 15988 18086
rect 15936 18022 15988 18028
rect 15658 17912 15714 17921
rect 15658 17847 15714 17856
rect 15672 17814 15700 17847
rect 15660 17808 15712 17814
rect 15660 17750 15712 17756
rect 15672 17490 15700 17750
rect 15752 17672 15804 17678
rect 15752 17614 15804 17620
rect 15580 17462 15700 17490
rect 15580 17134 15608 17462
rect 15658 17368 15714 17377
rect 15764 17338 15792 17614
rect 15658 17303 15714 17312
rect 15752 17332 15804 17338
rect 15568 17128 15620 17134
rect 15568 17070 15620 17076
rect 15568 16992 15620 16998
rect 15568 16934 15620 16940
rect 15580 16590 15608 16934
rect 15568 16584 15620 16590
rect 15568 16526 15620 16532
rect 15580 15706 15608 16526
rect 15568 15700 15620 15706
rect 15568 15642 15620 15648
rect 15672 14550 15700 17303
rect 15752 17274 15804 17280
rect 15764 16776 15792 17274
rect 15948 16998 15976 18022
rect 15936 16992 15988 16998
rect 15936 16934 15988 16940
rect 15844 16788 15896 16794
rect 15764 16748 15844 16776
rect 15844 16730 15896 16736
rect 15844 15972 15896 15978
rect 15844 15914 15896 15920
rect 15856 15706 15884 15914
rect 15844 15700 15896 15706
rect 15844 15642 15896 15648
rect 15660 14544 15712 14550
rect 15660 14486 15712 14492
rect 15672 14006 15700 14486
rect 15752 14476 15804 14482
rect 15752 14418 15804 14424
rect 15764 14074 15792 14418
rect 15936 14408 15988 14414
rect 15936 14350 15988 14356
rect 15752 14068 15804 14074
rect 15752 14010 15804 14016
rect 15660 14000 15712 14006
rect 15660 13942 15712 13948
rect 15948 13938 15976 14350
rect 15476 13932 15528 13938
rect 15476 13874 15528 13880
rect 15936 13932 15988 13938
rect 15936 13874 15988 13880
rect 15488 13530 15516 13874
rect 16040 13802 16068 18924
rect 16132 15162 16160 22442
rect 16396 21344 16448 21350
rect 16396 21286 16448 21292
rect 16210 19816 16266 19825
rect 16210 19751 16266 19760
rect 16120 15156 16172 15162
rect 16120 15098 16172 15104
rect 16028 13796 16080 13802
rect 16028 13738 16080 13744
rect 15476 13524 15528 13530
rect 15476 13466 15528 13472
rect 15382 13288 15438 13297
rect 15382 13223 15438 13232
rect 15292 13184 15344 13190
rect 15292 13126 15344 13132
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 14660 12838 14964 12866
rect 14648 12708 14700 12714
rect 14648 12650 14700 12656
rect 14660 12442 14688 12650
rect 14648 12436 14700 12442
rect 14648 12378 14700 12384
rect 14660 12102 14688 12378
rect 14936 12322 14964 12838
rect 15016 12640 15068 12646
rect 15016 12582 15068 12588
rect 15200 12640 15252 12646
rect 15200 12582 15252 12588
rect 15028 12442 15056 12582
rect 15016 12436 15068 12442
rect 15016 12378 15068 12384
rect 15212 12356 15240 12582
rect 15212 12328 15332 12356
rect 14936 12294 15056 12322
rect 14740 12232 14792 12238
rect 15028 12209 15056 12294
rect 14740 12174 14792 12180
rect 15014 12200 15070 12209
rect 14648 12096 14700 12102
rect 14648 12038 14700 12044
rect 14660 11898 14688 12038
rect 14648 11892 14700 11898
rect 14648 11834 14700 11840
rect 14648 11008 14700 11014
rect 14648 10950 14700 10956
rect 14660 10810 14688 10950
rect 14648 10804 14700 10810
rect 14648 10746 14700 10752
rect 14556 10668 14608 10674
rect 14556 10610 14608 10616
rect 14752 10606 14780 12174
rect 15014 12135 15070 12144
rect 14832 12096 14884 12102
rect 14832 12038 14884 12044
rect 14844 11898 14872 12038
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 14832 11892 14884 11898
rect 14832 11834 14884 11840
rect 15304 11830 15332 12328
rect 15292 11824 15344 11830
rect 14830 11792 14886 11801
rect 15292 11766 15344 11772
rect 14830 11727 14886 11736
rect 14740 10600 14792 10606
rect 14740 10542 14792 10548
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14752 9897 14780 10406
rect 14738 9888 14794 9897
rect 14738 9823 14794 9832
rect 14556 9580 14608 9586
rect 14556 9522 14608 9528
rect 14568 5778 14596 9522
rect 14738 8800 14794 8809
rect 14738 8735 14794 8744
rect 14752 8401 14780 8735
rect 14738 8392 14794 8401
rect 14738 8327 14794 8336
rect 14648 8288 14700 8294
rect 14648 8230 14700 8236
rect 14660 7342 14688 8230
rect 14740 7948 14792 7954
rect 14740 7890 14792 7896
rect 14752 7721 14780 7890
rect 14738 7712 14794 7721
rect 14738 7647 14794 7656
rect 14648 7336 14700 7342
rect 14648 7278 14700 7284
rect 14844 6882 14872 11727
rect 15488 11268 15516 13466
rect 15568 13388 15620 13394
rect 15568 13330 15620 13336
rect 15580 12646 15608 13330
rect 15660 13184 15712 13190
rect 15660 13126 15712 13132
rect 15568 12640 15620 12646
rect 15568 12582 15620 12588
rect 15568 11280 15620 11286
rect 15488 11240 15568 11268
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15304 10470 15332 11086
rect 15488 10538 15516 11240
rect 15568 11222 15620 11228
rect 15568 11076 15620 11082
rect 15568 11018 15620 11024
rect 15476 10532 15528 10538
rect 15476 10474 15528 10480
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15304 9110 15332 10202
rect 15476 9920 15528 9926
rect 15476 9862 15528 9868
rect 15382 9752 15438 9761
rect 15382 9687 15384 9696
rect 15436 9687 15438 9696
rect 15384 9658 15436 9664
rect 15488 9382 15516 9862
rect 15580 9654 15608 11018
rect 15568 9648 15620 9654
rect 15568 9590 15620 9596
rect 15476 9376 15528 9382
rect 15476 9318 15528 9324
rect 15292 9104 15344 9110
rect 15292 9046 15344 9052
rect 15384 8832 15436 8838
rect 15384 8774 15436 8780
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15106 8120 15162 8129
rect 15106 8055 15108 8064
rect 15160 8055 15162 8064
rect 15108 8026 15160 8032
rect 15396 7886 15424 8774
rect 15384 7880 15436 7886
rect 15384 7822 15436 7828
rect 15292 7744 15344 7750
rect 15396 7721 15424 7822
rect 15292 7686 15344 7692
rect 15382 7712 15438 7721
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14752 6854 14872 6882
rect 14752 6390 14780 6854
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 14740 6384 14792 6390
rect 14740 6326 14792 6332
rect 14844 6322 14872 6598
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 14832 6316 14884 6322
rect 14832 6258 14884 6264
rect 14844 6225 14872 6258
rect 14830 6216 14886 6225
rect 15304 6202 15332 7686
rect 15382 7647 15438 7656
rect 15384 7200 15436 7206
rect 15384 7142 15436 7148
rect 15396 6322 15424 7142
rect 15384 6316 15436 6322
rect 15384 6258 15436 6264
rect 15304 6174 15424 6202
rect 14830 6151 14886 6160
rect 15292 6112 15344 6118
rect 15292 6054 15344 6060
rect 15304 5778 15332 6054
rect 15396 5914 15424 6174
rect 15384 5908 15436 5914
rect 15384 5850 15436 5856
rect 14556 5772 14608 5778
rect 14556 5714 14608 5720
rect 15292 5772 15344 5778
rect 15292 5714 15344 5720
rect 14476 5630 14780 5658
rect 14648 5568 14700 5574
rect 14648 5510 14700 5516
rect 14554 5128 14610 5137
rect 14554 5063 14556 5072
rect 14608 5063 14610 5072
rect 14556 5034 14608 5040
rect 14464 4752 14516 4758
rect 14462 4720 14464 4729
rect 14516 4720 14518 4729
rect 14462 4655 14518 4664
rect 14372 4072 14424 4078
rect 14200 4032 14320 4060
rect 14096 4004 14148 4010
rect 14096 3946 14148 3952
rect 14292 2666 14320 4032
rect 14372 4014 14424 4020
rect 14556 3392 14608 3398
rect 14556 3334 14608 3340
rect 14568 2990 14596 3334
rect 14556 2984 14608 2990
rect 14556 2926 14608 2932
rect 14292 2638 14596 2666
rect 14568 480 14596 2638
rect 14660 2378 14688 5510
rect 14648 2372 14700 2378
rect 14648 2314 14700 2320
rect 14752 1306 14780 5630
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 15396 5370 15424 5850
rect 15384 5364 15436 5370
rect 15384 5306 15436 5312
rect 15488 5302 15516 9318
rect 15568 8832 15620 8838
rect 15568 8774 15620 8780
rect 15580 5710 15608 8774
rect 15568 5704 15620 5710
rect 15568 5646 15620 5652
rect 15476 5296 15528 5302
rect 15476 5238 15528 5244
rect 15384 5092 15436 5098
rect 15384 5034 15436 5040
rect 14924 5024 14976 5030
rect 14924 4966 14976 4972
rect 14936 4758 14964 4966
rect 14924 4752 14976 4758
rect 14924 4694 14976 4700
rect 15292 4548 15344 4554
rect 15292 4490 15344 4496
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 15200 3936 15252 3942
rect 15200 3878 15252 3884
rect 15212 3670 15240 3878
rect 15200 3664 15252 3670
rect 15200 3606 15252 3612
rect 15304 3602 15332 4490
rect 15396 4457 15424 5034
rect 15382 4448 15438 4457
rect 15382 4383 15438 4392
rect 15292 3596 15344 3602
rect 15292 3538 15344 3544
rect 14832 3392 14884 3398
rect 14832 3334 14884 3340
rect 15476 3392 15528 3398
rect 15476 3334 15528 3340
rect 14844 2922 14872 3334
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 15488 3058 15516 3334
rect 15476 3052 15528 3058
rect 15476 2994 15528 3000
rect 14832 2916 14884 2922
rect 14832 2858 14884 2864
rect 15108 2848 15160 2854
rect 15108 2790 15160 2796
rect 15120 2632 15148 2790
rect 15200 2644 15252 2650
rect 15120 2604 15200 2632
rect 15200 2586 15252 2592
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 14752 1278 15148 1306
rect 15120 480 15148 1278
rect 15672 480 15700 13126
rect 15752 12776 15804 12782
rect 15752 12718 15804 12724
rect 15764 12442 15792 12718
rect 16118 12608 16174 12617
rect 16118 12543 16174 12552
rect 15752 12436 15804 12442
rect 15752 12378 15804 12384
rect 15752 12300 15804 12306
rect 15752 12242 15804 12248
rect 15764 11354 15792 12242
rect 16132 11898 16160 12543
rect 16120 11892 16172 11898
rect 16120 11834 16172 11840
rect 15934 11656 15990 11665
rect 15934 11591 15936 11600
rect 15988 11591 15990 11600
rect 15936 11562 15988 11568
rect 15752 11348 15804 11354
rect 15752 11290 15804 11296
rect 15764 10266 15792 11290
rect 15844 11008 15896 11014
rect 15844 10950 15896 10956
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 15856 10130 15884 10950
rect 15844 10124 15896 10130
rect 15844 10066 15896 10072
rect 15936 10056 15988 10062
rect 15936 9998 15988 10004
rect 15948 9722 15976 9998
rect 15936 9716 15988 9722
rect 15936 9658 15988 9664
rect 16224 9568 16252 19751
rect 16408 18630 16436 21286
rect 16670 20496 16726 20505
rect 16670 20431 16672 20440
rect 16724 20431 16726 20440
rect 16672 20402 16724 20408
rect 17420 20058 17448 27520
rect 17500 24268 17552 24274
rect 17500 24210 17552 24216
rect 17512 23526 17540 24210
rect 17972 24154 18000 27520
rect 18144 24744 18196 24750
rect 18144 24686 18196 24692
rect 17880 24138 18000 24154
rect 17868 24132 18000 24138
rect 17920 24126 18000 24132
rect 18050 24168 18106 24177
rect 18050 24103 18106 24112
rect 17868 24074 17920 24080
rect 18064 23662 18092 24103
rect 18052 23656 18104 23662
rect 18052 23598 18104 23604
rect 17500 23520 17552 23526
rect 17500 23462 17552 23468
rect 17408 20052 17460 20058
rect 17408 19994 17460 20000
rect 16580 19916 16632 19922
rect 16580 19858 16632 19864
rect 16592 19514 16620 19858
rect 16580 19508 16632 19514
rect 16580 19450 16632 19456
rect 16672 19236 16724 19242
rect 16672 19178 16724 19184
rect 16684 18970 16712 19178
rect 16764 19168 16816 19174
rect 16764 19110 16816 19116
rect 16672 18964 16724 18970
rect 16672 18906 16724 18912
rect 16776 18737 16804 19110
rect 18052 18896 18104 18902
rect 18156 18873 18184 24686
rect 18236 24608 18288 24614
rect 18236 24550 18288 24556
rect 18248 24313 18276 24550
rect 18524 24410 18552 27520
rect 18786 24712 18842 24721
rect 18786 24647 18842 24656
rect 18800 24410 18828 24647
rect 18512 24404 18564 24410
rect 18512 24346 18564 24352
rect 18788 24404 18840 24410
rect 18788 24346 18840 24352
rect 18234 24304 18290 24313
rect 18234 24239 18290 24248
rect 18512 24268 18564 24274
rect 18512 24210 18564 24216
rect 18420 23656 18472 23662
rect 18420 23598 18472 23604
rect 18236 23180 18288 23186
rect 18236 23122 18288 23128
rect 18248 22438 18276 23122
rect 18236 22432 18288 22438
rect 18236 22374 18288 22380
rect 18248 19417 18276 22374
rect 18234 19408 18290 19417
rect 18234 19343 18290 19352
rect 18052 18838 18104 18844
rect 18142 18864 18198 18873
rect 18064 18748 18092 18838
rect 18198 18822 18276 18850
rect 18142 18799 18198 18808
rect 16762 18728 16818 18737
rect 16762 18663 16818 18672
rect 17130 18728 17186 18737
rect 18064 18720 18184 18748
rect 17130 18663 17186 18672
rect 16396 18624 16448 18630
rect 16396 18566 16448 18572
rect 16408 18086 16436 18566
rect 16396 18080 16448 18086
rect 16396 18022 16448 18028
rect 16408 17542 16436 18022
rect 16764 17672 16816 17678
rect 16764 17614 16816 17620
rect 16396 17536 16448 17542
rect 16396 17478 16448 17484
rect 16672 17536 16724 17542
rect 16672 17478 16724 17484
rect 16408 17105 16436 17478
rect 16394 17096 16450 17105
rect 16394 17031 16450 17040
rect 16408 16046 16436 17031
rect 16684 16998 16712 17478
rect 16776 17134 16804 17614
rect 16856 17536 16908 17542
rect 16856 17478 16908 17484
rect 16764 17128 16816 17134
rect 16764 17070 16816 17076
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 16488 16448 16540 16454
rect 16488 16390 16540 16396
rect 16396 16040 16448 16046
rect 16396 15982 16448 15988
rect 16304 15632 16356 15638
rect 16304 15574 16356 15580
rect 16316 15094 16344 15574
rect 16500 15434 16528 16390
rect 16776 16250 16804 17070
rect 16764 16244 16816 16250
rect 16764 16186 16816 16192
rect 16868 15745 16896 17478
rect 17144 16794 17172 18663
rect 17408 17740 17460 17746
rect 17408 17682 17460 17688
rect 17420 17377 17448 17682
rect 17500 17672 17552 17678
rect 17500 17614 17552 17620
rect 17406 17368 17462 17377
rect 17512 17338 17540 17614
rect 17406 17303 17408 17312
rect 17460 17303 17462 17312
rect 17500 17332 17552 17338
rect 17408 17274 17460 17280
rect 17500 17274 17552 17280
rect 17684 17128 17736 17134
rect 17684 17070 17736 17076
rect 17696 16794 17724 17070
rect 17868 16992 17920 16998
rect 17868 16934 17920 16940
rect 17132 16788 17184 16794
rect 17132 16730 17184 16736
rect 17684 16788 17736 16794
rect 17684 16730 17736 16736
rect 16948 16448 17000 16454
rect 16948 16390 17000 16396
rect 16854 15736 16910 15745
rect 16854 15671 16910 15680
rect 16960 15638 16988 16390
rect 17144 16250 17172 16730
rect 17316 16584 17368 16590
rect 17314 16552 17316 16561
rect 17500 16584 17552 16590
rect 17368 16552 17370 16561
rect 17500 16526 17552 16532
rect 17880 16538 17908 16934
rect 17314 16487 17370 16496
rect 17132 16244 17184 16250
rect 17132 16186 17184 16192
rect 17328 15638 17356 16487
rect 17512 15978 17540 16526
rect 17880 16510 18000 16538
rect 17500 15972 17552 15978
rect 17500 15914 17552 15920
rect 17972 15910 18000 16510
rect 17868 15904 17920 15910
rect 17868 15846 17920 15852
rect 17960 15904 18012 15910
rect 17960 15846 18012 15852
rect 16948 15632 17000 15638
rect 16948 15574 17000 15580
rect 17316 15632 17368 15638
rect 17316 15574 17368 15580
rect 17224 15496 17276 15502
rect 17224 15438 17276 15444
rect 16488 15428 16540 15434
rect 16488 15370 16540 15376
rect 16500 15314 16528 15370
rect 16500 15286 16620 15314
rect 16304 15088 16356 15094
rect 16304 15030 16356 15036
rect 16592 15026 16620 15286
rect 16580 15020 16632 15026
rect 16580 14962 16632 14968
rect 16764 14816 16816 14822
rect 16764 14758 16816 14764
rect 16670 14376 16726 14385
rect 16670 14311 16726 14320
rect 16488 14272 16540 14278
rect 16488 14214 16540 14220
rect 16500 13462 16528 14214
rect 16684 13530 16712 14311
rect 16776 14074 16804 14758
rect 17236 14482 17264 15438
rect 17880 15366 17908 15846
rect 17960 15632 18012 15638
rect 17960 15574 18012 15580
rect 17868 15360 17920 15366
rect 17868 15302 17920 15308
rect 17500 15156 17552 15162
rect 17500 15098 17552 15104
rect 17512 14793 17540 15098
rect 17592 15088 17644 15094
rect 17592 15030 17644 15036
rect 17498 14784 17554 14793
rect 17498 14719 17554 14728
rect 17224 14476 17276 14482
rect 17224 14418 17276 14424
rect 16764 14068 16816 14074
rect 16764 14010 16816 14016
rect 16762 13968 16818 13977
rect 16762 13903 16764 13912
rect 16816 13903 16818 13912
rect 16764 13874 16816 13880
rect 17236 13870 17264 14418
rect 17224 13864 17276 13870
rect 17224 13806 17276 13812
rect 17224 13728 17276 13734
rect 17224 13670 17276 13676
rect 16672 13524 16724 13530
rect 16672 13466 16724 13472
rect 16488 13456 16540 13462
rect 16488 13398 16540 13404
rect 16500 12322 16528 13398
rect 17236 13190 17264 13670
rect 17500 13388 17552 13394
rect 17500 13330 17552 13336
rect 17224 13184 17276 13190
rect 17224 13126 17276 13132
rect 17236 12782 17264 13126
rect 17512 12986 17540 13330
rect 17500 12980 17552 12986
rect 17500 12922 17552 12928
rect 17224 12776 17276 12782
rect 16762 12744 16818 12753
rect 17224 12718 17276 12724
rect 16762 12679 16764 12688
rect 16816 12679 16818 12688
rect 16764 12650 16816 12656
rect 16500 12306 16620 12322
rect 16500 12300 16632 12306
rect 16500 12294 16580 12300
rect 16580 12242 16632 12248
rect 16304 12096 16356 12102
rect 16304 12038 16356 12044
rect 16316 11558 16344 12038
rect 16396 11620 16448 11626
rect 16396 11562 16448 11568
rect 16304 11552 16356 11558
rect 16304 11494 16356 11500
rect 16316 11150 16344 11494
rect 16408 11354 16436 11562
rect 16396 11348 16448 11354
rect 16396 11290 16448 11296
rect 16672 11348 16724 11354
rect 16672 11290 16724 11296
rect 16304 11144 16356 11150
rect 16304 11086 16356 11092
rect 16408 10810 16436 11290
rect 16396 10804 16448 10810
rect 16396 10746 16448 10752
rect 16684 10606 16712 11290
rect 16776 10674 16804 12650
rect 16856 12640 16908 12646
rect 16856 12582 16908 12588
rect 16868 12306 16896 12582
rect 16856 12300 16908 12306
rect 16856 12242 16908 12248
rect 16868 11762 16896 12242
rect 16856 11756 16908 11762
rect 16856 11698 16908 11704
rect 17408 11280 17460 11286
rect 17408 11222 17460 11228
rect 17132 11212 17184 11218
rect 17132 11154 17184 11160
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 16948 10668 17000 10674
rect 16948 10610 17000 10616
rect 16672 10600 16724 10606
rect 16672 10542 16724 10548
rect 16304 10464 16356 10470
rect 16304 10406 16356 10412
rect 15856 9540 16252 9568
rect 15752 7948 15804 7954
rect 15752 7890 15804 7896
rect 15764 7002 15792 7890
rect 15752 6996 15804 7002
rect 15752 6938 15804 6944
rect 15856 5930 15884 9540
rect 16316 9518 16344 10406
rect 16960 10130 16988 10610
rect 17144 10198 17172 11154
rect 17420 11082 17448 11222
rect 17604 11121 17632 15030
rect 17880 12646 17908 15302
rect 17972 15162 18000 15574
rect 18052 15564 18104 15570
rect 18052 15506 18104 15512
rect 17960 15156 18012 15162
rect 17960 15098 18012 15104
rect 18064 15094 18092 15506
rect 18052 15088 18104 15094
rect 18052 15030 18104 15036
rect 17960 14068 18012 14074
rect 17960 14010 18012 14016
rect 17972 12986 18000 14010
rect 17960 12980 18012 12986
rect 17960 12922 18012 12928
rect 17868 12640 17920 12646
rect 17868 12582 17920 12588
rect 18156 12594 18184 18720
rect 18248 15570 18276 18822
rect 18432 17921 18460 23598
rect 18524 23594 18552 24210
rect 19076 23866 19104 27520
rect 19628 25786 19656 27520
rect 19536 25758 19656 25786
rect 19536 23866 19564 25758
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 20272 24721 20300 27520
rect 20258 24712 20314 24721
rect 20258 24647 20314 24656
rect 20442 24712 20498 24721
rect 20442 24647 20498 24656
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 20456 24041 20484 24647
rect 20824 24426 20852 27520
rect 20640 24398 20852 24426
rect 20442 24032 20498 24041
rect 20442 23967 20498 23976
rect 19064 23860 19116 23866
rect 19064 23802 19116 23808
rect 19524 23860 19576 23866
rect 19524 23802 19576 23808
rect 18512 23588 18564 23594
rect 18512 23530 18564 23536
rect 18418 17912 18474 17921
rect 18418 17847 18474 17856
rect 18236 15564 18288 15570
rect 18236 15506 18288 15512
rect 18328 14884 18380 14890
rect 18328 14826 18380 14832
rect 18340 14618 18368 14826
rect 18328 14612 18380 14618
rect 18328 14554 18380 14560
rect 18236 13320 18288 13326
rect 18236 13262 18288 13268
rect 18328 13320 18380 13326
rect 18328 13262 18380 13268
rect 18248 12714 18276 13262
rect 18236 12708 18288 12714
rect 18236 12650 18288 12656
rect 18340 12646 18368 13262
rect 18432 12866 18460 17847
rect 18524 15706 18552 23530
rect 20076 23520 20128 23526
rect 20076 23462 20128 23468
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19432 23180 19484 23186
rect 19432 23122 19484 23128
rect 19444 22778 19472 23122
rect 19432 22772 19484 22778
rect 19432 22714 19484 22720
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 20088 18193 20116 23462
rect 20166 23352 20222 23361
rect 20640 23322 20668 24398
rect 20812 24268 20864 24274
rect 20812 24210 20864 24216
rect 20824 23526 20852 24210
rect 21376 23866 21404 27520
rect 21928 23866 21956 27520
rect 22008 24268 22060 24274
rect 22008 24210 22060 24216
rect 21364 23860 21416 23866
rect 21364 23802 21416 23808
rect 21916 23860 21968 23866
rect 21916 23802 21968 23808
rect 21364 23656 21416 23662
rect 21364 23598 21416 23604
rect 20812 23520 20864 23526
rect 20812 23462 20864 23468
rect 21180 23520 21232 23526
rect 21180 23462 21232 23468
rect 20166 23287 20222 23296
rect 20628 23316 20680 23322
rect 20180 22137 20208 23287
rect 20628 23258 20680 23264
rect 20166 22128 20222 22137
rect 20166 22063 20222 22072
rect 20824 20369 20852 23462
rect 21192 23254 21220 23462
rect 21180 23248 21232 23254
rect 20902 23216 20958 23225
rect 21180 23190 21232 23196
rect 20902 23151 20904 23160
rect 20956 23151 20958 23160
rect 20904 23122 20956 23128
rect 20916 22778 20944 23122
rect 20904 22772 20956 22778
rect 20904 22714 20956 22720
rect 21376 20913 21404 23598
rect 22020 23526 22048 24210
rect 22480 24138 22508 27520
rect 23124 24410 23152 27520
rect 23294 24440 23350 24449
rect 23112 24404 23164 24410
rect 23294 24375 23296 24384
rect 23112 24346 23164 24352
rect 23348 24375 23350 24384
rect 23296 24346 23348 24352
rect 23296 24268 23348 24274
rect 23296 24210 23348 24216
rect 22468 24132 22520 24138
rect 22468 24074 22520 24080
rect 22376 23656 22428 23662
rect 22376 23598 22428 23604
rect 22008 23520 22060 23526
rect 22008 23462 22060 23468
rect 22388 21457 22416 23598
rect 23308 23526 23336 24210
rect 23676 23866 23704 27520
rect 23664 23860 23716 23866
rect 23664 23802 23716 23808
rect 24228 23769 24256 27520
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24780 24449 24808 27520
rect 24766 24440 24822 24449
rect 24766 24375 24822 24384
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 25332 23866 25360 27520
rect 25976 24313 26004 27520
rect 26528 25158 26556 27520
rect 26516 25152 26568 25158
rect 26516 25094 26568 25100
rect 27080 24721 27108 27520
rect 27066 24712 27122 24721
rect 27066 24647 27122 24656
rect 25962 24304 26018 24313
rect 25962 24239 26018 24248
rect 25320 23860 25372 23866
rect 25320 23802 25372 23808
rect 24214 23760 24270 23769
rect 24214 23695 24270 23704
rect 23480 23656 23532 23662
rect 23480 23598 23532 23604
rect 23296 23520 23348 23526
rect 23296 23462 23348 23468
rect 22468 23180 22520 23186
rect 22468 23122 22520 23128
rect 22480 22574 22508 23122
rect 22468 22568 22520 22574
rect 22466 22536 22468 22545
rect 22520 22536 22522 22545
rect 22466 22471 22522 22480
rect 22374 21448 22430 21457
rect 22374 21383 22430 21392
rect 21362 20904 21418 20913
rect 21362 20839 21418 20848
rect 20810 20360 20866 20369
rect 20810 20295 20866 20304
rect 23308 19961 23336 23462
rect 23492 23338 23520 23598
rect 23400 23310 23520 23338
rect 23400 23254 23428 23310
rect 23388 23248 23440 23254
rect 23388 23190 23440 23196
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 23294 19952 23350 19961
rect 23294 19887 23350 19896
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 27632 18737 27660 27520
rect 27618 18728 27674 18737
rect 27618 18663 27674 18672
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 20074 18184 20130 18193
rect 20074 18119 20130 18128
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 18696 15904 18748 15910
rect 18696 15846 18748 15852
rect 18512 15700 18564 15706
rect 18512 15642 18564 15648
rect 18708 14958 18736 15846
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 20626 15464 20682 15473
rect 20626 15399 20682 15408
rect 18696 14952 18748 14958
rect 18696 14894 18748 14900
rect 18708 14278 18736 14894
rect 19432 14816 19484 14822
rect 19432 14758 19484 14764
rect 18696 14272 18748 14278
rect 18696 14214 18748 14220
rect 18708 13870 18736 14214
rect 19444 13977 19472 14758
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19430 13968 19486 13977
rect 19430 13903 19486 13912
rect 18696 13864 18748 13870
rect 18694 13832 18696 13841
rect 18748 13832 18750 13841
rect 18512 13796 18564 13802
rect 18694 13767 18750 13776
rect 18512 13738 18564 13744
rect 18524 13682 18552 13738
rect 18524 13654 18644 13682
rect 18432 12838 18552 12866
rect 18616 12850 18644 13654
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 18788 13184 18840 13190
rect 18788 13126 18840 13132
rect 18328 12640 18380 12646
rect 18156 12566 18276 12594
rect 18420 12640 18472 12646
rect 18328 12582 18380 12588
rect 18418 12608 18420 12617
rect 18472 12608 18474 12617
rect 17960 11620 18012 11626
rect 17960 11562 18012 11568
rect 17684 11212 17736 11218
rect 17684 11154 17736 11160
rect 17590 11112 17646 11121
rect 17408 11076 17460 11082
rect 17590 11047 17646 11056
rect 17408 11018 17460 11024
rect 17132 10192 17184 10198
rect 17420 10169 17448 11018
rect 17696 10810 17724 11154
rect 17972 11132 18000 11562
rect 18052 11552 18104 11558
rect 18052 11494 18104 11500
rect 18064 11354 18092 11494
rect 18052 11348 18104 11354
rect 18052 11290 18104 11296
rect 18052 11144 18104 11150
rect 17972 11112 18052 11132
rect 18104 11112 18106 11121
rect 17972 11104 18050 11112
rect 18050 11047 18106 11056
rect 17684 10804 17736 10810
rect 17684 10746 17736 10752
rect 18142 10704 18198 10713
rect 18142 10639 18198 10648
rect 18052 10600 18104 10606
rect 18052 10542 18104 10548
rect 17960 10464 18012 10470
rect 17880 10412 17960 10418
rect 17880 10406 18012 10412
rect 17880 10390 18000 10406
rect 17132 10134 17184 10140
rect 17406 10160 17462 10169
rect 16948 10124 17000 10130
rect 16948 10066 17000 10072
rect 16580 9920 16632 9926
rect 16580 9862 16632 9868
rect 16592 9586 16620 9862
rect 17040 9648 17092 9654
rect 17040 9590 17092 9596
rect 16580 9580 16632 9586
rect 16580 9522 16632 9528
rect 16304 9512 16356 9518
rect 16304 9454 16356 9460
rect 16028 9376 16080 9382
rect 16028 9318 16080 9324
rect 16040 8634 16068 9318
rect 16316 9178 16344 9454
rect 16304 9172 16356 9178
rect 16304 9114 16356 9120
rect 16592 8838 16620 9522
rect 17052 9518 17080 9590
rect 17040 9512 17092 9518
rect 17040 9454 17092 9460
rect 16854 9208 16910 9217
rect 16854 9143 16910 9152
rect 16868 9110 16896 9143
rect 17052 9110 17080 9454
rect 16856 9104 16908 9110
rect 16856 9046 16908 9052
rect 17040 9104 17092 9110
rect 17040 9046 17092 9052
rect 16580 8832 16632 8838
rect 16580 8774 16632 8780
rect 16868 8634 16896 9046
rect 16028 8628 16080 8634
rect 16028 8570 16080 8576
rect 16856 8628 16908 8634
rect 16856 8570 16908 8576
rect 16040 8430 16068 8570
rect 16028 8424 16080 8430
rect 16028 8366 16080 8372
rect 16672 8356 16724 8362
rect 16672 8298 16724 8304
rect 16212 8288 16264 8294
rect 16212 8230 16264 8236
rect 16028 7744 16080 7750
rect 16028 7686 16080 7692
rect 15936 6724 15988 6730
rect 15936 6666 15988 6672
rect 15764 5902 15884 5930
rect 15948 5914 15976 6666
rect 15936 5908 15988 5914
rect 15764 4672 15792 5902
rect 15936 5850 15988 5856
rect 15844 5772 15896 5778
rect 15844 5714 15896 5720
rect 15856 5250 15884 5714
rect 15948 5409 15976 5850
rect 16040 5574 16068 7686
rect 16118 7168 16174 7177
rect 16118 7103 16174 7112
rect 16132 6866 16160 7103
rect 16224 6905 16252 8230
rect 16396 7812 16448 7818
rect 16396 7754 16448 7760
rect 16210 6896 16266 6905
rect 16120 6860 16172 6866
rect 16266 6854 16344 6882
rect 16210 6831 16266 6840
rect 16120 6802 16172 6808
rect 16132 6662 16160 6802
rect 16212 6792 16264 6798
rect 16212 6734 16264 6740
rect 16120 6656 16172 6662
rect 16120 6598 16172 6604
rect 16224 6458 16252 6734
rect 16212 6452 16264 6458
rect 16212 6394 16264 6400
rect 16212 6248 16264 6254
rect 16212 6190 16264 6196
rect 16120 5704 16172 5710
rect 16120 5646 16172 5652
rect 16028 5568 16080 5574
rect 16028 5510 16080 5516
rect 15934 5400 15990 5409
rect 16132 5370 16160 5646
rect 15934 5335 15990 5344
rect 16120 5364 16172 5370
rect 16120 5306 16172 5312
rect 16224 5250 16252 6190
rect 15856 5222 16068 5250
rect 15764 4644 15976 4672
rect 15750 4584 15806 4593
rect 15750 4519 15806 4528
rect 15764 4078 15792 4519
rect 15844 4480 15896 4486
rect 15844 4422 15896 4428
rect 15856 4214 15884 4422
rect 15844 4208 15896 4214
rect 15844 4150 15896 4156
rect 15948 4146 15976 4644
rect 15936 4140 15988 4146
rect 15936 4082 15988 4088
rect 15752 4072 15804 4078
rect 15752 4014 15804 4020
rect 15750 3904 15806 3913
rect 15750 3839 15806 3848
rect 15764 1873 15792 3839
rect 15936 3664 15988 3670
rect 15936 3606 15988 3612
rect 15948 3194 15976 3606
rect 15936 3188 15988 3194
rect 15936 3130 15988 3136
rect 15842 2544 15898 2553
rect 15842 2479 15844 2488
rect 15896 2479 15898 2488
rect 15844 2450 15896 2456
rect 16040 2145 16068 5222
rect 16132 5222 16252 5250
rect 16132 2582 16160 5222
rect 16316 5166 16344 6854
rect 16304 5160 16356 5166
rect 16304 5102 16356 5108
rect 16408 5030 16436 7754
rect 16684 7750 16712 8298
rect 17052 8022 17080 9046
rect 17040 8016 17092 8022
rect 17040 7958 17092 7964
rect 16764 7948 16816 7954
rect 16764 7890 16816 7896
rect 16672 7744 16724 7750
rect 16672 7686 16724 7692
rect 16672 7540 16724 7546
rect 16672 7482 16724 7488
rect 16580 7268 16632 7274
rect 16580 7210 16632 7216
rect 16592 6746 16620 7210
rect 16500 6730 16620 6746
rect 16488 6724 16620 6730
rect 16540 6718 16620 6724
rect 16488 6666 16540 6672
rect 16684 6497 16712 7482
rect 16776 7206 16804 7890
rect 17052 7342 17080 7958
rect 17040 7336 17092 7342
rect 17040 7278 17092 7284
rect 17052 7206 17080 7278
rect 16764 7200 16816 7206
rect 16764 7142 16816 7148
rect 17040 7200 17092 7206
rect 17040 7142 17092 7148
rect 16948 6860 17000 6866
rect 16948 6802 17000 6808
rect 16856 6792 16908 6798
rect 16856 6734 16908 6740
rect 16670 6488 16726 6497
rect 16670 6423 16726 6432
rect 16868 6322 16896 6734
rect 16960 6458 16988 6802
rect 17052 6730 17080 7142
rect 17040 6724 17092 6730
rect 17040 6666 17092 6672
rect 16948 6452 17000 6458
rect 16948 6394 17000 6400
rect 16580 6316 16632 6322
rect 16580 6258 16632 6264
rect 16856 6316 16908 6322
rect 16856 6258 16908 6264
rect 16592 5914 16620 6258
rect 17052 6254 17080 6666
rect 17040 6248 17092 6254
rect 17040 6190 17092 6196
rect 16856 6180 16908 6186
rect 16856 6122 16908 6128
rect 16764 6112 16816 6118
rect 16762 6080 16764 6089
rect 16816 6080 16818 6089
rect 16762 6015 16818 6024
rect 16868 5914 16896 6122
rect 16580 5908 16632 5914
rect 16580 5850 16632 5856
rect 16856 5908 16908 5914
rect 16856 5850 16908 5856
rect 17052 5710 17080 6190
rect 16580 5704 16632 5710
rect 16580 5646 16632 5652
rect 17040 5704 17092 5710
rect 17040 5646 17092 5652
rect 16396 5024 16448 5030
rect 16396 4966 16448 4972
rect 16394 4856 16450 4865
rect 16394 4791 16450 4800
rect 16304 4752 16356 4758
rect 16304 4694 16356 4700
rect 16212 4684 16264 4690
rect 16212 4626 16264 4632
rect 16224 4486 16252 4626
rect 16316 4593 16344 4694
rect 16302 4584 16358 4593
rect 16302 4519 16358 4528
rect 16212 4480 16264 4486
rect 16212 4422 16264 4428
rect 16224 3398 16252 4422
rect 16408 4282 16436 4791
rect 16592 4486 16620 5646
rect 16762 5536 16818 5545
rect 16762 5471 16818 5480
rect 16776 5234 16804 5471
rect 16764 5228 16816 5234
rect 16764 5170 16816 5176
rect 16856 5024 16908 5030
rect 16856 4966 16908 4972
rect 16580 4480 16632 4486
rect 16580 4422 16632 4428
rect 16396 4276 16448 4282
rect 16396 4218 16448 4224
rect 16764 4004 16816 4010
rect 16764 3946 16816 3952
rect 16776 3777 16804 3946
rect 16762 3768 16818 3777
rect 16762 3703 16818 3712
rect 16316 3534 16344 3565
rect 16304 3528 16356 3534
rect 16302 3496 16304 3505
rect 16356 3496 16358 3505
rect 16302 3431 16358 3440
rect 16580 3460 16632 3466
rect 16212 3392 16264 3398
rect 16212 3334 16264 3340
rect 16316 3194 16344 3431
rect 16580 3402 16632 3408
rect 16304 3188 16356 3194
rect 16304 3130 16356 3136
rect 16210 3088 16266 3097
rect 16210 3023 16266 3032
rect 16120 2576 16172 2582
rect 16120 2518 16172 2524
rect 16026 2136 16082 2145
rect 16026 2071 16082 2080
rect 15750 1864 15806 1873
rect 15750 1799 15806 1808
rect 16224 480 16252 3023
rect 16592 2938 16620 3402
rect 16762 3360 16818 3369
rect 16762 3295 16818 3304
rect 16776 3058 16804 3295
rect 16764 3052 16816 3058
rect 16764 2994 16816 3000
rect 16500 2910 16620 2938
rect 16500 2378 16528 2910
rect 16580 2848 16632 2854
rect 16580 2790 16632 2796
rect 16592 2650 16620 2790
rect 16868 2666 16896 4966
rect 17144 4146 17172 10134
rect 17406 10095 17462 10104
rect 17880 9654 17908 10390
rect 17972 10266 18000 10390
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 18064 10198 18092 10542
rect 18052 10192 18104 10198
rect 18052 10134 18104 10140
rect 18156 9994 18184 10639
rect 18144 9988 18196 9994
rect 18144 9930 18196 9936
rect 17868 9648 17920 9654
rect 17868 9590 17920 9596
rect 17958 9480 18014 9489
rect 17958 9415 18014 9424
rect 17224 9376 17276 9382
rect 17224 9318 17276 9324
rect 17236 9178 17264 9318
rect 17972 9178 18000 9415
rect 17224 9172 17276 9178
rect 17224 9114 17276 9120
rect 17960 9172 18012 9178
rect 17960 9114 18012 9120
rect 17236 8809 17264 9114
rect 17222 8800 17278 8809
rect 17222 8735 17278 8744
rect 17682 8664 17738 8673
rect 17682 8599 17738 8608
rect 17406 8120 17462 8129
rect 17406 8055 17462 8064
rect 17420 7342 17448 8055
rect 17408 7336 17460 7342
rect 17408 7278 17460 7284
rect 17314 6896 17370 6905
rect 17314 6831 17370 6840
rect 17328 6798 17356 6831
rect 17316 6792 17368 6798
rect 17316 6734 17368 6740
rect 17224 5840 17276 5846
rect 17224 5782 17276 5788
rect 17236 5030 17264 5782
rect 17224 5024 17276 5030
rect 17224 4966 17276 4972
rect 17236 4826 17264 4966
rect 17224 4820 17276 4826
rect 17224 4762 17276 4768
rect 17236 4214 17264 4762
rect 17224 4208 17276 4214
rect 17696 4185 17724 8599
rect 17960 8560 18012 8566
rect 17960 8502 18012 8508
rect 17972 8265 18000 8502
rect 18052 8288 18104 8294
rect 17958 8256 18014 8265
rect 18052 8230 18104 8236
rect 17958 8191 18014 8200
rect 18064 7290 18092 8230
rect 18144 7744 18196 7750
rect 18144 7686 18196 7692
rect 17972 7262 18092 7290
rect 17972 7041 18000 7262
rect 18052 7200 18104 7206
rect 18052 7142 18104 7148
rect 17958 7032 18014 7041
rect 17958 6967 18014 6976
rect 17958 6624 18014 6633
rect 17958 6559 18014 6568
rect 17224 4150 17276 4156
rect 17682 4176 17738 4185
rect 17132 4140 17184 4146
rect 17682 4111 17738 4120
rect 17868 4140 17920 4146
rect 17132 4082 17184 4088
rect 17868 4082 17920 4088
rect 17880 3913 17908 4082
rect 17972 3942 18000 6559
rect 18064 5681 18092 7142
rect 18156 6866 18184 7686
rect 18144 6860 18196 6866
rect 18144 6802 18196 6808
rect 18156 6458 18184 6802
rect 18144 6452 18196 6458
rect 18144 6394 18196 6400
rect 18050 5672 18106 5681
rect 18050 5607 18106 5616
rect 18050 5400 18106 5409
rect 18050 5335 18052 5344
rect 18104 5335 18106 5344
rect 18052 5306 18104 5312
rect 18142 4448 18198 4457
rect 18142 4383 18198 4392
rect 17960 3936 18012 3942
rect 17866 3904 17922 3913
rect 17960 3878 18012 3884
rect 17866 3839 17922 3848
rect 17406 3496 17462 3505
rect 17406 3431 17462 3440
rect 16580 2644 16632 2650
rect 16580 2586 16632 2592
rect 16776 2638 16896 2666
rect 16488 2372 16540 2378
rect 16488 2314 16540 2320
rect 16776 480 16804 2638
rect 17040 2440 17092 2446
rect 17038 2408 17040 2417
rect 17092 2408 17094 2417
rect 17038 2343 17094 2352
rect 17314 2408 17370 2417
rect 17314 2343 17316 2352
rect 17368 2343 17370 2352
rect 17316 2314 17368 2320
rect 17420 480 17448 3431
rect 17592 3392 17644 3398
rect 17592 3334 17644 3340
rect 17604 3097 17632 3334
rect 17590 3088 17646 3097
rect 17590 3023 17646 3032
rect 17958 2952 18014 2961
rect 17868 2916 17920 2922
rect 17958 2887 18014 2896
rect 17868 2858 17920 2864
rect 17880 2825 17908 2858
rect 17866 2816 17922 2825
rect 17866 2751 17922 2760
rect 17972 480 18000 2887
rect 18052 2848 18104 2854
rect 18052 2790 18104 2796
rect 18064 2582 18092 2790
rect 18156 2650 18184 4383
rect 18248 3992 18276 12566
rect 18418 12543 18474 12552
rect 18524 12458 18552 12838
rect 18604 12844 18656 12850
rect 18604 12786 18656 12792
rect 18340 12430 18552 12458
rect 18616 12442 18644 12786
rect 18800 12782 18828 13126
rect 18788 12776 18840 12782
rect 18788 12718 18840 12724
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 18604 12436 18656 12442
rect 18340 5658 18368 12430
rect 18604 12378 18656 12384
rect 18512 12368 18564 12374
rect 18512 12310 18564 12316
rect 18524 11898 18552 12310
rect 18512 11892 18564 11898
rect 18512 11834 18564 11840
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 18604 11144 18656 11150
rect 18604 11086 18656 11092
rect 18512 11008 18564 11014
rect 18512 10950 18564 10956
rect 18418 10568 18474 10577
rect 18418 10503 18420 10512
rect 18472 10503 18474 10512
rect 18420 10474 18472 10480
rect 18524 10198 18552 10950
rect 18616 10674 18644 11086
rect 18604 10668 18656 10674
rect 18604 10610 18656 10616
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 18512 10192 18564 10198
rect 18512 10134 18564 10140
rect 19340 10192 19392 10198
rect 19340 10134 19392 10140
rect 18972 10056 19024 10062
rect 18970 10024 18972 10033
rect 19024 10024 19026 10033
rect 18970 9959 19026 9968
rect 18878 9344 18934 9353
rect 18878 9279 18934 9288
rect 18604 8900 18656 8906
rect 18604 8842 18656 8848
rect 18616 8498 18644 8842
rect 18788 8832 18840 8838
rect 18788 8774 18840 8780
rect 18604 8492 18656 8498
rect 18604 8434 18656 8440
rect 18800 8362 18828 8774
rect 18788 8356 18840 8362
rect 18788 8298 18840 8304
rect 18696 8288 18748 8294
rect 18696 8230 18748 8236
rect 18708 7750 18736 8230
rect 18696 7744 18748 7750
rect 18696 7686 18748 7692
rect 18420 7404 18472 7410
rect 18420 7346 18472 7352
rect 18432 7002 18460 7346
rect 18512 7200 18564 7206
rect 18512 7142 18564 7148
rect 18420 6996 18472 7002
rect 18420 6938 18472 6944
rect 18432 6458 18460 6938
rect 18524 6934 18552 7142
rect 18512 6928 18564 6934
rect 18708 6905 18736 7686
rect 18512 6870 18564 6876
rect 18694 6896 18750 6905
rect 18694 6831 18750 6840
rect 18420 6452 18472 6458
rect 18420 6394 18472 6400
rect 18512 6248 18564 6254
rect 18512 6190 18564 6196
rect 18524 5914 18552 6190
rect 18512 5908 18564 5914
rect 18512 5850 18564 5856
rect 18340 5630 18460 5658
rect 18328 5568 18380 5574
rect 18328 5510 18380 5516
rect 18340 5234 18368 5510
rect 18328 5228 18380 5234
rect 18328 5170 18380 5176
rect 18340 4826 18368 5170
rect 18328 4820 18380 4826
rect 18328 4762 18380 4768
rect 18432 4146 18460 5630
rect 18512 5568 18564 5574
rect 18512 5510 18564 5516
rect 18524 5030 18552 5510
rect 18602 5128 18658 5137
rect 18602 5063 18658 5072
rect 18512 5024 18564 5030
rect 18512 4966 18564 4972
rect 18524 4865 18552 4966
rect 18510 4856 18566 4865
rect 18616 4826 18644 5063
rect 18800 4826 18828 8298
rect 18892 8022 18920 9279
rect 18984 9178 19012 9959
rect 19352 9654 19380 10134
rect 19432 9920 19484 9926
rect 19432 9862 19484 9868
rect 19340 9648 19392 9654
rect 19340 9590 19392 9596
rect 19444 9466 19472 9862
rect 19982 9752 20038 9761
rect 19982 9687 20038 9696
rect 19352 9450 19472 9466
rect 19340 9444 19472 9450
rect 19392 9438 19472 9444
rect 19340 9386 19392 9392
rect 19432 9376 19484 9382
rect 19432 9318 19484 9324
rect 19444 9217 19472 9318
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19430 9208 19486 9217
rect 18972 9172 19024 9178
rect 19622 9200 19918 9220
rect 19430 9143 19486 9152
rect 18972 9114 19024 9120
rect 19432 9036 19484 9042
rect 19432 8978 19484 8984
rect 19340 8968 19392 8974
rect 19340 8910 19392 8916
rect 19064 8832 19116 8838
rect 19064 8774 19116 8780
rect 19076 8430 19104 8774
rect 19352 8566 19380 8910
rect 19340 8560 19392 8566
rect 19340 8502 19392 8508
rect 19444 8498 19472 8978
rect 19524 8832 19576 8838
rect 19524 8774 19576 8780
rect 19432 8492 19484 8498
rect 19432 8434 19484 8440
rect 19064 8424 19116 8430
rect 19064 8366 19116 8372
rect 19076 8090 19104 8366
rect 19340 8356 19392 8362
rect 19340 8298 19392 8304
rect 19352 8106 19380 8298
rect 19260 8090 19380 8106
rect 19064 8084 19116 8090
rect 19064 8026 19116 8032
rect 19248 8084 19380 8090
rect 19300 8078 19380 8084
rect 19248 8026 19300 8032
rect 18880 8016 18932 8022
rect 19444 7993 19472 8434
rect 19536 8294 19564 8774
rect 19616 8560 19668 8566
rect 19616 8502 19668 8508
rect 19628 8401 19656 8502
rect 19614 8392 19670 8401
rect 19614 8327 19670 8336
rect 19524 8288 19576 8294
rect 19524 8230 19576 8236
rect 18880 7958 18932 7964
rect 19430 7984 19486 7993
rect 18892 7546 18920 7958
rect 19430 7919 19486 7928
rect 19536 7818 19564 8230
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19996 8090 20024 9687
rect 20074 8936 20130 8945
rect 20074 8871 20076 8880
rect 20128 8871 20130 8880
rect 20076 8842 20128 8848
rect 20088 8566 20116 8842
rect 20444 8832 20496 8838
rect 20258 8800 20314 8809
rect 20444 8774 20496 8780
rect 20258 8735 20314 8744
rect 20076 8560 20128 8566
rect 20076 8502 20128 8508
rect 19984 8084 20036 8090
rect 19984 8026 20036 8032
rect 19614 7848 19670 7857
rect 19524 7812 19576 7818
rect 19614 7783 19670 7792
rect 19524 7754 19576 7760
rect 18880 7540 18932 7546
rect 18880 7482 18932 7488
rect 19536 7410 19564 7754
rect 19628 7546 19656 7783
rect 19616 7540 19668 7546
rect 19616 7482 19668 7488
rect 19524 7404 19576 7410
rect 19524 7346 19576 7352
rect 18970 7304 19026 7313
rect 18970 7239 19026 7248
rect 18984 5234 19012 7239
rect 19536 7002 19564 7346
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19524 6996 19576 7002
rect 19524 6938 19576 6944
rect 19996 6934 20024 8026
rect 20076 7744 20128 7750
rect 20076 7686 20128 7692
rect 20088 7206 20116 7686
rect 20168 7268 20220 7274
rect 20168 7210 20220 7216
rect 20076 7200 20128 7206
rect 20076 7142 20128 7148
rect 19984 6928 20036 6934
rect 19984 6870 20036 6876
rect 19982 6488 20038 6497
rect 19982 6423 20038 6432
rect 19340 6112 19392 6118
rect 19340 6054 19392 6060
rect 19352 5273 19380 6054
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19524 5772 19576 5778
rect 19524 5714 19576 5720
rect 19432 5568 19484 5574
rect 19536 5545 19564 5714
rect 19432 5510 19484 5516
rect 19522 5536 19578 5545
rect 19338 5264 19394 5273
rect 18972 5228 19024 5234
rect 19338 5199 19394 5208
rect 18972 5170 19024 5176
rect 18510 4791 18566 4800
rect 18604 4820 18656 4826
rect 18604 4762 18656 4768
rect 18788 4820 18840 4826
rect 18788 4762 18840 4768
rect 18616 4214 18644 4762
rect 18984 4554 19012 5170
rect 19248 5160 19300 5166
rect 19248 5102 19300 5108
rect 19064 5024 19116 5030
rect 19062 4992 19064 5001
rect 19116 4992 19118 5001
rect 19062 4927 19118 4936
rect 19154 4720 19210 4729
rect 19154 4655 19156 4664
rect 19208 4655 19210 4664
rect 19156 4626 19208 4632
rect 18972 4548 19024 4554
rect 18972 4490 19024 4496
rect 18604 4208 18656 4214
rect 18510 4176 18566 4185
rect 18420 4140 18472 4146
rect 18604 4150 18656 4156
rect 18510 4111 18566 4120
rect 18420 4082 18472 4088
rect 18248 3964 18368 3992
rect 18340 3738 18368 3964
rect 18328 3732 18380 3738
rect 18328 3674 18380 3680
rect 18340 3194 18368 3674
rect 18328 3188 18380 3194
rect 18328 3130 18380 3136
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 18052 2576 18104 2582
rect 18050 2544 18052 2553
rect 18104 2544 18106 2553
rect 18050 2479 18106 2488
rect 18328 2304 18380 2310
rect 18328 2246 18380 2252
rect 18340 2009 18368 2246
rect 18326 2000 18382 2009
rect 18326 1935 18382 1944
rect 18524 480 18552 4111
rect 18984 3738 19012 4490
rect 19168 4282 19196 4626
rect 19260 4622 19288 5102
rect 19340 5024 19392 5030
rect 19340 4966 19392 4972
rect 19248 4616 19300 4622
rect 19248 4558 19300 4564
rect 19156 4276 19208 4282
rect 19156 4218 19208 4224
rect 19260 3942 19288 4558
rect 19352 4457 19380 4966
rect 19338 4448 19394 4457
rect 19338 4383 19394 4392
rect 19444 4185 19472 5510
rect 19522 5471 19578 5480
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19430 4176 19486 4185
rect 19430 4111 19486 4120
rect 19996 4078 20024 6423
rect 20088 5370 20116 7142
rect 20076 5364 20128 5370
rect 20076 5306 20128 5312
rect 20180 4593 20208 7210
rect 20166 4584 20222 4593
rect 20166 4519 20222 4528
rect 20272 4486 20300 8735
rect 20456 8430 20484 8774
rect 20444 8424 20496 8430
rect 20444 8366 20496 8372
rect 20536 7744 20588 7750
rect 20350 7712 20406 7721
rect 20536 7686 20588 7692
rect 20350 7647 20406 7656
rect 20260 4480 20312 4486
rect 20260 4422 20312 4428
rect 20364 4078 20392 7647
rect 20548 6662 20576 7686
rect 20640 7528 20668 15399
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 25502 15056 25558 15065
rect 25502 14991 25558 15000
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 25516 14074 25544 14991
rect 25504 14068 25556 14074
rect 25504 14010 25556 14016
rect 24398 13968 24454 13977
rect 24398 13903 24454 13912
rect 24412 13870 24440 13903
rect 24124 13864 24176 13870
rect 24122 13832 24124 13841
rect 24400 13864 24452 13870
rect 24176 13832 24178 13841
rect 24400 13806 24452 13812
rect 24122 13767 24178 13776
rect 24136 13530 24164 13767
rect 24124 13524 24176 13530
rect 24124 13466 24176 13472
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 21914 12880 21970 12889
rect 21914 12815 21970 12824
rect 20810 12200 20866 12209
rect 20810 12135 20866 12144
rect 20718 11112 20774 11121
rect 20718 11047 20774 11056
rect 20732 8634 20760 11047
rect 20720 8628 20772 8634
rect 20720 8570 20772 8576
rect 20720 7540 20772 7546
rect 20640 7500 20720 7528
rect 20720 7482 20772 7488
rect 20536 6656 20588 6662
rect 20536 6598 20588 6604
rect 20442 6488 20498 6497
rect 20442 6423 20444 6432
rect 20496 6423 20498 6432
rect 20444 6394 20496 6400
rect 20548 5914 20576 6598
rect 20824 6390 20852 12135
rect 21180 8832 21232 8838
rect 21180 8774 21232 8780
rect 20994 8664 21050 8673
rect 20994 8599 21050 8608
rect 21008 8566 21036 8599
rect 20996 8560 21048 8566
rect 21192 8537 21220 8774
rect 20996 8502 21048 8508
rect 21178 8528 21234 8537
rect 21178 8463 21180 8472
rect 21232 8463 21234 8472
rect 21180 8434 21232 8440
rect 21192 8403 21220 8434
rect 21640 8288 21692 8294
rect 21640 8230 21692 8236
rect 21652 7954 21680 8230
rect 21640 7948 21692 7954
rect 21640 7890 21692 7896
rect 20994 7440 21050 7449
rect 20994 7375 20996 7384
rect 21048 7375 21050 7384
rect 20996 7346 21048 7352
rect 21180 7268 21232 7274
rect 21180 7210 21232 7216
rect 20994 6896 21050 6905
rect 20994 6831 21050 6840
rect 21008 6390 21036 6831
rect 21192 6798 21220 7210
rect 21548 7200 21600 7206
rect 21548 7142 21600 7148
rect 21180 6792 21232 6798
rect 21178 6760 21180 6769
rect 21232 6760 21234 6769
rect 21178 6695 21234 6704
rect 21560 6662 21588 7142
rect 21548 6656 21600 6662
rect 21548 6598 21600 6604
rect 20812 6384 20864 6390
rect 20812 6326 20864 6332
rect 20996 6384 21048 6390
rect 20996 6326 21048 6332
rect 20536 5908 20588 5914
rect 20536 5850 20588 5856
rect 20548 5370 20576 5850
rect 21560 5817 21588 6598
rect 21652 6474 21680 7890
rect 21652 6446 21772 6474
rect 21640 6316 21692 6322
rect 21640 6258 21692 6264
rect 21546 5808 21602 5817
rect 21546 5743 21602 5752
rect 21178 5672 21234 5681
rect 21178 5607 21234 5616
rect 20720 5568 20772 5574
rect 20720 5510 20772 5516
rect 20536 5364 20588 5370
rect 20536 5306 20588 5312
rect 20548 4826 20576 5306
rect 20732 5234 20760 5510
rect 20720 5228 20772 5234
rect 20720 5170 20772 5176
rect 21192 5166 21220 5607
rect 21652 5574 21680 6258
rect 21640 5568 21692 5574
rect 21640 5510 21692 5516
rect 21180 5160 21232 5166
rect 21180 5102 21232 5108
rect 21456 5092 21508 5098
rect 21456 5034 21508 5040
rect 21364 5024 21416 5030
rect 21364 4966 21416 4972
rect 21376 4826 21404 4966
rect 20536 4820 20588 4826
rect 20536 4762 20588 4768
rect 21364 4820 21416 4826
rect 21364 4762 21416 4768
rect 20628 4480 20680 4486
rect 20680 4440 20760 4468
rect 20628 4422 20680 4428
rect 19984 4072 20036 4078
rect 19984 4014 20036 4020
rect 20352 4072 20404 4078
rect 20352 4014 20404 4020
rect 20260 4004 20312 4010
rect 20260 3946 20312 3952
rect 19248 3936 19300 3942
rect 19248 3878 19300 3884
rect 19524 3936 19576 3942
rect 20076 3936 20128 3942
rect 19524 3878 19576 3884
rect 20074 3904 20076 3913
rect 20128 3904 20130 3913
rect 18972 3732 19024 3738
rect 18972 3674 19024 3680
rect 19154 3632 19210 3641
rect 19154 3567 19156 3576
rect 19208 3567 19210 3576
rect 19156 3538 19208 3544
rect 18604 3528 18656 3534
rect 18604 3470 18656 3476
rect 18616 3058 18644 3470
rect 19064 3188 19116 3194
rect 19064 3130 19116 3136
rect 18604 3052 18656 3058
rect 18604 2994 18656 3000
rect 18616 2378 18644 2994
rect 19076 2553 19104 3130
rect 19260 2990 19288 3878
rect 19338 3768 19394 3777
rect 19338 3703 19394 3712
rect 19352 3602 19380 3703
rect 19536 3641 19564 3878
rect 19622 3836 19918 3856
rect 20074 3839 20130 3848
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 20168 3732 20220 3738
rect 20168 3674 20220 3680
rect 19522 3632 19578 3641
rect 19340 3596 19392 3602
rect 19522 3567 19578 3576
rect 19340 3538 19392 3544
rect 19352 3194 19380 3538
rect 19524 3392 19576 3398
rect 19524 3334 19576 3340
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 19536 3097 19564 3334
rect 19522 3088 19578 3097
rect 19522 3023 19578 3032
rect 19248 2984 19300 2990
rect 19248 2926 19300 2932
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 19522 2952 19578 2961
rect 19352 2689 19380 2926
rect 19522 2887 19578 2896
rect 19338 2680 19394 2689
rect 19338 2615 19394 2624
rect 19062 2544 19118 2553
rect 19062 2479 19118 2488
rect 18604 2372 18656 2378
rect 18604 2314 18656 2320
rect 19062 1592 19118 1601
rect 19062 1527 19118 1536
rect 19076 480 19104 1527
rect 19536 1442 19564 2887
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 20180 2689 20208 3674
rect 20166 2680 20222 2689
rect 20166 2615 20222 2624
rect 19892 2508 19944 2514
rect 19892 2450 19944 2456
rect 19904 2145 19932 2450
rect 19890 2136 19946 2145
rect 19890 2071 19946 2080
rect 19536 1414 19656 1442
rect 19628 480 19656 1414
rect 20272 480 20300 3946
rect 20364 3738 20392 4014
rect 20732 3738 20760 4440
rect 21376 3738 21404 4762
rect 21468 4690 21496 5034
rect 21456 4684 21508 4690
rect 21456 4626 21508 4632
rect 21468 4282 21496 4626
rect 21456 4276 21508 4282
rect 21456 4218 21508 4224
rect 20352 3732 20404 3738
rect 20352 3674 20404 3680
rect 20720 3732 20772 3738
rect 20720 3674 20772 3680
rect 21364 3732 21416 3738
rect 21364 3674 21416 3680
rect 20904 3596 20956 3602
rect 20904 3538 20956 3544
rect 20812 3392 20864 3398
rect 20812 3334 20864 3340
rect 20718 3224 20774 3233
rect 20718 3159 20774 3168
rect 20732 2990 20760 3159
rect 20720 2984 20772 2990
rect 20720 2926 20772 2932
rect 20720 2304 20772 2310
rect 20718 2272 20720 2281
rect 20772 2272 20774 2281
rect 20718 2207 20774 2216
rect 20824 480 20852 3334
rect 20916 3194 20944 3538
rect 21744 3194 21772 6446
rect 21928 4729 21956 12815
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 22008 6248 22060 6254
rect 22060 6196 22324 6202
rect 22008 6190 22324 6196
rect 22020 6174 22324 6190
rect 22100 6112 22152 6118
rect 22100 6054 22152 6060
rect 22112 5030 22140 6054
rect 22100 5024 22152 5030
rect 22100 4966 22152 4972
rect 21914 4720 21970 4729
rect 21914 4655 21970 4664
rect 21824 4072 21876 4078
rect 21824 4014 21876 4020
rect 21836 3398 21864 4014
rect 22008 3936 22060 3942
rect 22008 3878 22060 3884
rect 22020 3505 22048 3878
rect 22006 3496 22062 3505
rect 22006 3431 22062 3440
rect 22100 3460 22152 3466
rect 22100 3402 22152 3408
rect 21824 3392 21876 3398
rect 21822 3360 21824 3369
rect 21876 3360 21878 3369
rect 21822 3295 21878 3304
rect 22112 3194 22140 3402
rect 22192 3392 22244 3398
rect 22192 3334 22244 3340
rect 20904 3188 20956 3194
rect 20904 3130 20956 3136
rect 21732 3188 21784 3194
rect 21732 3130 21784 3136
rect 22100 3188 22152 3194
rect 22100 3130 22152 3136
rect 21364 3120 21416 3126
rect 21364 3062 21416 3068
rect 21178 2544 21234 2553
rect 21178 2479 21180 2488
rect 21232 2479 21234 2488
rect 21180 2450 21232 2456
rect 21376 480 21404 3062
rect 21744 2990 21772 3130
rect 21732 2984 21784 2990
rect 22204 2961 22232 3334
rect 21732 2926 21784 2932
rect 22190 2952 22246 2961
rect 22190 2887 22246 2896
rect 22006 2816 22062 2825
rect 22006 2751 22062 2760
rect 22020 2650 22048 2751
rect 22098 2680 22154 2689
rect 22008 2644 22060 2650
rect 22098 2615 22100 2624
rect 22008 2586 22060 2592
rect 22152 2615 22154 2624
rect 22100 2586 22152 2592
rect 22296 2514 22324 6174
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 22374 5128 22430 5137
rect 22374 5063 22430 5072
rect 22388 4690 22416 5063
rect 22376 4684 22428 4690
rect 22376 4626 22428 4632
rect 22388 4282 22416 4626
rect 23480 4616 23532 4622
rect 23480 4558 23532 4564
rect 23112 4480 23164 4486
rect 23112 4422 23164 4428
rect 22376 4276 22428 4282
rect 22376 4218 22428 4224
rect 22468 2916 22520 2922
rect 22468 2858 22520 2864
rect 22284 2508 22336 2514
rect 22284 2450 22336 2456
rect 21916 2372 21968 2378
rect 21916 2314 21968 2320
rect 21928 480 21956 2314
rect 22480 480 22508 2858
rect 23124 480 23152 4422
rect 23492 4078 23520 4558
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 23480 4072 23532 4078
rect 23480 4014 23532 4020
rect 25320 3936 25372 3942
rect 25320 3878 25372 3884
rect 26514 3904 26570 3913
rect 24122 3768 24178 3777
rect 24122 3703 24178 3712
rect 24032 2508 24084 2514
rect 24032 2450 24084 2456
rect 23664 2372 23716 2378
rect 23664 2314 23716 2320
rect 23480 2304 23532 2310
rect 23480 2246 23532 2252
rect 23492 1601 23520 2246
rect 23478 1592 23534 1601
rect 23478 1527 23534 1536
rect 23676 480 23704 2314
rect 24044 1873 24072 2450
rect 24030 1864 24086 1873
rect 24030 1799 24086 1808
rect 24136 1442 24164 3703
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24766 2816 24822 2825
rect 24766 2751 24822 2760
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24136 1414 24256 1442
rect 24228 480 24256 1414
rect 24780 480 24808 2751
rect 25332 480 25360 3878
rect 26514 3839 26570 3848
rect 25962 3088 26018 3097
rect 25962 3023 26018 3032
rect 25976 480 26004 3023
rect 26528 480 26556 3839
rect 27618 3632 27674 3641
rect 27618 3567 27674 3576
rect 27066 2408 27122 2417
rect 27066 2343 27122 2352
rect 27080 480 27108 2343
rect 27632 480 27660 3567
rect 294 0 350 480
rect 846 0 902 480
rect 1398 0 1454 480
rect 1950 0 2006 480
rect 2502 0 2558 480
rect 3146 0 3202 480
rect 3698 0 3754 480
rect 4250 0 4306 480
rect 4802 0 4858 480
rect 5354 0 5410 480
rect 5998 0 6054 480
rect 6550 0 6606 480
rect 7102 0 7158 480
rect 7654 0 7710 480
rect 8206 0 8262 480
rect 8850 0 8906 480
rect 9402 0 9458 480
rect 9954 0 10010 480
rect 10506 0 10562 480
rect 11058 0 11114 480
rect 11702 0 11758 480
rect 12254 0 12310 480
rect 12806 0 12862 480
rect 13358 0 13414 480
rect 13910 0 13966 480
rect 14554 0 14610 480
rect 15106 0 15162 480
rect 15658 0 15714 480
rect 16210 0 16266 480
rect 16762 0 16818 480
rect 17406 0 17462 480
rect 17958 0 18014 480
rect 18510 0 18566 480
rect 19062 0 19118 480
rect 19614 0 19670 480
rect 20258 0 20314 480
rect 20810 0 20866 480
rect 21362 0 21418 480
rect 21914 0 21970 480
rect 22466 0 22522 480
rect 23110 0 23166 480
rect 23662 0 23718 480
rect 24214 0 24270 480
rect 24766 0 24822 480
rect 25318 0 25374 480
rect 25962 0 26018 480
rect 26514 0 26570 480
rect 27066 0 27122 480
rect 27618 0 27674 480
<< via2 >>
rect 3514 27648 3570 27704
rect 294 20984 350 21040
rect 1766 24676 1822 24712
rect 1766 24656 1768 24676
rect 1768 24656 1820 24676
rect 1820 24656 1822 24676
rect 1766 24248 1822 24304
rect 1582 21936 1638 21992
rect 1674 20848 1730 20904
rect 1766 20440 1822 20496
rect 1490 19216 1546 19272
rect 1950 24520 2006 24576
rect 2042 21528 2098 21584
rect 2134 21392 2190 21448
rect 2226 19796 2228 19816
rect 2228 19796 2280 19816
rect 2280 19796 2282 19816
rect 2226 19760 2282 19796
rect 1582 16360 1638 16416
rect 1398 13232 1454 13288
rect 1582 13096 1638 13152
rect 2042 15544 2098 15600
rect 2410 23860 2466 23896
rect 2410 23840 2412 23860
rect 2412 23840 2464 23860
rect 2464 23840 2466 23860
rect 2686 23704 2742 23760
rect 2502 20304 2558 20360
rect 2870 20712 2926 20768
rect 2686 20168 2742 20224
rect 2594 17992 2650 18048
rect 2502 16088 2558 16144
rect 2410 15136 2466 15192
rect 2502 13912 2558 13968
rect 2042 13388 2098 13424
rect 2042 13368 2044 13388
rect 2044 13368 2096 13388
rect 2096 13368 2098 13388
rect 1858 13096 1914 13152
rect 1398 9460 1400 9480
rect 1400 9460 1452 9480
rect 1452 9460 1454 9480
rect 1398 9424 1454 9460
rect 1122 4392 1178 4448
rect 846 2080 902 2136
rect 294 1672 350 1728
rect 1582 9560 1638 9616
rect 1490 9016 1546 9072
rect 2410 13640 2466 13696
rect 2042 10412 2044 10432
rect 2044 10412 2096 10432
rect 2096 10412 2098 10432
rect 2042 10376 2098 10412
rect 1858 10240 1914 10296
rect 1950 8608 2006 8664
rect 1766 7384 1822 7440
rect 1858 4936 1914 4992
rect 1398 3304 1454 3360
rect 1306 856 1362 912
rect 2686 16360 2742 16416
rect 2778 15816 2834 15872
rect 2686 15408 2742 15464
rect 3514 27104 3570 27160
rect 3330 25336 3386 25392
rect 3146 21800 3202 21856
rect 3514 24112 3570 24168
rect 3606 22636 3662 22672
rect 3606 22616 3608 22636
rect 3608 22616 3660 22636
rect 3660 22616 3662 22636
rect 3238 21256 3294 21312
rect 3330 20984 3386 21040
rect 3054 19488 3110 19544
rect 3238 18944 3294 19000
rect 2962 17584 3018 17640
rect 2962 17176 3018 17232
rect 2870 13912 2926 13968
rect 2962 13640 3018 13696
rect 2686 12688 2742 12744
rect 3238 13812 3240 13832
rect 3240 13812 3292 13832
rect 3292 13812 3294 13832
rect 3238 13776 3294 13812
rect 4066 26580 4122 26616
rect 4066 26560 4068 26580
rect 4068 26560 4120 26580
rect 4120 26560 4122 26580
rect 4066 25880 4122 25936
rect 4066 24792 4122 24848
rect 4066 23568 4122 23624
rect 3974 22480 4030 22536
rect 3514 17312 3570 17368
rect 4250 19080 4306 19136
rect 3698 16632 3754 16688
rect 2410 8356 2466 8392
rect 2410 8336 2412 8356
rect 2412 8336 2464 8356
rect 2464 8336 2466 8356
rect 3422 13368 3478 13424
rect 3606 13504 3662 13560
rect 3514 13096 3570 13152
rect 3422 12416 3478 12472
rect 2962 10648 3018 10704
rect 3054 9016 3110 9072
rect 2410 5752 2466 5808
rect 1950 4120 2006 4176
rect 2042 3984 2098 4040
rect 2318 5072 2374 5128
rect 2318 4120 2374 4176
rect 3054 5480 3110 5536
rect 2594 3304 2650 3360
rect 2870 3032 2926 3088
rect 2318 2896 2374 2952
rect 2502 2760 2558 2816
rect 3054 3712 3110 3768
rect 3146 3032 3202 3088
rect 4158 16496 4214 16552
rect 3882 15680 3938 15736
rect 3790 15408 3846 15464
rect 3974 15000 4030 15056
rect 3882 14864 3938 14920
rect 3698 13368 3754 13424
rect 4526 21256 4582 21312
rect 4802 20204 4804 20224
rect 4804 20204 4856 20224
rect 4856 20204 4858 20224
rect 4802 20168 4858 20204
rect 5170 23840 5226 23896
rect 4986 23296 5042 23352
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5814 23160 5870 23216
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5170 20984 5226 21040
rect 4618 17992 4674 18048
rect 4342 15680 4398 15736
rect 3882 12824 3938 12880
rect 4434 15544 4490 15600
rect 4526 15136 4582 15192
rect 4710 15852 4712 15872
rect 4712 15852 4764 15872
rect 4764 15852 4766 15872
rect 4710 15816 4766 15852
rect 4526 13232 4582 13288
rect 3974 11192 4030 11248
rect 3790 10920 3846 10976
rect 3330 7928 3386 7984
rect 4066 10376 4122 10432
rect 3974 10104 4030 10160
rect 3790 7792 3846 7848
rect 3974 7792 4030 7848
rect 3330 4936 3386 4992
rect 3238 2488 3294 2544
rect 3606 5228 3662 5264
rect 3606 5208 3608 5228
rect 3608 5208 3660 5228
rect 3660 5208 3662 5228
rect 3422 3884 3424 3904
rect 3424 3884 3476 3904
rect 3476 3884 3478 3904
rect 3422 3848 3478 3884
rect 3974 6840 4030 6896
rect 3882 4528 3938 4584
rect 3882 3984 3938 4040
rect 3790 3712 3846 3768
rect 3698 3168 3754 3224
rect 3698 2896 3754 2952
rect 3606 2352 3662 2408
rect 4066 5888 4122 5944
rect 4066 5636 4122 5672
rect 4066 5616 4068 5636
rect 4068 5616 4120 5636
rect 4120 5616 4122 5636
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5446 18400 5502 18456
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 6182 23568 6238 23624
rect 6090 21528 6146 21584
rect 6918 24656 6974 24712
rect 6550 23296 6606 23352
rect 6458 23024 6514 23080
rect 6274 22616 6330 22672
rect 6274 21528 6330 21584
rect 6182 20984 6238 21040
rect 6734 23296 6790 23352
rect 6550 20168 6606 20224
rect 6642 19508 6698 19544
rect 6642 19488 6644 19508
rect 6644 19488 6696 19508
rect 6696 19488 6698 19508
rect 6550 18672 6606 18728
rect 5814 16768 5870 16824
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5170 15952 5226 16008
rect 5078 14884 5134 14920
rect 5078 14864 5080 14884
rect 5080 14864 5132 14884
rect 5132 14864 5134 14884
rect 5262 14184 5318 14240
rect 5170 12144 5226 12200
rect 4342 7928 4398 7984
rect 4618 8200 4674 8256
rect 4526 7384 4582 7440
rect 4526 4664 4582 4720
rect 4342 1944 4398 2000
rect 4710 3304 4766 3360
rect 5078 9580 5134 9616
rect 5078 9560 5080 9580
rect 5080 9560 5132 9580
rect 5132 9560 5134 9580
rect 5170 7420 5172 7440
rect 5172 7420 5224 7440
rect 5224 7420 5226 7440
rect 5170 7384 5226 7420
rect 5078 5752 5134 5808
rect 5998 15444 6000 15464
rect 6000 15444 6052 15464
rect 6052 15444 6054 15464
rect 5998 15408 6054 15444
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5998 15136 6054 15192
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5630 13776 5686 13832
rect 5538 13640 5594 13696
rect 5814 13368 5870 13424
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5814 10684 5816 10704
rect 5816 10684 5868 10704
rect 5868 10684 5870 10704
rect 5814 10648 5870 10684
rect 5630 10260 5686 10296
rect 5630 10240 5632 10260
rect 5632 10240 5684 10260
rect 5684 10240 5686 10260
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 6090 15000 6146 15056
rect 6182 14320 6238 14376
rect 6090 10140 6092 10160
rect 6092 10140 6144 10160
rect 6144 10140 6146 10160
rect 6090 10104 6146 10140
rect 5998 8508 6000 8528
rect 6000 8508 6052 8528
rect 6052 8508 6054 8528
rect 5998 8472 6054 8508
rect 5538 8336 5594 8392
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5998 6704 6054 6760
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 6090 5772 6146 5808
rect 6090 5752 6092 5772
rect 6092 5752 6144 5772
rect 6144 5752 6146 5772
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5998 4392 6054 4448
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 6090 3712 6146 3768
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5630 3068 5632 3088
rect 5632 3068 5684 3088
rect 5684 3068 5686 3088
rect 5630 3032 5686 3068
rect 5262 2488 5318 2544
rect 5354 2352 5410 2408
rect 5170 2080 5226 2136
rect 4894 1400 4950 1456
rect 6090 2216 6146 2272
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 6458 16632 6514 16688
rect 6918 23976 6974 24032
rect 6918 23024 6974 23080
rect 7746 24384 7802 24440
rect 7838 24248 7894 24304
rect 7010 20304 7066 20360
rect 6826 18400 6882 18456
rect 7010 19116 7012 19136
rect 7012 19116 7064 19136
rect 7064 19116 7066 19136
rect 7010 19080 7066 19116
rect 6642 15680 6698 15736
rect 6550 15000 6606 15056
rect 6642 13640 6698 13696
rect 6274 8780 6276 8800
rect 6276 8780 6328 8800
rect 6328 8780 6330 8800
rect 6274 8744 6330 8780
rect 7102 15136 7158 15192
rect 7102 13812 7104 13832
rect 7104 13812 7156 13832
rect 7156 13812 7158 13832
rect 7102 13776 7158 13812
rect 6826 13640 6882 13696
rect 7286 15544 7342 15600
rect 6734 12552 6790 12608
rect 6458 8064 6514 8120
rect 6642 8372 6644 8392
rect 6644 8372 6696 8392
rect 6696 8372 6698 8392
rect 6642 8336 6698 8372
rect 6642 7520 6698 7576
rect 6826 12416 6882 12472
rect 6826 10532 6882 10568
rect 6826 10512 6828 10532
rect 6828 10512 6880 10532
rect 6880 10512 6882 10532
rect 7378 13096 7434 13152
rect 7010 11192 7066 11248
rect 7194 10648 7250 10704
rect 7102 9988 7158 10024
rect 7102 9968 7104 9988
rect 7104 9968 7156 9988
rect 7156 9968 7158 9988
rect 7194 9424 7250 9480
rect 7102 8200 7158 8256
rect 6826 7248 6882 7304
rect 6826 6332 6828 6352
rect 6828 6332 6880 6352
rect 6880 6332 6882 6352
rect 6826 6296 6882 6332
rect 6918 5908 6974 5944
rect 6918 5888 6920 5908
rect 6920 5888 6972 5908
rect 6972 5888 6974 5908
rect 6366 2388 6368 2408
rect 6368 2388 6420 2408
rect 6420 2388 6422 2408
rect 6366 2352 6422 2388
rect 6826 3984 6882 4040
rect 7102 7656 7158 7712
rect 7286 6432 7342 6488
rect 7286 6024 7342 6080
rect 7378 3848 7434 3904
rect 6734 3440 6790 3496
rect 7654 21392 7710 21448
rect 7654 18128 7710 18184
rect 7746 17992 7802 18048
rect 7838 17176 7894 17232
rect 8666 24148 8668 24168
rect 8668 24148 8720 24168
rect 8720 24148 8722 24168
rect 8666 24112 8722 24148
rect 8022 22108 8024 22128
rect 8024 22108 8076 22128
rect 8076 22108 8078 22128
rect 8022 22072 8078 22108
rect 8482 22480 8538 22536
rect 8390 20032 8446 20088
rect 8022 19760 8078 19816
rect 8206 18964 8262 19000
rect 8206 18944 8208 18964
rect 8208 18944 8260 18964
rect 8260 18944 8262 18964
rect 8850 24384 8906 24440
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 9034 23860 9090 23896
rect 9678 24248 9734 24304
rect 9034 23840 9036 23860
rect 9036 23840 9088 23860
rect 9088 23840 9090 23860
rect 9494 23704 9550 23760
rect 8942 23160 8998 23216
rect 8850 19760 8906 19816
rect 8482 18128 8538 18184
rect 8850 18808 8906 18864
rect 8850 18536 8906 18592
rect 8758 18264 8814 18320
rect 8482 16768 8538 16824
rect 8666 16632 8722 16688
rect 8206 13232 8262 13288
rect 9126 21120 9182 21176
rect 9678 23296 9734 23352
rect 9494 20576 9550 20632
rect 9126 20168 9182 20224
rect 8942 17992 8998 18048
rect 9494 19488 9550 19544
rect 9218 19352 9274 19408
rect 9770 21292 9772 21312
rect 9772 21292 9824 21312
rect 9824 21292 9826 21312
rect 9770 21256 9826 21292
rect 9770 17720 9826 17776
rect 9586 17076 9588 17096
rect 9588 17076 9640 17096
rect 9640 17076 9642 17096
rect 9586 17040 9642 17076
rect 8942 16652 8998 16688
rect 8942 16632 8944 16652
rect 8944 16632 8996 16652
rect 8996 16632 8998 16652
rect 7562 7384 7618 7440
rect 7838 7928 7894 7984
rect 9770 15544 9826 15600
rect 8482 10104 8538 10160
rect 8114 9424 8170 9480
rect 8206 8508 8208 8528
rect 8208 8508 8260 8528
rect 8260 8508 8262 8528
rect 8206 8472 8262 8508
rect 8850 8336 8906 8392
rect 8666 7828 8668 7848
rect 8668 7828 8720 7848
rect 8720 7828 8722 7848
rect 8666 7792 8722 7828
rect 8666 7540 8722 7576
rect 8666 7520 8668 7540
rect 8668 7520 8720 7540
rect 8720 7520 8722 7540
rect 8206 6840 8262 6896
rect 8022 6160 8078 6216
rect 7746 4392 7802 4448
rect 7470 3032 7526 3088
rect 7930 4972 7932 4992
rect 7932 4972 7984 4992
rect 7984 4972 7986 4992
rect 7930 4936 7986 4972
rect 7838 2352 7894 2408
rect 7654 1808 7710 1864
rect 8850 4120 8906 4176
rect 8390 2896 8446 2952
rect 8758 3168 8814 3224
rect 8758 2796 8760 2816
rect 8760 2796 8812 2816
rect 8812 2796 8814 2816
rect 8758 2760 8814 2796
rect 9218 9288 9274 9344
rect 9494 8880 9550 8936
rect 9310 7812 9366 7848
rect 9310 7792 9312 7812
rect 9312 7792 9364 7812
rect 9364 7792 9366 7812
rect 9678 7948 9734 7984
rect 9678 7928 9680 7948
rect 9680 7928 9732 7948
rect 9732 7928 9734 7948
rect 9586 6996 9642 7032
rect 9586 6976 9588 6996
rect 9588 6976 9640 6996
rect 9640 6976 9642 6996
rect 9678 6024 9734 6080
rect 9034 5636 9090 5672
rect 9034 5616 9036 5636
rect 9036 5616 9088 5636
rect 9088 5616 9090 5636
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10230 21800 10286 21856
rect 10046 20440 10102 20496
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10138 18944 10194 19000
rect 9954 18400 10010 18456
rect 11242 24112 11298 24168
rect 11058 23840 11114 23896
rect 11702 23840 11758 23896
rect 11242 22616 11298 22672
rect 11058 22072 11114 22128
rect 11242 22072 11298 22128
rect 10874 19488 10930 19544
rect 11794 20304 11850 20360
rect 11242 19488 11298 19544
rect 11150 19236 11206 19272
rect 11150 19216 11152 19236
rect 11152 19216 11204 19236
rect 11204 19216 11206 19236
rect 11242 18944 11298 19000
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 11242 18536 11298 18592
rect 10874 17856 10930 17912
rect 10782 17720 10838 17776
rect 10874 16788 10930 16824
rect 10874 16768 10876 16788
rect 10876 16768 10928 16788
rect 10928 16768 10930 16788
rect 11242 17584 11298 17640
rect 11242 16768 11298 16824
rect 10782 15700 10838 15736
rect 10782 15680 10784 15700
rect 10784 15680 10836 15700
rect 10836 15680 10838 15700
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10138 12416 10194 12472
rect 10046 11328 10102 11384
rect 10782 13776 10838 13832
rect 11242 15272 11298 15328
rect 11702 15952 11758 16008
rect 11702 15564 11758 15600
rect 11702 15544 11704 15564
rect 11704 15544 11756 15564
rect 11756 15544 11758 15564
rect 11610 14864 11666 14920
rect 11334 14728 11390 14784
rect 10690 12144 10746 12200
rect 11334 13232 11390 13288
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10138 11056 10194 11112
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10598 9560 10654 9616
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10138 9016 10194 9072
rect 10046 8744 10102 8800
rect 9954 8200 10010 8256
rect 10690 8236 10692 8256
rect 10692 8236 10744 8256
rect 10744 8236 10746 8256
rect 10690 8200 10746 8236
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10138 7112 10194 7168
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10690 6316 10746 6352
rect 10690 6296 10692 6316
rect 10692 6296 10744 6316
rect 10744 6296 10746 6316
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10690 5788 10692 5808
rect 10692 5788 10744 5808
rect 10744 5788 10746 5808
rect 10690 5752 10746 5788
rect 9862 4664 9918 4720
rect 9402 3576 9458 3632
rect 9310 3440 9366 3496
rect 8942 2896 8998 2952
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10690 3984 10746 4040
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 11426 11736 11482 11792
rect 11610 10804 11666 10840
rect 11610 10784 11612 10804
rect 11612 10784 11664 10804
rect 11664 10784 11666 10804
rect 11242 9560 11298 9616
rect 11334 9424 11390 9480
rect 11242 9324 11244 9344
rect 11244 9324 11296 9344
rect 11296 9324 11298 9344
rect 11242 9288 11298 9324
rect 11150 8880 11206 8936
rect 11150 6432 11206 6488
rect 11242 5616 11298 5672
rect 11426 8200 11482 8256
rect 11518 6024 11574 6080
rect 11334 5480 11390 5536
rect 11334 4528 11390 4584
rect 11150 2896 11206 2952
rect 11242 2372 11298 2408
rect 11242 2352 11244 2372
rect 11244 2352 11296 2372
rect 11296 2352 11298 2372
rect 11518 3304 11574 3360
rect 11610 3032 11666 3088
rect 11426 2896 11482 2952
rect 11334 2216 11390 2272
rect 11610 1672 11666 1728
rect 12070 24656 12126 24712
rect 11978 19624 12034 19680
rect 12162 21564 12164 21584
rect 12164 21564 12216 21584
rect 12216 21564 12218 21584
rect 12162 21528 12218 21564
rect 12622 23740 12624 23760
rect 12624 23740 12676 23760
rect 12676 23740 12678 23760
rect 12622 23704 12678 23740
rect 13358 24656 13414 24712
rect 13450 23468 13452 23488
rect 13452 23468 13504 23488
rect 13504 23468 13506 23488
rect 12530 20868 12586 20904
rect 12530 20848 12532 20868
rect 12532 20848 12584 20868
rect 12584 20848 12586 20868
rect 12254 18944 12310 19000
rect 13450 23432 13506 23468
rect 12806 20440 12862 20496
rect 12898 19760 12954 19816
rect 12806 19352 12862 19408
rect 12622 18844 12624 18864
rect 12624 18844 12676 18864
rect 12676 18844 12678 18864
rect 12622 18808 12678 18844
rect 12714 17876 12770 17912
rect 12714 17856 12716 17876
rect 12716 17856 12768 17876
rect 12768 17856 12770 17876
rect 12346 17584 12402 17640
rect 12254 17176 12310 17232
rect 11978 17040 12034 17096
rect 11886 12416 11942 12472
rect 11978 11736 12034 11792
rect 11886 11056 11942 11112
rect 11794 8608 11850 8664
rect 12070 6160 12126 6216
rect 11886 4936 11942 4992
rect 11978 2488 12034 2544
rect 12162 3848 12218 3904
rect 11886 1536 11942 1592
rect 12622 17740 12678 17776
rect 12622 17720 12624 17740
rect 12624 17720 12676 17740
rect 12676 17720 12678 17740
rect 12530 16496 12586 16552
rect 12622 16124 12624 16144
rect 12624 16124 12676 16144
rect 12676 16124 12678 16144
rect 12622 16088 12678 16124
rect 12346 7248 12402 7304
rect 13174 19896 13230 19952
rect 12990 19216 13046 19272
rect 12990 18808 13046 18864
rect 13174 18264 13230 18320
rect 12990 16632 13046 16688
rect 13726 23432 13782 23488
rect 13910 22636 13966 22672
rect 13910 22616 13912 22636
rect 13912 22616 13964 22636
rect 13964 22616 13966 22636
rect 14002 21800 14058 21856
rect 13358 19352 13414 19408
rect 13266 15272 13322 15328
rect 13542 19216 13598 19272
rect 13450 19080 13506 19136
rect 13450 18264 13506 18320
rect 13910 19080 13966 19136
rect 14094 20576 14150 20632
rect 13726 16632 13782 16688
rect 13634 16496 13690 16552
rect 12898 13232 12954 13288
rect 12898 12436 12954 12472
rect 12898 12416 12900 12436
rect 12900 12416 12952 12436
rect 12952 12416 12954 12436
rect 12714 10920 12770 10976
rect 13174 13776 13230 13832
rect 13358 13096 13414 13152
rect 14370 23840 14426 23896
rect 14278 19760 14334 19816
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 15566 23432 15622 23488
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14830 21392 14886 21448
rect 14738 20848 14794 20904
rect 14646 19216 14702 19272
rect 14738 18944 14794 19000
rect 15382 21936 15438 21992
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14278 14356 14280 14376
rect 14280 14356 14332 14376
rect 14332 14356 14334 14376
rect 14278 14320 14334 14356
rect 14462 14456 14518 14512
rect 13634 12980 13690 13016
rect 13634 12960 13636 12980
rect 13636 12960 13688 12980
rect 13688 12960 13690 12980
rect 13818 12824 13874 12880
rect 13450 10784 13506 10840
rect 12898 6296 12954 6352
rect 12714 3712 12770 3768
rect 12714 3476 12716 3496
rect 12716 3476 12768 3496
rect 12768 3476 12770 3496
rect 12714 3440 12770 3476
rect 12438 2796 12440 2816
rect 12440 2796 12492 2816
rect 12492 2796 12494 2816
rect 12438 2760 12494 2796
rect 12990 3168 13046 3224
rect 13542 8628 13598 8664
rect 13542 8608 13544 8628
rect 13544 8608 13596 8628
rect 13596 8608 13598 8628
rect 14094 9696 14150 9752
rect 14094 8064 14150 8120
rect 13358 3848 13414 3904
rect 13082 2624 13138 2680
rect 12990 2488 13046 2544
rect 12898 1944 12954 2000
rect 13634 3712 13690 3768
rect 13634 3596 13690 3632
rect 13634 3576 13636 3596
rect 13636 3576 13688 3596
rect 13688 3576 13690 3596
rect 13542 2352 13598 2408
rect 14278 12280 14334 12336
rect 14370 11056 14426 11112
rect 14278 10920 14334 10976
rect 14278 9444 14334 9480
rect 14278 9424 14280 9444
rect 14280 9424 14332 9444
rect 14332 9424 14334 9444
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 15014 17076 15016 17096
rect 15016 17076 15068 17096
rect 15068 17076 15070 17096
rect 15014 17040 15070 17076
rect 15290 16768 15346 16824
rect 14922 16668 14924 16688
rect 14924 16668 14976 16688
rect 14976 16668 14978 16688
rect 14922 16632 14978 16668
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 16394 24268 16450 24304
rect 16394 24248 16396 24268
rect 16396 24248 16448 24268
rect 16448 24248 16450 24268
rect 16486 23976 16542 24032
rect 16854 22652 16856 22672
rect 16856 22652 16908 22672
rect 16908 22652 16910 22672
rect 16854 22616 16910 22652
rect 15658 19080 15714 19136
rect 15474 18128 15530 18184
rect 15658 17856 15714 17912
rect 15658 17312 15714 17368
rect 16210 19760 16266 19816
rect 15382 13232 15438 13288
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 15014 12144 15070 12200
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14830 11736 14886 11792
rect 14738 9832 14794 9888
rect 14738 8744 14794 8800
rect 14738 8336 14794 8392
rect 14738 7656 14794 7712
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 15382 9716 15438 9752
rect 15382 9696 15384 9716
rect 15384 9696 15436 9716
rect 15436 9696 15438 9716
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 15106 8084 15162 8120
rect 15106 8064 15108 8084
rect 15108 8064 15160 8084
rect 15160 8064 15162 8084
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14830 6160 14886 6216
rect 15382 7656 15438 7712
rect 14554 5092 14610 5128
rect 14554 5072 14556 5092
rect 14556 5072 14608 5092
rect 14608 5072 14610 5092
rect 14462 4700 14464 4720
rect 14464 4700 14516 4720
rect 14516 4700 14518 4720
rect 14462 4664 14518 4700
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 15382 4392 15438 4448
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 16118 12552 16174 12608
rect 15934 11620 15990 11656
rect 15934 11600 15936 11620
rect 15936 11600 15988 11620
rect 15988 11600 15990 11620
rect 16670 20460 16726 20496
rect 16670 20440 16672 20460
rect 16672 20440 16724 20460
rect 16724 20440 16726 20460
rect 18050 24112 18106 24168
rect 18786 24656 18842 24712
rect 18234 24248 18290 24304
rect 18234 19352 18290 19408
rect 18142 18808 18198 18864
rect 16762 18672 16818 18728
rect 17130 18672 17186 18728
rect 16394 17040 16450 17096
rect 17406 17332 17462 17368
rect 17406 17312 17408 17332
rect 17408 17312 17460 17332
rect 17460 17312 17462 17332
rect 16854 15680 16910 15736
rect 17314 16532 17316 16552
rect 17316 16532 17368 16552
rect 17368 16532 17370 16552
rect 17314 16496 17370 16532
rect 16670 14320 16726 14376
rect 17498 14728 17554 14784
rect 16762 13932 16818 13968
rect 16762 13912 16764 13932
rect 16764 13912 16816 13932
rect 16816 13912 16818 13932
rect 16762 12708 16818 12744
rect 16762 12688 16764 12708
rect 16764 12688 16816 12708
rect 16816 12688 16818 12708
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 20258 24656 20314 24712
rect 20442 24656 20498 24712
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 20442 23976 20498 24032
rect 18418 17856 18474 17912
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 20166 23296 20222 23352
rect 20166 22072 20222 22128
rect 20902 23180 20958 23216
rect 20902 23160 20904 23180
rect 20904 23160 20956 23180
rect 20956 23160 20958 23180
rect 23294 24404 23350 24440
rect 23294 24384 23296 24404
rect 23296 24384 23348 24404
rect 23348 24384 23350 24404
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24766 24384 24822 24440
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 27066 24656 27122 24712
rect 25962 24248 26018 24304
rect 24214 23704 24270 23760
rect 22466 22516 22468 22536
rect 22468 22516 22520 22536
rect 22520 22516 22522 22536
rect 22466 22480 22522 22516
rect 22374 21392 22430 21448
rect 21362 20848 21418 20904
rect 20810 20304 20866 20360
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 23294 19896 23350 19952
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 27618 18672 27674 18728
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 20074 18128 20130 18184
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 20626 15408 20682 15464
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19430 13912 19486 13968
rect 18694 13812 18696 13832
rect 18696 13812 18748 13832
rect 18748 13812 18750 13832
rect 18694 13776 18750 13812
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 18418 12588 18420 12608
rect 18420 12588 18472 12608
rect 18472 12588 18474 12608
rect 17590 11056 17646 11112
rect 18050 11092 18052 11112
rect 18052 11092 18104 11112
rect 18104 11092 18106 11112
rect 18050 11056 18106 11092
rect 18142 10648 18198 10704
rect 16854 9152 16910 9208
rect 16118 7112 16174 7168
rect 16210 6840 16266 6896
rect 15934 5344 15990 5400
rect 15750 4528 15806 4584
rect 15750 3848 15806 3904
rect 15842 2508 15898 2544
rect 15842 2488 15844 2508
rect 15844 2488 15896 2508
rect 15896 2488 15898 2508
rect 16670 6432 16726 6488
rect 16762 6060 16764 6080
rect 16764 6060 16816 6080
rect 16816 6060 16818 6080
rect 16762 6024 16818 6060
rect 16394 4800 16450 4856
rect 16302 4528 16358 4584
rect 16762 5480 16818 5536
rect 16762 3712 16818 3768
rect 16302 3476 16304 3496
rect 16304 3476 16356 3496
rect 16356 3476 16358 3496
rect 16302 3440 16358 3476
rect 16210 3032 16266 3088
rect 16026 2080 16082 2136
rect 15750 1808 15806 1864
rect 16762 3304 16818 3360
rect 17406 10104 17462 10160
rect 17958 9424 18014 9480
rect 17222 8744 17278 8800
rect 17682 8608 17738 8664
rect 17406 8064 17462 8120
rect 17314 6840 17370 6896
rect 17958 8200 18014 8256
rect 17958 6976 18014 7032
rect 17958 6568 18014 6624
rect 17682 4120 17738 4176
rect 18050 5616 18106 5672
rect 18050 5364 18106 5400
rect 18050 5344 18052 5364
rect 18052 5344 18104 5364
rect 18104 5344 18106 5364
rect 18142 4392 18198 4448
rect 17866 3848 17922 3904
rect 17406 3440 17462 3496
rect 17038 2388 17040 2408
rect 17040 2388 17092 2408
rect 17092 2388 17094 2408
rect 17038 2352 17094 2388
rect 17314 2372 17370 2408
rect 17314 2352 17316 2372
rect 17316 2352 17368 2372
rect 17368 2352 17370 2372
rect 17590 3032 17646 3088
rect 17958 2896 18014 2952
rect 17866 2760 17922 2816
rect 18418 12552 18474 12588
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 18418 10532 18474 10568
rect 18418 10512 18420 10532
rect 18420 10512 18472 10532
rect 18472 10512 18474 10532
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 18970 10004 18972 10024
rect 18972 10004 19024 10024
rect 19024 10004 19026 10024
rect 18970 9968 19026 10004
rect 18878 9288 18934 9344
rect 18694 6840 18750 6896
rect 18602 5072 18658 5128
rect 18510 4800 18566 4856
rect 19982 9696 20038 9752
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19430 9152 19486 9208
rect 19614 8336 19670 8392
rect 19430 7928 19486 7984
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 20074 8900 20130 8936
rect 20074 8880 20076 8900
rect 20076 8880 20128 8900
rect 20128 8880 20130 8900
rect 20258 8744 20314 8800
rect 19614 7792 19670 7848
rect 18970 7248 19026 7304
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19982 6432 20038 6488
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19338 5208 19394 5264
rect 19062 4972 19064 4992
rect 19064 4972 19116 4992
rect 19116 4972 19118 4992
rect 19062 4936 19118 4972
rect 19154 4684 19210 4720
rect 19154 4664 19156 4684
rect 19156 4664 19208 4684
rect 19208 4664 19210 4684
rect 18510 4120 18566 4176
rect 18050 2524 18052 2544
rect 18052 2524 18104 2544
rect 18104 2524 18106 2544
rect 18050 2488 18106 2524
rect 18326 1944 18382 2000
rect 19338 4392 19394 4448
rect 19522 5480 19578 5536
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19430 4120 19486 4176
rect 20166 4528 20222 4584
rect 20350 7656 20406 7712
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 25502 15000 25558 15056
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24398 13912 24454 13968
rect 24122 13812 24124 13832
rect 24124 13812 24176 13832
rect 24176 13812 24178 13832
rect 24122 13776 24178 13812
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 21914 12824 21970 12880
rect 20810 12144 20866 12200
rect 20718 11056 20774 11112
rect 20442 6452 20498 6488
rect 20442 6432 20444 6452
rect 20444 6432 20496 6452
rect 20496 6432 20498 6452
rect 20994 8608 21050 8664
rect 21178 8492 21234 8528
rect 21178 8472 21180 8492
rect 21180 8472 21232 8492
rect 21232 8472 21234 8492
rect 20994 7404 21050 7440
rect 20994 7384 20996 7404
rect 20996 7384 21048 7404
rect 21048 7384 21050 7404
rect 20994 6840 21050 6896
rect 21178 6740 21180 6760
rect 21180 6740 21232 6760
rect 21232 6740 21234 6760
rect 21178 6704 21234 6740
rect 21546 5752 21602 5808
rect 21178 5616 21234 5672
rect 20074 3884 20076 3904
rect 20076 3884 20128 3904
rect 20128 3884 20130 3904
rect 19154 3596 19210 3632
rect 19154 3576 19156 3596
rect 19156 3576 19208 3596
rect 19208 3576 19210 3596
rect 19338 3712 19394 3768
rect 20074 3848 20130 3884
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19522 3576 19578 3632
rect 19522 3032 19578 3088
rect 19522 2896 19578 2952
rect 19338 2624 19394 2680
rect 19062 2488 19118 2544
rect 19062 1536 19118 1592
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 20166 2624 20222 2680
rect 19890 2080 19946 2136
rect 20718 3168 20774 3224
rect 20718 2252 20720 2272
rect 20720 2252 20772 2272
rect 20772 2252 20774 2272
rect 20718 2216 20774 2252
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 21914 4664 21970 4720
rect 22006 3440 22062 3496
rect 21822 3340 21824 3360
rect 21824 3340 21876 3360
rect 21876 3340 21878 3360
rect 21822 3304 21878 3340
rect 21178 2508 21234 2544
rect 21178 2488 21180 2508
rect 21180 2488 21232 2508
rect 21232 2488 21234 2508
rect 22190 2896 22246 2952
rect 22006 2760 22062 2816
rect 22098 2644 22154 2680
rect 22098 2624 22100 2644
rect 22100 2624 22152 2644
rect 22152 2624 22154 2644
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 22374 5072 22430 5128
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24122 3712 24178 3768
rect 23478 1536 23534 1592
rect 24030 1808 24086 1864
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24766 2760 24822 2816
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 26514 3848 26570 3904
rect 25962 3032 26018 3088
rect 27618 3576 27674 3632
rect 27066 2352 27122 2408
<< metal3 >>
rect 0 27706 480 27736
rect 3509 27706 3575 27709
rect 0 27704 3575 27706
rect 0 27648 3514 27704
rect 3570 27648 3575 27704
rect 0 27646 3575 27648
rect 0 27616 480 27646
rect 3509 27643 3575 27646
rect 0 27162 480 27192
rect 3509 27162 3575 27165
rect 0 27160 3575 27162
rect 0 27104 3514 27160
rect 3570 27104 3575 27160
rect 0 27102 3575 27104
rect 0 27072 480 27102
rect 3509 27099 3575 27102
rect 0 26618 480 26648
rect 4061 26618 4127 26621
rect 0 26616 4127 26618
rect 0 26560 4066 26616
rect 4122 26560 4127 26616
rect 0 26558 4127 26560
rect 0 26528 480 26558
rect 4061 26555 4127 26558
rect 0 25938 480 25968
rect 4061 25938 4127 25941
rect 0 25936 4127 25938
rect 0 25880 4066 25936
rect 4122 25880 4127 25936
rect 0 25878 4127 25880
rect 0 25848 480 25878
rect 4061 25875 4127 25878
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 0 25394 480 25424
rect 3325 25394 3391 25397
rect 0 25392 3391 25394
rect 0 25336 3330 25392
rect 3386 25336 3391 25392
rect 0 25334 3391 25336
rect 0 25304 480 25334
rect 3325 25331 3391 25334
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 0 24850 480 24880
rect 4061 24850 4127 24853
rect 0 24848 4127 24850
rect 0 24792 4066 24848
rect 4122 24792 4127 24848
rect 0 24790 4127 24792
rect 0 24760 480 24790
rect 4061 24787 4127 24790
rect 1761 24714 1827 24717
rect 6913 24714 6979 24717
rect 1761 24712 6979 24714
rect 1761 24656 1766 24712
rect 1822 24656 6918 24712
rect 6974 24656 6979 24712
rect 1761 24654 6979 24656
rect 1761 24651 1827 24654
rect 6913 24651 6979 24654
rect 12065 24714 12131 24717
rect 13353 24714 13419 24717
rect 12065 24712 13419 24714
rect 12065 24656 12070 24712
rect 12126 24656 13358 24712
rect 13414 24656 13419 24712
rect 12065 24654 13419 24656
rect 12065 24651 12131 24654
rect 13353 24651 13419 24654
rect 18781 24714 18847 24717
rect 20253 24714 20319 24717
rect 18781 24712 20319 24714
rect 18781 24656 18786 24712
rect 18842 24656 20258 24712
rect 20314 24656 20319 24712
rect 18781 24654 20319 24656
rect 18781 24651 18847 24654
rect 20253 24651 20319 24654
rect 20437 24714 20503 24717
rect 27061 24714 27127 24717
rect 20437 24712 27127 24714
rect 20437 24656 20442 24712
rect 20498 24656 27066 24712
rect 27122 24656 27127 24712
rect 20437 24654 27127 24656
rect 20437 24651 20503 24654
rect 27061 24651 27127 24654
rect 1945 24578 2011 24581
rect 1945 24576 6194 24578
rect 1945 24520 1950 24576
rect 2006 24520 6194 24576
rect 1945 24518 6194 24520
rect 1945 24515 2011 24518
rect 6134 24442 6194 24518
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 7741 24442 7807 24445
rect 8845 24442 8911 24445
rect 6134 24440 8911 24442
rect 6134 24384 7746 24440
rect 7802 24384 8850 24440
rect 8906 24384 8911 24440
rect 6134 24382 8911 24384
rect 7741 24379 7807 24382
rect 8845 24379 8911 24382
rect 23289 24442 23355 24445
rect 24761 24442 24827 24445
rect 23289 24440 24827 24442
rect 23289 24384 23294 24440
rect 23350 24384 24766 24440
rect 24822 24384 24827 24440
rect 23289 24382 24827 24384
rect 23289 24379 23355 24382
rect 24761 24379 24827 24382
rect 1761 24306 1827 24309
rect 7833 24306 7899 24309
rect 1761 24304 7899 24306
rect 1761 24248 1766 24304
rect 1822 24248 7838 24304
rect 7894 24248 7899 24304
rect 1761 24246 7899 24248
rect 1761 24243 1827 24246
rect 7833 24243 7899 24246
rect 9673 24306 9739 24309
rect 16389 24306 16455 24309
rect 9673 24304 16455 24306
rect 9673 24248 9678 24304
rect 9734 24248 16394 24304
rect 16450 24248 16455 24304
rect 9673 24246 16455 24248
rect 9673 24243 9739 24246
rect 16389 24243 16455 24246
rect 18229 24306 18295 24309
rect 25957 24306 26023 24309
rect 18229 24304 26023 24306
rect 18229 24248 18234 24304
rect 18290 24248 25962 24304
rect 26018 24248 26023 24304
rect 18229 24246 26023 24248
rect 18229 24243 18295 24246
rect 25957 24243 26023 24246
rect 0 24170 480 24200
rect 3509 24170 3575 24173
rect 0 24168 3575 24170
rect 0 24112 3514 24168
rect 3570 24112 3575 24168
rect 0 24110 3575 24112
rect 0 24080 480 24110
rect 3509 24107 3575 24110
rect 8661 24170 8727 24173
rect 11237 24170 11303 24173
rect 18045 24170 18111 24173
rect 8661 24168 11303 24170
rect 8661 24112 8666 24168
rect 8722 24112 11242 24168
rect 11298 24112 11303 24168
rect 8661 24110 11303 24112
rect 8661 24107 8727 24110
rect 11237 24107 11303 24110
rect 11470 24168 18111 24170
rect 11470 24112 18050 24168
rect 18106 24112 18111 24168
rect 11470 24110 18111 24112
rect 6913 24034 6979 24037
rect 11470 24034 11530 24110
rect 18045 24107 18111 24110
rect 6913 24032 11530 24034
rect 6913 23976 6918 24032
rect 6974 23976 11530 24032
rect 6913 23974 11530 23976
rect 16481 24034 16547 24037
rect 20437 24034 20503 24037
rect 16481 24032 20503 24034
rect 16481 23976 16486 24032
rect 16542 23976 20442 24032
rect 20498 23976 20503 24032
rect 16481 23974 20503 23976
rect 6913 23971 6979 23974
rect 16481 23971 16547 23974
rect 20437 23971 20503 23974
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 2405 23898 2471 23901
rect 5165 23898 5231 23901
rect 2405 23896 5231 23898
rect 2405 23840 2410 23896
rect 2466 23840 5170 23896
rect 5226 23840 5231 23896
rect 2405 23838 5231 23840
rect 2405 23835 2471 23838
rect 5165 23835 5231 23838
rect 9029 23898 9095 23901
rect 11053 23898 11119 23901
rect 9029 23896 11119 23898
rect 9029 23840 9034 23896
rect 9090 23840 11058 23896
rect 11114 23840 11119 23896
rect 9029 23838 11119 23840
rect 9029 23835 9095 23838
rect 11053 23835 11119 23838
rect 11697 23898 11763 23901
rect 14365 23898 14431 23901
rect 11697 23896 14431 23898
rect 11697 23840 11702 23896
rect 11758 23840 14370 23896
rect 14426 23840 14431 23896
rect 11697 23838 14431 23840
rect 11697 23835 11763 23838
rect 14365 23835 14431 23838
rect 2681 23762 2747 23765
rect 9489 23762 9555 23765
rect 2681 23760 9555 23762
rect 2681 23704 2686 23760
rect 2742 23704 9494 23760
rect 9550 23704 9555 23760
rect 2681 23702 9555 23704
rect 2681 23699 2747 23702
rect 9489 23699 9555 23702
rect 12617 23762 12683 23765
rect 24209 23762 24275 23765
rect 12617 23760 24275 23762
rect 12617 23704 12622 23760
rect 12678 23704 24214 23760
rect 24270 23704 24275 23760
rect 12617 23702 24275 23704
rect 12617 23699 12683 23702
rect 24209 23699 24275 23702
rect 0 23626 480 23656
rect 4061 23626 4127 23629
rect 0 23624 4127 23626
rect 0 23568 4066 23624
rect 4122 23568 4127 23624
rect 0 23566 4127 23568
rect 0 23536 480 23566
rect 4061 23563 4127 23566
rect 6177 23626 6243 23629
rect 6177 23624 10794 23626
rect 6177 23568 6182 23624
rect 6238 23568 10794 23624
rect 6177 23566 10794 23568
rect 6177 23563 6243 23566
rect 10734 23490 10794 23566
rect 13445 23490 13511 23493
rect 10734 23488 13511 23490
rect 10734 23432 13450 23488
rect 13506 23432 13511 23488
rect 10734 23430 13511 23432
rect 13445 23427 13511 23430
rect 13721 23490 13787 23493
rect 15561 23490 15627 23493
rect 13721 23488 15627 23490
rect 13721 23432 13726 23488
rect 13782 23432 15566 23488
rect 15622 23432 15627 23488
rect 13721 23430 15627 23432
rect 13721 23427 13787 23430
rect 15561 23427 15627 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 4981 23354 5047 23357
rect 6545 23354 6611 23357
rect 4981 23352 6611 23354
rect 4981 23296 4986 23352
rect 5042 23296 6550 23352
rect 6606 23296 6611 23352
rect 4981 23294 6611 23296
rect 4981 23291 5047 23294
rect 6545 23291 6611 23294
rect 6729 23354 6795 23357
rect 9673 23354 9739 23357
rect 6729 23352 9739 23354
rect 6729 23296 6734 23352
rect 6790 23296 9678 23352
rect 9734 23296 9739 23352
rect 6729 23294 9739 23296
rect 6729 23291 6795 23294
rect 9673 23291 9739 23294
rect 20161 23354 20227 23357
rect 27520 23354 28000 23384
rect 20161 23352 28000 23354
rect 20161 23296 20166 23352
rect 20222 23296 28000 23352
rect 20161 23294 28000 23296
rect 20161 23291 20227 23294
rect 27520 23264 28000 23294
rect 5809 23218 5875 23221
rect 2638 23216 5875 23218
rect 2638 23160 5814 23216
rect 5870 23160 5875 23216
rect 2638 23158 5875 23160
rect 0 23082 480 23112
rect 2638 23082 2698 23158
rect 5809 23155 5875 23158
rect 8937 23218 9003 23221
rect 20897 23218 20963 23221
rect 8937 23216 20963 23218
rect 8937 23160 8942 23216
rect 8998 23160 20902 23216
rect 20958 23160 20963 23216
rect 8937 23158 20963 23160
rect 8937 23155 9003 23158
rect 20897 23155 20963 23158
rect 0 23022 2698 23082
rect 6453 23082 6519 23085
rect 6913 23082 6979 23085
rect 6453 23080 6979 23082
rect 6453 23024 6458 23080
rect 6514 23024 6918 23080
rect 6974 23024 6979 23080
rect 6453 23022 6979 23024
rect 0 22992 480 23022
rect 6453 23019 6519 23022
rect 6913 23019 6979 23022
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 3601 22674 3667 22677
rect 6269 22674 6335 22677
rect 11237 22674 11303 22677
rect 3601 22672 11303 22674
rect 3601 22616 3606 22672
rect 3662 22616 6274 22672
rect 6330 22616 11242 22672
rect 11298 22616 11303 22672
rect 3601 22614 11303 22616
rect 3601 22611 3667 22614
rect 6269 22611 6335 22614
rect 11237 22611 11303 22614
rect 13905 22674 13971 22677
rect 16849 22674 16915 22677
rect 13905 22672 16915 22674
rect 13905 22616 13910 22672
rect 13966 22616 16854 22672
rect 16910 22616 16915 22672
rect 13905 22614 16915 22616
rect 13905 22611 13971 22614
rect 16849 22611 16915 22614
rect 0 22538 480 22568
rect 3969 22538 4035 22541
rect 0 22536 4035 22538
rect 0 22480 3974 22536
rect 4030 22480 4035 22536
rect 0 22478 4035 22480
rect 0 22448 480 22478
rect 3969 22475 4035 22478
rect 8477 22538 8543 22541
rect 22461 22538 22527 22541
rect 8477 22536 22527 22538
rect 8477 22480 8482 22536
rect 8538 22480 22466 22536
rect 22522 22480 22527 22536
rect 8477 22478 22527 22480
rect 8477 22475 8543 22478
rect 22461 22475 22527 22478
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 8017 22130 8083 22133
rect 11053 22130 11119 22133
rect 8017 22128 11119 22130
rect 8017 22072 8022 22128
rect 8078 22072 11058 22128
rect 11114 22072 11119 22128
rect 8017 22070 11119 22072
rect 8017 22067 8083 22070
rect 11053 22067 11119 22070
rect 11237 22130 11303 22133
rect 20161 22130 20227 22133
rect 11237 22128 20227 22130
rect 11237 22072 11242 22128
rect 11298 22072 20166 22128
rect 20222 22072 20227 22128
rect 11237 22070 20227 22072
rect 11237 22067 11303 22070
rect 20161 22067 20227 22070
rect 1577 21994 1643 21997
rect 15377 21994 15443 21997
rect 1577 21992 15443 21994
rect 1577 21936 1582 21992
rect 1638 21936 15382 21992
rect 15438 21936 15443 21992
rect 1577 21934 15443 21936
rect 1577 21931 1643 21934
rect 15377 21931 15443 21934
rect 0 21858 480 21888
rect 3141 21858 3207 21861
rect 0 21856 3207 21858
rect 0 21800 3146 21856
rect 3202 21800 3207 21856
rect 0 21798 3207 21800
rect 0 21768 480 21798
rect 3141 21795 3207 21798
rect 10225 21858 10291 21861
rect 13997 21858 14063 21861
rect 10225 21856 14063 21858
rect 10225 21800 10230 21856
rect 10286 21800 14002 21856
rect 14058 21800 14063 21856
rect 10225 21798 14063 21800
rect 10225 21795 10291 21798
rect 13997 21795 14063 21798
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 2037 21586 2103 21589
rect 6085 21586 6151 21589
rect 2037 21584 6151 21586
rect 2037 21528 2042 21584
rect 2098 21528 6090 21584
rect 6146 21528 6151 21584
rect 2037 21526 6151 21528
rect 2037 21523 2103 21526
rect 6085 21523 6151 21526
rect 6269 21586 6335 21589
rect 12157 21586 12223 21589
rect 6269 21584 12223 21586
rect 6269 21528 6274 21584
rect 6330 21528 12162 21584
rect 12218 21528 12223 21584
rect 6269 21526 12223 21528
rect 6269 21523 6335 21526
rect 12157 21523 12223 21526
rect 2129 21450 2195 21453
rect 7649 21450 7715 21453
rect 2129 21448 7715 21450
rect 2129 21392 2134 21448
rect 2190 21392 7654 21448
rect 7710 21392 7715 21448
rect 2129 21390 7715 21392
rect 2129 21387 2195 21390
rect 7649 21387 7715 21390
rect 14825 21450 14891 21453
rect 22369 21450 22435 21453
rect 14825 21448 22435 21450
rect 14825 21392 14830 21448
rect 14886 21392 22374 21448
rect 22430 21392 22435 21448
rect 14825 21390 22435 21392
rect 14825 21387 14891 21390
rect 22369 21387 22435 21390
rect 0 21314 480 21344
rect 3233 21314 3299 21317
rect 0 21312 3299 21314
rect 0 21256 3238 21312
rect 3294 21256 3299 21312
rect 0 21254 3299 21256
rect 0 21224 480 21254
rect 3233 21251 3299 21254
rect 4521 21314 4587 21317
rect 9765 21314 9831 21317
rect 4521 21312 9831 21314
rect 4521 21256 4526 21312
rect 4582 21256 9770 21312
rect 9826 21256 9831 21312
rect 4521 21254 9831 21256
rect 4521 21251 4587 21254
rect 9765 21251 9831 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 9121 21178 9187 21181
rect 5030 21176 9187 21178
rect 5030 21120 9126 21176
rect 9182 21120 9187 21176
rect 5030 21118 9187 21120
rect 289 21042 355 21045
rect 3325 21042 3391 21045
rect 5030 21042 5090 21118
rect 9121 21115 9187 21118
rect 289 21040 5090 21042
rect 289 20984 294 21040
rect 350 20984 3330 21040
rect 3386 20984 5090 21040
rect 289 20982 5090 20984
rect 5165 21042 5231 21045
rect 6177 21042 6243 21045
rect 5165 21040 6243 21042
rect 5165 20984 5170 21040
rect 5226 20984 6182 21040
rect 6238 20984 6243 21040
rect 5165 20982 6243 20984
rect 289 20979 355 20982
rect 3325 20979 3391 20982
rect 5165 20979 5231 20982
rect 6177 20979 6243 20982
rect 1669 20906 1735 20909
rect 12525 20906 12591 20909
rect 1669 20904 12591 20906
rect 1669 20848 1674 20904
rect 1730 20848 12530 20904
rect 12586 20848 12591 20904
rect 1669 20846 12591 20848
rect 1669 20843 1735 20846
rect 12525 20843 12591 20846
rect 14733 20906 14799 20909
rect 21357 20906 21423 20909
rect 14733 20904 21423 20906
rect 14733 20848 14738 20904
rect 14794 20848 21362 20904
rect 21418 20848 21423 20904
rect 14733 20846 21423 20848
rect 14733 20843 14799 20846
rect 21357 20843 21423 20846
rect 0 20770 480 20800
rect 2865 20770 2931 20773
rect 0 20768 2931 20770
rect 0 20712 2870 20768
rect 2926 20712 2931 20768
rect 0 20710 2931 20712
rect 0 20680 480 20710
rect 2865 20707 2931 20710
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 9489 20634 9555 20637
rect 14089 20634 14155 20637
rect 9489 20632 14155 20634
rect 9489 20576 9494 20632
rect 9550 20576 14094 20632
rect 14150 20576 14155 20632
rect 9489 20574 14155 20576
rect 9489 20571 9555 20574
rect 14089 20571 14155 20574
rect 1761 20498 1827 20501
rect 10041 20498 10107 20501
rect 1761 20496 10107 20498
rect 1761 20440 1766 20496
rect 1822 20440 10046 20496
rect 10102 20440 10107 20496
rect 1761 20438 10107 20440
rect 1761 20435 1827 20438
rect 10041 20435 10107 20438
rect 12801 20498 12867 20501
rect 16665 20498 16731 20501
rect 12801 20496 16731 20498
rect 12801 20440 12806 20496
rect 12862 20440 16670 20496
rect 16726 20440 16731 20496
rect 12801 20438 16731 20440
rect 12801 20435 12867 20438
rect 16665 20435 16731 20438
rect 2497 20362 2563 20365
rect 7005 20362 7071 20365
rect 2497 20360 7071 20362
rect 2497 20304 2502 20360
rect 2558 20304 7010 20360
rect 7066 20304 7071 20360
rect 2497 20302 7071 20304
rect 2497 20299 2563 20302
rect 7005 20299 7071 20302
rect 11789 20362 11855 20365
rect 20805 20362 20871 20365
rect 11789 20360 20871 20362
rect 11789 20304 11794 20360
rect 11850 20304 20810 20360
rect 20866 20304 20871 20360
rect 11789 20302 20871 20304
rect 11789 20299 11855 20302
rect 20805 20299 20871 20302
rect 2681 20226 2747 20229
rect 4797 20226 4863 20229
rect 2681 20224 4863 20226
rect 2681 20168 2686 20224
rect 2742 20168 4802 20224
rect 4858 20168 4863 20224
rect 2681 20166 4863 20168
rect 2681 20163 2747 20166
rect 4797 20163 4863 20166
rect 6545 20226 6611 20229
rect 9121 20226 9187 20229
rect 6545 20224 9187 20226
rect 6545 20168 6550 20224
rect 6606 20168 9126 20224
rect 9182 20168 9187 20224
rect 6545 20166 9187 20168
rect 6545 20163 6611 20166
rect 9121 20163 9187 20166
rect 10277 20160 10597 20161
rect 0 20090 480 20120
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 8385 20090 8451 20093
rect 0 20088 8451 20090
rect 0 20032 8390 20088
rect 8446 20032 8451 20088
rect 0 20030 8451 20032
rect 0 20000 480 20030
rect 8385 20027 8451 20030
rect 13169 19954 13235 19957
rect 23289 19954 23355 19957
rect 13169 19952 23355 19954
rect 13169 19896 13174 19952
rect 13230 19896 23294 19952
rect 23350 19896 23355 19952
rect 13169 19894 23355 19896
rect 13169 19891 13235 19894
rect 23289 19891 23355 19894
rect 2221 19818 2287 19821
rect 8017 19818 8083 19821
rect 2221 19816 8083 19818
rect 2221 19760 2226 19816
rect 2282 19760 8022 19816
rect 8078 19760 8083 19816
rect 2221 19758 8083 19760
rect 2221 19755 2287 19758
rect 8017 19755 8083 19758
rect 8845 19818 8911 19821
rect 12893 19818 12959 19821
rect 8845 19816 12959 19818
rect 8845 19760 8850 19816
rect 8906 19760 12898 19816
rect 12954 19760 12959 19816
rect 8845 19758 12959 19760
rect 8845 19755 8911 19758
rect 12893 19755 12959 19758
rect 14273 19818 14339 19821
rect 16205 19818 16271 19821
rect 14273 19816 16271 19818
rect 14273 19760 14278 19816
rect 14334 19760 16210 19816
rect 16266 19760 16271 19816
rect 14273 19758 16271 19760
rect 14273 19755 14339 19758
rect 11973 19682 12039 19685
rect 10734 19680 12039 19682
rect 10734 19624 11978 19680
rect 12034 19624 12039 19680
rect 10734 19622 12039 19624
rect 5610 19616 5930 19617
rect 0 19546 480 19576
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 3049 19546 3115 19549
rect 0 19544 3115 19546
rect 0 19488 3054 19544
rect 3110 19488 3115 19544
rect 0 19486 3115 19488
rect 0 19456 480 19486
rect 3049 19483 3115 19486
rect 6637 19546 6703 19549
rect 9489 19546 9555 19549
rect 10734 19546 10794 19622
rect 11973 19619 12039 19622
rect 6637 19544 10794 19546
rect 6637 19488 6642 19544
rect 6698 19488 9494 19544
rect 9550 19488 10794 19544
rect 6637 19486 10794 19488
rect 10869 19546 10935 19549
rect 11237 19546 11303 19549
rect 14414 19546 14474 19758
rect 16205 19755 16271 19758
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 10869 19544 14474 19546
rect 10869 19488 10874 19544
rect 10930 19488 11242 19544
rect 11298 19488 14474 19544
rect 10869 19486 14474 19488
rect 6637 19483 6703 19486
rect 9489 19483 9555 19486
rect 10869 19483 10935 19486
rect 11237 19483 11303 19486
rect 9213 19410 9279 19413
rect 12801 19410 12867 19413
rect 9213 19408 12867 19410
rect 9213 19352 9218 19408
rect 9274 19352 12806 19408
rect 12862 19352 12867 19408
rect 9213 19350 12867 19352
rect 9213 19347 9279 19350
rect 12801 19347 12867 19350
rect 13353 19410 13419 19413
rect 18229 19410 18295 19413
rect 13353 19408 18295 19410
rect 13353 19352 13358 19408
rect 13414 19352 18234 19408
rect 18290 19352 18295 19408
rect 13353 19350 18295 19352
rect 13353 19347 13419 19350
rect 18229 19347 18295 19350
rect 1485 19274 1551 19277
rect 11145 19274 11211 19277
rect 12985 19274 13051 19277
rect 1485 19272 10794 19274
rect 1485 19216 1490 19272
rect 1546 19216 10794 19272
rect 1485 19214 10794 19216
rect 1485 19211 1551 19214
rect 4245 19138 4311 19141
rect 7005 19138 7071 19141
rect 4245 19136 7071 19138
rect 4245 19080 4250 19136
rect 4306 19080 7010 19136
rect 7066 19080 7071 19136
rect 4245 19078 7071 19080
rect 10734 19138 10794 19214
rect 11145 19272 13051 19274
rect 11145 19216 11150 19272
rect 11206 19216 12990 19272
rect 13046 19216 13051 19272
rect 11145 19214 13051 19216
rect 11145 19211 11211 19214
rect 12985 19211 13051 19214
rect 13537 19274 13603 19277
rect 14641 19274 14707 19277
rect 13537 19272 14707 19274
rect 13537 19216 13542 19272
rect 13598 19216 14646 19272
rect 14702 19216 14707 19272
rect 13537 19214 14707 19216
rect 13537 19211 13603 19214
rect 14641 19211 14707 19214
rect 13445 19138 13511 19141
rect 10734 19136 13511 19138
rect 10734 19080 13450 19136
rect 13506 19080 13511 19136
rect 10734 19078 13511 19080
rect 4245 19075 4311 19078
rect 7005 19075 7071 19078
rect 13445 19075 13511 19078
rect 13905 19138 13971 19141
rect 15653 19138 15719 19141
rect 13905 19136 15719 19138
rect 13905 19080 13910 19136
rect 13966 19080 15658 19136
rect 15714 19080 15719 19136
rect 13905 19078 15719 19080
rect 13905 19075 13971 19078
rect 15653 19075 15719 19078
rect 10277 19072 10597 19073
rect 0 19002 480 19032
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 3233 19002 3299 19005
rect 0 19000 3299 19002
rect 0 18944 3238 19000
rect 3294 18944 3299 19000
rect 0 18942 3299 18944
rect 0 18912 480 18942
rect 3233 18939 3299 18942
rect 8201 19002 8267 19005
rect 10133 19002 10199 19005
rect 8201 19000 10199 19002
rect 8201 18944 8206 19000
rect 8262 18944 10138 19000
rect 10194 18944 10199 19000
rect 8201 18942 10199 18944
rect 8201 18939 8267 18942
rect 10133 18939 10199 18942
rect 11237 19002 11303 19005
rect 12249 19002 12315 19005
rect 14733 19002 14799 19005
rect 11237 19000 14799 19002
rect 11237 18944 11242 19000
rect 11298 18944 12254 19000
rect 12310 18944 14738 19000
rect 14794 18944 14799 19000
rect 11237 18942 14799 18944
rect 11237 18939 11303 18942
rect 12249 18939 12315 18942
rect 14733 18939 14799 18942
rect 8845 18866 8911 18869
rect 12617 18866 12683 18869
rect 8845 18864 12683 18866
rect 8845 18808 8850 18864
rect 8906 18808 12622 18864
rect 12678 18808 12683 18864
rect 8845 18806 12683 18808
rect 8845 18803 8911 18806
rect 12617 18803 12683 18806
rect 12985 18866 13051 18869
rect 18137 18866 18203 18869
rect 12985 18864 18203 18866
rect 12985 18808 12990 18864
rect 13046 18808 18142 18864
rect 18198 18808 18203 18864
rect 12985 18806 18203 18808
rect 12985 18803 13051 18806
rect 18137 18803 18203 18806
rect 6545 18730 6611 18733
rect 16757 18730 16823 18733
rect 6545 18728 16823 18730
rect 6545 18672 6550 18728
rect 6606 18672 16762 18728
rect 16818 18672 16823 18728
rect 6545 18670 16823 18672
rect 6545 18667 6611 18670
rect 16757 18667 16823 18670
rect 17125 18730 17191 18733
rect 27613 18730 27679 18733
rect 17125 18728 27679 18730
rect 17125 18672 17130 18728
rect 17186 18672 27618 18728
rect 27674 18672 27679 18728
rect 17125 18670 27679 18672
rect 17125 18667 17191 18670
rect 27613 18667 27679 18670
rect 8845 18594 8911 18597
rect 11237 18594 11303 18597
rect 8845 18592 11303 18594
rect 8845 18536 8850 18592
rect 8906 18536 11242 18592
rect 11298 18536 11303 18592
rect 8845 18534 11303 18536
rect 8845 18531 8911 18534
rect 11237 18531 11303 18534
rect 5610 18528 5930 18529
rect 0 18458 480 18488
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 5441 18458 5507 18461
rect 0 18456 5507 18458
rect 0 18400 5446 18456
rect 5502 18400 5507 18456
rect 0 18398 5507 18400
rect 0 18368 480 18398
rect 5441 18395 5507 18398
rect 6821 18458 6887 18461
rect 9949 18458 10015 18461
rect 6821 18456 10015 18458
rect 6821 18400 6826 18456
rect 6882 18400 9954 18456
rect 10010 18400 10015 18456
rect 6821 18398 10015 18400
rect 6821 18395 6887 18398
rect 9949 18395 10015 18398
rect 8753 18322 8819 18325
rect 13169 18322 13235 18325
rect 13445 18322 13511 18325
rect 8753 18320 13511 18322
rect 8753 18264 8758 18320
rect 8814 18264 13174 18320
rect 13230 18264 13450 18320
rect 13506 18264 13511 18320
rect 8753 18262 13511 18264
rect 8753 18259 8819 18262
rect 13169 18259 13235 18262
rect 13445 18259 13511 18262
rect 7649 18186 7715 18189
rect 8477 18186 8543 18189
rect 7649 18184 8543 18186
rect 7649 18128 7654 18184
rect 7710 18128 8482 18184
rect 8538 18128 8543 18184
rect 7649 18126 8543 18128
rect 7649 18123 7715 18126
rect 8477 18123 8543 18126
rect 15469 18186 15535 18189
rect 20069 18186 20135 18189
rect 15469 18184 20135 18186
rect 15469 18128 15474 18184
rect 15530 18128 20074 18184
rect 20130 18128 20135 18184
rect 15469 18126 20135 18128
rect 15469 18123 15535 18126
rect 20069 18123 20135 18126
rect 2589 18050 2655 18053
rect 4613 18050 4679 18053
rect 2589 18048 4679 18050
rect 2589 17992 2594 18048
rect 2650 17992 4618 18048
rect 4674 17992 4679 18048
rect 2589 17990 4679 17992
rect 2589 17987 2655 17990
rect 4613 17987 4679 17990
rect 7741 18050 7807 18053
rect 8937 18050 9003 18053
rect 7741 18048 9003 18050
rect 7741 17992 7746 18048
rect 7802 17992 8942 18048
rect 8998 17992 9003 18048
rect 7741 17990 9003 17992
rect 7741 17987 7807 17990
rect 8937 17987 9003 17990
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 10869 17914 10935 17917
rect 12709 17914 12775 17917
rect 10869 17912 12775 17914
rect 10869 17856 10874 17912
rect 10930 17856 12714 17912
rect 12770 17856 12775 17912
rect 10869 17854 12775 17856
rect 10869 17851 10935 17854
rect 12709 17851 12775 17854
rect 15653 17914 15719 17917
rect 18413 17914 18479 17917
rect 15653 17912 18479 17914
rect 15653 17856 15658 17912
rect 15714 17856 18418 17912
rect 18474 17856 18479 17912
rect 15653 17854 18479 17856
rect 15653 17851 15719 17854
rect 18413 17851 18479 17854
rect 0 17778 480 17808
rect 9765 17778 9831 17781
rect 0 17776 9831 17778
rect 0 17720 9770 17776
rect 9826 17720 9831 17776
rect 0 17718 9831 17720
rect 0 17688 480 17718
rect 9765 17715 9831 17718
rect 10777 17778 10843 17781
rect 12617 17778 12683 17781
rect 10777 17776 12683 17778
rect 10777 17720 10782 17776
rect 10838 17720 12622 17776
rect 12678 17720 12683 17776
rect 10777 17718 12683 17720
rect 10777 17715 10843 17718
rect 12617 17715 12683 17718
rect 2957 17642 3023 17645
rect 11237 17642 11303 17645
rect 12341 17642 12407 17645
rect 2957 17640 12407 17642
rect 2957 17584 2962 17640
rect 3018 17584 11242 17640
rect 11298 17584 12346 17640
rect 12402 17584 12407 17640
rect 2957 17582 12407 17584
rect 2957 17579 3023 17582
rect 11237 17579 11303 17582
rect 12341 17579 12407 17582
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 3509 17372 3575 17373
rect 3509 17370 3556 17372
rect 3464 17368 3556 17370
rect 3464 17312 3514 17368
rect 3464 17310 3556 17312
rect 3509 17308 3556 17310
rect 3620 17308 3626 17372
rect 15653 17370 15719 17373
rect 16430 17370 16436 17372
rect 15653 17368 16436 17370
rect 15653 17312 15658 17368
rect 15714 17312 16436 17368
rect 15653 17310 16436 17312
rect 3509 17307 3575 17308
rect 15653 17307 15719 17310
rect 16430 17308 16436 17310
rect 16500 17370 16506 17372
rect 17401 17370 17467 17373
rect 16500 17368 17467 17370
rect 16500 17312 17406 17368
rect 17462 17312 17467 17368
rect 16500 17310 17467 17312
rect 16500 17308 16506 17310
rect 17401 17307 17467 17310
rect 0 17234 480 17264
rect 2957 17234 3023 17237
rect 0 17232 3023 17234
rect 0 17176 2962 17232
rect 3018 17176 3023 17232
rect 0 17174 3023 17176
rect 0 17144 480 17174
rect 2957 17171 3023 17174
rect 7833 17234 7899 17237
rect 12249 17234 12315 17237
rect 7833 17232 12315 17234
rect 7833 17176 7838 17232
rect 7894 17176 12254 17232
rect 12310 17176 12315 17232
rect 7833 17174 12315 17176
rect 7833 17171 7899 17174
rect 12249 17171 12315 17174
rect 9581 17098 9647 17101
rect 11973 17098 12039 17101
rect 9581 17096 12039 17098
rect 9581 17040 9586 17096
rect 9642 17040 11978 17096
rect 12034 17040 12039 17096
rect 9581 17038 12039 17040
rect 9581 17035 9647 17038
rect 11973 17035 12039 17038
rect 15009 17098 15075 17101
rect 16389 17098 16455 17101
rect 15009 17096 16455 17098
rect 15009 17040 15014 17096
rect 15070 17040 16394 17096
rect 16450 17040 16455 17096
rect 15009 17038 16455 17040
rect 15009 17035 15075 17038
rect 16389 17035 16455 17038
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 5809 16826 5875 16829
rect 8477 16826 8543 16829
rect 5809 16824 8543 16826
rect 5809 16768 5814 16824
rect 5870 16768 8482 16824
rect 8538 16768 8543 16824
rect 5809 16766 8543 16768
rect 5809 16763 5875 16766
rect 8477 16763 8543 16766
rect 10869 16826 10935 16829
rect 11237 16826 11303 16829
rect 15285 16826 15351 16829
rect 10869 16824 15351 16826
rect 10869 16768 10874 16824
rect 10930 16768 11242 16824
rect 11298 16768 15290 16824
rect 15346 16768 15351 16824
rect 10869 16766 15351 16768
rect 10869 16763 10935 16766
rect 11237 16763 11303 16766
rect 15285 16763 15351 16766
rect 0 16690 480 16720
rect 3693 16690 3759 16693
rect 0 16688 3759 16690
rect 0 16632 3698 16688
rect 3754 16632 3759 16688
rect 0 16630 3759 16632
rect 0 16600 480 16630
rect 3693 16627 3759 16630
rect 6453 16690 6519 16693
rect 8661 16690 8727 16693
rect 6453 16688 8727 16690
rect 6453 16632 6458 16688
rect 6514 16632 8666 16688
rect 8722 16632 8727 16688
rect 6453 16630 8727 16632
rect 6453 16627 6519 16630
rect 8661 16627 8727 16630
rect 8937 16690 9003 16693
rect 12985 16690 13051 16693
rect 8937 16688 13051 16690
rect 8937 16632 8942 16688
rect 8998 16632 12990 16688
rect 13046 16632 13051 16688
rect 8937 16630 13051 16632
rect 8937 16627 9003 16630
rect 12985 16627 13051 16630
rect 13721 16690 13787 16693
rect 14917 16690 14983 16693
rect 13721 16688 14983 16690
rect 13721 16632 13726 16688
rect 13782 16632 14922 16688
rect 14978 16632 14983 16688
rect 13721 16630 14983 16632
rect 13721 16627 13787 16630
rect 14917 16627 14983 16630
rect 4153 16554 4219 16557
rect 12525 16554 12591 16557
rect 4153 16552 12591 16554
rect 4153 16496 4158 16552
rect 4214 16496 12530 16552
rect 12586 16496 12591 16552
rect 4153 16494 12591 16496
rect 4153 16491 4219 16494
rect 12525 16491 12591 16494
rect 13629 16554 13695 16557
rect 17309 16554 17375 16557
rect 13629 16552 17375 16554
rect 13629 16496 13634 16552
rect 13690 16496 17314 16552
rect 17370 16496 17375 16552
rect 13629 16494 17375 16496
rect 13629 16491 13695 16494
rect 17309 16491 17375 16494
rect 1577 16418 1643 16421
rect 2681 16418 2747 16421
rect 1577 16416 2747 16418
rect 1577 16360 1582 16416
rect 1638 16360 2686 16416
rect 2742 16360 2747 16416
rect 1577 16358 2747 16360
rect 1577 16355 1643 16358
rect 2681 16355 2747 16358
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 2497 16146 2563 16149
rect 12617 16146 12683 16149
rect 2497 16144 12683 16146
rect 2497 16088 2502 16144
rect 2558 16088 12622 16144
rect 12678 16088 12683 16144
rect 2497 16086 12683 16088
rect 2497 16083 2563 16086
rect 12617 16083 12683 16086
rect 0 16010 480 16040
rect 5165 16010 5231 16013
rect 11697 16010 11763 16013
rect 0 15950 5090 16010
rect 0 15920 480 15950
rect 2773 15874 2839 15877
rect 4705 15874 4771 15877
rect 2773 15872 4771 15874
rect 2773 15816 2778 15872
rect 2834 15816 4710 15872
rect 4766 15816 4771 15872
rect 2773 15814 4771 15816
rect 5030 15874 5090 15950
rect 5165 16008 11763 16010
rect 5165 15952 5170 16008
rect 5226 15952 11702 16008
rect 11758 15952 11763 16008
rect 5165 15950 11763 15952
rect 5165 15947 5231 15950
rect 11697 15947 11763 15950
rect 5030 15814 10012 15874
rect 2773 15811 2839 15814
rect 4705 15811 4771 15814
rect 3877 15738 3943 15741
rect 4337 15738 4403 15741
rect 6637 15738 6703 15741
rect 3877 15736 6703 15738
rect 3877 15680 3882 15736
rect 3938 15680 4342 15736
rect 4398 15680 6642 15736
rect 6698 15680 6703 15736
rect 3877 15678 6703 15680
rect 3877 15675 3943 15678
rect 4337 15675 4403 15678
rect 6637 15675 6703 15678
rect 2037 15602 2103 15605
rect 4429 15602 4495 15605
rect 2037 15600 4495 15602
rect 2037 15544 2042 15600
rect 2098 15544 4434 15600
rect 4490 15544 4495 15600
rect 2037 15542 4495 15544
rect 2037 15539 2103 15542
rect 4429 15539 4495 15542
rect 7281 15602 7347 15605
rect 9765 15602 9831 15605
rect 7281 15600 9831 15602
rect 7281 15544 7286 15600
rect 7342 15544 9770 15600
rect 9826 15544 9831 15600
rect 7281 15542 9831 15544
rect 9952 15602 10012 15814
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 10777 15738 10843 15741
rect 16849 15738 16915 15741
rect 10777 15736 16915 15738
rect 10777 15680 10782 15736
rect 10838 15680 16854 15736
rect 16910 15680 16915 15736
rect 10777 15678 16915 15680
rect 10777 15675 10843 15678
rect 16849 15675 16915 15678
rect 11697 15602 11763 15605
rect 9952 15600 11763 15602
rect 9952 15544 11702 15600
rect 11758 15544 11763 15600
rect 9952 15542 11763 15544
rect 7281 15539 7347 15542
rect 9765 15539 9831 15542
rect 11697 15539 11763 15542
rect 0 15466 480 15496
rect 2681 15466 2747 15469
rect 0 15464 2747 15466
rect 0 15408 2686 15464
rect 2742 15408 2747 15464
rect 0 15406 2747 15408
rect 0 15376 480 15406
rect 2681 15403 2747 15406
rect 3785 15466 3851 15469
rect 5993 15466 6059 15469
rect 20621 15466 20687 15469
rect 3785 15464 20687 15466
rect 3785 15408 3790 15464
rect 3846 15408 5998 15464
rect 6054 15408 20626 15464
rect 20682 15408 20687 15464
rect 3785 15406 20687 15408
rect 3785 15403 3851 15406
rect 5993 15403 6059 15406
rect 20621 15403 20687 15406
rect 11237 15330 11303 15333
rect 13261 15330 13327 15333
rect 11237 15328 13327 15330
rect 11237 15272 11242 15328
rect 11298 15272 13266 15328
rect 13322 15272 13327 15328
rect 11237 15270 13327 15272
rect 11237 15267 11303 15270
rect 13261 15267 13327 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 2405 15194 2471 15197
rect 4521 15194 4587 15197
rect 2405 15192 4587 15194
rect 2405 15136 2410 15192
rect 2466 15136 4526 15192
rect 4582 15136 4587 15192
rect 2405 15134 4587 15136
rect 2405 15131 2471 15134
rect 4521 15131 4587 15134
rect 5993 15194 6059 15197
rect 7097 15194 7163 15197
rect 5993 15192 7163 15194
rect 5993 15136 5998 15192
rect 6054 15136 7102 15192
rect 7158 15136 7163 15192
rect 5993 15134 7163 15136
rect 5993 15131 6059 15134
rect 7097 15131 7163 15134
rect 3969 15058 4035 15061
rect 6085 15058 6151 15061
rect 3969 15056 6151 15058
rect 3969 15000 3974 15056
rect 4030 15000 6090 15056
rect 6146 15000 6151 15056
rect 3969 14998 6151 15000
rect 3969 14995 4035 14998
rect 6085 14995 6151 14998
rect 6545 15058 6611 15061
rect 25497 15058 25563 15061
rect 6545 15056 25563 15058
rect 6545 15000 6550 15056
rect 6606 15000 25502 15056
rect 25558 15000 25563 15056
rect 6545 14998 25563 15000
rect 6545 14995 6611 14998
rect 25497 14995 25563 14998
rect 0 14922 480 14952
rect 3877 14922 3943 14925
rect 0 14920 3943 14922
rect 0 14864 3882 14920
rect 3938 14864 3943 14920
rect 0 14862 3943 14864
rect 0 14832 480 14862
rect 3877 14859 3943 14862
rect 5073 14922 5139 14925
rect 11605 14922 11671 14925
rect 5073 14920 11671 14922
rect 5073 14864 5078 14920
rect 5134 14864 11610 14920
rect 11666 14864 11671 14920
rect 5073 14862 11671 14864
rect 5073 14859 5139 14862
rect 11605 14859 11671 14862
rect 11329 14786 11395 14789
rect 17493 14786 17559 14789
rect 11329 14784 17559 14786
rect 11329 14728 11334 14784
rect 11390 14728 17498 14784
rect 17554 14728 17559 14784
rect 11329 14726 17559 14728
rect 11329 14723 11395 14726
rect 17493 14723 17559 14726
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 14457 14514 14523 14517
rect 14590 14514 14596 14516
rect 14457 14512 14596 14514
rect 14457 14456 14462 14512
rect 14518 14456 14596 14512
rect 14457 14454 14596 14456
rect 14457 14451 14523 14454
rect 14590 14452 14596 14454
rect 14660 14452 14666 14516
rect 0 14378 480 14408
rect 6177 14378 6243 14381
rect 0 14376 6243 14378
rect 0 14320 6182 14376
rect 6238 14320 6243 14376
rect 0 14318 6243 14320
rect 0 14288 480 14318
rect 5214 14245 5274 14318
rect 6177 14315 6243 14318
rect 14273 14378 14339 14381
rect 16665 14378 16731 14381
rect 14273 14376 16731 14378
rect 14273 14320 14278 14376
rect 14334 14320 16670 14376
rect 16726 14320 16731 14376
rect 14273 14318 16731 14320
rect 14273 14315 14339 14318
rect 16665 14315 16731 14318
rect 5214 14240 5323 14245
rect 5214 14184 5262 14240
rect 5318 14184 5323 14240
rect 5214 14182 5323 14184
rect 5257 14179 5323 14182
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 2497 13970 2563 13973
rect 2865 13970 2931 13973
rect 2497 13968 2931 13970
rect 2497 13912 2502 13968
rect 2558 13912 2870 13968
rect 2926 13912 2931 13968
rect 2497 13910 2931 13912
rect 2497 13907 2563 13910
rect 2865 13907 2931 13910
rect 16757 13970 16823 13973
rect 19425 13970 19491 13973
rect 16757 13968 19491 13970
rect 16757 13912 16762 13968
rect 16818 13912 19430 13968
rect 19486 13912 19491 13968
rect 16757 13910 19491 13912
rect 16757 13907 16823 13910
rect 19425 13907 19491 13910
rect 24393 13970 24459 13973
rect 27520 13970 28000 14000
rect 24393 13968 28000 13970
rect 24393 13912 24398 13968
rect 24454 13912 28000 13968
rect 24393 13910 28000 13912
rect 24393 13907 24459 13910
rect 27520 13880 28000 13910
rect 3233 13834 3299 13837
rect 5625 13834 5691 13837
rect 3233 13832 5691 13834
rect 3233 13776 3238 13832
rect 3294 13776 5630 13832
rect 5686 13776 5691 13832
rect 3233 13774 5691 13776
rect 3233 13771 3299 13774
rect 5625 13771 5691 13774
rect 7097 13834 7163 13837
rect 10777 13834 10843 13837
rect 13169 13834 13235 13837
rect 7097 13832 13235 13834
rect 7097 13776 7102 13832
rect 7158 13776 10782 13832
rect 10838 13776 13174 13832
rect 13230 13776 13235 13832
rect 7097 13774 13235 13776
rect 7097 13771 7163 13774
rect 10777 13771 10843 13774
rect 13169 13771 13235 13774
rect 18689 13834 18755 13837
rect 24117 13834 24183 13837
rect 18689 13832 24183 13834
rect 18689 13776 18694 13832
rect 18750 13776 24122 13832
rect 24178 13776 24183 13832
rect 18689 13774 24183 13776
rect 18689 13771 18755 13774
rect 24117 13771 24183 13774
rect 0 13698 480 13728
rect 2405 13698 2471 13701
rect 2957 13698 3023 13701
rect 5533 13698 5599 13701
rect 0 13638 1410 13698
rect 0 13608 480 13638
rect 1350 13562 1410 13638
rect 2405 13696 5599 13698
rect 2405 13640 2410 13696
rect 2466 13640 2962 13696
rect 3018 13640 5538 13696
rect 5594 13640 5599 13696
rect 2405 13638 5599 13640
rect 2405 13635 2471 13638
rect 2957 13635 3023 13638
rect 5533 13635 5599 13638
rect 6637 13698 6703 13701
rect 6821 13698 6887 13701
rect 6637 13696 6887 13698
rect 6637 13640 6642 13696
rect 6698 13640 6826 13696
rect 6882 13640 6887 13696
rect 6637 13638 6887 13640
rect 6637 13635 6703 13638
rect 6821 13635 6887 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 3601 13562 3667 13565
rect 1350 13560 3667 13562
rect 1350 13504 3606 13560
rect 3662 13504 3667 13560
rect 1350 13502 3667 13504
rect 3601 13499 3667 13502
rect 2037 13426 2103 13429
rect 3417 13426 3483 13429
rect 2037 13424 3483 13426
rect 2037 13368 2042 13424
rect 2098 13368 3422 13424
rect 3478 13368 3483 13424
rect 2037 13366 3483 13368
rect 2037 13363 2103 13366
rect 3417 13363 3483 13366
rect 3693 13426 3759 13429
rect 5809 13426 5875 13429
rect 3693 13424 5875 13426
rect 3693 13368 3698 13424
rect 3754 13368 5814 13424
rect 5870 13368 5875 13424
rect 3693 13366 5875 13368
rect 3693 13363 3759 13366
rect 5809 13363 5875 13366
rect 1393 13290 1459 13293
rect 4521 13290 4587 13293
rect 1393 13288 4587 13290
rect 1393 13232 1398 13288
rect 1454 13232 4526 13288
rect 4582 13232 4587 13288
rect 1393 13230 4587 13232
rect 1393 13227 1459 13230
rect 4521 13227 4587 13230
rect 8201 13290 8267 13293
rect 11329 13290 11395 13293
rect 8201 13288 11395 13290
rect 8201 13232 8206 13288
rect 8262 13232 11334 13288
rect 11390 13232 11395 13288
rect 8201 13230 11395 13232
rect 8201 13227 8267 13230
rect 11329 13227 11395 13230
rect 12893 13290 12959 13293
rect 15377 13290 15443 13293
rect 12893 13288 15443 13290
rect 12893 13232 12898 13288
rect 12954 13232 15382 13288
rect 15438 13232 15443 13288
rect 12893 13230 15443 13232
rect 12893 13227 12959 13230
rect 15377 13227 15443 13230
rect 0 13154 480 13184
rect 1577 13154 1643 13157
rect 1853 13154 1919 13157
rect 0 13152 1919 13154
rect 0 13096 1582 13152
rect 1638 13096 1858 13152
rect 1914 13096 1919 13152
rect 0 13094 1919 13096
rect 0 13064 480 13094
rect 1577 13091 1643 13094
rect 1853 13091 1919 13094
rect 3366 13092 3372 13156
rect 3436 13154 3442 13156
rect 3509 13154 3575 13157
rect 3436 13152 3575 13154
rect 3436 13096 3514 13152
rect 3570 13096 3575 13152
rect 3436 13094 3575 13096
rect 3436 13092 3442 13094
rect 3509 13091 3575 13094
rect 7373 13154 7439 13157
rect 13353 13154 13419 13157
rect 7373 13152 13419 13154
rect 7373 13096 7378 13152
rect 7434 13096 13358 13152
rect 13414 13096 13419 13152
rect 7373 13094 13419 13096
rect 7373 13091 7439 13094
rect 13353 13091 13419 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 13629 13018 13695 13021
rect 13629 13016 14106 13018
rect 13629 12960 13634 13016
rect 13690 12960 14106 13016
rect 13629 12958 14106 12960
rect 13629 12955 13695 12958
rect 3877 12882 3943 12885
rect 13813 12882 13879 12885
rect 3877 12880 13879 12882
rect 3877 12824 3882 12880
rect 3938 12824 13818 12880
rect 13874 12824 13879 12880
rect 3877 12822 13879 12824
rect 14046 12882 14106 12958
rect 21909 12882 21975 12885
rect 14046 12880 21975 12882
rect 14046 12824 21914 12880
rect 21970 12824 21975 12880
rect 14046 12822 21975 12824
rect 3877 12819 3943 12822
rect 13813 12819 13879 12822
rect 21909 12819 21975 12822
rect 2681 12746 2747 12749
rect 16757 12746 16823 12749
rect 2681 12744 16823 12746
rect 2681 12688 2686 12744
rect 2742 12688 16762 12744
rect 16818 12688 16823 12744
rect 2681 12686 16823 12688
rect 2681 12683 2747 12686
rect 16757 12683 16823 12686
rect 0 12610 480 12640
rect 6729 12610 6795 12613
rect 0 12608 6795 12610
rect 0 12552 6734 12608
rect 6790 12552 6795 12608
rect 0 12550 6795 12552
rect 0 12520 480 12550
rect 6729 12547 6795 12550
rect 16113 12610 16179 12613
rect 18413 12610 18479 12613
rect 16113 12608 18479 12610
rect 16113 12552 16118 12608
rect 16174 12552 18418 12608
rect 18474 12552 18479 12608
rect 16113 12550 18479 12552
rect 16113 12547 16179 12550
rect 18413 12547 18479 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 3417 12474 3483 12477
rect 6821 12474 6887 12477
rect 10133 12474 10199 12477
rect 3417 12472 10199 12474
rect 3417 12416 3422 12472
rect 3478 12416 6826 12472
rect 6882 12416 10138 12472
rect 10194 12416 10199 12472
rect 3417 12414 10199 12416
rect 3417 12411 3483 12414
rect 6821 12411 6887 12414
rect 10133 12411 10199 12414
rect 11881 12474 11947 12477
rect 12893 12474 12959 12477
rect 11881 12472 12959 12474
rect 11881 12416 11886 12472
rect 11942 12416 12898 12472
rect 12954 12416 12959 12472
rect 11881 12414 12959 12416
rect 11881 12411 11947 12414
rect 12893 12411 12959 12414
rect 14273 12340 14339 12341
rect 14222 12338 14228 12340
rect 14182 12278 14228 12338
rect 14292 12336 14339 12340
rect 14334 12280 14339 12336
rect 14222 12276 14228 12278
rect 14292 12276 14339 12280
rect 14273 12275 14339 12276
rect 5165 12202 5231 12205
rect 10685 12202 10751 12205
rect 5165 12200 10751 12202
rect 5165 12144 5170 12200
rect 5226 12144 10690 12200
rect 10746 12144 10751 12200
rect 5165 12142 10751 12144
rect 5165 12139 5231 12142
rect 10685 12139 10751 12142
rect 15009 12202 15075 12205
rect 20805 12202 20871 12205
rect 15009 12200 20871 12202
rect 15009 12144 15014 12200
rect 15070 12144 20810 12200
rect 20866 12144 20871 12200
rect 15009 12142 20871 12144
rect 15009 12139 15075 12142
rect 20805 12139 20871 12142
rect 5610 12000 5930 12001
rect 0 11930 480 11960
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 0 11870 4906 11930
rect 0 11840 480 11870
rect 4846 11794 4906 11870
rect 11421 11794 11487 11797
rect 11973 11794 12039 11797
rect 4846 11792 12039 11794
rect 4846 11736 11426 11792
rect 11482 11736 11978 11792
rect 12034 11736 12039 11792
rect 4846 11734 12039 11736
rect 11421 11731 11487 11734
rect 11973 11731 12039 11734
rect 14590 11732 14596 11796
rect 14660 11794 14666 11796
rect 14825 11794 14891 11797
rect 14660 11792 14891 11794
rect 14660 11736 14830 11792
rect 14886 11736 14891 11792
rect 14660 11734 14891 11736
rect 14660 11732 14666 11734
rect 14825 11731 14891 11734
rect 15929 11658 15995 11661
rect 4846 11656 15995 11658
rect 4846 11600 15934 11656
rect 15990 11600 15995 11656
rect 4846 11598 15995 11600
rect 0 11386 480 11416
rect 4846 11386 4906 11598
rect 15929 11595 15995 11598
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 10041 11386 10107 11389
rect 0 11326 4906 11386
rect 9998 11384 10107 11386
rect 9998 11328 10046 11384
rect 10102 11328 10107 11384
rect 0 11296 480 11326
rect 9998 11323 10107 11328
rect 3969 11250 4035 11253
rect 7005 11250 7071 11253
rect 9998 11250 10058 11323
rect 3969 11248 10058 11250
rect 3969 11192 3974 11248
rect 4030 11192 7010 11248
rect 7066 11192 10058 11248
rect 3969 11190 10058 11192
rect 3969 11187 4035 11190
rect 7005 11187 7071 11190
rect 10133 11114 10199 11117
rect 11094 11114 11100 11116
rect 5398 11054 6194 11114
rect 3785 10978 3851 10981
rect 5398 10978 5458 11054
rect 3785 10976 5458 10978
rect 3785 10920 3790 10976
rect 3846 10920 5458 10976
rect 3785 10918 5458 10920
rect 6134 10978 6194 11054
rect 10133 11112 11100 11114
rect 10133 11056 10138 11112
rect 10194 11056 11100 11112
rect 10133 11054 11100 11056
rect 10133 11051 10199 11054
rect 11094 11052 11100 11054
rect 11164 11052 11170 11116
rect 11881 11114 11947 11117
rect 14365 11114 14431 11117
rect 17585 11114 17651 11117
rect 11881 11112 14290 11114
rect 11881 11056 11886 11112
rect 11942 11056 14290 11112
rect 11881 11054 14290 11056
rect 11881 11051 11947 11054
rect 14230 10981 14290 11054
rect 14365 11112 17651 11114
rect 14365 11056 14370 11112
rect 14426 11056 17590 11112
rect 17646 11056 17651 11112
rect 14365 11054 17651 11056
rect 14365 11051 14431 11054
rect 17585 11051 17651 11054
rect 18045 11114 18111 11117
rect 20713 11114 20779 11117
rect 18045 11112 20779 11114
rect 18045 11056 18050 11112
rect 18106 11056 20718 11112
rect 20774 11056 20779 11112
rect 18045 11054 20779 11056
rect 18045 11051 18111 11054
rect 20713 11051 20779 11054
rect 12709 10978 12775 10981
rect 6134 10976 12775 10978
rect 6134 10920 12714 10976
rect 12770 10920 12775 10976
rect 6134 10918 12775 10920
rect 14230 10976 14339 10981
rect 14230 10920 14278 10976
rect 14334 10920 14339 10976
rect 14230 10918 14339 10920
rect 3785 10915 3851 10918
rect 12709 10915 12775 10918
rect 14273 10915 14339 10918
rect 5610 10912 5930 10913
rect 0 10842 480 10872
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 11605 10842 11671 10845
rect 13445 10842 13511 10845
rect 0 10782 2882 10842
rect 0 10752 480 10782
rect 2822 10570 2882 10782
rect 5996 10840 13511 10842
rect 5996 10784 11610 10840
rect 11666 10784 13450 10840
rect 13506 10784 13511 10840
rect 5996 10782 13511 10784
rect 2957 10706 3023 10709
rect 5809 10706 5875 10709
rect 2957 10704 5875 10706
rect 2957 10648 2962 10704
rect 3018 10648 5814 10704
rect 5870 10648 5875 10704
rect 2957 10646 5875 10648
rect 2957 10643 3023 10646
rect 5809 10643 5875 10646
rect 5996 10570 6056 10782
rect 11605 10779 11671 10782
rect 13445 10779 13511 10782
rect 7189 10706 7255 10709
rect 18137 10706 18203 10709
rect 7189 10704 18203 10706
rect 7189 10648 7194 10704
rect 7250 10648 18142 10704
rect 18198 10648 18203 10704
rect 7189 10646 18203 10648
rect 7189 10643 7255 10646
rect 18137 10643 18203 10646
rect 2822 10510 6056 10570
rect 6821 10570 6887 10573
rect 18413 10570 18479 10573
rect 6821 10568 18479 10570
rect 6821 10512 6826 10568
rect 6882 10512 18418 10568
rect 18474 10512 18479 10568
rect 6821 10510 18479 10512
rect 6821 10507 6887 10510
rect 18413 10507 18479 10510
rect 2037 10434 2103 10437
rect 4061 10434 4127 10437
rect 2037 10432 4127 10434
rect 2037 10376 2042 10432
rect 2098 10376 4066 10432
rect 4122 10376 4127 10432
rect 2037 10374 4127 10376
rect 2037 10371 2103 10374
rect 4061 10371 4127 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 1853 10298 1919 10301
rect 5625 10298 5691 10301
rect 1853 10296 5691 10298
rect 1853 10240 1858 10296
rect 1914 10240 5630 10296
rect 5686 10240 5691 10296
rect 1853 10238 5691 10240
rect 1853 10235 1919 10238
rect 5625 10235 5691 10238
rect 0 10162 480 10192
rect 3969 10162 4035 10165
rect 0 10160 4035 10162
rect 0 10104 3974 10160
rect 4030 10104 4035 10160
rect 0 10102 4035 10104
rect 0 10072 480 10102
rect 3969 10099 4035 10102
rect 6085 10162 6151 10165
rect 8477 10162 8543 10165
rect 17401 10162 17467 10165
rect 6085 10160 17467 10162
rect 6085 10104 6090 10160
rect 6146 10104 8482 10160
rect 8538 10104 17406 10160
rect 17462 10104 17467 10160
rect 6085 10102 17467 10104
rect 6085 10099 6151 10102
rect 8477 10099 8543 10102
rect 17401 10099 17467 10102
rect 7097 10026 7163 10029
rect 18965 10026 19031 10029
rect 7097 10024 19031 10026
rect 7097 9968 7102 10024
rect 7158 9968 18970 10024
rect 19026 9968 19031 10024
rect 7097 9966 19031 9968
rect 7097 9963 7163 9966
rect 18965 9963 19031 9966
rect 14733 9890 14799 9893
rect 6134 9888 14799 9890
rect 6134 9832 14738 9888
rect 14794 9832 14799 9888
rect 6134 9830 14799 9832
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 3918 9692 3924 9756
rect 3988 9754 3994 9756
rect 3988 9694 5458 9754
rect 3988 9692 3994 9694
rect 0 9618 480 9648
rect 1577 9618 1643 9621
rect 5073 9618 5139 9621
rect 0 9558 1226 9618
rect 0 9528 480 9558
rect 1166 9346 1226 9558
rect 1577 9616 5139 9618
rect 1577 9560 1582 9616
rect 1638 9560 5078 9616
rect 5134 9560 5139 9616
rect 1577 9558 5139 9560
rect 5398 9618 5458 9694
rect 6134 9618 6194 9830
rect 14733 9827 14799 9830
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 14089 9754 14155 9757
rect 14222 9754 14228 9756
rect 14089 9752 14228 9754
rect 14089 9696 14094 9752
rect 14150 9696 14228 9752
rect 14089 9694 14228 9696
rect 14089 9691 14155 9694
rect 14222 9692 14228 9694
rect 14292 9692 14298 9756
rect 15377 9754 15443 9757
rect 19977 9754 20043 9757
rect 15377 9752 20043 9754
rect 15377 9696 15382 9752
rect 15438 9696 19982 9752
rect 20038 9696 20043 9752
rect 15377 9694 20043 9696
rect 15377 9691 15443 9694
rect 19977 9691 20043 9694
rect 5398 9558 6194 9618
rect 10593 9618 10659 9621
rect 11237 9618 11303 9621
rect 10593 9616 11303 9618
rect 10593 9560 10598 9616
rect 10654 9560 11242 9616
rect 11298 9560 11303 9616
rect 10593 9558 11303 9560
rect 1577 9555 1643 9558
rect 5073 9555 5139 9558
rect 10593 9555 10659 9558
rect 11237 9555 11303 9558
rect 1393 9482 1459 9485
rect 7189 9482 7255 9485
rect 1393 9480 7255 9482
rect 1393 9424 1398 9480
rect 1454 9424 7194 9480
rect 7250 9424 7255 9480
rect 1393 9422 7255 9424
rect 1393 9419 1459 9422
rect 7189 9419 7255 9422
rect 8109 9482 8175 9485
rect 11329 9482 11395 9485
rect 8109 9480 9874 9482
rect 8109 9424 8114 9480
rect 8170 9424 9874 9480
rect 10366 9480 11395 9482
rect 10366 9448 11334 9480
rect 8109 9422 9874 9424
rect 8109 9419 8175 9422
rect 9213 9346 9279 9349
rect 1166 9344 9279 9346
rect 1166 9288 9218 9344
rect 9274 9288 9279 9344
rect 1166 9286 9279 9288
rect 9814 9346 9874 9422
rect 10136 9424 11334 9448
rect 11390 9424 11395 9480
rect 10136 9422 11395 9424
rect 10136 9388 10426 9422
rect 11329 9419 11395 9422
rect 14273 9482 14339 9485
rect 17953 9482 18019 9485
rect 14273 9480 18019 9482
rect 14273 9424 14278 9480
rect 14334 9424 17958 9480
rect 18014 9424 18019 9480
rect 14273 9422 18019 9424
rect 14273 9419 14339 9422
rect 17953 9419 18019 9422
rect 10136 9346 10196 9388
rect 9814 9286 10196 9346
rect 11237 9346 11303 9349
rect 18873 9346 18939 9349
rect 11237 9344 18939 9346
rect 11237 9288 11242 9344
rect 11298 9288 18878 9344
rect 18934 9288 18939 9344
rect 11237 9286 18939 9288
rect 9213 9283 9279 9286
rect 11237 9283 11303 9286
rect 18873 9283 18939 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 16849 9210 16915 9213
rect 19425 9210 19491 9213
rect 16849 9208 19491 9210
rect 16849 9152 16854 9208
rect 16910 9152 19430 9208
rect 19486 9152 19491 9208
rect 16849 9150 19491 9152
rect 16849 9147 16915 9150
rect 19425 9147 19491 9150
rect 0 9074 480 9104
rect 1485 9074 1551 9077
rect 0 9072 1551 9074
rect 0 9016 1490 9072
rect 1546 9016 1551 9072
rect 0 9014 1551 9016
rect 0 8984 480 9014
rect 1485 9011 1551 9014
rect 3049 9074 3115 9077
rect 10133 9074 10199 9077
rect 12198 9074 12204 9076
rect 3049 9072 10199 9074
rect 3049 9016 3054 9072
rect 3110 9016 10138 9072
rect 10194 9016 10199 9072
rect 3049 9014 10199 9016
rect 3049 9011 3115 9014
rect 10133 9011 10199 9014
rect 10918 9014 12204 9074
rect 9489 8938 9555 8941
rect 10918 8938 10978 9014
rect 12198 9012 12204 9014
rect 12268 9012 12274 9076
rect 9489 8936 10978 8938
rect 9489 8880 9494 8936
rect 9550 8880 10978 8936
rect 9489 8878 10978 8880
rect 11145 8938 11211 8941
rect 20069 8938 20135 8941
rect 11145 8936 20135 8938
rect 11145 8880 11150 8936
rect 11206 8880 20074 8936
rect 20130 8880 20135 8936
rect 11145 8878 20135 8880
rect 9489 8875 9555 8878
rect 11145 8875 11211 8878
rect 20069 8875 20135 8878
rect 6269 8804 6335 8805
rect 6269 8802 6316 8804
rect 6224 8800 6316 8802
rect 6224 8744 6274 8800
rect 6224 8742 6316 8744
rect 6269 8740 6316 8742
rect 6380 8740 6386 8804
rect 10041 8802 10107 8805
rect 14733 8802 14799 8805
rect 10041 8800 14799 8802
rect 10041 8744 10046 8800
rect 10102 8744 14738 8800
rect 14794 8744 14799 8800
rect 10041 8742 14799 8744
rect 6269 8739 6335 8740
rect 10041 8739 10107 8742
rect 14733 8739 14799 8742
rect 17217 8802 17283 8805
rect 20253 8802 20319 8805
rect 17217 8800 20319 8802
rect 17217 8744 17222 8800
rect 17278 8744 20258 8800
rect 20314 8744 20319 8800
rect 17217 8742 20319 8744
rect 17217 8739 17283 8742
rect 20253 8739 20319 8742
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 1945 8666 2011 8669
rect 11789 8666 11855 8669
rect 13537 8666 13603 8669
rect 1945 8664 2514 8666
rect 1945 8608 1950 8664
rect 2006 8608 2514 8664
rect 1945 8606 2514 8608
rect 1945 8603 2011 8606
rect 0 8530 480 8560
rect 2454 8530 2514 8606
rect 11789 8664 13603 8666
rect 11789 8608 11794 8664
rect 11850 8608 13542 8664
rect 13598 8608 13603 8664
rect 11789 8606 13603 8608
rect 11789 8603 11855 8606
rect 13537 8603 13603 8606
rect 17677 8666 17743 8669
rect 20989 8666 21055 8669
rect 17677 8664 21055 8666
rect 17677 8608 17682 8664
rect 17738 8608 20994 8664
rect 21050 8608 21055 8664
rect 17677 8606 21055 8608
rect 17677 8603 17743 8606
rect 20989 8603 21055 8606
rect 5993 8530 6059 8533
rect 0 8470 2330 8530
rect 2454 8528 6059 8530
rect 2454 8472 5998 8528
rect 6054 8472 6059 8528
rect 2454 8470 6059 8472
rect 0 8440 480 8470
rect 2270 8122 2330 8470
rect 5993 8467 6059 8470
rect 8201 8530 8267 8533
rect 21173 8530 21239 8533
rect 8201 8528 21239 8530
rect 8201 8472 8206 8528
rect 8262 8472 21178 8528
rect 21234 8472 21239 8528
rect 8201 8470 21239 8472
rect 8201 8467 8267 8470
rect 21173 8467 21239 8470
rect 2405 8394 2471 8397
rect 5533 8394 5599 8397
rect 2405 8392 5599 8394
rect 2405 8336 2410 8392
rect 2466 8336 5538 8392
rect 5594 8336 5599 8392
rect 2405 8334 5599 8336
rect 2405 8331 2471 8334
rect 5533 8331 5599 8334
rect 6637 8394 6703 8397
rect 8845 8394 8911 8397
rect 6637 8392 8911 8394
rect 6637 8336 6642 8392
rect 6698 8336 8850 8392
rect 8906 8336 8911 8392
rect 6637 8334 8911 8336
rect 6637 8331 6703 8334
rect 8845 8331 8911 8334
rect 14733 8394 14799 8397
rect 19609 8394 19675 8397
rect 14733 8392 19675 8394
rect 14733 8336 14738 8392
rect 14794 8336 19614 8392
rect 19670 8336 19675 8392
rect 14733 8334 19675 8336
rect 14733 8331 14799 8334
rect 19609 8331 19675 8334
rect 4613 8258 4679 8261
rect 7097 8258 7163 8261
rect 9949 8258 10015 8261
rect 4613 8256 10015 8258
rect 4613 8200 4618 8256
rect 4674 8200 7102 8256
rect 7158 8200 9954 8256
rect 10010 8200 10015 8256
rect 4613 8198 10015 8200
rect 4613 8195 4679 8198
rect 7097 8195 7163 8198
rect 9949 8195 10015 8198
rect 10685 8258 10751 8261
rect 11421 8258 11487 8261
rect 10685 8256 11487 8258
rect 10685 8200 10690 8256
rect 10746 8200 11426 8256
rect 11482 8200 11487 8256
rect 10685 8198 11487 8200
rect 10685 8195 10751 8198
rect 11421 8195 11487 8198
rect 12198 8196 12204 8260
rect 12268 8258 12274 8260
rect 17953 8258 18019 8261
rect 12268 8256 18019 8258
rect 12268 8200 17958 8256
rect 18014 8200 18019 8256
rect 12268 8198 18019 8200
rect 12268 8196 12274 8198
rect 17953 8195 18019 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 6453 8122 6519 8125
rect 2270 8120 6519 8122
rect 2270 8064 6458 8120
rect 6514 8064 6519 8120
rect 2270 8062 6519 8064
rect 6453 8059 6519 8062
rect 14089 8122 14155 8125
rect 15101 8122 15167 8125
rect 17401 8122 17467 8125
rect 14089 8120 17467 8122
rect 14089 8064 14094 8120
rect 14150 8064 15106 8120
rect 15162 8064 17406 8120
rect 17462 8064 17467 8120
rect 14089 8062 17467 8064
rect 14089 8059 14155 8062
rect 15101 8059 15167 8062
rect 17401 8059 17467 8062
rect 3325 7986 3391 7989
rect 4337 7986 4403 7989
rect 7833 7986 7899 7989
rect 3325 7984 7899 7986
rect 3325 7928 3330 7984
rect 3386 7928 4342 7984
rect 4398 7928 7838 7984
rect 7894 7928 7899 7984
rect 3325 7926 7899 7928
rect 3325 7923 3391 7926
rect 4337 7923 4403 7926
rect 7833 7923 7899 7926
rect 9673 7986 9739 7989
rect 19425 7986 19491 7989
rect 9673 7984 19491 7986
rect 9673 7928 9678 7984
rect 9734 7928 19430 7984
rect 19486 7928 19491 7984
rect 9673 7926 19491 7928
rect 9673 7923 9739 7926
rect 19425 7923 19491 7926
rect 0 7850 480 7880
rect 3785 7850 3851 7853
rect 0 7848 3851 7850
rect 0 7792 3790 7848
rect 3846 7792 3851 7848
rect 0 7790 3851 7792
rect 0 7760 480 7790
rect 3785 7787 3851 7790
rect 3969 7850 4035 7853
rect 8661 7850 8727 7853
rect 3969 7848 8727 7850
rect 3969 7792 3974 7848
rect 4030 7792 8666 7848
rect 8722 7792 8727 7848
rect 3969 7790 8727 7792
rect 3969 7787 4035 7790
rect 8661 7787 8727 7790
rect 9305 7850 9371 7853
rect 19609 7850 19675 7853
rect 9305 7848 19675 7850
rect 9305 7792 9310 7848
rect 9366 7792 19614 7848
rect 19670 7792 19675 7848
rect 9305 7790 19675 7792
rect 9305 7787 9371 7790
rect 19609 7787 19675 7790
rect 7097 7714 7163 7717
rect 14733 7714 14799 7717
rect 7097 7712 14799 7714
rect 7097 7656 7102 7712
rect 7158 7656 14738 7712
rect 14794 7656 14799 7712
rect 7097 7654 14799 7656
rect 7097 7651 7163 7654
rect 14733 7651 14799 7654
rect 15377 7714 15443 7717
rect 20345 7714 20411 7717
rect 15377 7712 20411 7714
rect 15377 7656 15382 7712
rect 15438 7656 20350 7712
rect 20406 7656 20411 7712
rect 15377 7654 20411 7656
rect 15377 7651 15443 7654
rect 20345 7651 20411 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 6637 7578 6703 7581
rect 8661 7578 8727 7581
rect 14774 7578 14780 7580
rect 6637 7576 8218 7578
rect 6637 7520 6642 7576
rect 6698 7520 8218 7576
rect 6637 7518 8218 7520
rect 6637 7515 6703 7518
rect 1761 7442 1827 7445
rect 4521 7442 4587 7445
rect 1761 7440 4587 7442
rect 1761 7384 1766 7440
rect 1822 7384 4526 7440
rect 4582 7384 4587 7440
rect 1761 7382 4587 7384
rect 1761 7379 1827 7382
rect 4521 7379 4587 7382
rect 5165 7442 5231 7445
rect 7557 7442 7623 7445
rect 5165 7440 7623 7442
rect 5165 7384 5170 7440
rect 5226 7384 7562 7440
rect 7618 7384 7623 7440
rect 5165 7382 7623 7384
rect 8158 7442 8218 7518
rect 8661 7576 14780 7578
rect 8661 7520 8666 7576
rect 8722 7520 14780 7576
rect 8661 7518 14780 7520
rect 8661 7515 8727 7518
rect 14774 7516 14780 7518
rect 14844 7516 14850 7580
rect 20989 7442 21055 7445
rect 8158 7440 21055 7442
rect 8158 7384 20994 7440
rect 21050 7384 21055 7440
rect 8158 7382 21055 7384
rect 5165 7379 5231 7382
rect 7557 7379 7623 7382
rect 20989 7379 21055 7382
rect 0 7306 480 7336
rect 3918 7306 3924 7308
rect 0 7246 3924 7306
rect 0 7216 480 7246
rect 3918 7244 3924 7246
rect 3988 7244 3994 7308
rect 6821 7306 6887 7309
rect 12341 7306 12407 7309
rect 18965 7306 19031 7309
rect 6821 7304 10794 7306
rect 6821 7248 6826 7304
rect 6882 7248 10794 7304
rect 6821 7246 10794 7248
rect 6821 7243 6887 7246
rect 10133 7170 10199 7173
rect 2776 7168 10199 7170
rect 2776 7112 10138 7168
rect 10194 7112 10199 7168
rect 2776 7110 10199 7112
rect 10734 7170 10794 7246
rect 12341 7304 19031 7306
rect 12341 7248 12346 7304
rect 12402 7248 18970 7304
rect 19026 7248 19031 7304
rect 12341 7246 19031 7248
rect 12341 7243 12407 7246
rect 18965 7243 19031 7246
rect 16113 7170 16179 7173
rect 10734 7168 16179 7170
rect 10734 7112 16118 7168
rect 16174 7112 16179 7168
rect 10734 7110 16179 7112
rect 2776 6898 2836 7110
rect 10133 7107 10199 7110
rect 16113 7107 16179 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 9581 7034 9647 7037
rect 17953 7034 18019 7037
rect 9581 7032 10196 7034
rect 9581 6976 9586 7032
rect 9642 6976 10196 7032
rect 9581 6974 10196 6976
rect 9581 6971 9647 6974
rect 2638 6838 2836 6898
rect 3969 6898 4035 6901
rect 8201 6898 8267 6901
rect 3969 6896 8267 6898
rect 3969 6840 3974 6896
rect 4030 6840 8206 6896
rect 8262 6840 8267 6896
rect 3969 6838 8267 6840
rect 10136 6898 10196 6974
rect 10734 7032 18019 7034
rect 10734 6976 17958 7032
rect 18014 6976 18019 7032
rect 10734 6974 18019 6976
rect 10734 6898 10794 6974
rect 17953 6971 18019 6974
rect 10136 6838 10794 6898
rect 16205 6898 16271 6901
rect 17309 6898 17375 6901
rect 16205 6896 17375 6898
rect 16205 6840 16210 6896
rect 16266 6840 17314 6896
rect 17370 6840 17375 6896
rect 16205 6838 17375 6840
rect 0 6762 480 6792
rect 2638 6762 2698 6838
rect 3969 6835 4035 6838
rect 8201 6835 8267 6838
rect 16205 6835 16271 6838
rect 17309 6835 17375 6838
rect 18689 6898 18755 6901
rect 20989 6898 21055 6901
rect 18689 6896 21055 6898
rect 18689 6840 18694 6896
rect 18750 6840 20994 6896
rect 21050 6840 21055 6896
rect 18689 6838 21055 6840
rect 18689 6835 18755 6838
rect 20989 6835 21055 6838
rect 0 6702 2698 6762
rect 5993 6762 6059 6765
rect 21173 6762 21239 6765
rect 5993 6760 21239 6762
rect 5993 6704 5998 6760
rect 6054 6704 21178 6760
rect 21234 6704 21239 6760
rect 5993 6702 21239 6704
rect 0 6672 480 6702
rect 5993 6699 6059 6702
rect 21173 6699 21239 6702
rect 16614 6564 16620 6628
rect 16684 6626 16690 6628
rect 17953 6626 18019 6629
rect 16684 6624 18019 6626
rect 16684 6568 17958 6624
rect 18014 6568 18019 6624
rect 16684 6566 18019 6568
rect 16684 6564 16690 6566
rect 17953 6563 18019 6566
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 7281 6490 7347 6493
rect 11145 6490 11211 6493
rect 7281 6488 11211 6490
rect 7281 6432 7286 6488
rect 7342 6432 11150 6488
rect 11206 6432 11211 6488
rect 7281 6430 11211 6432
rect 7281 6427 7347 6430
rect 11145 6427 11211 6430
rect 16665 6490 16731 6493
rect 19977 6490 20043 6493
rect 16665 6488 20043 6490
rect 16665 6432 16670 6488
rect 16726 6432 19982 6488
rect 20038 6432 20043 6488
rect 16665 6430 20043 6432
rect 16665 6427 16731 6430
rect 19977 6427 20043 6430
rect 20294 6428 20300 6492
rect 20364 6490 20370 6492
rect 20437 6490 20503 6493
rect 20364 6488 20503 6490
rect 20364 6432 20442 6488
rect 20498 6432 20503 6488
rect 20364 6430 20503 6432
rect 20364 6428 20370 6430
rect 20437 6427 20503 6430
rect 6821 6354 6887 6357
rect 10685 6354 10751 6357
rect 12893 6354 12959 6357
rect 6821 6352 10751 6354
rect 6821 6296 6826 6352
rect 6882 6296 10690 6352
rect 10746 6296 10751 6352
rect 6821 6294 10751 6296
rect 6821 6291 6887 6294
rect 10685 6291 10751 6294
rect 10918 6352 12959 6354
rect 10918 6296 12898 6352
rect 12954 6296 12959 6352
rect 10918 6294 12959 6296
rect 8017 6218 8083 6221
rect 10918 6218 10978 6294
rect 12893 6291 12959 6294
rect 8017 6216 10978 6218
rect 8017 6160 8022 6216
rect 8078 6160 10978 6216
rect 8017 6158 10978 6160
rect 12065 6218 12131 6221
rect 14825 6218 14891 6221
rect 12065 6216 14891 6218
rect 12065 6160 12070 6216
rect 12126 6160 14830 6216
rect 14886 6160 14891 6216
rect 12065 6158 14891 6160
rect 8017 6155 8083 6158
rect 12065 6155 12131 6158
rect 14825 6155 14891 6158
rect 0 6082 480 6112
rect 7281 6082 7347 6085
rect 9673 6082 9739 6085
rect 0 6080 9739 6082
rect 0 6024 7286 6080
rect 7342 6024 9678 6080
rect 9734 6024 9739 6080
rect 0 6022 9739 6024
rect 0 5992 480 6022
rect 7281 6019 7347 6022
rect 9673 6019 9739 6022
rect 11513 6082 11579 6085
rect 16757 6082 16823 6085
rect 11513 6080 16823 6082
rect 11513 6024 11518 6080
rect 11574 6024 16762 6080
rect 16818 6024 16823 6080
rect 11513 6022 16823 6024
rect 11513 6019 11579 6022
rect 16757 6019 16823 6022
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 4061 5946 4127 5949
rect 6913 5946 6979 5949
rect 4061 5944 6979 5946
rect 4061 5888 4066 5944
rect 4122 5888 6918 5944
rect 6974 5888 6979 5944
rect 4061 5886 6979 5888
rect 4061 5883 4127 5886
rect 6913 5883 6979 5886
rect 2405 5810 2471 5813
rect 5073 5810 5139 5813
rect 5390 5810 5396 5812
rect 2405 5808 4906 5810
rect 2405 5752 2410 5808
rect 2466 5752 4906 5808
rect 2405 5750 4906 5752
rect 2405 5747 2471 5750
rect 3918 5612 3924 5676
rect 3988 5674 3994 5676
rect 4061 5674 4127 5677
rect 3988 5672 4127 5674
rect 3988 5616 4066 5672
rect 4122 5616 4127 5672
rect 3988 5614 4127 5616
rect 4846 5674 4906 5750
rect 5073 5808 5396 5810
rect 5073 5752 5078 5808
rect 5134 5752 5396 5808
rect 5073 5750 5396 5752
rect 5073 5747 5139 5750
rect 5390 5748 5396 5750
rect 5460 5748 5466 5812
rect 6085 5810 6151 5813
rect 10685 5810 10751 5813
rect 6085 5808 10751 5810
rect 6085 5752 6090 5808
rect 6146 5752 10690 5808
rect 10746 5752 10751 5808
rect 6085 5750 10751 5752
rect 6085 5747 6151 5750
rect 10685 5747 10751 5750
rect 21398 5748 21404 5812
rect 21468 5810 21474 5812
rect 21541 5810 21607 5813
rect 21468 5808 21607 5810
rect 21468 5752 21546 5808
rect 21602 5752 21607 5808
rect 21468 5750 21607 5752
rect 21468 5748 21474 5750
rect 21541 5747 21607 5750
rect 9029 5674 9095 5677
rect 4846 5672 9095 5674
rect 4846 5616 9034 5672
rect 9090 5616 9095 5672
rect 4846 5614 9095 5616
rect 3988 5612 3994 5614
rect 4061 5611 4127 5614
rect 9029 5611 9095 5614
rect 11094 5612 11100 5676
rect 11164 5674 11170 5676
rect 11237 5674 11303 5677
rect 11164 5672 11303 5674
rect 11164 5616 11242 5672
rect 11298 5616 11303 5672
rect 11164 5614 11303 5616
rect 11164 5612 11170 5614
rect 11237 5611 11303 5614
rect 18045 5674 18111 5677
rect 21173 5674 21239 5677
rect 18045 5672 21239 5674
rect 18045 5616 18050 5672
rect 18106 5616 21178 5672
rect 21234 5616 21239 5672
rect 18045 5614 21239 5616
rect 18045 5611 18111 5614
rect 21173 5611 21239 5614
rect 0 5538 480 5568
rect 3049 5538 3115 5541
rect 0 5536 3115 5538
rect 0 5480 3054 5536
rect 3110 5480 3115 5536
rect 0 5478 3115 5480
rect 0 5448 480 5478
rect 3049 5475 3115 5478
rect 11094 5476 11100 5540
rect 11164 5538 11170 5540
rect 11329 5538 11395 5541
rect 11164 5536 11395 5538
rect 11164 5480 11334 5536
rect 11390 5480 11395 5536
rect 11164 5478 11395 5480
rect 11164 5476 11170 5478
rect 11329 5475 11395 5478
rect 16757 5538 16823 5541
rect 19517 5538 19583 5541
rect 16757 5536 19583 5538
rect 16757 5480 16762 5536
rect 16818 5480 19522 5536
rect 19578 5480 19583 5536
rect 16757 5478 19583 5480
rect 16757 5475 16823 5478
rect 19517 5475 19583 5478
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 15929 5402 15995 5405
rect 18045 5402 18111 5405
rect 15929 5400 18111 5402
rect 15929 5344 15934 5400
rect 15990 5344 18050 5400
rect 18106 5344 18111 5400
rect 15929 5342 18111 5344
rect 15929 5339 15995 5342
rect 18045 5339 18111 5342
rect 3601 5266 3667 5269
rect 19333 5266 19399 5269
rect 3601 5264 19399 5266
rect 3601 5208 3606 5264
rect 3662 5208 19338 5264
rect 19394 5208 19399 5264
rect 3601 5206 19399 5208
rect 3601 5203 3667 5206
rect 19333 5203 19399 5206
rect 2313 5130 2379 5133
rect 14549 5130 14615 5133
rect 1534 5128 2379 5130
rect 1534 5072 2318 5128
rect 2374 5072 2379 5128
rect 1534 5070 2379 5072
rect 0 4994 480 5024
rect 1534 4994 1594 5070
rect 2313 5067 2379 5070
rect 2454 5128 14615 5130
rect 2454 5072 14554 5128
rect 14610 5072 14615 5128
rect 2454 5070 14615 5072
rect 0 4934 1594 4994
rect 1853 4994 1919 4997
rect 2454 4994 2514 5070
rect 14549 5067 14615 5070
rect 14774 5068 14780 5132
rect 14844 5130 14850 5132
rect 18597 5130 18663 5133
rect 22369 5132 22435 5133
rect 14844 5128 18663 5130
rect 14844 5072 18602 5128
rect 18658 5072 18663 5128
rect 14844 5070 18663 5072
rect 14844 5068 14850 5070
rect 18597 5067 18663 5070
rect 22318 5068 22324 5132
rect 22388 5130 22435 5132
rect 22388 5128 22480 5130
rect 22430 5072 22480 5128
rect 22388 5070 22480 5072
rect 22388 5068 22435 5070
rect 22369 5067 22435 5068
rect 1853 4992 2514 4994
rect 1853 4936 1858 4992
rect 1914 4936 2514 4992
rect 1853 4934 2514 4936
rect 3325 4994 3391 4997
rect 7925 4994 7991 4997
rect 3325 4992 7991 4994
rect 3325 4936 3330 4992
rect 3386 4936 7930 4992
rect 7986 4936 7991 4992
rect 3325 4934 7991 4936
rect 0 4904 480 4934
rect 1853 4931 1919 4934
rect 3325 4931 3391 4934
rect 7925 4931 7991 4934
rect 11881 4994 11947 4997
rect 19057 4994 19123 4997
rect 11881 4992 19123 4994
rect 11881 4936 11886 4992
rect 11942 4936 19062 4992
rect 19118 4936 19123 4992
rect 11881 4934 19123 4936
rect 11881 4931 11947 4934
rect 19057 4931 19123 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 16389 4858 16455 4861
rect 18505 4858 18571 4861
rect 16389 4856 18571 4858
rect 16389 4800 16394 4856
rect 16450 4800 18510 4856
rect 18566 4800 18571 4856
rect 16389 4798 18571 4800
rect 16389 4795 16455 4798
rect 18505 4795 18571 4798
rect 4521 4722 4587 4725
rect 9857 4722 9923 4725
rect 14457 4722 14523 4725
rect 19149 4722 19215 4725
rect 4521 4720 14523 4722
rect 4521 4664 4526 4720
rect 4582 4664 9862 4720
rect 9918 4664 14462 4720
rect 14518 4664 14523 4720
rect 4521 4662 14523 4664
rect 4521 4659 4587 4662
rect 9857 4659 9923 4662
rect 14457 4659 14523 4662
rect 14598 4720 19215 4722
rect 14598 4664 19154 4720
rect 19210 4664 19215 4720
rect 14598 4662 19215 4664
rect 3877 4586 3943 4589
rect 11094 4586 11100 4588
rect 3877 4584 11100 4586
rect 3877 4528 3882 4584
rect 3938 4528 11100 4584
rect 3877 4526 11100 4528
rect 3877 4523 3943 4526
rect 11094 4524 11100 4526
rect 11164 4524 11170 4588
rect 11329 4586 11395 4589
rect 14598 4586 14658 4662
rect 19149 4659 19215 4662
rect 21909 4722 21975 4725
rect 27520 4722 28000 4752
rect 21909 4720 28000 4722
rect 21909 4664 21914 4720
rect 21970 4664 28000 4720
rect 21909 4662 28000 4664
rect 21909 4659 21975 4662
rect 27520 4632 28000 4662
rect 15745 4586 15811 4589
rect 11329 4584 14658 4586
rect 11329 4528 11334 4584
rect 11390 4528 14658 4584
rect 11329 4526 14658 4528
rect 14782 4584 15811 4586
rect 14782 4528 15750 4584
rect 15806 4528 15811 4584
rect 14782 4526 15811 4528
rect 11329 4523 11395 4526
rect 0 4450 480 4480
rect 1117 4450 1183 4453
rect 0 4448 1183 4450
rect 0 4392 1122 4448
rect 1178 4392 1183 4448
rect 0 4390 1183 4392
rect 0 4360 480 4390
rect 1117 4387 1183 4390
rect 5993 4450 6059 4453
rect 7741 4450 7807 4453
rect 14782 4450 14842 4526
rect 15745 4523 15811 4526
rect 16297 4586 16363 4589
rect 20161 4586 20227 4589
rect 16297 4584 20227 4586
rect 16297 4528 16302 4584
rect 16358 4528 20166 4584
rect 20222 4528 20227 4584
rect 16297 4526 20227 4528
rect 16297 4523 16363 4526
rect 20161 4523 20227 4526
rect 5993 4448 14842 4450
rect 5993 4392 5998 4448
rect 6054 4392 7746 4448
rect 7802 4392 14842 4448
rect 5993 4390 14842 4392
rect 15377 4450 15443 4453
rect 18137 4450 18203 4453
rect 19333 4450 19399 4453
rect 15377 4448 19399 4450
rect 15377 4392 15382 4448
rect 15438 4392 18142 4448
rect 18198 4392 19338 4448
rect 19394 4392 19399 4448
rect 15377 4390 19399 4392
rect 5993 4387 6059 4390
rect 7741 4387 7807 4390
rect 15377 4387 15443 4390
rect 18137 4387 18203 4390
rect 19333 4387 19399 4390
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 1945 4178 2011 4181
rect 2313 4178 2379 4181
rect 1945 4176 2379 4178
rect 1945 4120 1950 4176
rect 2006 4120 2318 4176
rect 2374 4120 2379 4176
rect 1945 4118 2379 4120
rect 1945 4115 2011 4118
rect 2313 4115 2379 4118
rect 8845 4178 8911 4181
rect 17677 4178 17743 4181
rect 8845 4176 17743 4178
rect 8845 4120 8850 4176
rect 8906 4120 17682 4176
rect 17738 4120 17743 4176
rect 8845 4118 17743 4120
rect 8845 4115 8911 4118
rect 17677 4115 17743 4118
rect 18505 4178 18571 4181
rect 19425 4178 19491 4181
rect 18505 4176 19491 4178
rect 18505 4120 18510 4176
rect 18566 4120 19430 4176
rect 19486 4120 19491 4176
rect 18505 4118 19491 4120
rect 18505 4115 18571 4118
rect 19425 4115 19491 4118
rect 2037 4042 2103 4045
rect 3877 4042 3943 4045
rect 2037 4040 3943 4042
rect 2037 3984 2042 4040
rect 2098 3984 3882 4040
rect 3938 3984 3943 4040
rect 2037 3982 3943 3984
rect 2037 3979 2103 3982
rect 3877 3979 3943 3982
rect 6821 4042 6887 4045
rect 10685 4042 10751 4045
rect 6821 4040 10751 4042
rect 6821 3984 6826 4040
rect 6882 3984 10690 4040
rect 10746 3984 10751 4040
rect 6821 3982 10751 3984
rect 6821 3979 6887 3982
rect 10685 3979 10751 3982
rect 3417 3906 3483 3909
rect 7373 3906 7439 3909
rect 3417 3904 7439 3906
rect 3417 3848 3422 3904
rect 3478 3848 7378 3904
rect 7434 3848 7439 3904
rect 3417 3846 7439 3848
rect 3417 3843 3483 3846
rect 7373 3843 7439 3846
rect 12157 3906 12223 3909
rect 13353 3906 13419 3909
rect 12157 3904 13419 3906
rect 12157 3848 12162 3904
rect 12218 3848 13358 3904
rect 13414 3848 13419 3904
rect 12157 3846 13419 3848
rect 12157 3843 12223 3846
rect 13353 3843 13419 3846
rect 15745 3906 15811 3909
rect 17861 3906 17927 3909
rect 15745 3904 17927 3906
rect 15745 3848 15750 3904
rect 15806 3848 17866 3904
rect 17922 3848 17927 3904
rect 15745 3846 17927 3848
rect 15745 3843 15811 3846
rect 17861 3843 17927 3846
rect 20069 3906 20135 3909
rect 26509 3906 26575 3909
rect 20069 3904 26575 3906
rect 20069 3848 20074 3904
rect 20130 3848 26514 3904
rect 26570 3848 26575 3904
rect 20069 3846 26575 3848
rect 20069 3843 20135 3846
rect 26509 3843 26575 3846
rect 10277 3840 10597 3841
rect 0 3770 480 3800
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 3049 3770 3115 3773
rect 0 3768 3115 3770
rect 0 3712 3054 3768
rect 3110 3712 3115 3768
rect 0 3710 3115 3712
rect 0 3680 480 3710
rect 3049 3707 3115 3710
rect 3785 3770 3851 3773
rect 6085 3770 6151 3773
rect 3785 3768 6151 3770
rect 3785 3712 3790 3768
rect 3846 3712 6090 3768
rect 6146 3712 6151 3768
rect 3785 3710 6151 3712
rect 3785 3707 3851 3710
rect 6085 3707 6151 3710
rect 12709 3768 12775 3773
rect 12709 3712 12714 3768
rect 12770 3712 12775 3768
rect 12709 3707 12775 3712
rect 13629 3772 13695 3773
rect 13629 3768 13676 3772
rect 13740 3770 13746 3772
rect 16757 3770 16823 3773
rect 19333 3770 19399 3773
rect 13629 3712 13634 3768
rect 13629 3708 13676 3712
rect 13740 3710 13786 3770
rect 16757 3768 19399 3770
rect 16757 3712 16762 3768
rect 16818 3712 19338 3768
rect 19394 3712 19399 3768
rect 16757 3710 19399 3712
rect 13740 3708 13746 3710
rect 13629 3707 13695 3708
rect 16757 3707 16823 3710
rect 19333 3707 19399 3710
rect 23422 3708 23428 3772
rect 23492 3770 23498 3772
rect 24117 3770 24183 3773
rect 23492 3768 24183 3770
rect 23492 3712 24122 3768
rect 24178 3712 24183 3768
rect 23492 3710 24183 3712
rect 23492 3708 23498 3710
rect 24117 3707 24183 3710
rect 9397 3634 9463 3637
rect 12712 3634 12772 3707
rect 9397 3632 12772 3634
rect 9397 3576 9402 3632
rect 9458 3576 12772 3632
rect 9397 3574 12772 3576
rect 13629 3634 13695 3637
rect 19149 3634 19215 3637
rect 13629 3632 19215 3634
rect 13629 3576 13634 3632
rect 13690 3576 19154 3632
rect 19210 3576 19215 3632
rect 13629 3574 19215 3576
rect 9397 3571 9463 3574
rect 13629 3571 13695 3574
rect 19149 3571 19215 3574
rect 19517 3634 19583 3637
rect 27613 3634 27679 3637
rect 19517 3632 27679 3634
rect 19517 3576 19522 3632
rect 19578 3576 27618 3632
rect 27674 3576 27679 3632
rect 19517 3574 27679 3576
rect 19517 3571 19583 3574
rect 27613 3571 27679 3574
rect 6729 3498 6795 3501
rect 9305 3498 9371 3501
rect 4708 3438 6562 3498
rect 4708 3365 4768 3438
rect 1393 3362 1459 3365
rect 2589 3362 2655 3365
rect 4705 3362 4771 3365
rect 1393 3360 4771 3362
rect 1393 3304 1398 3360
rect 1454 3304 2594 3360
rect 2650 3304 4710 3360
rect 4766 3304 4771 3360
rect 1393 3302 4771 3304
rect 6502 3362 6562 3438
rect 6729 3496 9371 3498
rect 6729 3440 6734 3496
rect 6790 3440 9310 3496
rect 9366 3440 9371 3496
rect 6729 3438 9371 3440
rect 6729 3435 6795 3438
rect 9305 3435 9371 3438
rect 12709 3498 12775 3501
rect 16297 3498 16363 3501
rect 12709 3496 16363 3498
rect 12709 3440 12714 3496
rect 12770 3440 16302 3496
rect 16358 3440 16363 3496
rect 12709 3438 16363 3440
rect 12709 3435 12775 3438
rect 16297 3435 16363 3438
rect 17401 3498 17467 3501
rect 22001 3498 22067 3501
rect 17401 3496 22067 3498
rect 17401 3440 17406 3496
rect 17462 3440 22006 3496
rect 22062 3440 22067 3496
rect 17401 3438 22067 3440
rect 17401 3435 17467 3438
rect 22001 3435 22067 3438
rect 11513 3362 11579 3365
rect 6502 3360 11579 3362
rect 6502 3304 11518 3360
rect 11574 3304 11579 3360
rect 6502 3302 11579 3304
rect 1393 3299 1459 3302
rect 2589 3299 2655 3302
rect 4705 3299 4771 3302
rect 11513 3299 11579 3302
rect 16757 3362 16823 3365
rect 21817 3362 21883 3365
rect 16757 3360 21883 3362
rect 16757 3304 16762 3360
rect 16818 3304 21822 3360
rect 21878 3304 21883 3360
rect 16757 3302 21883 3304
rect 16757 3299 16823 3302
rect 21817 3299 21883 3302
rect 5610 3296 5930 3297
rect 0 3226 480 3256
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 3693 3226 3759 3229
rect 0 3224 3759 3226
rect 0 3168 3698 3224
rect 3754 3168 3759 3224
rect 0 3166 3759 3168
rect 0 3136 480 3166
rect 3693 3163 3759 3166
rect 8753 3226 8819 3229
rect 12985 3226 13051 3229
rect 20713 3228 20779 3229
rect 8753 3224 13051 3226
rect 8753 3168 8758 3224
rect 8814 3168 12990 3224
rect 13046 3168 13051 3224
rect 8753 3166 13051 3168
rect 8753 3163 8819 3166
rect 12985 3163 13051 3166
rect 20662 3164 20668 3228
rect 20732 3226 20779 3228
rect 20732 3224 20824 3226
rect 20774 3168 20824 3224
rect 20732 3166 20824 3168
rect 20732 3164 20779 3166
rect 20713 3163 20779 3164
rect 2865 3090 2931 3093
rect 2998 3090 3004 3092
rect 2865 3088 3004 3090
rect 2865 3032 2870 3088
rect 2926 3032 3004 3088
rect 2865 3030 3004 3032
rect 2865 3027 2931 3030
rect 2998 3028 3004 3030
rect 3068 3028 3074 3092
rect 3141 3090 3207 3093
rect 5625 3090 5691 3093
rect 7465 3092 7531 3093
rect 3141 3088 5691 3090
rect 3141 3032 3146 3088
rect 3202 3032 5630 3088
rect 5686 3032 5691 3088
rect 3141 3030 5691 3032
rect 3141 3027 3207 3030
rect 5625 3027 5691 3030
rect 7414 3028 7420 3092
rect 7484 3090 7531 3092
rect 11605 3090 11671 3093
rect 16205 3090 16271 3093
rect 17585 3092 17651 3093
rect 7484 3088 7576 3090
rect 7526 3032 7576 3088
rect 7484 3030 7576 3032
rect 11605 3088 16271 3090
rect 11605 3032 11610 3088
rect 11666 3032 16210 3088
rect 16266 3032 16271 3088
rect 11605 3030 16271 3032
rect 7484 3028 7531 3030
rect 7465 3027 7531 3028
rect 11605 3027 11671 3030
rect 16205 3027 16271 3030
rect 17534 3028 17540 3092
rect 17604 3090 17651 3092
rect 19517 3090 19583 3093
rect 25957 3090 26023 3093
rect 17604 3088 17696 3090
rect 17646 3032 17696 3088
rect 17604 3030 17696 3032
rect 19517 3088 26023 3090
rect 19517 3032 19522 3088
rect 19578 3032 25962 3088
rect 26018 3032 26023 3088
rect 19517 3030 26023 3032
rect 17604 3028 17651 3030
rect 17585 3027 17651 3028
rect 19517 3027 19583 3030
rect 25957 3027 26023 3030
rect 2313 2954 2379 2957
rect 3693 2954 3759 2957
rect 8385 2954 8451 2957
rect 2313 2952 8451 2954
rect 2313 2896 2318 2952
rect 2374 2896 3698 2952
rect 3754 2896 8390 2952
rect 8446 2896 8451 2952
rect 2313 2894 8451 2896
rect 2313 2891 2379 2894
rect 3693 2891 3759 2894
rect 8385 2891 8451 2894
rect 8937 2954 9003 2957
rect 11145 2954 11211 2957
rect 8937 2952 11211 2954
rect 8937 2896 8942 2952
rect 8998 2896 11150 2952
rect 11206 2896 11211 2952
rect 8937 2894 11211 2896
rect 8937 2891 9003 2894
rect 11145 2891 11211 2894
rect 11421 2954 11487 2957
rect 17953 2954 18019 2957
rect 11421 2952 18019 2954
rect 11421 2896 11426 2952
rect 11482 2896 17958 2952
rect 18014 2896 18019 2952
rect 11421 2894 18019 2896
rect 11421 2891 11487 2894
rect 17953 2891 18019 2894
rect 19517 2954 19583 2957
rect 22185 2954 22251 2957
rect 19517 2952 22251 2954
rect 19517 2896 19522 2952
rect 19578 2896 22190 2952
rect 22246 2896 22251 2952
rect 19517 2894 22251 2896
rect 19517 2891 19583 2894
rect 22185 2891 22251 2894
rect 2497 2818 2563 2821
rect 8753 2818 8819 2821
rect 2497 2816 8819 2818
rect 2497 2760 2502 2816
rect 2558 2760 8758 2816
rect 8814 2760 8819 2816
rect 2497 2758 8819 2760
rect 2497 2755 2563 2758
rect 8753 2755 8819 2758
rect 12433 2818 12499 2821
rect 17861 2818 17927 2821
rect 12433 2816 17927 2818
rect 12433 2760 12438 2816
rect 12494 2760 17866 2816
rect 17922 2760 17927 2816
rect 12433 2758 17927 2760
rect 12433 2755 12499 2758
rect 17861 2755 17927 2758
rect 22001 2818 22067 2821
rect 24761 2818 24827 2821
rect 22001 2816 24827 2818
rect 22001 2760 22006 2816
rect 22062 2760 24766 2816
rect 24822 2760 24827 2816
rect 22001 2758 24827 2760
rect 22001 2755 22067 2758
rect 24761 2755 24827 2758
rect 10277 2752 10597 2753
rect 0 2682 480 2712
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 13077 2682 13143 2685
rect 19333 2682 19399 2685
rect 0 2622 674 2682
rect 0 2592 480 2622
rect 614 2546 674 2622
rect 13077 2680 19399 2682
rect 13077 2624 13082 2680
rect 13138 2624 19338 2680
rect 19394 2624 19399 2680
rect 13077 2622 19399 2624
rect 13077 2619 13143 2622
rect 19333 2619 19399 2622
rect 20161 2682 20227 2685
rect 22093 2682 22159 2685
rect 20161 2680 22159 2682
rect 20161 2624 20166 2680
rect 20222 2624 22098 2680
rect 22154 2624 22159 2680
rect 20161 2622 22159 2624
rect 20161 2619 20227 2622
rect 22093 2619 22159 2622
rect 3233 2546 3299 2549
rect 614 2544 3299 2546
rect 614 2488 3238 2544
rect 3294 2488 3299 2544
rect 614 2486 3299 2488
rect 3233 2483 3299 2486
rect 5257 2546 5323 2549
rect 11973 2546 12039 2549
rect 5257 2544 12039 2546
rect 5257 2488 5262 2544
rect 5318 2488 11978 2544
rect 12034 2488 12039 2544
rect 5257 2486 12039 2488
rect 5257 2483 5323 2486
rect 11973 2483 12039 2486
rect 12985 2546 13051 2549
rect 15837 2546 15903 2549
rect 18045 2546 18111 2549
rect 12985 2544 15762 2546
rect 12985 2488 12990 2544
rect 13046 2488 15762 2544
rect 12985 2486 15762 2488
rect 12985 2483 13051 2486
rect 3601 2410 3667 2413
rect 5349 2410 5415 2413
rect 3601 2408 5415 2410
rect 3601 2352 3606 2408
rect 3662 2352 5354 2408
rect 5410 2352 5415 2408
rect 3601 2350 5415 2352
rect 3601 2347 3667 2350
rect 5349 2347 5415 2350
rect 6361 2410 6427 2413
rect 7833 2410 7899 2413
rect 11237 2410 11303 2413
rect 6361 2408 11303 2410
rect 6361 2352 6366 2408
rect 6422 2352 7838 2408
rect 7894 2352 11242 2408
rect 11298 2352 11303 2408
rect 6361 2350 11303 2352
rect 6361 2347 6427 2350
rect 7833 2347 7899 2350
rect 11237 2347 11303 2350
rect 13537 2410 13603 2413
rect 15702 2410 15762 2486
rect 15837 2544 18111 2546
rect 15837 2488 15842 2544
rect 15898 2488 18050 2544
rect 18106 2488 18111 2544
rect 15837 2486 18111 2488
rect 15837 2483 15903 2486
rect 18045 2483 18111 2486
rect 19057 2546 19123 2549
rect 21173 2546 21239 2549
rect 19057 2544 21239 2546
rect 19057 2488 19062 2544
rect 19118 2488 21178 2544
rect 21234 2488 21239 2544
rect 19057 2486 21239 2488
rect 19057 2483 19123 2486
rect 21173 2483 21239 2486
rect 17033 2410 17099 2413
rect 13537 2408 15394 2410
rect 13537 2352 13542 2408
rect 13598 2352 15394 2408
rect 13537 2350 15394 2352
rect 15702 2408 17099 2410
rect 15702 2352 17038 2408
rect 17094 2352 17099 2408
rect 15702 2350 17099 2352
rect 13537 2347 13603 2350
rect 6085 2274 6151 2277
rect 11329 2274 11395 2277
rect 6085 2272 11395 2274
rect 6085 2216 6090 2272
rect 6146 2216 11334 2272
rect 11390 2216 11395 2272
rect 6085 2214 11395 2216
rect 15334 2274 15394 2350
rect 17033 2347 17099 2350
rect 17309 2410 17375 2413
rect 27061 2410 27127 2413
rect 17309 2408 27127 2410
rect 17309 2352 17314 2408
rect 17370 2352 27066 2408
rect 27122 2352 27127 2408
rect 17309 2350 27127 2352
rect 17309 2347 17375 2350
rect 27061 2347 27127 2350
rect 20713 2274 20779 2277
rect 15334 2272 20779 2274
rect 15334 2216 20718 2272
rect 20774 2216 20779 2272
rect 15334 2214 20779 2216
rect 6085 2211 6151 2214
rect 11329 2211 11395 2214
rect 20713 2211 20779 2214
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 841 2138 907 2141
rect 5165 2138 5231 2141
rect 841 2136 5231 2138
rect 841 2080 846 2136
rect 902 2080 5170 2136
rect 5226 2080 5231 2136
rect 841 2078 5231 2080
rect 841 2075 907 2078
rect 5165 2075 5231 2078
rect 16021 2138 16087 2141
rect 19885 2138 19951 2141
rect 16021 2136 19951 2138
rect 16021 2080 16026 2136
rect 16082 2080 19890 2136
rect 19946 2080 19951 2136
rect 16021 2078 19951 2080
rect 16021 2075 16087 2078
rect 19885 2075 19951 2078
rect 0 2002 480 2032
rect 4337 2002 4403 2005
rect 0 2000 4403 2002
rect 0 1944 4342 2000
rect 4398 1944 4403 2000
rect 0 1942 4403 1944
rect 0 1912 480 1942
rect 4337 1939 4403 1942
rect 12893 2002 12959 2005
rect 18321 2002 18387 2005
rect 12893 2000 18387 2002
rect 12893 1944 12898 2000
rect 12954 1944 18326 2000
rect 18382 1944 18387 2000
rect 12893 1942 18387 1944
rect 12893 1939 12959 1942
rect 18321 1939 18387 1942
rect 7649 1866 7715 1869
rect 15745 1866 15811 1869
rect 24025 1866 24091 1869
rect 7649 1864 15811 1866
rect 7649 1808 7654 1864
rect 7710 1808 15750 1864
rect 15806 1808 15811 1864
rect 7649 1806 15811 1808
rect 7649 1803 7715 1806
rect 15745 1803 15811 1806
rect 17174 1864 24091 1866
rect 17174 1808 24030 1864
rect 24086 1808 24091 1864
rect 17174 1806 24091 1808
rect 289 1730 355 1733
rect 11605 1730 11671 1733
rect 289 1728 11671 1730
rect 289 1672 294 1728
rect 350 1672 11610 1728
rect 11666 1672 11671 1728
rect 289 1670 11671 1672
rect 289 1667 355 1670
rect 11605 1667 11671 1670
rect 11881 1594 11947 1597
rect 17174 1594 17234 1806
rect 24025 1803 24091 1806
rect 11881 1592 17234 1594
rect 11881 1536 11886 1592
rect 11942 1536 17234 1592
rect 11881 1534 17234 1536
rect 19057 1594 19123 1597
rect 23473 1594 23539 1597
rect 19057 1592 23539 1594
rect 19057 1536 19062 1592
rect 19118 1536 23478 1592
rect 23534 1536 23539 1592
rect 19057 1534 23539 1536
rect 11881 1531 11947 1534
rect 19057 1531 19123 1534
rect 23473 1531 23539 1534
rect 0 1458 480 1488
rect 4889 1458 4955 1461
rect 0 1456 4955 1458
rect 0 1400 4894 1456
rect 4950 1400 4955 1456
rect 0 1398 4955 1400
rect 0 1368 480 1398
rect 4889 1395 4955 1398
rect 0 914 480 944
rect 1301 914 1367 917
rect 0 912 1367 914
rect 0 856 1306 912
rect 1362 856 1367 912
rect 0 854 1367 856
rect 0 824 480 854
rect 1301 851 1367 854
rect 0 370 480 400
rect 3366 370 3372 372
rect 0 310 3372 370
rect 0 280 480 310
rect 3366 308 3372 310
rect 3436 308 3442 372
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 3556 17368 3620 17372
rect 3556 17312 3570 17368
rect 3570 17312 3620 17368
rect 3556 17308 3620 17312
rect 16436 17308 16500 17372
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 14596 14452 14660 14516
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 3372 13092 3436 13156
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 14228 12336 14292 12340
rect 14228 12280 14278 12336
rect 14278 12280 14292 12336
rect 14228 12276 14292 12280
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 14596 11732 14660 11796
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 11100 11052 11164 11116
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 3924 9692 3988 9756
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 14228 9692 14292 9756
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 12204 9012 12268 9076
rect 6316 8800 6380 8804
rect 6316 8744 6330 8800
rect 6330 8744 6380 8800
rect 6316 8740 6380 8744
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 12204 8196 12268 8260
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 14780 7516 14844 7580
rect 3924 7244 3988 7308
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 16620 6564 16684 6628
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 20300 6428 20364 6492
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 3924 5612 3988 5676
rect 5396 5748 5460 5812
rect 21404 5748 21468 5812
rect 11100 5612 11164 5676
rect 11100 5476 11164 5540
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 14780 5068 14844 5132
rect 22324 5128 22388 5132
rect 22324 5072 22374 5128
rect 22374 5072 22388 5128
rect 22324 5068 22388 5072
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 11100 4524 11164 4588
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 13676 3768 13740 3772
rect 13676 3712 13690 3768
rect 13690 3712 13740 3768
rect 13676 3708 13740 3712
rect 23428 3708 23492 3772
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 20668 3224 20732 3228
rect 20668 3168 20718 3224
rect 20718 3168 20732 3224
rect 20668 3164 20732 3168
rect 3004 3028 3068 3092
rect 7420 3088 7484 3092
rect 7420 3032 7470 3088
rect 7470 3032 7484 3088
rect 7420 3028 7484 3032
rect 17540 3088 17604 3092
rect 17540 3032 17590 3088
rect 17590 3032 17604 3088
rect 17540 3028 17604 3032
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
rect 3372 308 3436 372
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 3371 13156 3437 13157
rect 3371 13092 3372 13156
rect 3436 13092 3437 13156
rect 3371 13091 3437 13092
rect 3374 373 3434 13091
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 3923 9756 3989 9757
rect 3923 9692 3924 9756
rect 3988 9692 3989 9756
rect 3923 9691 3989 9692
rect 3926 7309 3986 9691
rect 5610 8736 5931 9760
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14595 14516 14661 14517
rect 14595 14452 14596 14516
rect 14660 14452 14661 14516
rect 14595 14451 14661 14452
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 14227 12340 14293 12341
rect 14227 12276 14228 12340
rect 14292 12276 14293 12340
rect 14227 12275 14293 12276
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 11099 11116 11165 11117
rect 11099 11052 11100 11116
rect 11164 11052 11165 11116
rect 11099 11051 11165 11052
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 6318 8805 6378 9062
rect 6315 8804 6381 8805
rect 6315 8740 6316 8804
rect 6380 8740 6381 8804
rect 6315 8739 6381 8740
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 3923 7308 3989 7309
rect 3923 7244 3924 7308
rect 3988 7244 3989 7308
rect 3923 7243 3989 7244
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 3923 5676 3989 5677
rect 3923 5612 3924 5676
rect 3988 5612 3989 5676
rect 3923 5611 3989 5612
rect 3926 5218 3986 5611
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 11102 6578 11162 11051
rect 14230 9757 14290 12275
rect 14598 11797 14658 14451
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14595 11796 14661 11797
rect 14595 11732 14596 11796
rect 14660 11732 14661 11796
rect 14595 11731 14661 11732
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14227 9756 14293 9757
rect 14227 9692 14228 9756
rect 14292 9692 14293 9756
rect 14227 9691 14293 9692
rect 12203 9076 12269 9077
rect 12203 9012 12204 9076
rect 12268 9012 12269 9076
rect 12203 9011 12269 9012
rect 12206 8261 12266 9011
rect 14944 8736 15264 9760
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 12203 8260 12269 8261
rect 12203 8196 12204 8260
rect 12268 8196 12269 8260
rect 12203 8195 12269 8196
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14779 7580 14845 7581
rect 14779 7516 14780 7580
rect 14844 7516 14845 7580
rect 14779 7515 14845 7516
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 11102 5677 11162 6342
rect 11099 5676 11165 5677
rect 11099 5612 11100 5676
rect 11164 5612 11165 5676
rect 11099 5611 11165 5612
rect 11099 5540 11165 5541
rect 11099 5476 11100 5540
rect 11164 5476 11165 5540
rect 11099 5475 11165 5476
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 11102 4589 11162 5475
rect 14782 5133 14842 7515
rect 14944 6560 15264 7584
rect 16622 6629 16682 9062
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 16619 6628 16685 6629
rect 16619 6564 16620 6628
rect 16684 6564 16685 6628
rect 16619 6563 16685 6564
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14779 5132 14845 5133
rect 14779 5068 14780 5132
rect 14844 5068 14845 5132
rect 14779 5067 14845 5068
rect 11099 4588 11165 4589
rect 11099 4538 11100 4588
rect 11164 4538 11165 4588
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 19610 6016 19930 7040
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 2752 19930 3776
rect 20670 3229 20730 4302
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 20667 3228 20733 3229
rect 20667 3164 20668 3228
rect 20732 3164 20733 3228
rect 20667 3163 20733 3164
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
rect 3371 372 3437 373
rect 3371 308 3372 372
rect 3436 308 3437 372
rect 3371 307 3437 308
<< via4 >>
rect 3470 17372 3706 17458
rect 3470 17308 3556 17372
rect 3556 17308 3620 17372
rect 3620 17308 3706 17372
rect 3470 17222 3706 17308
rect 2918 3092 3154 3178
rect 2918 3028 3004 3092
rect 3004 3028 3068 3092
rect 3068 3028 3154 3092
rect 2918 2942 3154 3028
rect 16350 17372 16586 17458
rect 16350 17308 16436 17372
rect 16436 17308 16500 17372
rect 16500 17308 16586 17372
rect 16350 17222 16586 17308
rect 6230 9062 6466 9298
rect 5310 5812 5546 5898
rect 5310 5748 5396 5812
rect 5396 5748 5460 5812
rect 5460 5748 5546 5812
rect 5310 5662 5546 5748
rect 3838 4982 4074 5218
rect 16534 9062 16770 9298
rect 11014 6342 11250 6578
rect 11014 4524 11100 4538
rect 11100 4524 11164 4538
rect 11164 4524 11250 4538
rect 11014 4302 11250 4524
rect 7334 3092 7570 3178
rect 7334 3028 7420 3092
rect 7420 3028 7484 3092
rect 7484 3028 7570 3092
rect 7334 2942 7570 3028
rect 13590 3772 13826 3858
rect 13590 3708 13676 3772
rect 13676 3708 13740 3772
rect 13740 3708 13826 3772
rect 13590 3622 13826 3708
rect 20214 6492 20450 6578
rect 20214 6428 20300 6492
rect 20300 6428 20364 6492
rect 20364 6428 20450 6492
rect 20214 6342 20450 6428
rect 21318 5812 21554 5898
rect 21318 5748 21404 5812
rect 21404 5748 21468 5812
rect 21468 5748 21554 5812
rect 21318 5662 21554 5748
rect 22238 5132 22474 5218
rect 22238 5068 22324 5132
rect 22324 5068 22388 5132
rect 22388 5068 22474 5132
rect 22238 4982 22474 5068
rect 20582 4302 20818 4538
rect 17454 3092 17690 3178
rect 17454 3028 17540 3092
rect 17540 3028 17604 3092
rect 17604 3028 17690 3092
rect 17454 2942 17690 3028
rect 23342 3772 23578 3858
rect 23342 3708 23428 3772
rect 23428 3708 23492 3772
rect 23492 3708 23578 3772
rect 23342 3622 23578 3708
<< metal5 >>
rect 3428 17458 16628 17500
rect 3428 17222 3470 17458
rect 3706 17222 16350 17458
rect 16586 17222 16628 17458
rect 3428 17180 16628 17222
rect 6188 9298 16812 9340
rect 6188 9062 6230 9298
rect 6466 9062 16534 9298
rect 16770 9062 16812 9298
rect 6188 9020 16812 9062
rect 10972 6578 20492 6620
rect 10972 6342 11014 6578
rect 11250 6342 20214 6578
rect 20450 6342 20492 6578
rect 10972 6300 20492 6342
rect 5268 5898 21596 5940
rect 5268 5662 5310 5898
rect 5546 5662 21318 5898
rect 21554 5662 21596 5898
rect 5268 5620 21596 5662
rect 3796 5218 22516 5260
rect 3796 4982 3838 5218
rect 4074 4982 22238 5218
rect 22474 4982 22516 5218
rect 3796 4940 22516 4982
rect 10972 4538 20860 4580
rect 10972 4302 11014 4538
rect 11250 4302 20582 4538
rect 20818 4302 20860 4538
rect 10972 4260 20860 4302
rect 13548 3858 23620 3900
rect 13548 3622 13590 3858
rect 13826 3622 23342 3858
rect 23578 3622 23620 3858
rect 13548 3580 23620 3622
rect 2876 3178 17732 3220
rect 2876 2942 2918 3178
rect 3154 2942 7334 3178
rect 7570 2942 17454 3178
rect 17690 2942 17732 3178
rect 2876 2900 17732 2942
use sky130_fd_sc_hd__decap_4  FILLER_1_10 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2024 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7
timestamp 1604681595
transform 1 0 1748 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1472 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_1_16
timestamp 1604681595
transform 1 0 2576 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 2392 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2852 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23
timestamp 1604681595
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27
timestamp 1604681595
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35
timestamp 1604681595
transform 1 0 4324 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _043_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_38
timestamp 1604681595
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41
timestamp 1604681595
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_46
timestamp 1604681595
transform 1 0 5336 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_42
timestamp 1604681595
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 5520 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 5152 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1604681595
transform 1 0 5244 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1604681595
transform 1 0 5704 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1604681595
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_53
timestamp 1604681595
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1604681595
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58
timestamp 1604681595
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 7176 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 8740 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_81
timestamp 1604681595
transform 1 0 8556 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_85
timestamp 1604681595
transform 1 0 8924 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1604681595
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1604681595
transform 1 0 8924 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 9108 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l4_in_0_
timestamp 1604681595
transform 1 0 9292 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_102
timestamp 1604681595
transform 1 0 10488 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_98
timestamp 1604681595
transform 1 0 10120 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 10672 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 10304 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9844 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_1_112
timestamp 1604681595
transform 1 0 11408 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_114
timestamp 1604681595
transform 1 0 11592 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 10856 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_118
timestamp 1604681595
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_116
timestamp 1604681595
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1604681595
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120
timestamp 1604681595
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_125
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13156 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 12972 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 14168 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_140
timestamp 1604681595
transform 1 0 13984 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_144
timestamp 1604681595
transform 1 0 14352 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_142
timestamp 1604681595
transform 1 0 14168 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_146
timestamp 1604681595
transform 1 0 14536 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_151
timestamp 1604681595
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_148
timestamp 1604681595
transform 1 0 14720 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 14720 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_0_
timestamp 1604681595
transform 1 0 14904 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_163
timestamp 1604681595
transform 1 0 16100 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_159
timestamp 1604681595
transform 1 0 15732 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_165
timestamp 1604681595
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 15916 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16284 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_173
timestamp 1604681595
transform 1 0 17020 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_169
timestamp 1604681595
transform 1 0 16652 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1604681595
transform 1 0 16928 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16468 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _086_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 17112 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_178
timestamp 1604681595
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_179
timestamp 1604681595
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_182
timestamp 1604681595
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_3_
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_193
timestamp 1604681595
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_197
timestamp 1604681595
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_200
timestamp 1604681595
transform 1 0 19504 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_196
timestamp 1604681595
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 19320 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1604681595
transform 1 0 19412 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19044 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19596 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_207
timestamp 1604681595
transform 1 0 20148 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_208
timestamp 1604681595
transform 1 0 20240 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 19688 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1604681595
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_211
timestamp 1604681595
transform 1 0 20516 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_212
timestamp 1604681595
transform 1 0 20608 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20332 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1604681595
transform 1 0 20700 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1604681595
transform 1 0 20424 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_216
timestamp 1604681595
transform 1 0 20976 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 20792 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1604681595
transform 1 0 20884 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_219
timestamp 1604681595
transform 1 0 21252 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1604681595
transform 1 0 21528 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1604681595
transform 1 0 21436 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_223
timestamp 1604681595
transform 1 0 21620 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_226
timestamp 1604681595
transform 1 0 21896 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1604681595
transform 1 0 21804 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1604681595
transform 1 0 21712 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1604681595
transform 1 0 21988 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 22080 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_235 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 22724 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_231
timestamp 1604681595
transform 1 0 22356 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_238
timestamp 1604681595
transform 1 0 23000 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_234
timestamp 1604681595
transform 1 0 22632 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1604681595
transform 1 0 22540 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1604681595
transform 1 0 22816 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1604681595
transform 1 0 22264 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_243
timestamp 1604681595
transform 1 0 23460 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_246
timestamp 1604681595
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1604681595
transform 1 0 24012 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_245 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1604681595
transform 1 0 24564 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1604681595
transform 1 0 24380 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_257
timestamp 1604681595
transform 1 0 24748 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_269
timestamp 1604681595
transform 1 0 25852 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_257
timestamp 1604681595
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_269
timestamp 1604681595
transform 1 0 25852 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 1840 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 2208 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_7
timestamp 1604681595
transform 1 0 1748 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_10
timestamp 1604681595
transform 1 0 2024 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_23
timestamp 1604681595
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27
timestamp 1604681595
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 6716 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 6532 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 5980 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_51
timestamp 1604681595
transform 1 0 5796 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_55
timestamp 1604681595
transform 1 0 6164 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 8004 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 7820 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_67
timestamp 1604681595
transform 1 0 7268 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_71
timestamp 1604681595
transform 1 0 7636 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_84
timestamp 1604681595
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_88
timestamp 1604681595
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_102
timestamp 1604681595
transform 1 0 10488 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 11224 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 12420 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 10856 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_108
timestamp 1604681595
transform 1 0 11040 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_119
timestamp 1604681595
transform 1 0 12052 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_125
timestamp 1604681595
transform 1 0 12604 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_1_
timestamp 1604681595
transform 1 0 13340 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 13156 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 12788 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_129
timestamp 1604681595
transform 1 0 12972 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_142
timestamp 1604681595
transform 1 0 14168 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 14904 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 14536 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_148
timestamp 1604681595
transform 1 0 14720 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_152
timestamp 1604681595
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 17756 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17572 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 17204 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_173
timestamp 1604681595
transform 1 0 17020 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_177
timestamp 1604681595
transform 1 0 17388 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1604681595
transform 1 0 19320 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 18768 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 19136 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 19872 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 20240 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_190
timestamp 1604681595
transform 1 0 18584 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1604681595
transform 1 0 18952 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_202
timestamp 1604681595
transform 1 0 19688 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_206
timestamp 1604681595
transform 1 0 20056 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1604681595
transform 1 0 21988 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1604681595
transform 1 0 21804 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 21436 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_210
timestamp 1604681595
transform 1 0 20424 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_219
timestamp 1604681595
transform 1 0 21252 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_223
timestamp 1604681595
transform 1 0 21620 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_231
timestamp 1604681595
transform 1 0 22356 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_243
timestamp 1604681595
transform 1 0 23460 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_255
timestamp 1604681595
transform 1 0 24564 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_267
timestamp 1604681595
transform 1 0 25668 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_276
timestamp 1604681595
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1604681595
transform 1 0 1840 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 1656 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 2852 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_17
timestamp 1604681595
transform 1 0 2668 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 3404 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3220 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_21
timestamp 1604681595
transform 1 0 3036 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_34
timestamp 1604681595
transform 1 0 4232 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_40
timestamp 1604681595
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_3_
timestamp 1604681595
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_53
timestamp 1604681595
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1604681595
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 8740 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 8556 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 7820 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_71
timestamp 1604681595
transform 1 0 7636 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_75
timestamp 1604681595
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_79
timestamp 1604681595
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10672 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_102
timestamp 1604681595
transform 1 0 10488 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1604681595
transform 1 0 11224 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1604681595
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 11040 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_106
timestamp 1604681595
transform 1 0 10856 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_114
timestamp 1604681595
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_118
timestamp 1604681595
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 13800 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1604681595
transform 1 0 12972 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 13340 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_127
timestamp 1604681595
transform 1 0 12788 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_131
timestamp 1604681595
transform 1 0 13156 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_135
timestamp 1604681595
transform 1 0 13524 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 16192 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15824 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_157
timestamp 1604681595
transform 1 0 15548 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_162
timestamp 1604681595
transform 1 0 16008 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_175
timestamp 1604681595
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_179
timestamp 1604681595
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1604681595
transform 1 0 19596 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1604681595
transform 1 0 20148 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_193
timestamp 1604681595
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_197
timestamp 1604681595
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_205
timestamp 1604681595
transform 1 0 19964 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1604681595
transform 1 0 20700 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1604681595
transform 1 0 21804 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A
timestamp 1604681595
transform 1 0 21252 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1604681595
transform 1 0 21620 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 20516 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_209
timestamp 1604681595
transform 1 0 20332 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_217
timestamp 1604681595
transform 1 0 21068 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_221
timestamp 1604681595
transform 1 0 21436 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_229
timestamp 1604681595
transform 1 0 22172 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1604681595
transform 1 0 23644 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 22356 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_233
timestamp 1604681595
transform 1 0 22540 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_241
timestamp 1604681595
transform 1 0 23276 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_249
timestamp 1604681595
transform 1 0 24012 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1604681595
transform 1 0 24196 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_253
timestamp 1604681595
transform 1 0 24380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_265
timestamp 1604681595
transform 1 0 25484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1604681595
transform 1 0 1840 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2944 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 1564 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7
timestamp 1604681595
transform 1 0 1748 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_17
timestamp 1604681595
transform 1 0 2668 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 4232 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 3312 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3680 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_22
timestamp 1604681595
transform 1 0 3128 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1604681595
transform 1 0 3496 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_30
timestamp 1604681595
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_32
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 6808 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6164 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_53
timestamp 1604681595
transform 1 0 5980 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_57
timestamp 1604681595
transform 1 0 6348 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_61
timestamp 1604681595
transform 1 0 6716 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 7544 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 8556 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 7176 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_64
timestamp 1604681595
transform 1 0 6992 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_68
timestamp 1604681595
transform 1 0 7360 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_79
timestamp 1604681595
transform 1 0 8372 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_83
timestamp 1604681595
transform 1 0 8740 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_88
timestamp 1604681595
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_102
timestamp 1604681595
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 11592 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1604681595
transform 1 0 11224 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 12604 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_106
timestamp 1604681595
transform 1 0 10856 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_112
timestamp 1604681595
transform 1 0 11408 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_123
timestamp 1604681595
transform 1 0 12420 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_3_
timestamp 1604681595
transform 1 0 13156 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 14168 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 12972 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_127
timestamp 1604681595
transform 1 0 12788 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_140
timestamp 1604681595
transform 1 0 13984 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_144
timestamp 1604681595
transform 1 0 14352 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_152
timestamp 1604681595
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_148
timestamp 1604681595
transform 1 0 14720 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 14536 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 14904 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_161
timestamp 1604681595
transform 1 0 15916 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_157
timestamp 1604681595
transform 1 0 15548 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 15732 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 16284 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 18216 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_184
timestamp 1604681595
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18768 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 19780 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 18584 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 20148 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_188
timestamp 1604681595
transform 1 0 18400 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_201
timestamp 1604681595
transform 1 0 19596 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_205
timestamp 1604681595
transform 1 0 19964 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 20516 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_209
timestamp 1604681595
transform 1 0 20332 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_213
timestamp 1604681595
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_219
timestamp 1604681595
transform 1 0 21252 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 22356 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_237
timestamp 1604681595
transform 1 0 22908 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_249
timestamp 1604681595
transform 1 0 24012 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_261
timestamp 1604681595
transform 1 0 25116 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_273
timestamp 1604681595
transform 1 0 26220 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_276
timestamp 1604681595
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2944 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_1_
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2760 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 2392 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_12
timestamp 1604681595
transform 1 0 2208 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_16
timestamp 1604681595
transform 1 0 2576 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4048 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_29
timestamp 1604681595
transform 1 0 3772 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_34
timestamp 1604681595
transform 1 0 4232 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_40
timestamp 1604681595
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_2_
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_53
timestamp 1604681595
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1604681595
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 8556 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 8372 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_71
timestamp 1604681595
transform 1 0 7636 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_77
timestamp 1604681595
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 10488 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_100
timestamp 1604681595
transform 1 0 10304 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_104
timestamp 1604681595
transform 1 0 10672 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1604681595
transform 1 0 11224 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_2_
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 11040 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_114
timestamp 1604681595
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_118
timestamp 1604681595
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_6__A1
timestamp 1604681595
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_6__A0
timestamp 1604681595
transform 1 0 13800 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_6__S
timestamp 1604681595
transform 1 0 14168 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_132
timestamp 1604681595
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_136
timestamp 1604681595
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_140
timestamp 1604681595
transform 1 0 13984 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_144
timestamp 1604681595
transform 1 0 14352 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 14904 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 14720 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 15916 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 16284 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_159
timestamp 1604681595
transform 1 0 15732 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_163
timestamp 1604681595
transform 1 0 16100 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16468 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_173
timestamp 1604681595
transform 1 0 17020 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_177
timestamp 1604681595
transform 1 0 17388 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1604681595
transform 1 0 19596 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_193
timestamp 1604681595
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_197
timestamp 1604681595
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 21160 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 21896 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 20608 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_210
timestamp 1604681595
transform 1 0 20424 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_214
timestamp 1604681595
transform 1 0 20792 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_224
timestamp 1604681595
transform 1 0 21712 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_228
timestamp 1604681595
transform 1 0 22080 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_240
timestamp 1604681595
transform 1 0 23184 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_245
timestamp 1604681595
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_257
timestamp 1604681595
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_269
timestamp 1604681595
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 1472 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 1564 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_28
timestamp 1604681595
transform 1 0 3680 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_24
timestamp 1604681595
transform 1 0 3312 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_27
timestamp 1604681595
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_23
timestamp 1604681595
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 3864 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 3496 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_39
timestamp 1604681595
transform 1 0 4692 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_35
timestamp 1604681595
transform 1 0 4324 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 4508 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1604681595
transform 1 0 4048 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_41
timestamp 1604681595
transform 1 0 4876 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 4876 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_46
timestamp 1604681595
transform 1 0 5336 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 5152 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1604681595
transform 1 0 5060 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5612 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1604681595
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_52
timestamp 1604681595
transform 1 0 5888 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_58
timestamp 1604681595
transform 1 0 6440 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_3_
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_71
timestamp 1604681595
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_71
timestamp 1604681595
transform 1 0 7636 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_68
timestamp 1604681595
transform 1 0 7360 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_64
timestamp 1604681595
transform 1 0 6992 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_75
timestamp 1604681595
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 7820 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 8188 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_4_
timestamp 1604681595
transform 1 0 8004 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 8372 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_6_88
timestamp 1604681595
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_84
timestamp 1604681595
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l4_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_102
timestamp 1604681595
transform 1 0 10488 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_98
timestamp 1604681595
transform 1 0 10120 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_102
timestamp 1604681595
transform 1 0 10488 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 10304 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10672 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10672 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_114
timestamp 1604681595
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1604681595
transform 1 0 11224 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_106
timestamp 1604681595
transform 1 0 10856 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_110
timestamp 1604681595
transform 1 0 11224 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_106
timestamp 1604681595
transform 1 0 10856 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11040 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 11316 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1604681595
transform 1 0 11500 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_7_123
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_118
timestamp 1604681595
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_122
timestamp 1604681595
transform 1 0 12328 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 12512 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_130
timestamp 1604681595
transform 1 0 13064 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_127
timestamp 1604681595
transform 1 0 12788 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_126
timestamp 1604681595
transform 1 0 12696 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 12880 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 12880 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_6_
timestamp 1604681595
transform 1 0 13064 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13248 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_141
timestamp 1604681595
transform 1 0 14076 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_143
timestamp 1604681595
transform 1 0 14260 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_139
timestamp 1604681595
transform 1 0 13892 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 14076 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 14260 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_145
timestamp 1604681595
transform 1 0 14444 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_154
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1604681595
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_147
timestamp 1604681595
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14628 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 14812 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_162
timestamp 1604681595
transform 1 0 16008 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_158
timestamp 1604681595
transform 1 0 15640 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_165
timestamp 1604681595
transform 1 0 16284 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 15824 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 16192 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 15456 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_175
timestamp 1604681595
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_169
timestamp 1604681595
transform 1 0 16652 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16836 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16468 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_184
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_179
timestamp 1604681595
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 18308 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 17020 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_6_196
timestamp 1604681595
transform 1 0 19136 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_192
timestamp 1604681595
transform 1 0 18768 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 18952 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_208
timestamp 1604681595
transform 1 0 20240 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_208
timestamp 1604681595
transform 1 0 20240 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_204
timestamp 1604681595
transform 1 0 19872 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 19320 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1604681595
transform 1 0 20056 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1604681595
transform 1 0 19504 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 18492 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_7_212
timestamp 1604681595
transform 1 0 20608 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_215
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_212
timestamp 1604681595
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 20424 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21068 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 20424 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20792 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20976 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1604681595
transform 1 0 21804 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 21988 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_229
timestamp 1604681595
transform 1 0 22172 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_219
timestamp 1604681595
transform 1 0 21252 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_231
timestamp 1604681595
transform 1 0 22356 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_243
timestamp 1604681595
transform 1 0 23460 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_241
timestamp 1604681595
transform 1 0 23276 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_245
timestamp 1604681595
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_255
timestamp 1604681595
transform 1 0 24564 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_267
timestamp 1604681595
transform 1 0 25668 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_257
timestamp 1604681595
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_269
timestamp 1604681595
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_276
timestamp 1604681595
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1604681595
transform 1 0 2944 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_2_
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 2392 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 2760 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_12
timestamp 1604681595
transform 1 0 2208 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_16
timestamp 1604681595
transform 1 0 2576 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_23
timestamp 1604681595
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_27
timestamp 1604681595
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_39
timestamp 1604681595
transform 1 0 4692 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_36
timestamp 1604681595
transform 1 0 4416 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 4508 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 4876 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 5060 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_8_62
timestamp 1604681595
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1604681595
transform 1 0 7544 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 8556 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 6992 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 7360 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_66
timestamp 1604681595
transform 1 0 7176 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_79
timestamp 1604681595
transform 1 0 8372 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_83
timestamp 1604681595
transform 1 0 8740 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_87
timestamp 1604681595
transform 1 0 9108 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1604681595
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 12328 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 11592 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11960 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_112
timestamp 1604681595
transform 1 0 11408 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_116
timestamp 1604681595
transform 1 0 11776 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_120
timestamp 1604681595
transform 1 0 12144 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_124
timestamp 1604681595
transform 1 0 12512 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12880 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13892 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12696 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 14444 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_137
timestamp 1604681595
transform 1 0 13708 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_141
timestamp 1604681595
transform 1 0 14076 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_151
timestamp 1604681595
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_147
timestamp 1604681595
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14812 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_161
timestamp 1604681595
transform 1 0 15916 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_157
timestamp 1604681595
transform 1 0 15548 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1604681595
transform 1 0 15732 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1604681595
transform 1 0 16284 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 17848 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 17664 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17296 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_174
timestamp 1604681595
transform 1 0 17112 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_178
timestamp 1604681595
transform 1 0 17480 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 19780 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 20148 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_201
timestamp 1604681595
transform 1 0 19596 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_205
timestamp 1604681595
transform 1 0 19964 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 21160 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 21528 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 20516 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_209
timestamp 1604681595
transform 1 0 20332 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1604681595
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_215
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_220
timestamp 1604681595
transform 1 0 21344 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_224
timestamp 1604681595
transform 1 0 21712 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_236
timestamp 1604681595
transform 1 0 22816 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_248
timestamp 1604681595
transform 1 0 23920 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_260
timestamp 1604681595
transform 1 0 25024 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_272
timestamp 1604681595
transform 1 0 26128 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_276
timestamp 1604681595
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 2208 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 1564 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 2024 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_7
timestamp 1604681595
transform 1 0 1748 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 4140 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_31
timestamp 1604681595
transform 1 0 3956 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_35
timestamp 1604681595
transform 1 0 4324 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_40
timestamp 1604681595
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_2_
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_2_
timestamp 1604681595
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_53
timestamp 1604681595
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1604681595
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 8556 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_71
timestamp 1604681595
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_75
timestamp 1604681595
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_79
timestamp 1604681595
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_83
timestamp 1604681595
transform 1 0 8740 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 9200 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_5__A1
timestamp 1604681595
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 9016 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_5__S
timestamp 1604681595
transform 1 0 10212 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_97
timestamp 1604681595
transform 1 0 10028 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_101
timestamp 1604681595
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_5_
timestamp 1604681595
transform 1 0 10764 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12604 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_114
timestamp 1604681595
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_118
timestamp 1604681595
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_123
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13156 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14168 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12972 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_127
timestamp 1604681595
transform 1 0 12788 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_140
timestamp 1604681595
transform 1 0 13984 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_144
timestamp 1604681595
transform 1 0 14352 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 14720 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 14536 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 17204 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 16652 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 17020 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_167
timestamp 1604681595
transform 1 0 16468 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_171
timestamp 1604681595
transform 1 0 16836 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_178
timestamp 1604681595
transform 1 0 17480 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 19596 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_193
timestamp 1604681595
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_197
timestamp 1604681595
transform 1 0 19228 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1604681595
transform 1 0 21160 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 20608 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 20976 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_210
timestamp 1604681595
transform 1 0 20424 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_214
timestamp 1604681595
transform 1 0 20792 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_227
timestamp 1604681595
transform 1 0 21988 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_239
timestamp 1604681595
transform 1 0 23092 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_243
timestamp 1604681595
transform 1 0 23460 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_245
timestamp 1604681595
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_257
timestamp 1604681595
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_269
timestamp 1604681595
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_3_
timestamp 1604681595
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 1564 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_7
timestamp 1604681595
transform 1 0 1748 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_11
timestamp 1604681595
transform 1 0 2116 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_23
timestamp 1604681595
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1604681595
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_35
timestamp 1604681595
transform 1 0 4324 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_39
timestamp 1604681595
transform 1 0 4692 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4508 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 5244 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_10_43
timestamp 1604681595
transform 1 0 5060 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1604681595
transform 1 0 7728 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 7176 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 7544 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 8740 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_64
timestamp 1604681595
transform 1 0 6992 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_68
timestamp 1604681595
transform 1 0 7360 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_81
timestamp 1604681595
transform 1 0 8556 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10120 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_85
timestamp 1604681595
transform 1 0 8924 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1604681595
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_96
timestamp 1604681595
transform 1 0 9936 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_100
timestamp 1604681595
transform 1 0 10304 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_104
timestamp 1604681595
transform 1 0 10672 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11132 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_5__A0
timestamp 1604681595
transform 1 0 10764 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_107
timestamp 1604681595
transform 1 0 10948 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 13432 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13064 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_128
timestamp 1604681595
transform 1 0 12880 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_132
timestamp 1604681595
transform 1 0 13248 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_145
timestamp 1604681595
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_149
timestamp 1604681595
transform 1 0 14812 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_prog_clk_A
timestamp 1604681595
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_158
timestamp 1604681595
transform 1 0 15640 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 15824 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_162
timestamp 1604681595
transform 1 0 16008 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 16192 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_166
timestamp 1604681595
transform 1 0 16376 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 16652 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_2_
timestamp 1604681595
transform 1 0 19136 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 18584 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 20148 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 18952 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_188
timestamp 1604681595
transform 1 0 18400 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_192
timestamp 1604681595
transform 1 0 18768 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_205
timestamp 1604681595
transform 1 0 19964 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21160 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 20516 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_209
timestamp 1604681595
transform 1 0 20332 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_213
timestamp 1604681595
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_215
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_220
timestamp 1604681595
transform 1 0 21344 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_232
timestamp 1604681595
transform 1 0 22448 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_244
timestamp 1604681595
transform 1 0 23552 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_256
timestamp 1604681595
transform 1 0 24656 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_268 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 25760 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_274
timestamp 1604681595
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_276
timestamp 1604681595
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 1472 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 2484 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2852 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_13
timestamp 1604681595
transform 1 0 2300 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_17
timestamp 1604681595
transform 1 0 2668 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 4600 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 3036 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 4416 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_30
timestamp 1604681595
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_34
timestamp 1604681595
transform 1 0 4232 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1604681595
transform 1 0 6440 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 5612 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_47
timestamp 1604681595
transform 1 0 5428 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_51
timestamp 1604681595
transform 1 0 5796 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_55
timestamp 1604681595
transform 1 0 6164 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 8740 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_81
timestamp 1604681595
transform 1 0 8556 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9936 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 9752 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 9384 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_85
timestamp 1604681595
transform 1 0 8924 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_89
timestamp 1604681595
transform 1 0 9292 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_92
timestamp 1604681595
transform 1 0 9568 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1604681595
transform 1 0 12052 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_prog_clk_A
timestamp 1604681595
transform 1 0 11868 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 11500 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_105
timestamp 1604681595
transform 1 0 10764 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_111
timestamp 1604681595
transform 1 0 11316 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_115
timestamp 1604681595
transform 1 0 11684 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_123
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1604681595
transform 1 0 12696 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 13708 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 13524 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 13156 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_129
timestamp 1604681595
transform 1 0 12972 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_133
timestamp 1604681595
transform 1 0 13340 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l4_in_0_
timestamp 1604681595
transform 1 0 16192 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 16008 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 15640 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_156
timestamp 1604681595
transform 1 0 15456 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_160
timestamp 1604681595
transform 1 0 15824 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_173
timestamp 1604681595
transform 1 0 17020 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_177
timestamp 1604681595
transform 1 0 17388 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_1_
timestamp 1604681595
transform 1 0 19596 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 19044 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 19412 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_193
timestamp 1604681595
transform 1 0 18860 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_197
timestamp 1604681595
transform 1 0 19228 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21160 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20976 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 20608 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_210
timestamp 1604681595
transform 1 0 20424 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_214
timestamp 1604681595
transform 1 0 20792 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_227
timestamp 1604681595
transform 1 0 21988 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_239
timestamp 1604681595
transform 1 0 23092 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_243
timestamp 1604681595
transform 1 0 23460 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_245
timestamp 1604681595
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_257
timestamp 1604681595
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_269
timestamp 1604681595
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 3312 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3680 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_22
timestamp 1604681595
transform 1 0 3128 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1604681595
transform 1 0 3496 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_30
timestamp 1604681595
transform 1 0 3864 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_41
timestamp 1604681595
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_45
timestamp 1604681595
transform 1 0 5244 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 5060 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 5428 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk
timestamp 1604681595
transform 1 0 5612 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_52
timestamp 1604681595
transform 1 0 5888 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_56
timestamp 1604681595
transform 1 0 6256 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6072 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_60
timestamp 1604681595
transform 1 0 6624 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6440 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 7084 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_12_64
timestamp 1604681595
transform 1 0 6992 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1604681595
transform 1 0 10028 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 9108 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 9844 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_84
timestamp 1604681595
transform 1 0 8832 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_89
timestamp 1604681595
transform 1 0 9292 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_93
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_100
timestamp 1604681595
transform 1 0 10304 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 11132 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_12_106
timestamp 1604681595
transform 1 0 10856 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_3_
timestamp 1604681595
transform 1 0 13616 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 13432 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 13064 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_128
timestamp 1604681595
transform 1 0 12880 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_132
timestamp 1604681595
transform 1 0 13248 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_145
timestamp 1604681595
transform 1 0 14444 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_149
timestamp 1604681595
transform 1 0 14812 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_154
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_158
timestamp 1604681595
transform 1 0 15640 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 15456 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_164
timestamp 1604681595
transform 1 0 16192 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 16008 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 16376 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 16560 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_12_187
timestamp 1604681595
transform 1 0 18308 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_3_
timestamp 1604681595
transform 1 0 19044 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 20056 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 18492 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 18860 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_191
timestamp 1604681595
transform 1 0 18676 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_204
timestamp 1604681595
transform 1 0 19872 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_208
timestamp 1604681595
transform 1 0 20240 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21160 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 20424 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_212
timestamp 1604681595
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_215
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_220
timestamp 1604681595
transform 1 0 21344 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_232
timestamp 1604681595
transform 1 0 22448 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_244
timestamp 1604681595
transform 1 0 23552 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_256
timestamp 1604681595
transform 1 0 24656 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_268
timestamp 1604681595
transform 1 0 25760 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_274
timestamp 1604681595
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_276
timestamp 1604681595
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_7
timestamp 1604681595
transform 1 0 1748 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_9
timestamp 1604681595
transform 1 0 1932 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 1564 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_11
timestamp 1604681595
transform 1 0 2116 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_16
timestamp 1604681595
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_13
timestamp 1604681595
transform 1 0 2300 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_2_
timestamp 1604681595
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 2760 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_14_27
timestamp 1604681595
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_23
timestamp 1604681595
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_37
timestamp 1604681595
transform 1 0 4508 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4692 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_41
timestamp 1604681595
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_41
timestamp 1604681595
transform 1 0 4876 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_49
timestamp 1604681595
transform 1 0 5612 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_45
timestamp 1604681595
transform 1 0 5244 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_51
timestamp 1604681595
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 5060 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 5428 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 5060 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 5244 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_62
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1604681595
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_55
timestamp 1604681595
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 5704 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_14_69
timestamp 1604681595
transform 1 0 7452 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_66
timestamp 1604681595
transform 1 0 7176 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 7636 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 6992 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 7360 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1604681595
transform 1 0 7544 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_81
timestamp 1604681595
transform 1 0 8556 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_77
timestamp 1604681595
transform 1 0 8188 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_73
timestamp 1604681595
transform 1 0 7820 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_79
timestamp 1604681595
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 8372 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8004 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_83
timestamp 1604681595
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 8740 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_93
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_89
timestamp 1604681595
transform 1 0 9292 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1604681595
transform 1 0 8924 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 9108 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_2_
timestamp 1604681595
transform 1 0 9108 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_101
timestamp 1604681595
transform 1 0 10396 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_97
timestamp 1604681595
transform 1 0 10028 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_100
timestamp 1604681595
transform 1 0 10304 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_96
timestamp 1604681595
transform 1 0 9936 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10212 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9844 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 10120 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 10488 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10672 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 10488 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 11684 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1604681595
transform 1 0 11500 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_117
timestamp 1604681595
transform 1 0 11868 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_123
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_121
timestamp 1604681595
transform 1 0 12236 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_125
timestamp 1604681595
transform 1 0 12604 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_128
timestamp 1604681595
transform 1 0 12880 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 12696 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 13064 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 12788 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12972 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_142
timestamp 1604681595
transform 1 0 14168 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1604681595
transform 1 0 13800 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 14352 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 13984 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 13248 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_14_154
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_150
timestamp 1604681595
transform 1 0 14904 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_146
timestamp 1604681595
transform 1 0 14536 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_155
timestamp 1604681595
transform 1 0 15364 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_151
timestamp 1604681595
transform 1 0 14996 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14720 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_158
timestamp 1604681595
transform 1 0 15640 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_158
timestamp 1604681595
transform 1 0 15640 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 15824 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 15732 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_1_
timestamp 1604681595
transform 1 0 16008 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 15916 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_13_175
timestamp 1604681595
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_171
timestamp 1604681595
transform 1 0 16836 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 17020 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_186
timestamp 1604681595
transform 1 0 18216 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_180
timestamp 1604681595
transform 1 0 17664 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_179
timestamp 1604681595
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18400 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 19964 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 19412 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 19780 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_203
timestamp 1604681595
transform 1 0 19780 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_207
timestamp 1604681595
transform 1 0 20148 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1604681595
transform 1 0 19228 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_201
timestamp 1604681595
transform 1 0 19596 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_205
timestamp 1604681595
transform 1 0 19964 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_219
timestamp 1604681595
transform 1 0 21252 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1604681595
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_215
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_227
timestamp 1604681595
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_231
timestamp 1604681595
transform 1 0 22356 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_243
timestamp 1604681595
transform 1 0 23460 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_245
timestamp 1604681595
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_239
timestamp 1604681595
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_257
timestamp 1604681595
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_269
timestamp 1604681595
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_251
timestamp 1604681595
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_263
timestamp 1604681595
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_276
timestamp 1604681595
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 1564 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 2576 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 2944 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_14
timestamp 1604681595
transform 1 0 2392 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_18
timestamp 1604681595
transform 1 0 2760 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 3128 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_15_41
timestamp 1604681595
transform 1 0 4876 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_45
timestamp 1604681595
transform 1 0 5244 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 5060 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 5428 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1604681595
transform 1 0 5612 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_53
timestamp 1604681595
transform 1 0 5980 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_60
timestamp 1604681595
transform 1 0 6624 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_57
timestamp 1604681595
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6440 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8004 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7452 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_65
timestamp 1604681595
transform 1 0 7084 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_71
timestamp 1604681595
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 9660 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 9476 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9108 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_84
timestamp 1604681595
transform 1 0 8832 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_89
timestamp 1604681595
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_2_
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 11684 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_112
timestamp 1604681595
transform 1 0 11408 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_117
timestamp 1604681595
transform 1 0 11868 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_3_
timestamp 1604681595
transform 1 0 13984 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 13800 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_132
timestamp 1604681595
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_136
timestamp 1604681595
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_3_
timestamp 1604681595
transform 1 0 16284 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 15272 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_149
timestamp 1604681595
transform 1 0 14812 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_153
timestamp 1604681595
transform 1 0 15180 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_156
timestamp 1604681595
transform 1 0 15456 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_160
timestamp 1604681595
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_164
timestamp 1604681595
transform 1 0 16192 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_174
timestamp 1604681595
transform 1 0 17112 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_178
timestamp 1604681595
transform 1 0 17480 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1604681595
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_193
timestamp 1604681595
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_197
timestamp 1604681595
transform 1 0 19228 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_209
timestamp 1604681595
transform 1 0 20332 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_221
timestamp 1604681595
transform 1 0 21436 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_233
timestamp 1604681595
transform 1 0 22540 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_241
timestamp 1604681595
transform 1 0 23276 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_245
timestamp 1604681595
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_257
timestamp 1604681595
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_269
timestamp 1604681595
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1604681595
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 1564 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 1932 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_7
timestamp 1604681595
transform 1 0 1748 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_11
timestamp 1604681595
transform 1 0 2116 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_23
timestamp 1604681595
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1604681595
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_41
timestamp 1604681595
transform 1 0 4876 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 6440 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 5060 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1604681595
transform 1 0 5612 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 5980 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_45
timestamp 1604681595
transform 1 0 5244 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_51
timestamp 1604681595
transform 1 0 5796 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_55
timestamp 1604681595
transform 1 0 6164 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 8372 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 8740 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_77
timestamp 1604681595
transform 1 0 8188 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_81
timestamp 1604681595
transform 1 0 8556 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10672 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_85
timestamp 1604681595
transform 1 0 8924 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_89
timestamp 1604681595
transform 1 0 9292 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_102
timestamp 1604681595
transform 1 0 10488 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_2_
timestamp 1604681595
transform 1 0 11684 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 11500 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11132 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_106
timestamp 1604681595
transform 1 0 10856 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_111
timestamp 1604681595
transform 1 0 11316 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_124
timestamp 1604681595
transform 1 0 12512 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1604681595
transform 1 0 13248 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 12696 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 13064 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14260 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_128
timestamp 1604681595
transform 1 0 12880 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1604681595
transform 1 0 14076 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_145
timestamp 1604681595
transform 1 0 14444 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_2_
timestamp 1604681595
transform 1 0 16008 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 15824 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 14628 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 15456 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_149
timestamp 1604681595
transform 1 0 14812 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_154
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_158
timestamp 1604681595
transform 1 0 15640 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 17572 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 17020 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17388 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_171
timestamp 1604681595
transform 1 0 16836 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_175
timestamp 1604681595
transform 1 0 17204 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 18584 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_188
timestamp 1604681595
transform 1 0 18400 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_192
timestamp 1604681595
transform 1 0 18768 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_204
timestamp 1604681595
transform 1 0 19872 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_212
timestamp 1604681595
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_215
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_227
timestamp 1604681595
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_239
timestamp 1604681595
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_251
timestamp 1604681595
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_263
timestamp 1604681595
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_276
timestamp 1604681595
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 2024 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 1840 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_7
timestamp 1604681595
transform 1 0 1748 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_3_
timestamp 1604681595
transform 1 0 4508 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 4324 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 3956 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_29
timestamp 1604681595
transform 1 0 3772 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_33
timestamp 1604681595
transform 1 0 4140 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 5520 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_46
timestamp 1604681595
transform 1 0 5336 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_50
timestamp 1604681595
transform 1 0 5704 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_54
timestamp 1604681595
transform 1 0 6072 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1604681595
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_62
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 7452 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 6992 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_66
timestamp 1604681595
transform 1 0 7176 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9936 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_88
timestamp 1604681595
transform 1 0 9200 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_92
timestamp 1604681595
transform 1 0 9568 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_95
timestamp 1604681595
transform 1 0 9844 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_105
timestamp 1604681595
transform 1 0 10764 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 10948 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_109
timestamp 1604681595
transform 1 0 11132 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11316 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1604681595
transform 1 0 11500 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_117
timestamp 1604681595
transform 1 0 11868 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12052 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_123
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1604681595
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 13248 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 13064 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 12696 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_128
timestamp 1604681595
transform 1 0 12880 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_2_
timestamp 1604681595
transform 1 0 16100 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 15916 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 15548 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 15180 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_151
timestamp 1604681595
transform 1 0 14996 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_155
timestamp 1604681595
transform 1 0 15364 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_159
timestamp 1604681595
transform 1 0 15732 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 17112 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_172
timestamp 1604681595
transform 1 0 16928 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_176
timestamp 1604681595
transform 1 0 17296 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1604681595
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_187
timestamp 1604681595
transform 1 0 18308 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 18492 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_191
timestamp 1604681595
transform 1 0 18676 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_203
timestamp 1604681595
transform 1 0 19780 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_215
timestamp 1604681595
transform 1 0 20884 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_227
timestamp 1604681595
transform 1 0 21988 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_239
timestamp 1604681595
transform 1 0 23092 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_243
timestamp 1604681595
transform 1 0 23460 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_245
timestamp 1604681595
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_257
timestamp 1604681595
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_269
timestamp 1604681595
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 1472 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_23
timestamp 1604681595
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1604681595
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_41
timestamp 1604681595
transform 1 0 4876 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_45
timestamp 1604681595
transform 1 0 5244 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 5060 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 5428 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1604681595
transform 1 0 5612 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_52
timestamp 1604681595
transform 1 0 5888 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_56
timestamp 1604681595
transform 1 0 6256 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 6072 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_60
timestamp 1604681595
transform 1 0 6624 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 6440 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6992 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 8004 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 8372 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 8740 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_73
timestamp 1604681595
transform 1 0 7820 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_77
timestamp 1604681595
transform 1 0 8188 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_81
timestamp 1604681595
transform 1 0 8556 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_2_
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_85
timestamp 1604681595
transform 1 0 8924 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_89
timestamp 1604681595
transform 1 0 9292 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_102
timestamp 1604681595
transform 1 0 10488 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1604681595
transform 1 0 11316 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12420 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10764 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11132 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_107
timestamp 1604681595
transform 1 0 10948 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_120
timestamp 1604681595
transform 1 0 12144 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13432 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_132
timestamp 1604681595
transform 1 0 13248 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_145
timestamp 1604681595
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_149
timestamp 1604681595
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_157
timestamp 1604681595
transform 1 0 15548 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_161
timestamp 1604681595
transform 1 0 15916 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 15732 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_165
timestamp 1604681595
transform 1 0 16284 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 16560 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_18_187
timestamp 1604681595
transform 1 0 18308 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 18492 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 18860 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_191
timestamp 1604681595
transform 1 0 18676 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_195
timestamp 1604681595
transform 1 0 19044 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_207
timestamp 1604681595
transform 1 0 20148 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_213
timestamp 1604681595
transform 1 0 20700 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_215
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_227
timestamp 1604681595
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_239
timestamp 1604681595
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_251
timestamp 1604681595
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_263
timestamp 1604681595
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_276
timestamp 1604681595
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_7
timestamp 1604681595
transform 1 0 1748 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 1932 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 1564 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_11
timestamp 1604681595
transform 1 0 2116 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_16
timestamp 1604681595
transform 1 0 2576 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_12
timestamp 1604681595
transform 1 0 2208 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 2760 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2392 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 2944 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4876 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_39
timestamp 1604681595
transform 1 0 4692 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_23
timestamp 1604681595
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_27
timestamp 1604681595
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_41
timestamp 1604681595
transform 1 0 4876 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_45
timestamp 1604681595
transform 1 0 5244 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_43
timestamp 1604681595
transform 1 0 5060 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 5060 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 5244 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_47
timestamp 1604681595
transform 1 0 5428 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 5428 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1604681595
transform 1 0 5612 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1604681595
transform 1 0 5704 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_53
timestamp 1604681595
transform 1 0 5980 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_53
timestamp 1604681595
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1604681595
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_61
timestamp 1604681595
transform 1 0 6716 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_57
timestamp 1604681595
transform 1 0 6348 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1604681595
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 6532 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_62
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_71
timestamp 1604681595
transform 1 0 7636 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_67
timestamp 1604681595
transform 1 0 7268 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6900 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 7452 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l3_in_0_
timestamp 1604681595
transform 1 0 7084 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1604681595
transform 1 0 6992 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1604681595
transform 1 0 8648 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_78
timestamp 1604681595
transform 1 0 8280 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_74
timestamp 1604681595
transform 1 0 7912 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 8464 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 8096 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 7912 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 8096 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_20_90
timestamp 1604681595
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_86
timestamp 1604681595
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_99
timestamp 1604681595
transform 1 0 10212 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_95
timestamp 1604681595
transform 1 0 9844 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 10028 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_20_112
timestamp 1604681595
transform 1 0 11408 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_114
timestamp 1604681595
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 11592 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_125
timestamp 1604681595
transform 1 0 12604 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_120
timestamp 1604681595
transform 1 0 12144 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_116
timestamp 1604681595
transform 1 0 11776 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_118
timestamp 1604681595
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11960 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 14168 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 12788 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 14904 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 16100 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_161
timestamp 1604681595
transform 1 0 15916 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_165
timestamp 1604681595
transform 1 0 16284 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_147
timestamp 1604681595
transform 1 0 14628 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_152
timestamp 1604681595
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_173
timestamp 1604681595
transform 1 0 17020 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_175
timestamp 1604681595
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_171
timestamp 1604681595
transform 1 0 16836 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 17204 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 17020 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1604681595
transform 1 0 16560 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_177
timestamp 1604681595
transform 1 0 17388 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_179
timestamp 1604681595
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 17572 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_3_
timestamp 1604681595
transform 1 0 17756 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 18768 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_193
timestamp 1604681595
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_197
timestamp 1604681595
transform 1 0 19228 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_190
timestamp 1604681595
transform 1 0 18584 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_194
timestamp 1604681595
transform 1 0 18952 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_206
timestamp 1604681595
transform 1 0 20056 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_209
timestamp 1604681595
transform 1 0 20332 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_221
timestamp 1604681595
transform 1 0 21436 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_215
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_227
timestamp 1604681595
transform 1 0 21988 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 24104 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_233
timestamp 1604681595
transform 1 0 22540 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_241
timestamp 1604681595
transform 1 0 23276 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_245
timestamp 1604681595
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_239
timestamp 1604681595
transform 1 0 23092 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_247
timestamp 1604681595
transform 1 0 23828 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_257
timestamp 1604681595
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_269
timestamp 1604681595
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_252
timestamp 1604681595
transform 1 0 24288 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_264
timestamp 1604681595
transform 1 0 25392 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_272
timestamp 1604681595
transform 1 0 26128 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_276
timestamp 1604681595
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2944 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2392 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2760 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_12
timestamp 1604681595
transform 1 0 2208 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_16
timestamp 1604681595
transform 1 0 2576 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 4232 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 4048 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 3680 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_26
timestamp 1604681595
transform 1 0 3496 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_30
timestamp 1604681595
transform 1 0 3864 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_43
timestamp 1604681595
transform 1 0 5060 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_47
timestamp 1604681595
transform 1 0 5428 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 5244 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 5612 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_51
timestamp 1604681595
transform 1 0 5796 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_55
timestamp 1604681595
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1604681595
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_62
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 7544 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 6992 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 7360 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_66
timestamp 1604681595
transform 1 0 7176 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10580 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 9752 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_89
timestamp 1604681595
transform 1 0 9292 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_93
timestamp 1604681595
transform 1 0 9660 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_96
timestamp 1604681595
transform 1 0 9936 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_101
timestamp 1604681595
transform 1 0 10396 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10764 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_114
timestamp 1604681595
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1604681595
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 14352 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_142
timestamp 1604681595
transform 1 0 14168 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1604681595
transform 1 0 14904 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 14720 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15916 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 16284 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_146
timestamp 1604681595
transform 1 0 14536 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_159
timestamp 1604681595
transform 1 0 15732 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_163
timestamp 1604681595
transform 1 0 16100 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_167
timestamp 1604681595
transform 1 0 16468 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16652 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_171
timestamp 1604681595
transform 1 0 16836 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_175
timestamp 1604681595
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 17020 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_179
timestamp 1604681595
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_184
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 18216 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 18584 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_188
timestamp 1604681595
transform 1 0 18400 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_192
timestamp 1604681595
transform 1 0 18768 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_204
timestamp 1604681595
transform 1 0 19872 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_216
timestamp 1604681595
transform 1 0 20976 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_228
timestamp 1604681595
transform 1 0 22080 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 24104 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 23920 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_240
timestamp 1604681595
transform 1 0 23184 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_245
timestamp 1604681595
transform 1 0 23644 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_269
timestamp 1604681595
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 1840 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 2208 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_6
timestamp 1604681595
transform 1 0 1656 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_10
timestamp 1604681595
transform 1 0 2024 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 4140 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_23
timestamp 1604681595
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1604681595
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_32
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 6624 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6072 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6440 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_52
timestamp 1604681595
transform 1 0 5888 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_56
timestamp 1604681595
transform 1 0 6256 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 8556 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_79
timestamp 1604681595
transform 1 0 8372 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_83
timestamp 1604681595
transform 1 0 8740 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9752 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 8924 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9292 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_87
timestamp 1604681595
transform 1 0 9108 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_91
timestamp 1604681595
transform 1 0 9476 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_93
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_100
timestamp 1604681595
transform 1 0 10304 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_104
timestamp 1604681595
transform 1 0 10672 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1604681595
transform 1 0 12604 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l3_in_0_
timestamp 1604681595
transform 1 0 11040 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10764 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 12052 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 12420 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_107
timestamp 1604681595
transform 1 0 10948 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_117
timestamp 1604681595
transform 1 0 11868 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_121
timestamp 1604681595
transform 1 0 12236 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1604681595
transform 1 0 13616 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 13432 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 13064 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_128
timestamp 1604681595
transform 1 0 12880 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_132
timestamp 1604681595
transform 1 0 13248 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_145
timestamp 1604681595
transform 1 0 14444 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 14904 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_149
timestamp 1604681595
transform 1 0 14812 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_152
timestamp 1604681595
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_163
timestamp 1604681595
transform 1 0 16100 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 16928 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 16468 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_169
timestamp 1604681595
transform 1 0 16652 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 18860 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_191
timestamp 1604681595
transform 1 0 18676 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_195
timestamp 1604681595
transform 1 0 19044 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_207
timestamp 1604681595
transform 1 0 20148 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_213
timestamp 1604681595
transform 1 0 20700 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_215
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_227
timestamp 1604681595
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_239
timestamp 1604681595
transform 1 0 23092 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_251
timestamp 1604681595
transform 1 0 24196 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_263
timestamp 1604681595
transform 1 0 25300 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_276
timestamp 1604681595
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 1656 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4692 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 4508 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 4140 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3772 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_25
timestamp 1604681595
transform 1 0 3404 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_31
timestamp 1604681595
transform 1 0 3956 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_35
timestamp 1604681595
transform 1 0 4324 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 5796 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_48
timestamp 1604681595
transform 1 0 5520 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_53
timestamp 1604681595
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1604681595
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 8740 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 8556 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_71
timestamp 1604681595
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_75
timestamp 1604681595
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_79
timestamp 1604681595
transform 1 0 8372 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10672 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_102
timestamp 1604681595
transform 1 0 10488 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_106
timestamp 1604681595
transform 1 0 10856 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 11040 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1604681595
transform 1 0 11224 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_6__A1
timestamp 1604681595
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_114
timestamp 1604681595
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_118
timestamp 1604681595
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_6__A0
timestamp 1604681595
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_6__S
timestamp 1604681595
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_123
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_5__S
timestamp 1604681595
transform 1 0 12604 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 13616 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_5__A0
timestamp 1604681595
transform 1 0 12972 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_5__A1
timestamp 1604681595
transform 1 0 13340 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_127
timestamp 1604681595
transform 1 0 12788 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_131
timestamp 1604681595
transform 1 0 13156 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_135
timestamp 1604681595
transform 1 0 13524 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l4_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 16192 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 15824 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_155
timestamp 1604681595
transform 1 0 15364 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_159
timestamp 1604681595
transform 1 0 15732 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_162
timestamp 1604681595
transform 1 0 16008 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_175
timestamp 1604681595
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_179
timestamp 1604681595
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_203
timestamp 1604681595
transform 1 0 19780 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_215
timestamp 1604681595
transform 1 0 20884 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_227
timestamp 1604681595
transform 1 0 21988 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_239
timestamp 1604681595
transform 1 0 23092 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_243
timestamp 1604681595
transform 1 0 23460 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_245
timestamp 1604681595
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_257
timestamp 1604681595
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_269
timestamp 1604681595
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 2024 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 1656 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_8
timestamp 1604681595
transform 1 0 1840 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_12
timestamp 1604681595
transform 1 0 2208 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_23
timestamp 1604681595
transform 1 0 3220 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1604681595
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_41
timestamp 1604681595
transform 1 0 4876 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_3_
timestamp 1604681595
transform 1 0 6164 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 5152 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 5520 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 5888 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_46
timestamp 1604681595
transform 1 0 5336 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_50
timestamp 1604681595
transform 1 0 5704 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_54
timestamp 1604681595
transform 1 0 6072 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1604681595
transform 1 0 7728 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7176 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7544 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8740 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_64
timestamp 1604681595
transform 1 0 6992 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_68
timestamp 1604681595
transform 1 0 7360 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_81
timestamp 1604681595
transform 1 0 8556 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 9108 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1604681595
transform 1 0 8924 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_89
timestamp 1604681595
transform 1 0 9292 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_102
timestamp 1604681595
transform 1 0 10488 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_6_
timestamp 1604681595
transform 1 0 11408 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 11132 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 12420 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_106
timestamp 1604681595
transform 1 0 10856 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_111
timestamp 1604681595
transform 1 0 11316 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_121
timestamp 1604681595
transform 1 0 12236 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_125
timestamp 1604681595
transform 1 0 12604 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_5_
timestamp 1604681595
transform 1 0 12972 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13984 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 14352 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_prog_clk_A
timestamp 1604681595
transform 1 0 12788 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1604681595
transform 1 0 13800 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_142
timestamp 1604681595
transform 1 0 14168 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_150
timestamp 1604681595
transform 1 0 14904 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_146
timestamp 1604681595
transform 1 0 14536 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_154
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_158
timestamp 1604681595
transform 1 0 15640 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 15824 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15456 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_162
timestamp 1604681595
transform 1 0 16008 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 16284 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18032 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16468 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 17848 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 17480 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_176
timestamp 1604681595
transform 1 0 17296 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_180
timestamp 1604681595
transform 1 0 17664 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_193
timestamp 1604681595
transform 1 0 18860 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_205
timestamp 1604681595
transform 1 0 19964 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_213
timestamp 1604681595
transform 1 0 20700 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_215
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_227
timestamp 1604681595
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_239
timestamp 1604681595
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_251
timestamp 1604681595
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_263
timestamp 1604681595
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_276
timestamp 1604681595
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 2024 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 1840 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_7
timestamp 1604681595
transform 1 0 1748 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_19
timestamp 1604681595
transform 1 0 2852 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 3588 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 3404 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 3036 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 4600 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_23
timestamp 1604681595
transform 1 0 3220 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_36
timestamp 1604681595
transform 1 0 4416 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_40
timestamp 1604681595
transform 1 0 4784 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 5152 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 4968 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_53
timestamp 1604681595
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1604681595
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_62
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6992 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8556 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8372 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_73
timestamp 1604681595
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_77
timestamp 1604681595
transform 1 0 8188 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9568 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1604681595
transform 1 0 9936 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_90
timestamp 1604681595
transform 1 0 9384 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_94
timestamp 1604681595
transform 1 0 9752 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_98
timestamp 1604681595
transform 1 0 10120 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_102
timestamp 1604681595
transform 1 0 10488 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_2_
timestamp 1604681595
transform 1 0 10764 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_114
timestamp 1604681595
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_118
timestamp 1604681595
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_123
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13616 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13432 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13064 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12696 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_128
timestamp 1604681595
transform 1 0 12880 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_132
timestamp 1604681595
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_145
timestamp 1604681595
transform 1 0 14444 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 15180 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14628 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_149
timestamp 1604681595
transform 1 0 14812 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17112 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17480 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 18216 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_172
timestamp 1604681595
transform 1 0 16928 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_176
timestamp 1604681595
transform 1 0 17296 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_180
timestamp 1604681595
transform 1 0 17664 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_184
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_188
timestamp 1604681595
transform 1 0 18400 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_200
timestamp 1604681595
transform 1 0 19504 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_212
timestamp 1604681595
transform 1 0 20608 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_224
timestamp 1604681595
transform 1 0 21712 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_236
timestamp 1604681595
transform 1 0 22816 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_245
timestamp 1604681595
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_257
timestamp 1604681595
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_269
timestamp 1604681595
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_20
timestamp 1604681595
transform 1 0 2944 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_16
timestamp 1604681595
transform 1 0 2576 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_12
timestamp 1604681595
transform 1 0 2208 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2760 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2392 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 1472 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1604681595
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_23
timestamp 1604681595
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 3128 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_35
timestamp 1604681595
transform 1 0 4324 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_31
timestamp 1604681595
transform 1 0 3956 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_38
timestamp 1604681595
transform 1 0 4600 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4784 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 4508 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 4140 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4692 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_48
timestamp 1604681595
transform 1 0 5520 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_46
timestamp 1604681595
transform 1 0 5336 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_42
timestamp 1604681595
transform 1 0 4968 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 5704 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 5152 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_3_
timestamp 1604681595
transform 1 0 5428 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1604681595
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_52
timestamp 1604681595
transform 1 0 5888 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_60
timestamp 1604681595
transform 1 0 6624 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_56
timestamp 1604681595
transform 1 0 6256 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6440 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_2_
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_71
timestamp 1604681595
transform 1 0 7636 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_72
timestamp 1604681595
transform 1 0 7728 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_68
timestamp 1604681595
transform 1 0 7360 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_64
timestamp 1604681595
transform 1 0 6992 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 7544 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 7176 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_79
timestamp 1604681595
transform 1 0 8372 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_75
timestamp 1604681595
transform 1 0 8004 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1604681595
transform 1 0 8648 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8188 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 8556 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7820 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 8740 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_26_86
timestamp 1604681595
transform 1 0 9016 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9200 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_90
timestamp 1604681595
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_97
timestamp 1604681595
transform 1 0 10028 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_102
timestamp 1604681595
transform 1 0 10488 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_101
timestamp 1604681595
transform 1 0 10396 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10212 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1604681595
transform 1 0 11500 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_107
timestamp 1604681595
transform 1 0 10948 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_107
timestamp 1604681595
transform 1 0 10948 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 10764 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 10764 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_3_
timestamp 1604681595
transform 1 0 11132 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1604681595
transform 1 0 11224 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_123
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_117
timestamp 1604681595
transform 1 0 11868 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_122
timestamp 1604681595
transform 1 0 12328 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_118
timestamp 1604681595
transform 1 0 11960 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 12144 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11684 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 12604 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12512 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 13156 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 14444 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12972 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_127
timestamp 1604681595
transform 1 0 12788 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_134
timestamp 1604681595
transform 1 0 13432 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_145
timestamp 1604681595
transform 1 0 14444 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_143
timestamp 1604681595
transform 1 0 14260 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_147
timestamp 1604681595
transform 1 0 14628 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_149
timestamp 1604681595
transform 1 0 14812 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 14628 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 14812 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_26_163
timestamp 1604681595
transform 1 0 16100 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 16376 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 14996 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_27_174
timestamp 1604681595
transform 1 0 17112 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_170
timestamp 1604681595
transform 1 0 16744 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_168
timestamp 1604681595
transform 1 0 16560 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 17296 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 16928 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16836 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_184
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_181
timestamp 1604681595
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_180
timestamp 1604681595
transform 1 0 17664 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_prog_clk_A
timestamp 1604681595
transform 1 0 17848 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 18216 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 17480 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_184
timestamp 1604681595
transform 1 0 18032 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_196
timestamp 1604681595
transform 1 0 19136 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_208
timestamp 1604681595
transform 1 0 20240 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_188
timestamp 1604681595
transform 1 0 18400 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_200
timestamp 1604681595
transform 1 0 19504 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_215
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_227
timestamp 1604681595
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_212
timestamp 1604681595
transform 1 0 20608 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_224
timestamp 1604681595
transform 1 0 21712 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_239
timestamp 1604681595
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_236
timestamp 1604681595
transform 1 0 22816 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_245
timestamp 1604681595
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_251
timestamp 1604681595
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_263
timestamp 1604681595
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_257
timestamp 1604681595
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_269
timestamp 1604681595
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_276
timestamp 1604681595
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 1564 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 1932 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_7
timestamp 1604681595
transform 1 0 1748 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_11
timestamp 1604681595
transform 1 0 2116 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 4416 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 4232 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_23
timestamp 1604681595
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_27
timestamp 1604681595
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_32
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6348 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 6716 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_55
timestamp 1604681595
transform 1 0 6164 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_59
timestamp 1604681595
transform 1 0 6532 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1604681595
transform 1 0 8464 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_1_
timestamp 1604681595
transform 1 0 6900 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 7912 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 8280 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_72
timestamp 1604681595
transform 1 0 7728 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_76
timestamp 1604681595
transform 1 0 8096 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_83
timestamp 1604681595
transform 1 0 8740 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_87
timestamp 1604681595
transform 1 0 9108 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 8924 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_91
timestamp 1604681595
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9292 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_96
timestamp 1604681595
transform 1 0 9936 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 10120 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_100
timestamp 1604681595
transform 1 0 10304 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 10580 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 10764 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_28_124
timestamp 1604681595
transform 1 0 12512 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_0_
timestamp 1604681595
transform 1 0 13248 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 13064 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 14260 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 12696 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_128
timestamp 1604681595
transform 1 0 12880 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1604681595
transform 1 0 14076 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_145
timestamp 1604681595
transform 1 0 14444 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_4_
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 14904 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 16284 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_149
timestamp 1604681595
transform 1 0 14812 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_152
timestamp 1604681595
transform 1 0 15088 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_163
timestamp 1604681595
transform 1 0 16100 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 16836 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 16652 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_167
timestamp 1604681595
transform 1 0 16468 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_180
timestamp 1604681595
transform 1 0 17664 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_192
timestamp 1604681595
transform 1 0 18768 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_204
timestamp 1604681595
transform 1 0 19872 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_212
timestamp 1604681595
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_215
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_227
timestamp 1604681595
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_239
timestamp 1604681595
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_251
timestamp 1604681595
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_263
timestamp 1604681595
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_276
timestamp 1604681595
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 2024 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 1840 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_7
timestamp 1604681595
transform 1 0 1748 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 4140 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 4508 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_29
timestamp 1604681595
transform 1 0 3772 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_35
timestamp 1604681595
transform 1 0 4324 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_39
timestamp 1604681595
transform 1 0 4692 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l4_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 4968 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_53
timestamp 1604681595
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1604681595
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_62
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 7084 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1604681595
transform 1 0 9660 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 10120 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1604681595
transform 1 0 9016 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 9476 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_84
timestamp 1604681595
transform 1 0 8832 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_88
timestamp 1604681595
transform 1 0 9200 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_96
timestamp 1604681595
transform 1 0 9936 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_100
timestamp 1604681595
transform 1 0 10304 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_1_
timestamp 1604681595
transform 1 0 10764 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_114
timestamp 1604681595
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_118
timestamp 1604681595
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 14352 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_142
timestamp 1604681595
transform 1 0 14168 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_1_
timestamp 1604681595
transform 1 0 14904 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 14720 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 15916 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 16284 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_146
timestamp 1604681595
transform 1 0 14536 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_159
timestamp 1604681595
transform 1 0 15732 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_163
timestamp 1604681595
transform 1 0 16100 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1604681595
transform 1 0 16468 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_170
timestamp 1604681595
transform 1 0 16744 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_182
timestamp 1604681595
transform 1 0 17848 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1604681595
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1604681595
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_220
timestamp 1604681595
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_232
timestamp 1604681595
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_245
timestamp 1604681595
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_257
timestamp 1604681595
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_269
timestamp 1604681595
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1604681595
transform 1 0 2944 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 2392 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2760 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_12
timestamp 1604681595
transform 1 0 2208 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_16
timestamp 1604681595
transform 1 0 2576 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4140 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 3404 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_23
timestamp 1604681595
transform 1 0 3220 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_27
timestamp 1604681595
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_32
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 5704 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 5152 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1604681595
transform 1 0 5520 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_42
timestamp 1604681595
transform 1 0 4968 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_46
timestamp 1604681595
transform 1 0 5336 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1604681595
transform 1 0 8188 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7636 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 8004 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8740 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_69
timestamp 1604681595
transform 1 0 7452 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_73
timestamp 1604681595
transform 1 0 7820 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_81
timestamp 1604681595
transform 1 0 8556 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10028 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9844 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 9108 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1604681595
transform 1 0 8924 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_89
timestamp 1604681595
transform 1 0 9292 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_93
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 11592 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11408 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 11040 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 12604 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_106
timestamp 1604681595
transform 1 0 10856 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_110
timestamp 1604681595
transform 1 0 11224 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_123
timestamp 1604681595
transform 1 0 12420 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12972 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 13432 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_127
timestamp 1604681595
transform 1 0 12788 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_131
timestamp 1604681595
transform 1 0 13156 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_145
timestamp 1604681595
transform 1 0 14444 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 14904 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_149
timestamp 1604681595
transform 1 0 14812 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_152
timestamp 1604681595
transform 1 0 15088 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_173
timestamp 1604681595
transform 1 0 17020 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_185
timestamp 1604681595
transform 1 0 18124 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_197
timestamp 1604681595
transform 1 0 19228 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_209
timestamp 1604681595
transform 1 0 20332 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_213
timestamp 1604681595
transform 1 0 20700 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_215
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_227
timestamp 1604681595
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_239
timestamp 1604681595
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_251
timestamp 1604681595
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_263
timestamp 1604681595
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_276
timestamp 1604681595
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 1472 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 2484 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 2852 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_13
timestamp 1604681595
transform 1 0 2300 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_17
timestamp 1604681595
transform 1 0 2668 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 3036 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_31_40
timestamp 1604681595
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_44
timestamp 1604681595
transform 1 0 5152 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 5336 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 4968 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1604681595
transform 1 0 5520 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_60
timestamp 1604681595
transform 1 0 6624 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_56
timestamp 1604681595
transform 1 0 6256 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_52
timestamp 1604681595
transform 1 0 5888 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6440 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6072 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_3_
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8372 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8188 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_71
timestamp 1604681595
transform 1 0 7636 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_75
timestamp 1604681595
transform 1 0 8004 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10580 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9752 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10212 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_88
timestamp 1604681595
transform 1 0 9200 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_92
timestamp 1604681595
transform 1 0 9568 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_96
timestamp 1604681595
transform 1 0 9936 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_101
timestamp 1604681595
transform 1 0 10396 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_114
timestamp 1604681595
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_118
timestamp 1604681595
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_123
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12972 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12788 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 13984 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14444 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_138
timestamp 1604681595
transform 1 0 13800 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_142
timestamp 1604681595
transform 1 0 14168 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 15364 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 15180 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14812 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_147
timestamp 1604681595
transform 1 0 14628 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_151
timestamp 1604681595
transform 1 0 14996 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1604681595
transform 1 0 17296 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_174
timestamp 1604681595
transform 1 0 17112 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_178
timestamp 1604681595
transform 1 0 17480 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_182
timestamp 1604681595
transform 1 0 17848 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1604681595
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1604681595
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_220
timestamp 1604681595
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_232
timestamp 1604681595
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_245
timestamp 1604681595
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_257
timestamp 1604681595
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_269
timestamp 1604681595
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2668 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2116 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 2484 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_9
timestamp 1604681595
transform 1 0 1932 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_13
timestamp 1604681595
transform 1 0 2300 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1604681595
transform 1 0 4324 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_23
timestamp 1604681595
transform 1 0 3220 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_27
timestamp 1604681595
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_32
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5888 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 5704 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 5336 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_44
timestamp 1604681595
transform 1 0 5152 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_48
timestamp 1604681595
transform 1 0 5520 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_61
timestamp 1604681595
transform 1 0 6716 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7452 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 6900 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 7268 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8464 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_65
timestamp 1604681595
transform 1 0 7084 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_78
timestamp 1604681595
transform 1 0 8280 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1604681595
transform 1 0 8648 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9752 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 9016 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 8832 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_89
timestamp 1604681595
transform 1 0 9292 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_93
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_103
timestamp 1604681595
transform 1 0 10580 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 11316 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10764 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11132 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_107
timestamp 1604681595
transform 1 0 10948 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13800 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13248 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_130
timestamp 1604681595
transform 1 0 13064 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_134
timestamp 1604681595
transform 1 0 13432 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_144
timestamp 1604681595
transform 1 0 14352 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16008 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_150
timestamp 1604681595
transform 1 0 14904 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_160
timestamp 1604681595
transform 1 0 15824 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_164
timestamp 1604681595
transform 1 0 16192 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _123_
timestamp 1604681595
transform 1 0 16560 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_172
timestamp 1604681595
transform 1 0 16928 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_184
timestamp 1604681595
transform 1 0 18032 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_196
timestamp 1604681595
transform 1 0 19136 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_208
timestamp 1604681595
transform 1 0 20240 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_215
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_227
timestamp 1604681595
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_239
timestamp 1604681595
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_251
timestamp 1604681595
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_263
timestamp 1604681595
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_276
timestamp 1604681595
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_7
timestamp 1604681595
transform 1 0 1748 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_13
timestamp 1604681595
transform 1 0 2300 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1748 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1932 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_19
timestamp 1604681595
transform 1 0 2852 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_15
timestamp 1604681595
transform 1 0 2484 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_17
timestamp 1604681595
transform 1 0 2668 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 2668 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1604681595
transform 1 0 2852 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2484 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_23
timestamp 1604681595
transform 1 0 3220 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_29
timestamp 1604681595
transform 1 0 3772 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_25
timestamp 1604681595
transform 1 0 3404 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 3036 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3864 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1604681595
transform 1 0 3036 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_36
timestamp 1604681595
transform 1 0 4416 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_32
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_36
timestamp 1604681595
transform 1 0 4416 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_32
timestamp 1604681595
transform 1 0 4048 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 4692 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 4232 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 4232 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4600 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4784 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 4876 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_33_49
timestamp 1604681595
transform 1 0 5612 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 5796 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_60
timestamp 1604681595
transform 1 0 6624 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_60
timestamp 1604681595
transform 1 0 6624 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_53
timestamp 1604681595
transform 1 0 5980 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6808 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1604681595
transform 1 0 6348 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_1_
timestamp 1604681595
transform 1 0 7360 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 8740 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 7176 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8372 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_81
timestamp 1604681595
transform 1 0 8556 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_64
timestamp 1604681595
transform 1 0 6992 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_77
timestamp 1604681595
transform 1 0 8188 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_81
timestamp 1604681595
transform 1 0 8556 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_93
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_91
timestamp 1604681595
transform 1 0 9476 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_87
timestamp 1604681595
transform 1 0 9108 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_85
timestamp 1604681595
transform 1 0 8924 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 8924 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9292 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 9108 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9844 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10028 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9292 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_33_112
timestamp 1604681595
transform 1 0 11408 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_108
timestamp 1604681595
transform 1 0 11040 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11224 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11960 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_118
timestamp 1604681595
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_116
timestamp 1604681595
transform 1 0 11776 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12328 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_123
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_120
timestamp 1604681595
transform 1 0 12144 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12512 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 12604 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1604681595
transform 1 0 14168 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 13524 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 13984 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_144
timestamp 1604681595
transform 1 0 14352 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_133
timestamp 1604681595
transform 1 0 13340 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_137
timestamp 1604681595
transform 1 0 13708 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_145
timestamp 1604681595
transform 1 0 14444 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_148
timestamp 1604681595
transform 1 0 14720 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 14536 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 14904 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604681595
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1604681595
transform 1 0 15088 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_33_165
timestamp 1604681595
transform 1 0 16284 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_161
timestamp 1604681595
transform 1 0 15916 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16100 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_163
timestamp 1604681595
transform 1 0 16100 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1604681595
transform 1 0 16652 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 16468 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_172
timestamp 1604681595
transform 1 0 16928 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_180
timestamp 1604681595
transform 1 0 17664 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1604681595
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_175
timestamp 1604681595
transform 1 0 17204 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_187
timestamp 1604681595
transform 1 0 18308 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_196
timestamp 1604681595
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_208
timestamp 1604681595
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_199
timestamp 1604681595
transform 1 0 19412 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604681595
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_220
timestamp 1604681595
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_211
timestamp 1604681595
transform 1 0 20516 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_215
timestamp 1604681595
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_227
timestamp 1604681595
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_232
timestamp 1604681595
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_245
timestamp 1604681595
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_239
timestamp 1604681595
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_257
timestamp 1604681595
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_269
timestamp 1604681595
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_251
timestamp 1604681595
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_263
timestamp 1604681595
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604681595
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_276
timestamp 1604681595
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1840 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1604681595
transform 1 0 2852 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1656 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_3
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_14
timestamp 1604681595
transform 1 0 2392 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_18
timestamp 1604681595
transform 1 0 2760 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1604681595
transform 1 0 3128 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4140 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 3956 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 3588 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_21
timestamp 1604681595
transform 1 0 3036 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_25
timestamp 1604681595
transform 1 0 3404 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_29
timestamp 1604681595
transform 1 0 3772 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_46
timestamp 1604681595
transform 1 0 5336 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_42
timestamp 1604681595
transform 1 0 4968 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 5152 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 5520 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1604681595
transform 1 0 5704 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_53
timestamp 1604681595
transform 1 0 5980 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 6164 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1604681595
transform 1 0 6348 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604681595
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_62
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 7452 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7268 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_66
timestamp 1604681595
transform 1 0 7176 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9936 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 9752 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_88
timestamp 1604681595
transform 1 0 9200 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_92
timestamp 1604681595
transform 1 0 9568 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_113
timestamp 1604681595
transform 1 0 11500 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_109
timestamp 1604681595
transform 1 0 11132 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_105
timestamp 1604681595
transform 1 0 10764 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11316 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 10948 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_118
timestamp 1604681595
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604681595
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 13984 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 13800 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 13432 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_132
timestamp 1604681595
transform 1 0 13248 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_136
timestamp 1604681595
transform 1 0 13616 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 15916 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 16284 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_159
timestamp 1604681595
transform 1 0 15732 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_163
timestamp 1604681595
transform 1 0 16100 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604681595
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_167
timestamp 1604681595
transform 1 0 16468 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_179
timestamp 1604681595
transform 1 0 17572 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1604681595
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_196
timestamp 1604681595
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_208
timestamp 1604681595
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_220
timestamp 1604681595
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604681595
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_232
timestamp 1604681595
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_245
timestamp 1604681595
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_257
timestamp 1604681595
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_269
timestamp 1604681595
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1604681595
transform 1 0 2852 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1564 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604681595
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2392 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1604681595
transform 1 0 1380 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_11
timestamp 1604681595
transform 1 0 2116 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_16
timestamp 1604681595
transform 1 0 2576 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_27
timestamp 1604681595
transform 1 0 3588 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_23
timestamp 1604681595
transform 1 0 3220 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604681595
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_39
timestamp 1604681595
transform 1 0 4692 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_36
timestamp 1604681595
transform 1 0 4416 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_32
timestamp 1604681595
transform 1 0 4048 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4508 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_39.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 4876 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_36_60
timestamp 1604681595
transform 1 0 6624 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7636 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6992 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 7452 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 8648 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_66
timestamp 1604681595
transform 1 0 7176 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_80
timestamp 1604681595
transform 1 0 8464 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9752 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604681595
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_84
timestamp 1604681595
transform 1 0 8832 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_88
timestamp 1604681595
transform 1 0 9200 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_93
timestamp 1604681595
transform 1 0 9660 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_103
timestamp 1604681595
transform 1 0 10580 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1604681595
transform 1 0 12604 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1604681595
transform 1 0 11316 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 12420 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 10764 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_107
timestamp 1604681595
transform 1 0 10948 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_114
timestamp 1604681595
transform 1 0 11592 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_122
timestamp 1604681595
transform 1 0 12328 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13800 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13248 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13616 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_128
timestamp 1604681595
transform 1 0 12880 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_134
timestamp 1604681595
transform 1 0 13432 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_144
timestamp 1604681595
transform 1 0 14352 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 15364 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604681595
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14996 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_150
timestamp 1604681595
transform 1 0 14904 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_154
timestamp 1604681595
transform 1 0 15272 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_174
timestamp 1604681595
transform 1 0 17112 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_186
timestamp 1604681595
transform 1 0 18216 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_198
timestamp 1604681595
transform 1 0 19320 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604681595
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_210
timestamp 1604681595
transform 1 0 20424 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_215
timestamp 1604681595
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_227
timestamp 1604681595
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_239
timestamp 1604681595
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_251
timestamp 1604681595
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_263
timestamp 1604681595
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604681595
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604681595
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_276
timestamp 1604681595
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2944 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1656 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604681595
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2760 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 2392 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_3
timestamp 1604681595
transform 1 0 1380 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_12
timestamp 1604681595
transform 1 0 2208 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_16
timestamp 1604681595
transform 1 0 2576 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4508 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4324 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 3956 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_29
timestamp 1604681595
transform 1 0 3772 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_33
timestamp 1604681595
transform 1 0 4140 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604681595
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 5520 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_46
timestamp 1604681595
transform 1 0 5336 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_50
timestamp 1604681595
transform 1 0 5704 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_54
timestamp 1604681595
transform 1 0 6072 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1604681595
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_62
timestamp 1604681595
transform 1 0 6808 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 8556 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6992 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 8372 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8004 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_73
timestamp 1604681595
transform 1 0 7820 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_77
timestamp 1604681595
transform 1 0 8188 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 10488 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_100
timestamp 1604681595
transform 1 0 10304 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_104
timestamp 1604681595
transform 1 0 10672 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1604681595
transform 1 0 11040 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604681595
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 10856 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_111
timestamp 1604681595
transform 1 0 11316 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_119
timestamp 1604681595
transform 1 0 12052 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_123
timestamp 1604681595
transform 1 0 12420 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13248 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13064 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12696 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_128
timestamp 1604681595
transform 1 0 12880 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_141
timestamp 1604681595
transform 1 0 14076 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_145
timestamp 1604681595
transform 1 0 14444 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_29.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 15456 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 15272 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 14904 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 14536 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_148
timestamp 1604681595
transform 1 0 14720 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_152
timestamp 1604681595
transform 1 0 15088 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604681595
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 18216 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17388 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_175
timestamp 1604681595
transform 1 0 17204 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_179
timestamp 1604681595
transform 1 0 17572 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_184
timestamp 1604681595
transform 1 0 18032 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1604681595
transform 1 0 19412 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_188
timestamp 1604681595
transform 1 0 18400 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_196
timestamp 1604681595
transform 1 0 19136 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_201
timestamp 1604681595
transform 1 0 19596 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20884 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_213
timestamp 1604681595
transform 1 0 20700 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_217
timestamp 1604681595
transform 1 0 21068 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_229
timestamp 1604681595
transform 1 0 22172 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604681595
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 22448 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_234
timestamp 1604681595
transform 1 0 22632 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_242
timestamp 1604681595
transform 1 0 23368 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_245
timestamp 1604681595
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_257
timestamp 1604681595
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_269
timestamp 1604681595
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604681595
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1604681595
transform 1 0 1380 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604681595
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 2208 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1840 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_6
timestamp 1604681595
transform 1 0 1656 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_10
timestamp 1604681595
transform 1 0 2024 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_39.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 4048 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604681595
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_23
timestamp 1604681595
transform 1 0 3220 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_27
timestamp 1604681595
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 5980 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_51
timestamp 1604681595
transform 1 0 5796 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_55
timestamp 1604681595
transform 1 0 6164 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_35.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 7084 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 6900 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_31.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10212 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604681595
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9936 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9384 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_84
timestamp 1604681595
transform 1 0 8832 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_88
timestamp 1604681595
transform 1 0 9200 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_93
timestamp 1604681595
transform 1 0 9660 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_38_98
timestamp 1604681595
transform 1 0 10120 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12144 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12512 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_118
timestamp 1604681595
transform 1 0 11960 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_122
timestamp 1604681595
transform 1 0 12328 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_31.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12696 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_38_145
timestamp 1604681595
transform 1 0 14444 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604681595
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 16284 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_163
timestamp 1604681595
transform 1 0 16100 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18124 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16836 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_167
timestamp 1604681595
transform 1 0 16468 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_177
timestamp 1604681595
transform 1 0 17388 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1604681595
transform 1 0 19412 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_191
timestamp 1604681595
transform 1 0 18676 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_203
timestamp 1604681595
transform 1 0 19780 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20884 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604681595
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_211
timestamp 1604681595
transform 1 0 20516 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_221
timestamp 1604681595
transform 1 0 21436 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_229
timestamp 1604681595
transform 1 0 22172 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 22448 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_38_238
timestamp 1604681595
transform 1 0 23000 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_250
timestamp 1604681595
transform 1 0 24104 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_262
timestamp 1604681595
transform 1 0 25208 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604681595
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1604681595
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_274
timestamp 1604681595
transform 1 0 26312 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_276
timestamp 1604681595
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_3
timestamp 1604681595
transform 1 0 1380 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_39_3
timestamp 1604681595
transform 1 0 1380 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604681595
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604681595
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1656 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1472 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_12
timestamp 1604681595
transform 1 0 2208 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_14
timestamp 1604681595
transform 1 0 2392 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_10
timestamp 1604681595
transform 1 0 2024 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2576 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2208 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_20
timestamp 1604681595
transform 1 0 2944 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_18
timestamp 1604681595
transform 1 0 2760 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 2944 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_30
timestamp 1604681595
transform 1 0 3864 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_24
timestamp 1604681595
transform 1 0 3312 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 3128 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1604681595
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_40
timestamp 1604681595
transform 1 0 4784 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_36
timestamp 1604681595
transform 1 0 4416 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_41
timestamp 1604681595
transform 1 0 4876 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1604681595
transform 1 0 4600 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1604681595
transform 1 0 4048 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_37.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 3128 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_40_44
timestamp 1604681595
transform 1 0 5152 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_47
timestamp 1604681595
transform 1 0 5428 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 5244 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1604681595
transform 1 0 5612 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_62
timestamp 1604681595
transform 1 0 6808 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1604681595
transform 1 0 6348 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_53
timestamp 1604681595
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1604681595
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1604681595
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_37.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 5244 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_35.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 6992 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7820 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 7176 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_83
timestamp 1604681595
transform 1 0 8740 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_64
timestamp 1604681595
transform 1 0 6992 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_68
timestamp 1604681595
transform 1 0 7360 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_72
timestamp 1604681595
transform 1 0 7728 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_93
timestamp 1604681595
transform 1 0 9660 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_84
timestamp 1604681595
transform 1 0 8832 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_91
timestamp 1604681595
transform 1 0 9476 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_87
timestamp 1604681595
transform 1 0 9108 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9660 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9292 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8924 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1604681595
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9936 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9844 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1604681595
transform 1 0 12420 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1604681595
transform 1 0 11500 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1604681595
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 11776 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_114
timestamp 1604681595
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_118
timestamp 1604681595
transform 1 0 11960 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_105
timestamp 1604681595
transform 1 0 10764 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_40_122
timestamp 1604681595
transform 1 0 12328 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_131
timestamp 1604681595
transform 1 0 13156 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_127
timestamp 1604681595
transform 1 0 12788 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12880 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13340 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1604681595
transform 1 0 12972 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13064 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_40_143
timestamp 1604681595
transform 1 0 14260 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_139
timestamp 1604681595
transform 1 0 13892 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 14076 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_29.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 13524 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_40_151
timestamp 1604681595
transform 1 0 14996 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_154
timestamp 1604681595
transform 1 0 15272 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1604681595
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _125_
timestamp 1604681595
transform 1 0 15272 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_158
timestamp 1604681595
transform 1 0 15640 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_158
timestamp 1604681595
transform 1 0 15640 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 15824 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1604681595
transform 1 0 15456 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16008 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _122_
timestamp 1604681595
transform 1 0 16376 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_170
timestamp 1604681595
transform 1 0 16744 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_39_172
timestamp 1604681595
transform 1 0 16928 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_168
timestamp 1604681595
transform 1 0 16560 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__A
timestamp 1604681595
transform 1 0 16744 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_182
timestamp 1604681595
transform 1 0 17848 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_180
timestamp 1604681595
transform 1 0 17664 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1604681595
transform 1 0 17480 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1604681595
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _121_
timestamp 1604681595
transform 1 0 17480 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _120_
timestamp 1604681595
transform 1 0 18032 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_192
timestamp 1604681595
transform 1 0 18768 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_188
timestamp 1604681595
transform 1 0 18400 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A
timestamp 1604681595
transform 1 0 18952 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A
timestamp 1604681595
transform 1 0 18584 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _119_
timestamp 1604681595
transform 1 0 19136 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1604681595
transform 1 0 18584 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_206
timestamp 1604681595
transform 1 0 20056 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_204
timestamp 1604681595
transform 1 0 19872 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_200
timestamp 1604681595
transform 1 0 19504 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1604681595
transform 1 0 20056 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1604681595
transform 1 0 19688 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1604681595
transform 1 0 20240 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_194
timestamp 1604681595
transform 1 0 18952 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_217
timestamp 1604681595
transform 1 0 21068 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_212
timestamp 1604681595
transform 1 0 20608 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1604681595
transform 1 0 20884 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1604681595
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1604681595
transform 1 0 20884 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_219
timestamp 1604681595
transform 1 0 21252 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_224
timestamp 1604681595
transform 1 0 21712 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1604681595
transform 1 0 21896 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1604681595
transform 1 0 21344 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_228
timestamp 1604681595
transform 1 0 22080 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1604681595
transform 1 0 21988 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_231
timestamp 1604681595
transform 1 0 22356 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_236
timestamp 1604681595
transform 1 0 22816 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1604681595
transform 1 0 22264 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1604681595
transform 1 0 23000 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1604681595
transform 1 0 22448 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1604681595
transform 1 0 23092 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_249
timestamp 1604681595
transform 1 0 24012 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_240
timestamp 1604681595
transform 1 0 23184 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1604681595
transform 1 0 23368 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1604681595
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1604681595
transform 1 0 23644 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_243
timestamp 1604681595
transform 1 0 23460 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1604681595
transform 1 0 24196 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_253
timestamp 1604681595
transform 1 0 24380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_265
timestamp 1604681595
transform 1 0 25484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_255
timestamp 1604681595
transform 1 0 24564 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_267
timestamp 1604681595
transform 1 0 25668 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604681595
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604681595
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1604681595
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_276
timestamp 1604681595
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1604681595
transform 1 0 2760 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1472 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604681595
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A
timestamp 1604681595
transform 1 0 2208 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1604681595
transform 1 0 2576 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_3
timestamp 1604681595
transform 1 0 1380 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_10
timestamp 1604681595
transform 1 0 2024 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_14
timestamp 1604681595
transform 1 0 2392 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1604681595
transform 1 0 3864 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1604681595
transform 1 0 4416 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A
timestamp 1604681595
transform 1 0 3312 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1604681595
transform 1 0 3680 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_22
timestamp 1604681595
transform 1 0 3128 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_26
timestamp 1604681595
transform 1 0 3496 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_34
timestamp 1604681595
transform 1 0 4232 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_38
timestamp 1604681595
transform 1 0 4600 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1604681595
transform 1 0 6808 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1604681595
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4968 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6164 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_53
timestamp 1604681595
transform 1 0 5980 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_57
timestamp 1604681595
transform 1 0 6348 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1604681595
transform 1 0 7912 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1604681595
transform 1 0 7360 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A
timestamp 1604681595
transform 1 0 7728 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A
timestamp 1604681595
transform 1 0 8464 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_66
timestamp 1604681595
transform 1 0 7176 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_70
timestamp 1604681595
transform 1 0 7544 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_78
timestamp 1604681595
transform 1 0 8280 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_82
timestamp 1604681595
transform 1 0 8648 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9568 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 10304 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1604681595
transform 1 0 8832 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1604681595
transform 1 0 9384 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_86
timestamp 1604681595
transform 1 0 9016 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_98
timestamp 1604681595
transform 1 0 10120 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_102
timestamp 1604681595
transform 1 0 10488 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12420 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1604681595
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_114
timestamp 1604681595
transform 1 0 11592 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 13156 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 13524 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_129
timestamp 1604681595
transform 1 0 12972 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_133
timestamp 1604681595
transform 1 0 13340 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_137
timestamp 1604681595
transform 1 0 13708 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1604681595
transform 1 0 16192 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _124_
timestamp 1604681595
transform 1 0 15088 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1604681595
transform 1 0 15640 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1604681595
transform 1 0 14904 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_149
timestamp 1604681595
transform 1 0 14812 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_156
timestamp 1604681595
transform 1 0 15456 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_160
timestamp 1604681595
transform 1 0 15824 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1604681595
transform 1 0 18032 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1604681595
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1604681595
transform 1 0 16744 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_168
timestamp 1604681595
transform 1 0 16560 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_172
timestamp 1604681595
transform 1 0 16928 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_180
timestamp 1604681595
transform 1 0 17664 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A
timestamp 1604681595
transform 1 0 18584 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_188
timestamp 1604681595
transform 1 0 18400 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_192
timestamp 1604681595
transform 1 0 18768 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_204
timestamp 1604681595
transform 1 0 19872 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_216
timestamp 1604681595
transform 1 0 20976 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_228
timestamp 1604681595
transform 1 0 22080 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1604681595
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_240
timestamp 1604681595
transform 1 0 23184 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_245
timestamp 1604681595
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_257
timestamp 1604681595
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_269
timestamp 1604681595
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604681595
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1604681595
transform 1 0 2484 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1604681595
transform 1 0 1380 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604681595
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1932 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_7
timestamp 1604681595
transform 1 0 1748 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_11
timestamp 1604681595
transform 1 0 2116 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_19
timestamp 1604681595
transform 1 0 2852 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1604681595
transform 1 0 4048 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1604681595
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_36
timestamp 1604681595
transform 1 0 4416 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1604681595
transform 1 0 5152 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1604681595
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1604681595
transform 1 0 5704 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_48
timestamp 1604681595
transform 1 0 5520 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_52
timestamp 1604681595
transform 1 0 5888 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_60
timestamp 1604681595
transform 1 0 6624 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1604681595
transform 1 0 8004 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1604681595
transform 1 0 6900 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_67
timestamp 1604681595
transform 1 0 7268 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_79
timestamp 1604681595
transform 1 0 8372 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1604681595
transform 1 0 9752 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1604681595
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_91
timestamp 1604681595
transform 1 0 9476 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_98
timestamp 1604681595
transform 1 0 10120 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1604681595
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_110
timestamp 1604681595
transform 1 0 11224 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_122
timestamp 1604681595
transform 1 0 12328 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_125
timestamp 1604681595
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_137
timestamp 1604681595
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1604681595
transform 1 0 15456 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1604681595
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_149
timestamp 1604681595
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_160
timestamp 1604681595
transform 1 0 15824 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1604681595
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_172
timestamp 1604681595
transform 1 0 16928 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_184
timestamp 1604681595
transform 1 0 18032 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_187
timestamp 1604681595
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_199
timestamp 1604681595
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1604681595
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_211
timestamp 1604681595
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_218
timestamp 1604681595
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1604681595
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_230
timestamp 1604681595
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_242
timestamp 1604681595
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_249
timestamp 1604681595
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_261
timestamp 1604681595
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604681595
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_273
timestamp 1604681595
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 294 0 350 480 6 bottom_left_grid_pin_42_
port 0 nsew default input
rlabel metal2 s 846 0 902 480 6 bottom_left_grid_pin_43_
port 1 nsew default input
rlabel metal2 s 1398 0 1454 480 6 bottom_left_grid_pin_44_
port 2 nsew default input
rlabel metal2 s 1950 0 2006 480 6 bottom_left_grid_pin_45_
port 3 nsew default input
rlabel metal2 s 2502 0 2558 480 6 bottom_left_grid_pin_46_
port 4 nsew default input
rlabel metal2 s 3146 0 3202 480 6 bottom_left_grid_pin_47_
port 5 nsew default input
rlabel metal2 s 3698 0 3754 480 6 bottom_left_grid_pin_48_
port 6 nsew default input
rlabel metal2 s 4250 0 4306 480 6 bottom_left_grid_pin_49_
port 7 nsew default input
rlabel metal2 s 27618 0 27674 480 6 bottom_right_grid_pin_1_
port 8 nsew default input
rlabel metal3 s 27520 13880 28000 14000 6 ccff_head
port 9 nsew default input
rlabel metal3 s 27520 23264 28000 23384 6 ccff_tail
port 10 nsew default tristate
rlabel metal3 s 0 4904 480 5024 6 chanx_left_in[0]
port 11 nsew default input
rlabel metal3 s 0 10752 480 10872 6 chanx_left_in[10]
port 12 nsew default input
rlabel metal3 s 0 11296 480 11416 6 chanx_left_in[11]
port 13 nsew default input
rlabel metal3 s 0 11840 480 11960 6 chanx_left_in[12]
port 14 nsew default input
rlabel metal3 s 0 12520 480 12640 6 chanx_left_in[13]
port 15 nsew default input
rlabel metal3 s 0 13064 480 13184 6 chanx_left_in[14]
port 16 nsew default input
rlabel metal3 s 0 13608 480 13728 6 chanx_left_in[15]
port 17 nsew default input
rlabel metal3 s 0 14288 480 14408 6 chanx_left_in[16]
port 18 nsew default input
rlabel metal3 s 0 14832 480 14952 6 chanx_left_in[17]
port 19 nsew default input
rlabel metal3 s 0 15376 480 15496 6 chanx_left_in[18]
port 20 nsew default input
rlabel metal3 s 0 15920 480 16040 6 chanx_left_in[19]
port 21 nsew default input
rlabel metal3 s 0 5448 480 5568 6 chanx_left_in[1]
port 22 nsew default input
rlabel metal3 s 0 5992 480 6112 6 chanx_left_in[2]
port 23 nsew default input
rlabel metal3 s 0 6672 480 6792 6 chanx_left_in[3]
port 24 nsew default input
rlabel metal3 s 0 7216 480 7336 6 chanx_left_in[4]
port 25 nsew default input
rlabel metal3 s 0 7760 480 7880 6 chanx_left_in[5]
port 26 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_left_in[6]
port 27 nsew default input
rlabel metal3 s 0 8984 480 9104 6 chanx_left_in[7]
port 28 nsew default input
rlabel metal3 s 0 9528 480 9648 6 chanx_left_in[8]
port 29 nsew default input
rlabel metal3 s 0 10072 480 10192 6 chanx_left_in[9]
port 30 nsew default input
rlabel metal3 s 0 16600 480 16720 6 chanx_left_out[0]
port 31 nsew default tristate
rlabel metal3 s 0 22448 480 22568 6 chanx_left_out[10]
port 32 nsew default tristate
rlabel metal3 s 0 22992 480 23112 6 chanx_left_out[11]
port 33 nsew default tristate
rlabel metal3 s 0 23536 480 23656 6 chanx_left_out[12]
port 34 nsew default tristate
rlabel metal3 s 0 24080 480 24200 6 chanx_left_out[13]
port 35 nsew default tristate
rlabel metal3 s 0 24760 480 24880 6 chanx_left_out[14]
port 36 nsew default tristate
rlabel metal3 s 0 25304 480 25424 6 chanx_left_out[15]
port 37 nsew default tristate
rlabel metal3 s 0 25848 480 25968 6 chanx_left_out[16]
port 38 nsew default tristate
rlabel metal3 s 0 26528 480 26648 6 chanx_left_out[17]
port 39 nsew default tristate
rlabel metal3 s 0 27072 480 27192 6 chanx_left_out[18]
port 40 nsew default tristate
rlabel metal3 s 0 27616 480 27736 6 chanx_left_out[19]
port 41 nsew default tristate
rlabel metal3 s 0 17144 480 17264 6 chanx_left_out[1]
port 42 nsew default tristate
rlabel metal3 s 0 17688 480 17808 6 chanx_left_out[2]
port 43 nsew default tristate
rlabel metal3 s 0 18368 480 18488 6 chanx_left_out[3]
port 44 nsew default tristate
rlabel metal3 s 0 18912 480 19032 6 chanx_left_out[4]
port 45 nsew default tristate
rlabel metal3 s 0 19456 480 19576 6 chanx_left_out[5]
port 46 nsew default tristate
rlabel metal3 s 0 20000 480 20120 6 chanx_left_out[6]
port 47 nsew default tristate
rlabel metal3 s 0 20680 480 20800 6 chanx_left_out[7]
port 48 nsew default tristate
rlabel metal3 s 0 21224 480 21344 6 chanx_left_out[8]
port 49 nsew default tristate
rlabel metal3 s 0 21768 480 21888 6 chanx_left_out[9]
port 50 nsew default tristate
rlabel metal2 s 4802 0 4858 480 6 chany_bottom_in[0]
port 51 nsew default input
rlabel metal2 s 10506 0 10562 480 6 chany_bottom_in[10]
port 52 nsew default input
rlabel metal2 s 11058 0 11114 480 6 chany_bottom_in[11]
port 53 nsew default input
rlabel metal2 s 11702 0 11758 480 6 chany_bottom_in[12]
port 54 nsew default input
rlabel metal2 s 12254 0 12310 480 6 chany_bottom_in[13]
port 55 nsew default input
rlabel metal2 s 12806 0 12862 480 6 chany_bottom_in[14]
port 56 nsew default input
rlabel metal2 s 13358 0 13414 480 6 chany_bottom_in[15]
port 57 nsew default input
rlabel metal2 s 13910 0 13966 480 6 chany_bottom_in[16]
port 58 nsew default input
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_in[17]
port 59 nsew default input
rlabel metal2 s 15106 0 15162 480 6 chany_bottom_in[18]
port 60 nsew default input
rlabel metal2 s 15658 0 15714 480 6 chany_bottom_in[19]
port 61 nsew default input
rlabel metal2 s 5354 0 5410 480 6 chany_bottom_in[1]
port 62 nsew default input
rlabel metal2 s 5998 0 6054 480 6 chany_bottom_in[2]
port 63 nsew default input
rlabel metal2 s 6550 0 6606 480 6 chany_bottom_in[3]
port 64 nsew default input
rlabel metal2 s 7102 0 7158 480 6 chany_bottom_in[4]
port 65 nsew default input
rlabel metal2 s 7654 0 7710 480 6 chany_bottom_in[5]
port 66 nsew default input
rlabel metal2 s 8206 0 8262 480 6 chany_bottom_in[6]
port 67 nsew default input
rlabel metal2 s 8850 0 8906 480 6 chany_bottom_in[7]
port 68 nsew default input
rlabel metal2 s 9402 0 9458 480 6 chany_bottom_in[8]
port 69 nsew default input
rlabel metal2 s 9954 0 10010 480 6 chany_bottom_in[9]
port 70 nsew default input
rlabel metal2 s 16210 0 16266 480 6 chany_bottom_out[0]
port 71 nsew default tristate
rlabel metal2 s 21914 0 21970 480 6 chany_bottom_out[10]
port 72 nsew default tristate
rlabel metal2 s 22466 0 22522 480 6 chany_bottom_out[11]
port 73 nsew default tristate
rlabel metal2 s 23110 0 23166 480 6 chany_bottom_out[12]
port 74 nsew default tristate
rlabel metal2 s 23662 0 23718 480 6 chany_bottom_out[13]
port 75 nsew default tristate
rlabel metal2 s 24214 0 24270 480 6 chany_bottom_out[14]
port 76 nsew default tristate
rlabel metal2 s 24766 0 24822 480 6 chany_bottom_out[15]
port 77 nsew default tristate
rlabel metal2 s 25318 0 25374 480 6 chany_bottom_out[16]
port 78 nsew default tristate
rlabel metal2 s 25962 0 26018 480 6 chany_bottom_out[17]
port 79 nsew default tristate
rlabel metal2 s 26514 0 26570 480 6 chany_bottom_out[18]
port 80 nsew default tristate
rlabel metal2 s 27066 0 27122 480 6 chany_bottom_out[19]
port 81 nsew default tristate
rlabel metal2 s 16762 0 16818 480 6 chany_bottom_out[1]
port 82 nsew default tristate
rlabel metal2 s 17406 0 17462 480 6 chany_bottom_out[2]
port 83 nsew default tristate
rlabel metal2 s 17958 0 18014 480 6 chany_bottom_out[3]
port 84 nsew default tristate
rlabel metal2 s 18510 0 18566 480 6 chany_bottom_out[4]
port 85 nsew default tristate
rlabel metal2 s 19062 0 19118 480 6 chany_bottom_out[5]
port 86 nsew default tristate
rlabel metal2 s 19614 0 19670 480 6 chany_bottom_out[6]
port 87 nsew default tristate
rlabel metal2 s 20258 0 20314 480 6 chany_bottom_out[7]
port 88 nsew default tristate
rlabel metal2 s 20810 0 20866 480 6 chany_bottom_out[8]
port 89 nsew default tristate
rlabel metal2 s 21362 0 21418 480 6 chany_bottom_out[9]
port 90 nsew default tristate
rlabel metal2 s 4802 27520 4858 28000 6 chany_top_in[0]
port 91 nsew default input
rlabel metal2 s 10506 27520 10562 28000 6 chany_top_in[10]
port 92 nsew default input
rlabel metal2 s 11058 27520 11114 28000 6 chany_top_in[11]
port 93 nsew default input
rlabel metal2 s 11702 27520 11758 28000 6 chany_top_in[12]
port 94 nsew default input
rlabel metal2 s 12254 27520 12310 28000 6 chany_top_in[13]
port 95 nsew default input
rlabel metal2 s 12806 27520 12862 28000 6 chany_top_in[14]
port 96 nsew default input
rlabel metal2 s 13358 27520 13414 28000 6 chany_top_in[15]
port 97 nsew default input
rlabel metal2 s 13910 27520 13966 28000 6 chany_top_in[16]
port 98 nsew default input
rlabel metal2 s 14554 27520 14610 28000 6 chany_top_in[17]
port 99 nsew default input
rlabel metal2 s 15106 27520 15162 28000 6 chany_top_in[18]
port 100 nsew default input
rlabel metal2 s 15658 27520 15714 28000 6 chany_top_in[19]
port 101 nsew default input
rlabel metal2 s 5354 27520 5410 28000 6 chany_top_in[1]
port 102 nsew default input
rlabel metal2 s 5998 27520 6054 28000 6 chany_top_in[2]
port 103 nsew default input
rlabel metal2 s 6550 27520 6606 28000 6 chany_top_in[3]
port 104 nsew default input
rlabel metal2 s 7102 27520 7158 28000 6 chany_top_in[4]
port 105 nsew default input
rlabel metal2 s 7654 27520 7710 28000 6 chany_top_in[5]
port 106 nsew default input
rlabel metal2 s 8206 27520 8262 28000 6 chany_top_in[6]
port 107 nsew default input
rlabel metal2 s 8850 27520 8906 28000 6 chany_top_in[7]
port 108 nsew default input
rlabel metal2 s 9402 27520 9458 28000 6 chany_top_in[8]
port 109 nsew default input
rlabel metal2 s 9954 27520 10010 28000 6 chany_top_in[9]
port 110 nsew default input
rlabel metal2 s 16210 27520 16266 28000 6 chany_top_out[0]
port 111 nsew default tristate
rlabel metal2 s 21914 27520 21970 28000 6 chany_top_out[10]
port 112 nsew default tristate
rlabel metal2 s 22466 27520 22522 28000 6 chany_top_out[11]
port 113 nsew default tristate
rlabel metal2 s 23110 27520 23166 28000 6 chany_top_out[12]
port 114 nsew default tristate
rlabel metal2 s 23662 27520 23718 28000 6 chany_top_out[13]
port 115 nsew default tristate
rlabel metal2 s 24214 27520 24270 28000 6 chany_top_out[14]
port 116 nsew default tristate
rlabel metal2 s 24766 27520 24822 28000 6 chany_top_out[15]
port 117 nsew default tristate
rlabel metal2 s 25318 27520 25374 28000 6 chany_top_out[16]
port 118 nsew default tristate
rlabel metal2 s 25962 27520 26018 28000 6 chany_top_out[17]
port 119 nsew default tristate
rlabel metal2 s 26514 27520 26570 28000 6 chany_top_out[18]
port 120 nsew default tristate
rlabel metal2 s 27066 27520 27122 28000 6 chany_top_out[19]
port 121 nsew default tristate
rlabel metal2 s 16762 27520 16818 28000 6 chany_top_out[1]
port 122 nsew default tristate
rlabel metal2 s 17406 27520 17462 28000 6 chany_top_out[2]
port 123 nsew default tristate
rlabel metal2 s 17958 27520 18014 28000 6 chany_top_out[3]
port 124 nsew default tristate
rlabel metal2 s 18510 27520 18566 28000 6 chany_top_out[4]
port 125 nsew default tristate
rlabel metal2 s 19062 27520 19118 28000 6 chany_top_out[5]
port 126 nsew default tristate
rlabel metal2 s 19614 27520 19670 28000 6 chany_top_out[6]
port 127 nsew default tristate
rlabel metal2 s 20258 27520 20314 28000 6 chany_top_out[7]
port 128 nsew default tristate
rlabel metal2 s 20810 27520 20866 28000 6 chany_top_out[8]
port 129 nsew default tristate
rlabel metal2 s 21362 27520 21418 28000 6 chany_top_out[9]
port 130 nsew default tristate
rlabel metal3 s 0 280 480 400 6 left_bottom_grid_pin_34_
port 131 nsew default input
rlabel metal3 s 0 824 480 944 6 left_bottom_grid_pin_35_
port 132 nsew default input
rlabel metal3 s 0 1368 480 1488 6 left_bottom_grid_pin_36_
port 133 nsew default input
rlabel metal3 s 0 1912 480 2032 6 left_bottom_grid_pin_37_
port 134 nsew default input
rlabel metal3 s 0 2592 480 2712 6 left_bottom_grid_pin_38_
port 135 nsew default input
rlabel metal3 s 0 3136 480 3256 6 left_bottom_grid_pin_39_
port 136 nsew default input
rlabel metal3 s 0 3680 480 3800 6 left_bottom_grid_pin_40_
port 137 nsew default input
rlabel metal3 s 0 4360 480 4480 6 left_bottom_grid_pin_41_
port 138 nsew default input
rlabel metal3 s 27520 4632 28000 4752 6 prog_clk
port 139 nsew default input
rlabel metal2 s 294 27520 350 28000 6 top_left_grid_pin_42_
port 140 nsew default input
rlabel metal2 s 846 27520 902 28000 6 top_left_grid_pin_43_
port 141 nsew default input
rlabel metal2 s 1398 27520 1454 28000 6 top_left_grid_pin_44_
port 142 nsew default input
rlabel metal2 s 1950 27520 2006 28000 6 top_left_grid_pin_45_
port 143 nsew default input
rlabel metal2 s 2502 27520 2558 28000 6 top_left_grid_pin_46_
port 144 nsew default input
rlabel metal2 s 3146 27520 3202 28000 6 top_left_grid_pin_47_
port 145 nsew default input
rlabel metal2 s 3698 27520 3754 28000 6 top_left_grid_pin_48_
port 146 nsew default input
rlabel metal2 s 4250 27520 4306 28000 6 top_left_grid_pin_49_
port 147 nsew default input
rlabel metal2 s 27618 27520 27674 28000 6 top_right_grid_pin_1_
port 148 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 VPWR
port 149 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 VGND
port 150 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
