magic
tech EFS8A
magscale 1 2
timestamp 1602539203
<< locali >>
rect 4807 231081 4813 231115
rect 4807 231013 4841 231081
rect 4807 226729 4813 226763
rect 4807 226661 4841 226729
rect 4807 225641 4813 225675
rect 4807 225573 4841 225641
rect 3979 214999 4013 215067
rect 3979 214965 3985 214999
<< viali >>
rect 2237 244681 2271 244715
rect 2053 244477 2087 244511
rect 2697 244341 2731 244375
rect 7665 241961 7699 241995
rect 7481 241825 7515 241859
rect 7481 241077 7515 241111
rect 7021 239241 7055 239275
rect 6837 239037 6871 239071
rect 7389 239037 7423 239071
rect 2513 237473 2547 237507
rect 2697 237405 2731 237439
rect 3157 237269 3191 237303
rect 2513 237065 2547 237099
rect 2973 236725 3007 236759
rect 4398 234277 4432 234311
rect 6745 234209 6779 234243
rect 4077 234141 4111 234175
rect 6929 234141 6963 234175
rect 4997 234005 5031 234039
rect 7389 234005 7423 234039
rect 7021 233801 7055 233835
rect 5089 233733 5123 233767
rect 4629 233665 4663 233699
rect 4445 233597 4479 233631
rect 3801 233461 3835 233495
rect 4169 233461 4203 233495
rect 7389 233461 7423 233495
rect 4537 233257 4571 233291
rect 4905 233257 4939 233291
rect 3801 232713 3835 232747
rect 2881 232509 2915 232543
rect 2789 232441 2823 232475
rect 3243 232441 3277 232475
rect 2973 231829 3007 231863
rect 4813 231081 4847 231115
rect 5365 231081 5399 231115
rect 4445 230877 4479 230911
rect 2973 230741 3007 230775
rect 2789 230469 2823 230503
rect 3157 230333 3191 230367
rect 3341 230333 3375 230367
rect 3709 230333 3743 230367
rect 4077 230333 4111 230367
rect 2421 230197 2455 230231
rect 4077 230197 4111 230231
rect 4721 230197 4755 230231
rect 4997 230197 5031 230231
rect 2973 229993 3007 230027
rect 4445 229925 4479 229959
rect 4077 229857 4111 229891
rect 4261 229857 4295 229891
rect 4353 229857 4387 229891
rect 4813 229789 4847 229823
rect 3249 229653 3283 229687
rect 2789 229449 2823 229483
rect 5365 229449 5399 229483
rect 5089 229381 5123 229415
rect 2053 229313 2087 229347
rect 4353 229313 4387 229347
rect 2881 229245 2915 229279
rect 3341 229245 3375 229279
rect 3709 229245 3743 229279
rect 4077 229245 4111 229279
rect 5733 229245 5767 229279
rect 2421 229109 2455 229143
rect 4721 229109 4755 229143
rect 2605 228905 2639 228939
rect 3433 228905 3467 228939
rect 2789 228837 2823 228871
rect 2697 228769 2731 228803
rect 4077 228769 4111 228803
rect 4721 228769 4755 228803
rect 2421 228701 2455 228735
rect 3157 228701 3191 228735
rect 2329 228565 2363 228599
rect 2053 228361 2087 228395
rect 2421 228293 2455 228327
rect 2881 228293 2915 228327
rect 3709 228225 3743 228259
rect 3325 228157 3359 228191
rect 2973 228089 3007 228123
rect 1777 228021 1811 228055
rect 3157 228021 3191 228055
rect 3249 228021 3283 228055
rect 4169 228021 4203 228055
rect 3065 227817 3099 227851
rect 2881 227681 2915 227715
rect 2513 227477 2547 227511
rect 3341 227477 3375 227511
rect 3709 227477 3743 227511
rect 2053 227273 2087 227307
rect 2329 227273 2363 227307
rect 2789 227069 2823 227103
rect 3157 227069 3191 227103
rect 3341 227069 3375 227103
rect 3709 227069 3743 227103
rect 4077 227069 4111 227103
rect 4077 226933 4111 226967
rect 3433 226729 3467 226763
rect 4813 226729 4847 226763
rect 2421 226661 2455 226695
rect 2513 226593 2547 226627
rect 4445 226593 4479 226627
rect 5365 226389 5399 226423
rect 2421 226185 2455 226219
rect 3525 226185 3559 226219
rect 5641 226185 5675 226219
rect 4445 226049 4479 226083
rect 3985 225981 4019 226015
rect 4353 225913 4387 225947
rect 4766 225913 4800 225947
rect 5365 225845 5399 225879
rect 4813 225641 4847 225675
rect 4445 225505 4479 225539
rect 6285 225505 6319 225539
rect 6469 225437 6503 225471
rect 5365 225301 5399 225335
rect 6653 225301 6687 225335
rect 4813 225097 4847 225131
rect 5917 225097 5951 225131
rect 6285 225097 6319 225131
rect 4537 225029 4571 225063
rect 6837 224961 6871 224995
rect 7021 224893 7055 224927
rect 7481 224757 7515 224791
rect 2605 224553 2639 224587
rect 6929 224553 6963 224587
rect 7205 224553 7239 224587
rect 5825 224417 5859 224451
rect 6009 224349 6043 224383
rect 6469 224213 6503 224247
rect 2421 224009 2455 224043
rect 5825 224009 5859 224043
rect 6285 224009 6319 224043
rect 2605 223805 2639 223839
rect 3249 223805 3283 223839
rect 3433 223805 3467 223839
rect 3801 223805 3835 223839
rect 2145 223737 2179 223771
rect 2881 223669 2915 223703
rect 2697 223465 2731 223499
rect 3065 222377 3099 222411
rect 2513 221833 2547 221867
rect 2881 221833 2915 221867
rect 2973 221697 3007 221731
rect 4537 221697 4571 221731
rect 3249 221629 3283 221663
rect 4445 221629 4479 221663
rect 4629 221629 4663 221663
rect 3157 221561 3191 221595
rect 3341 221561 3375 221595
rect 3709 221561 3743 221595
rect 2973 220949 3007 220983
rect 3617 215169 3651 215203
rect 3525 214965 3559 214999
rect 3985 214965 4019 214999
rect 4537 214965 4571 214999
rect 3709 214761 3743 214795
rect 7665 214217 7699 214251
rect 7481 214013 7515 214047
rect 8033 214013 8067 214047
rect 4261 212041 4295 212075
rect 4445 211905 4479 211939
rect 4629 211905 4663 211939
rect 5089 211701 5123 211735
rect 4537 211497 4571 211531
rect 7021 210953 7055 210987
rect 6837 210749 6871 210783
rect 7389 210749 7423 210783
rect 3341 209865 3375 209899
rect 2697 209661 2731 209695
rect 2881 209661 2915 209695
rect 2513 209525 2547 209559
rect 2789 208981 2823 209015
rect 3709 208777 3743 208811
rect 2789 208641 2823 208675
rect 2697 208505 2731 208539
rect 3151 208505 3185 208539
rect 2881 208233 2915 208267
rect 7665 172329 7699 172363
rect 7481 172193 7515 172227
rect 7481 171785 7515 171819
rect 4261 158185 4295 158219
rect 4065 158049 4099 158083
rect 4077 157641 4111 157675
rect 7021 50949 7055 50983
rect 6837 50813 6871 50847
rect 7389 50813 7423 50847
<< metal1 >>
rect 566 332528 572 332580
rect 624 332568 630 332580
rect 1210 332568 1216 332580
rect 624 332540 1216 332568
rect 624 332528 630 332540
rect 1210 332528 1216 332540
rect 1268 332528 1274 332580
rect 3050 332528 3056 332580
rect 3108 332568 3114 332580
rect 3878 332568 3884 332580
rect 3108 332540 3884 332568
rect 3108 332528 3114 332540
rect 3878 332528 3884 332540
rect 3936 332528 3942 332580
rect 4246 332528 4252 332580
rect 4304 332568 4310 332580
rect 5442 332568 5448 332580
rect 4304 332540 5448 332568
rect 4304 332528 4310 332540
rect 5442 332528 5448 332540
rect 5500 332528 5506 332580
rect 8294 332528 8300 332580
rect 8352 332568 8358 332580
rect 9306 332568 9312 332580
rect 8352 332540 9312 332568
rect 8352 332528 8358 332540
rect 9306 332528 9312 332540
rect 9364 332528 9370 332580
rect 1104 330778 8832 330800
rect 1104 330726 2648 330778
rect 2700 330726 2712 330778
rect 2764 330726 2776 330778
rect 2828 330726 2840 330778
rect 2892 330726 5982 330778
rect 6034 330726 6046 330778
rect 6098 330726 6110 330778
rect 6162 330726 6174 330778
rect 6226 330726 8832 330778
rect 1104 330704 8832 330726
rect 1104 330234 8832 330256
rect 1104 330182 4315 330234
rect 4367 330182 4379 330234
rect 4431 330182 4443 330234
rect 4495 330182 4507 330234
rect 4559 330182 7648 330234
rect 7700 330182 7712 330234
rect 7764 330182 7776 330234
rect 7828 330182 7840 330234
rect 7892 330182 8832 330234
rect 1104 330160 8832 330182
rect 1104 329690 8832 329712
rect 1104 329638 2648 329690
rect 2700 329638 2712 329690
rect 2764 329638 2776 329690
rect 2828 329638 2840 329690
rect 2892 329638 5982 329690
rect 6034 329638 6046 329690
rect 6098 329638 6110 329690
rect 6162 329638 6174 329690
rect 6226 329638 8832 329690
rect 1104 329616 8832 329638
rect 1104 329146 8832 329168
rect 1104 329094 4315 329146
rect 4367 329094 4379 329146
rect 4431 329094 4443 329146
rect 4495 329094 4507 329146
rect 4559 329094 7648 329146
rect 7700 329094 7712 329146
rect 7764 329094 7776 329146
rect 7828 329094 7840 329146
rect 7892 329094 8832 329146
rect 1104 329072 8832 329094
rect 1104 328602 8832 328624
rect 1104 328550 2648 328602
rect 2700 328550 2712 328602
rect 2764 328550 2776 328602
rect 2828 328550 2840 328602
rect 2892 328550 5982 328602
rect 6034 328550 6046 328602
rect 6098 328550 6110 328602
rect 6162 328550 6174 328602
rect 6226 328550 8832 328602
rect 1104 328528 8832 328550
rect 1104 328058 8832 328080
rect 1104 328006 4315 328058
rect 4367 328006 4379 328058
rect 4431 328006 4443 328058
rect 4495 328006 4507 328058
rect 4559 328006 7648 328058
rect 7700 328006 7712 328058
rect 7764 328006 7776 328058
rect 7828 328006 7840 328058
rect 7892 328006 8832 328058
rect 1104 327984 8832 328006
rect 1104 327514 8832 327536
rect 1104 327462 2648 327514
rect 2700 327462 2712 327514
rect 2764 327462 2776 327514
rect 2828 327462 2840 327514
rect 2892 327462 5982 327514
rect 6034 327462 6046 327514
rect 6098 327462 6110 327514
rect 6162 327462 6174 327514
rect 6226 327462 8832 327514
rect 1104 327440 8832 327462
rect 1104 326970 8832 326992
rect 1104 326918 4315 326970
rect 4367 326918 4379 326970
rect 4431 326918 4443 326970
rect 4495 326918 4507 326970
rect 4559 326918 7648 326970
rect 7700 326918 7712 326970
rect 7764 326918 7776 326970
rect 7828 326918 7840 326970
rect 7892 326918 8832 326970
rect 1104 326896 8832 326918
rect 1104 326426 8832 326448
rect 1104 326374 2648 326426
rect 2700 326374 2712 326426
rect 2764 326374 2776 326426
rect 2828 326374 2840 326426
rect 2892 326374 5982 326426
rect 6034 326374 6046 326426
rect 6098 326374 6110 326426
rect 6162 326374 6174 326426
rect 6226 326374 8832 326426
rect 1104 326352 8832 326374
rect 1104 325882 8832 325904
rect 1104 325830 4315 325882
rect 4367 325830 4379 325882
rect 4431 325830 4443 325882
rect 4495 325830 4507 325882
rect 4559 325830 7648 325882
rect 7700 325830 7712 325882
rect 7764 325830 7776 325882
rect 7828 325830 7840 325882
rect 7892 325830 8832 325882
rect 1104 325808 8832 325830
rect 1104 325338 8832 325360
rect 1104 325286 2648 325338
rect 2700 325286 2712 325338
rect 2764 325286 2776 325338
rect 2828 325286 2840 325338
rect 2892 325286 5982 325338
rect 6034 325286 6046 325338
rect 6098 325286 6110 325338
rect 6162 325286 6174 325338
rect 6226 325286 8832 325338
rect 1104 325264 8832 325286
rect 1104 324794 8832 324816
rect 1104 324742 4315 324794
rect 4367 324742 4379 324794
rect 4431 324742 4443 324794
rect 4495 324742 4507 324794
rect 4559 324742 7648 324794
rect 7700 324742 7712 324794
rect 7764 324742 7776 324794
rect 7828 324742 7840 324794
rect 7892 324742 8832 324794
rect 1104 324720 8832 324742
rect 1104 324250 8832 324272
rect 1104 324198 2648 324250
rect 2700 324198 2712 324250
rect 2764 324198 2776 324250
rect 2828 324198 2840 324250
rect 2892 324198 5982 324250
rect 6034 324198 6046 324250
rect 6098 324198 6110 324250
rect 6162 324198 6174 324250
rect 6226 324198 8832 324250
rect 1104 324176 8832 324198
rect 1104 323706 8832 323728
rect 1104 323654 4315 323706
rect 4367 323654 4379 323706
rect 4431 323654 4443 323706
rect 4495 323654 4507 323706
rect 4559 323654 7648 323706
rect 7700 323654 7712 323706
rect 7764 323654 7776 323706
rect 7828 323654 7840 323706
rect 7892 323654 8832 323706
rect 1104 323632 8832 323654
rect 1104 323162 8832 323184
rect 1104 323110 2648 323162
rect 2700 323110 2712 323162
rect 2764 323110 2776 323162
rect 2828 323110 2840 323162
rect 2892 323110 5982 323162
rect 6034 323110 6046 323162
rect 6098 323110 6110 323162
rect 6162 323110 6174 323162
rect 6226 323110 8832 323162
rect 1104 323088 8832 323110
rect 1104 322618 8832 322640
rect 1104 322566 4315 322618
rect 4367 322566 4379 322618
rect 4431 322566 4443 322618
rect 4495 322566 4507 322618
rect 4559 322566 7648 322618
rect 7700 322566 7712 322618
rect 7764 322566 7776 322618
rect 7828 322566 7840 322618
rect 7892 322566 8832 322618
rect 1104 322544 8832 322566
rect 1104 322074 8832 322096
rect 1104 322022 2648 322074
rect 2700 322022 2712 322074
rect 2764 322022 2776 322074
rect 2828 322022 2840 322074
rect 2892 322022 5982 322074
rect 6034 322022 6046 322074
rect 6098 322022 6110 322074
rect 6162 322022 6174 322074
rect 6226 322022 8832 322074
rect 1104 322000 8832 322022
rect 1104 321530 8832 321552
rect 1104 321478 4315 321530
rect 4367 321478 4379 321530
rect 4431 321478 4443 321530
rect 4495 321478 4507 321530
rect 4559 321478 7648 321530
rect 7700 321478 7712 321530
rect 7764 321478 7776 321530
rect 7828 321478 7840 321530
rect 7892 321478 8832 321530
rect 1104 321456 8832 321478
rect 1104 320986 8832 321008
rect 1104 320934 2648 320986
rect 2700 320934 2712 320986
rect 2764 320934 2776 320986
rect 2828 320934 2840 320986
rect 2892 320934 5982 320986
rect 6034 320934 6046 320986
rect 6098 320934 6110 320986
rect 6162 320934 6174 320986
rect 6226 320934 8832 320986
rect 1104 320912 8832 320934
rect 1104 320442 8832 320464
rect 1104 320390 4315 320442
rect 4367 320390 4379 320442
rect 4431 320390 4443 320442
rect 4495 320390 4507 320442
rect 4559 320390 7648 320442
rect 7700 320390 7712 320442
rect 7764 320390 7776 320442
rect 7828 320390 7840 320442
rect 7892 320390 8832 320442
rect 1104 320368 8832 320390
rect 1104 319898 8832 319920
rect 1104 319846 2648 319898
rect 2700 319846 2712 319898
rect 2764 319846 2776 319898
rect 2828 319846 2840 319898
rect 2892 319846 5982 319898
rect 6034 319846 6046 319898
rect 6098 319846 6110 319898
rect 6162 319846 6174 319898
rect 6226 319846 8832 319898
rect 1104 319824 8832 319846
rect 1104 319354 8832 319376
rect 1104 319302 4315 319354
rect 4367 319302 4379 319354
rect 4431 319302 4443 319354
rect 4495 319302 4507 319354
rect 4559 319302 7648 319354
rect 7700 319302 7712 319354
rect 7764 319302 7776 319354
rect 7828 319302 7840 319354
rect 7892 319302 8832 319354
rect 1104 319280 8832 319302
rect 1104 318810 8832 318832
rect 1104 318758 2648 318810
rect 2700 318758 2712 318810
rect 2764 318758 2776 318810
rect 2828 318758 2840 318810
rect 2892 318758 5982 318810
rect 6034 318758 6046 318810
rect 6098 318758 6110 318810
rect 6162 318758 6174 318810
rect 6226 318758 8832 318810
rect 1104 318736 8832 318758
rect 1104 318266 8832 318288
rect 1104 318214 4315 318266
rect 4367 318214 4379 318266
rect 4431 318214 4443 318266
rect 4495 318214 4507 318266
rect 4559 318214 7648 318266
rect 7700 318214 7712 318266
rect 7764 318214 7776 318266
rect 7828 318214 7840 318266
rect 7892 318214 8832 318266
rect 1104 318192 8832 318214
rect 1104 317722 8832 317744
rect 1104 317670 2648 317722
rect 2700 317670 2712 317722
rect 2764 317670 2776 317722
rect 2828 317670 2840 317722
rect 2892 317670 5982 317722
rect 6034 317670 6046 317722
rect 6098 317670 6110 317722
rect 6162 317670 6174 317722
rect 6226 317670 8832 317722
rect 1104 317648 8832 317670
rect 1104 317178 8832 317200
rect 1104 317126 4315 317178
rect 4367 317126 4379 317178
rect 4431 317126 4443 317178
rect 4495 317126 4507 317178
rect 4559 317126 7648 317178
rect 7700 317126 7712 317178
rect 7764 317126 7776 317178
rect 7828 317126 7840 317178
rect 7892 317126 8832 317178
rect 1104 317104 8832 317126
rect 1104 316634 8832 316656
rect 1104 316582 2648 316634
rect 2700 316582 2712 316634
rect 2764 316582 2776 316634
rect 2828 316582 2840 316634
rect 2892 316582 5982 316634
rect 6034 316582 6046 316634
rect 6098 316582 6110 316634
rect 6162 316582 6174 316634
rect 6226 316582 8832 316634
rect 1104 316560 8832 316582
rect 1104 316090 8832 316112
rect 1104 316038 4315 316090
rect 4367 316038 4379 316090
rect 4431 316038 4443 316090
rect 4495 316038 4507 316090
rect 4559 316038 7648 316090
rect 7700 316038 7712 316090
rect 7764 316038 7776 316090
rect 7828 316038 7840 316090
rect 7892 316038 8832 316090
rect 1104 316016 8832 316038
rect 1104 315546 8832 315568
rect 1104 315494 2648 315546
rect 2700 315494 2712 315546
rect 2764 315494 2776 315546
rect 2828 315494 2840 315546
rect 2892 315494 5982 315546
rect 6034 315494 6046 315546
rect 6098 315494 6110 315546
rect 6162 315494 6174 315546
rect 6226 315494 8832 315546
rect 1104 315472 8832 315494
rect 7374 315120 7380 315172
rect 7432 315160 7438 315172
rect 8018 315160 8024 315172
rect 7432 315132 8024 315160
rect 7432 315120 7438 315132
rect 8018 315120 8024 315132
rect 8076 315120 8082 315172
rect 1104 315002 8832 315024
rect 1104 314950 4315 315002
rect 4367 314950 4379 315002
rect 4431 314950 4443 315002
rect 4495 314950 4507 315002
rect 4559 314950 7648 315002
rect 7700 314950 7712 315002
rect 7764 314950 7776 315002
rect 7828 314950 7840 315002
rect 7892 314950 8832 315002
rect 1104 314928 8832 314950
rect 1104 314458 8832 314480
rect 1104 314406 2648 314458
rect 2700 314406 2712 314458
rect 2764 314406 2776 314458
rect 2828 314406 2840 314458
rect 2892 314406 5982 314458
rect 6034 314406 6046 314458
rect 6098 314406 6110 314458
rect 6162 314406 6174 314458
rect 6226 314406 8832 314458
rect 1104 314384 8832 314406
rect 1104 313914 8832 313936
rect 1104 313862 4315 313914
rect 4367 313862 4379 313914
rect 4431 313862 4443 313914
rect 4495 313862 4507 313914
rect 4559 313862 7648 313914
rect 7700 313862 7712 313914
rect 7764 313862 7776 313914
rect 7828 313862 7840 313914
rect 7892 313862 8832 313914
rect 1104 313840 8832 313862
rect 1104 313370 8832 313392
rect 1104 313318 2648 313370
rect 2700 313318 2712 313370
rect 2764 313318 2776 313370
rect 2828 313318 2840 313370
rect 2892 313318 5982 313370
rect 6034 313318 6046 313370
rect 6098 313318 6110 313370
rect 6162 313318 6174 313370
rect 6226 313318 8832 313370
rect 1104 313296 8832 313318
rect 1104 312826 8832 312848
rect 1104 312774 4315 312826
rect 4367 312774 4379 312826
rect 4431 312774 4443 312826
rect 4495 312774 4507 312826
rect 4559 312774 7648 312826
rect 7700 312774 7712 312826
rect 7764 312774 7776 312826
rect 7828 312774 7840 312826
rect 7892 312774 8832 312826
rect 1104 312752 8832 312774
rect 1104 312282 8832 312304
rect 1104 312230 2648 312282
rect 2700 312230 2712 312282
rect 2764 312230 2776 312282
rect 2828 312230 2840 312282
rect 2892 312230 5982 312282
rect 6034 312230 6046 312282
rect 6098 312230 6110 312282
rect 6162 312230 6174 312282
rect 6226 312230 8832 312282
rect 1104 312208 8832 312230
rect 1104 311738 8832 311760
rect 1104 311686 4315 311738
rect 4367 311686 4379 311738
rect 4431 311686 4443 311738
rect 4495 311686 4507 311738
rect 4559 311686 7648 311738
rect 7700 311686 7712 311738
rect 7764 311686 7776 311738
rect 7828 311686 7840 311738
rect 7892 311686 8832 311738
rect 1104 311664 8832 311686
rect 1104 311194 8832 311216
rect 1104 311142 2648 311194
rect 2700 311142 2712 311194
rect 2764 311142 2776 311194
rect 2828 311142 2840 311194
rect 2892 311142 5982 311194
rect 6034 311142 6046 311194
rect 6098 311142 6110 311194
rect 6162 311142 6174 311194
rect 6226 311142 8832 311194
rect 1104 311120 8832 311142
rect 1104 310650 8832 310672
rect 1104 310598 4315 310650
rect 4367 310598 4379 310650
rect 4431 310598 4443 310650
rect 4495 310598 4507 310650
rect 4559 310598 7648 310650
rect 7700 310598 7712 310650
rect 7764 310598 7776 310650
rect 7828 310598 7840 310650
rect 7892 310598 8832 310650
rect 1104 310576 8832 310598
rect 1104 310106 8832 310128
rect 1104 310054 2648 310106
rect 2700 310054 2712 310106
rect 2764 310054 2776 310106
rect 2828 310054 2840 310106
rect 2892 310054 5982 310106
rect 6034 310054 6046 310106
rect 6098 310054 6110 310106
rect 6162 310054 6174 310106
rect 6226 310054 8832 310106
rect 1104 310032 8832 310054
rect 1104 309562 8832 309584
rect 1104 309510 4315 309562
rect 4367 309510 4379 309562
rect 4431 309510 4443 309562
rect 4495 309510 4507 309562
rect 4559 309510 7648 309562
rect 7700 309510 7712 309562
rect 7764 309510 7776 309562
rect 7828 309510 7840 309562
rect 7892 309510 8832 309562
rect 1104 309488 8832 309510
rect 1104 309018 8832 309040
rect 1104 308966 2648 309018
rect 2700 308966 2712 309018
rect 2764 308966 2776 309018
rect 2828 308966 2840 309018
rect 2892 308966 5982 309018
rect 6034 308966 6046 309018
rect 6098 308966 6110 309018
rect 6162 308966 6174 309018
rect 6226 308966 8832 309018
rect 1104 308944 8832 308966
rect 1104 308474 8832 308496
rect 1104 308422 4315 308474
rect 4367 308422 4379 308474
rect 4431 308422 4443 308474
rect 4495 308422 4507 308474
rect 4559 308422 7648 308474
rect 7700 308422 7712 308474
rect 7764 308422 7776 308474
rect 7828 308422 7840 308474
rect 7892 308422 8832 308474
rect 1104 308400 8832 308422
rect 1104 307930 8832 307952
rect 1104 307878 2648 307930
rect 2700 307878 2712 307930
rect 2764 307878 2776 307930
rect 2828 307878 2840 307930
rect 2892 307878 5982 307930
rect 6034 307878 6046 307930
rect 6098 307878 6110 307930
rect 6162 307878 6174 307930
rect 6226 307878 8832 307930
rect 1104 307856 8832 307878
rect 1104 307386 8832 307408
rect 1104 307334 4315 307386
rect 4367 307334 4379 307386
rect 4431 307334 4443 307386
rect 4495 307334 4507 307386
rect 4559 307334 7648 307386
rect 7700 307334 7712 307386
rect 7764 307334 7776 307386
rect 7828 307334 7840 307386
rect 7892 307334 8832 307386
rect 1104 307312 8832 307334
rect 1104 306842 8832 306864
rect 1104 306790 2648 306842
rect 2700 306790 2712 306842
rect 2764 306790 2776 306842
rect 2828 306790 2840 306842
rect 2892 306790 5982 306842
rect 6034 306790 6046 306842
rect 6098 306790 6110 306842
rect 6162 306790 6174 306842
rect 6226 306790 8832 306842
rect 1104 306768 8832 306790
rect 1104 306298 8832 306320
rect 1104 306246 4315 306298
rect 4367 306246 4379 306298
rect 4431 306246 4443 306298
rect 4495 306246 4507 306298
rect 4559 306246 7648 306298
rect 7700 306246 7712 306298
rect 7764 306246 7776 306298
rect 7828 306246 7840 306298
rect 7892 306246 8832 306298
rect 1104 306224 8832 306246
rect 1104 305754 8832 305776
rect 1104 305702 2648 305754
rect 2700 305702 2712 305754
rect 2764 305702 2776 305754
rect 2828 305702 2840 305754
rect 2892 305702 5982 305754
rect 6034 305702 6046 305754
rect 6098 305702 6110 305754
rect 6162 305702 6174 305754
rect 6226 305702 8832 305754
rect 1104 305680 8832 305702
rect 1104 305210 8832 305232
rect 1104 305158 4315 305210
rect 4367 305158 4379 305210
rect 4431 305158 4443 305210
rect 4495 305158 4507 305210
rect 4559 305158 7648 305210
rect 7700 305158 7712 305210
rect 7764 305158 7776 305210
rect 7828 305158 7840 305210
rect 7892 305158 8832 305210
rect 1104 305136 8832 305158
rect 1104 304666 8832 304688
rect 1104 304614 2648 304666
rect 2700 304614 2712 304666
rect 2764 304614 2776 304666
rect 2828 304614 2840 304666
rect 2892 304614 5982 304666
rect 6034 304614 6046 304666
rect 6098 304614 6110 304666
rect 6162 304614 6174 304666
rect 6226 304614 8832 304666
rect 1104 304592 8832 304614
rect 1104 304122 8832 304144
rect 1104 304070 4315 304122
rect 4367 304070 4379 304122
rect 4431 304070 4443 304122
rect 4495 304070 4507 304122
rect 4559 304070 7648 304122
rect 7700 304070 7712 304122
rect 7764 304070 7776 304122
rect 7828 304070 7840 304122
rect 7892 304070 8832 304122
rect 1104 304048 8832 304070
rect 1104 303578 8832 303600
rect 1104 303526 2648 303578
rect 2700 303526 2712 303578
rect 2764 303526 2776 303578
rect 2828 303526 2840 303578
rect 2892 303526 5982 303578
rect 6034 303526 6046 303578
rect 6098 303526 6110 303578
rect 6162 303526 6174 303578
rect 6226 303526 8832 303578
rect 1104 303504 8832 303526
rect 1104 303034 8832 303056
rect 1104 302982 4315 303034
rect 4367 302982 4379 303034
rect 4431 302982 4443 303034
rect 4495 302982 4507 303034
rect 4559 302982 7648 303034
rect 7700 302982 7712 303034
rect 7764 302982 7776 303034
rect 7828 302982 7840 303034
rect 7892 302982 8832 303034
rect 1104 302960 8832 302982
rect 1104 302490 8832 302512
rect 1104 302438 2648 302490
rect 2700 302438 2712 302490
rect 2764 302438 2776 302490
rect 2828 302438 2840 302490
rect 2892 302438 5982 302490
rect 6034 302438 6046 302490
rect 6098 302438 6110 302490
rect 6162 302438 6174 302490
rect 6226 302438 8832 302490
rect 1104 302416 8832 302438
rect 1104 301946 8832 301968
rect 1104 301894 4315 301946
rect 4367 301894 4379 301946
rect 4431 301894 4443 301946
rect 4495 301894 4507 301946
rect 4559 301894 7648 301946
rect 7700 301894 7712 301946
rect 7764 301894 7776 301946
rect 7828 301894 7840 301946
rect 7892 301894 8832 301946
rect 1104 301872 8832 301894
rect 1104 301402 8832 301424
rect 1104 301350 2648 301402
rect 2700 301350 2712 301402
rect 2764 301350 2776 301402
rect 2828 301350 2840 301402
rect 2892 301350 5982 301402
rect 6034 301350 6046 301402
rect 6098 301350 6110 301402
rect 6162 301350 6174 301402
rect 6226 301350 8832 301402
rect 1104 301328 8832 301350
rect 1104 300858 8832 300880
rect 1104 300806 4315 300858
rect 4367 300806 4379 300858
rect 4431 300806 4443 300858
rect 4495 300806 4507 300858
rect 4559 300806 7648 300858
rect 7700 300806 7712 300858
rect 7764 300806 7776 300858
rect 7828 300806 7840 300858
rect 7892 300806 8832 300858
rect 1104 300784 8832 300806
rect 1104 300314 8832 300336
rect 1104 300262 2648 300314
rect 2700 300262 2712 300314
rect 2764 300262 2776 300314
rect 2828 300262 2840 300314
rect 2892 300262 5982 300314
rect 6034 300262 6046 300314
rect 6098 300262 6110 300314
rect 6162 300262 6174 300314
rect 6226 300262 8832 300314
rect 1104 300240 8832 300262
rect 1104 299770 8832 299792
rect 1104 299718 4315 299770
rect 4367 299718 4379 299770
rect 4431 299718 4443 299770
rect 4495 299718 4507 299770
rect 4559 299718 7648 299770
rect 7700 299718 7712 299770
rect 7764 299718 7776 299770
rect 7828 299718 7840 299770
rect 7892 299718 8832 299770
rect 1104 299696 8832 299718
rect 1104 299226 8832 299248
rect 1104 299174 2648 299226
rect 2700 299174 2712 299226
rect 2764 299174 2776 299226
rect 2828 299174 2840 299226
rect 2892 299174 5982 299226
rect 6034 299174 6046 299226
rect 6098 299174 6110 299226
rect 6162 299174 6174 299226
rect 6226 299174 8832 299226
rect 1104 299152 8832 299174
rect 1104 298682 8832 298704
rect 1104 298630 4315 298682
rect 4367 298630 4379 298682
rect 4431 298630 4443 298682
rect 4495 298630 4507 298682
rect 4559 298630 7648 298682
rect 7700 298630 7712 298682
rect 7764 298630 7776 298682
rect 7828 298630 7840 298682
rect 7892 298630 8832 298682
rect 1104 298608 8832 298630
rect 1104 298138 8832 298160
rect 1104 298086 2648 298138
rect 2700 298086 2712 298138
rect 2764 298086 2776 298138
rect 2828 298086 2840 298138
rect 2892 298086 5982 298138
rect 6034 298086 6046 298138
rect 6098 298086 6110 298138
rect 6162 298086 6174 298138
rect 6226 298086 8832 298138
rect 1104 298064 8832 298086
rect 1104 297594 8832 297616
rect 1104 297542 4315 297594
rect 4367 297542 4379 297594
rect 4431 297542 4443 297594
rect 4495 297542 4507 297594
rect 4559 297542 7648 297594
rect 7700 297542 7712 297594
rect 7764 297542 7776 297594
rect 7828 297542 7840 297594
rect 7892 297542 8832 297594
rect 1104 297520 8832 297542
rect 1104 297050 8832 297072
rect 1104 296998 2648 297050
rect 2700 296998 2712 297050
rect 2764 296998 2776 297050
rect 2828 296998 2840 297050
rect 2892 296998 5982 297050
rect 6034 296998 6046 297050
rect 6098 296998 6110 297050
rect 6162 296998 6174 297050
rect 6226 296998 8832 297050
rect 1104 296976 8832 296998
rect 1104 296506 8832 296528
rect 1104 296454 4315 296506
rect 4367 296454 4379 296506
rect 4431 296454 4443 296506
rect 4495 296454 4507 296506
rect 4559 296454 7648 296506
rect 7700 296454 7712 296506
rect 7764 296454 7776 296506
rect 7828 296454 7840 296506
rect 7892 296454 8832 296506
rect 1104 296432 8832 296454
rect 1104 295962 8832 295984
rect 1104 295910 2648 295962
rect 2700 295910 2712 295962
rect 2764 295910 2776 295962
rect 2828 295910 2840 295962
rect 2892 295910 5982 295962
rect 6034 295910 6046 295962
rect 6098 295910 6110 295962
rect 6162 295910 6174 295962
rect 6226 295910 8832 295962
rect 1104 295888 8832 295910
rect 1104 295418 8832 295440
rect 1104 295366 4315 295418
rect 4367 295366 4379 295418
rect 4431 295366 4443 295418
rect 4495 295366 4507 295418
rect 4559 295366 7648 295418
rect 7700 295366 7712 295418
rect 7764 295366 7776 295418
rect 7828 295366 7840 295418
rect 7892 295366 8832 295418
rect 1104 295344 8832 295366
rect 1104 294874 8832 294896
rect 1104 294822 2648 294874
rect 2700 294822 2712 294874
rect 2764 294822 2776 294874
rect 2828 294822 2840 294874
rect 2892 294822 5982 294874
rect 6034 294822 6046 294874
rect 6098 294822 6110 294874
rect 6162 294822 6174 294874
rect 6226 294822 8832 294874
rect 1104 294800 8832 294822
rect 1104 294330 8832 294352
rect 1104 294278 4315 294330
rect 4367 294278 4379 294330
rect 4431 294278 4443 294330
rect 4495 294278 4507 294330
rect 4559 294278 7648 294330
rect 7700 294278 7712 294330
rect 7764 294278 7776 294330
rect 7828 294278 7840 294330
rect 7892 294278 8832 294330
rect 1104 294256 8832 294278
rect 1104 293786 8832 293808
rect 1104 293734 2648 293786
rect 2700 293734 2712 293786
rect 2764 293734 2776 293786
rect 2828 293734 2840 293786
rect 2892 293734 5982 293786
rect 6034 293734 6046 293786
rect 6098 293734 6110 293786
rect 6162 293734 6174 293786
rect 6226 293734 8832 293786
rect 1104 293712 8832 293734
rect 1104 293242 8832 293264
rect 1104 293190 4315 293242
rect 4367 293190 4379 293242
rect 4431 293190 4443 293242
rect 4495 293190 4507 293242
rect 4559 293190 7648 293242
rect 7700 293190 7712 293242
rect 7764 293190 7776 293242
rect 7828 293190 7840 293242
rect 7892 293190 8832 293242
rect 1104 293168 8832 293190
rect 1104 292698 8832 292720
rect 1104 292646 2648 292698
rect 2700 292646 2712 292698
rect 2764 292646 2776 292698
rect 2828 292646 2840 292698
rect 2892 292646 5982 292698
rect 6034 292646 6046 292698
rect 6098 292646 6110 292698
rect 6162 292646 6174 292698
rect 6226 292646 8832 292698
rect 1104 292624 8832 292646
rect 1104 292154 8832 292176
rect 1104 292102 4315 292154
rect 4367 292102 4379 292154
rect 4431 292102 4443 292154
rect 4495 292102 4507 292154
rect 4559 292102 7648 292154
rect 7700 292102 7712 292154
rect 7764 292102 7776 292154
rect 7828 292102 7840 292154
rect 7892 292102 8832 292154
rect 1104 292080 8832 292102
rect 1104 291610 8832 291632
rect 1104 291558 2648 291610
rect 2700 291558 2712 291610
rect 2764 291558 2776 291610
rect 2828 291558 2840 291610
rect 2892 291558 5982 291610
rect 6034 291558 6046 291610
rect 6098 291558 6110 291610
rect 6162 291558 6174 291610
rect 6226 291558 8832 291610
rect 1104 291536 8832 291558
rect 1104 291066 8832 291088
rect 1104 291014 4315 291066
rect 4367 291014 4379 291066
rect 4431 291014 4443 291066
rect 4495 291014 4507 291066
rect 4559 291014 7648 291066
rect 7700 291014 7712 291066
rect 7764 291014 7776 291066
rect 7828 291014 7840 291066
rect 7892 291014 8832 291066
rect 1104 290992 8832 291014
rect 1104 290522 8832 290544
rect 1104 290470 2648 290522
rect 2700 290470 2712 290522
rect 2764 290470 2776 290522
rect 2828 290470 2840 290522
rect 2892 290470 5982 290522
rect 6034 290470 6046 290522
rect 6098 290470 6110 290522
rect 6162 290470 6174 290522
rect 6226 290470 8832 290522
rect 1104 290448 8832 290470
rect 1104 289978 8832 290000
rect 1104 289926 4315 289978
rect 4367 289926 4379 289978
rect 4431 289926 4443 289978
rect 4495 289926 4507 289978
rect 4559 289926 7648 289978
rect 7700 289926 7712 289978
rect 7764 289926 7776 289978
rect 7828 289926 7840 289978
rect 7892 289926 8832 289978
rect 1104 289904 8832 289926
rect 1104 289434 8832 289456
rect 1104 289382 2648 289434
rect 2700 289382 2712 289434
rect 2764 289382 2776 289434
rect 2828 289382 2840 289434
rect 2892 289382 5982 289434
rect 6034 289382 6046 289434
rect 6098 289382 6110 289434
rect 6162 289382 6174 289434
rect 6226 289382 8832 289434
rect 1104 289360 8832 289382
rect 1104 288890 8832 288912
rect 1104 288838 4315 288890
rect 4367 288838 4379 288890
rect 4431 288838 4443 288890
rect 4495 288838 4507 288890
rect 4559 288838 7648 288890
rect 7700 288838 7712 288890
rect 7764 288838 7776 288890
rect 7828 288838 7840 288890
rect 7892 288838 8832 288890
rect 1104 288816 8832 288838
rect 1104 288346 8832 288368
rect 1104 288294 2648 288346
rect 2700 288294 2712 288346
rect 2764 288294 2776 288346
rect 2828 288294 2840 288346
rect 2892 288294 5982 288346
rect 6034 288294 6046 288346
rect 6098 288294 6110 288346
rect 6162 288294 6174 288346
rect 6226 288294 8832 288346
rect 1104 288272 8832 288294
rect 1104 287802 8832 287824
rect 1104 287750 4315 287802
rect 4367 287750 4379 287802
rect 4431 287750 4443 287802
rect 4495 287750 4507 287802
rect 4559 287750 7648 287802
rect 7700 287750 7712 287802
rect 7764 287750 7776 287802
rect 7828 287750 7840 287802
rect 7892 287750 8832 287802
rect 1104 287728 8832 287750
rect 1104 287258 8832 287280
rect 1104 287206 2648 287258
rect 2700 287206 2712 287258
rect 2764 287206 2776 287258
rect 2828 287206 2840 287258
rect 2892 287206 5982 287258
rect 6034 287206 6046 287258
rect 6098 287206 6110 287258
rect 6162 287206 6174 287258
rect 6226 287206 8832 287258
rect 1104 287184 8832 287206
rect 1104 286714 8832 286736
rect 1104 286662 4315 286714
rect 4367 286662 4379 286714
rect 4431 286662 4443 286714
rect 4495 286662 4507 286714
rect 4559 286662 7648 286714
rect 7700 286662 7712 286714
rect 7764 286662 7776 286714
rect 7828 286662 7840 286714
rect 7892 286662 8832 286714
rect 1104 286640 8832 286662
rect 1104 286170 8832 286192
rect 1104 286118 2648 286170
rect 2700 286118 2712 286170
rect 2764 286118 2776 286170
rect 2828 286118 2840 286170
rect 2892 286118 5982 286170
rect 6034 286118 6046 286170
rect 6098 286118 6110 286170
rect 6162 286118 6174 286170
rect 6226 286118 8832 286170
rect 1104 286096 8832 286118
rect 1104 285626 8832 285648
rect 1104 285574 4315 285626
rect 4367 285574 4379 285626
rect 4431 285574 4443 285626
rect 4495 285574 4507 285626
rect 4559 285574 7648 285626
rect 7700 285574 7712 285626
rect 7764 285574 7776 285626
rect 7828 285574 7840 285626
rect 7892 285574 8832 285626
rect 1104 285552 8832 285574
rect 1104 285082 8832 285104
rect 1104 285030 2648 285082
rect 2700 285030 2712 285082
rect 2764 285030 2776 285082
rect 2828 285030 2840 285082
rect 2892 285030 5982 285082
rect 6034 285030 6046 285082
rect 6098 285030 6110 285082
rect 6162 285030 6174 285082
rect 6226 285030 8832 285082
rect 1104 285008 8832 285030
rect 1104 284538 8832 284560
rect 1104 284486 4315 284538
rect 4367 284486 4379 284538
rect 4431 284486 4443 284538
rect 4495 284486 4507 284538
rect 4559 284486 7648 284538
rect 7700 284486 7712 284538
rect 7764 284486 7776 284538
rect 7828 284486 7840 284538
rect 7892 284486 8832 284538
rect 1104 284464 8832 284486
rect 1104 283994 8832 284016
rect 1104 283942 2648 283994
rect 2700 283942 2712 283994
rect 2764 283942 2776 283994
rect 2828 283942 2840 283994
rect 2892 283942 5982 283994
rect 6034 283942 6046 283994
rect 6098 283942 6110 283994
rect 6162 283942 6174 283994
rect 6226 283942 8832 283994
rect 1104 283920 8832 283942
rect 1104 283450 8832 283472
rect 1104 283398 4315 283450
rect 4367 283398 4379 283450
rect 4431 283398 4443 283450
rect 4495 283398 4507 283450
rect 4559 283398 7648 283450
rect 7700 283398 7712 283450
rect 7764 283398 7776 283450
rect 7828 283398 7840 283450
rect 7892 283398 8832 283450
rect 1104 283376 8832 283398
rect 1104 282906 8832 282928
rect 1104 282854 2648 282906
rect 2700 282854 2712 282906
rect 2764 282854 2776 282906
rect 2828 282854 2840 282906
rect 2892 282854 5982 282906
rect 6034 282854 6046 282906
rect 6098 282854 6110 282906
rect 6162 282854 6174 282906
rect 6226 282854 8832 282906
rect 1104 282832 8832 282854
rect 1104 282362 8832 282384
rect 1104 282310 4315 282362
rect 4367 282310 4379 282362
rect 4431 282310 4443 282362
rect 4495 282310 4507 282362
rect 4559 282310 7648 282362
rect 7700 282310 7712 282362
rect 7764 282310 7776 282362
rect 7828 282310 7840 282362
rect 7892 282310 8832 282362
rect 1104 282288 8832 282310
rect 1104 281818 8832 281840
rect 1104 281766 2648 281818
rect 2700 281766 2712 281818
rect 2764 281766 2776 281818
rect 2828 281766 2840 281818
rect 2892 281766 5982 281818
rect 6034 281766 6046 281818
rect 6098 281766 6110 281818
rect 6162 281766 6174 281818
rect 6226 281766 8832 281818
rect 1104 281744 8832 281766
rect 1104 281274 8832 281296
rect 1104 281222 4315 281274
rect 4367 281222 4379 281274
rect 4431 281222 4443 281274
rect 4495 281222 4507 281274
rect 4559 281222 7648 281274
rect 7700 281222 7712 281274
rect 7764 281222 7776 281274
rect 7828 281222 7840 281274
rect 7892 281222 8832 281274
rect 1104 281200 8832 281222
rect 1104 280730 8832 280752
rect 1104 280678 2648 280730
rect 2700 280678 2712 280730
rect 2764 280678 2776 280730
rect 2828 280678 2840 280730
rect 2892 280678 5982 280730
rect 6034 280678 6046 280730
rect 6098 280678 6110 280730
rect 6162 280678 6174 280730
rect 6226 280678 8832 280730
rect 1104 280656 8832 280678
rect 1104 280186 8832 280208
rect 1104 280134 4315 280186
rect 4367 280134 4379 280186
rect 4431 280134 4443 280186
rect 4495 280134 4507 280186
rect 4559 280134 7648 280186
rect 7700 280134 7712 280186
rect 7764 280134 7776 280186
rect 7828 280134 7840 280186
rect 7892 280134 8832 280186
rect 1104 280112 8832 280134
rect 1104 279642 8832 279664
rect 1104 279590 2648 279642
rect 2700 279590 2712 279642
rect 2764 279590 2776 279642
rect 2828 279590 2840 279642
rect 2892 279590 5982 279642
rect 6034 279590 6046 279642
rect 6098 279590 6110 279642
rect 6162 279590 6174 279642
rect 6226 279590 8832 279642
rect 1104 279568 8832 279590
rect 1104 279098 8832 279120
rect 1104 279046 4315 279098
rect 4367 279046 4379 279098
rect 4431 279046 4443 279098
rect 4495 279046 4507 279098
rect 4559 279046 7648 279098
rect 7700 279046 7712 279098
rect 7764 279046 7776 279098
rect 7828 279046 7840 279098
rect 7892 279046 8832 279098
rect 1104 279024 8832 279046
rect 1104 278554 8832 278576
rect 1104 278502 2648 278554
rect 2700 278502 2712 278554
rect 2764 278502 2776 278554
rect 2828 278502 2840 278554
rect 2892 278502 5982 278554
rect 6034 278502 6046 278554
rect 6098 278502 6110 278554
rect 6162 278502 6174 278554
rect 6226 278502 8832 278554
rect 1104 278480 8832 278502
rect 1104 278010 8832 278032
rect 1104 277958 4315 278010
rect 4367 277958 4379 278010
rect 4431 277958 4443 278010
rect 4495 277958 4507 278010
rect 4559 277958 7648 278010
rect 7700 277958 7712 278010
rect 7764 277958 7776 278010
rect 7828 277958 7840 278010
rect 7892 277958 8832 278010
rect 1104 277936 8832 277958
rect 1104 277466 8832 277488
rect 1104 277414 2648 277466
rect 2700 277414 2712 277466
rect 2764 277414 2776 277466
rect 2828 277414 2840 277466
rect 2892 277414 5982 277466
rect 6034 277414 6046 277466
rect 6098 277414 6110 277466
rect 6162 277414 6174 277466
rect 6226 277414 8832 277466
rect 1104 277392 8832 277414
rect 1104 276922 8832 276944
rect 1104 276870 4315 276922
rect 4367 276870 4379 276922
rect 4431 276870 4443 276922
rect 4495 276870 4507 276922
rect 4559 276870 7648 276922
rect 7700 276870 7712 276922
rect 7764 276870 7776 276922
rect 7828 276870 7840 276922
rect 7892 276870 8832 276922
rect 1104 276848 8832 276870
rect 1104 276378 8832 276400
rect 1104 276326 2648 276378
rect 2700 276326 2712 276378
rect 2764 276326 2776 276378
rect 2828 276326 2840 276378
rect 2892 276326 5982 276378
rect 6034 276326 6046 276378
rect 6098 276326 6110 276378
rect 6162 276326 6174 276378
rect 6226 276326 8832 276378
rect 1104 276304 8832 276326
rect 1104 275834 8832 275856
rect 1104 275782 4315 275834
rect 4367 275782 4379 275834
rect 4431 275782 4443 275834
rect 4495 275782 4507 275834
rect 4559 275782 7648 275834
rect 7700 275782 7712 275834
rect 7764 275782 7776 275834
rect 7828 275782 7840 275834
rect 7892 275782 8832 275834
rect 1104 275760 8832 275782
rect 1104 275290 8832 275312
rect 1104 275238 2648 275290
rect 2700 275238 2712 275290
rect 2764 275238 2776 275290
rect 2828 275238 2840 275290
rect 2892 275238 5982 275290
rect 6034 275238 6046 275290
rect 6098 275238 6110 275290
rect 6162 275238 6174 275290
rect 6226 275238 8832 275290
rect 1104 275216 8832 275238
rect 1104 274746 8832 274768
rect 1104 274694 4315 274746
rect 4367 274694 4379 274746
rect 4431 274694 4443 274746
rect 4495 274694 4507 274746
rect 4559 274694 7648 274746
rect 7700 274694 7712 274746
rect 7764 274694 7776 274746
rect 7828 274694 7840 274746
rect 7892 274694 8832 274746
rect 1104 274672 8832 274694
rect 1104 274202 8832 274224
rect 1104 274150 2648 274202
rect 2700 274150 2712 274202
rect 2764 274150 2776 274202
rect 2828 274150 2840 274202
rect 2892 274150 5982 274202
rect 6034 274150 6046 274202
rect 6098 274150 6110 274202
rect 6162 274150 6174 274202
rect 6226 274150 8832 274202
rect 1104 274128 8832 274150
rect 1104 273658 8832 273680
rect 1104 273606 4315 273658
rect 4367 273606 4379 273658
rect 4431 273606 4443 273658
rect 4495 273606 4507 273658
rect 4559 273606 7648 273658
rect 7700 273606 7712 273658
rect 7764 273606 7776 273658
rect 7828 273606 7840 273658
rect 7892 273606 8832 273658
rect 1104 273584 8832 273606
rect 1104 273114 8832 273136
rect 1104 273062 2648 273114
rect 2700 273062 2712 273114
rect 2764 273062 2776 273114
rect 2828 273062 2840 273114
rect 2892 273062 5982 273114
rect 6034 273062 6046 273114
rect 6098 273062 6110 273114
rect 6162 273062 6174 273114
rect 6226 273062 8832 273114
rect 1104 273040 8832 273062
rect 1104 272570 8832 272592
rect 1104 272518 4315 272570
rect 4367 272518 4379 272570
rect 4431 272518 4443 272570
rect 4495 272518 4507 272570
rect 4559 272518 7648 272570
rect 7700 272518 7712 272570
rect 7764 272518 7776 272570
rect 7828 272518 7840 272570
rect 7892 272518 8832 272570
rect 1104 272496 8832 272518
rect 1104 272026 8832 272048
rect 1104 271974 2648 272026
rect 2700 271974 2712 272026
rect 2764 271974 2776 272026
rect 2828 271974 2840 272026
rect 2892 271974 5982 272026
rect 6034 271974 6046 272026
rect 6098 271974 6110 272026
rect 6162 271974 6174 272026
rect 6226 271974 8832 272026
rect 1104 271952 8832 271974
rect 1104 271482 8832 271504
rect 1104 271430 4315 271482
rect 4367 271430 4379 271482
rect 4431 271430 4443 271482
rect 4495 271430 4507 271482
rect 4559 271430 7648 271482
rect 7700 271430 7712 271482
rect 7764 271430 7776 271482
rect 7828 271430 7840 271482
rect 7892 271430 8832 271482
rect 1104 271408 8832 271430
rect 1104 270938 8832 270960
rect 1104 270886 2648 270938
rect 2700 270886 2712 270938
rect 2764 270886 2776 270938
rect 2828 270886 2840 270938
rect 2892 270886 5982 270938
rect 6034 270886 6046 270938
rect 6098 270886 6110 270938
rect 6162 270886 6174 270938
rect 6226 270886 8832 270938
rect 1104 270864 8832 270886
rect 1104 270394 8832 270416
rect 1104 270342 4315 270394
rect 4367 270342 4379 270394
rect 4431 270342 4443 270394
rect 4495 270342 4507 270394
rect 4559 270342 7648 270394
rect 7700 270342 7712 270394
rect 7764 270342 7776 270394
rect 7828 270342 7840 270394
rect 7892 270342 8832 270394
rect 1104 270320 8832 270342
rect 1104 269850 8832 269872
rect 1104 269798 2648 269850
rect 2700 269798 2712 269850
rect 2764 269798 2776 269850
rect 2828 269798 2840 269850
rect 2892 269798 5982 269850
rect 6034 269798 6046 269850
rect 6098 269798 6110 269850
rect 6162 269798 6174 269850
rect 6226 269798 8832 269850
rect 1104 269776 8832 269798
rect 1104 269306 8832 269328
rect 1104 269254 4315 269306
rect 4367 269254 4379 269306
rect 4431 269254 4443 269306
rect 4495 269254 4507 269306
rect 4559 269254 7648 269306
rect 7700 269254 7712 269306
rect 7764 269254 7776 269306
rect 7828 269254 7840 269306
rect 7892 269254 8832 269306
rect 1104 269232 8832 269254
rect 1104 268762 8832 268784
rect 1104 268710 2648 268762
rect 2700 268710 2712 268762
rect 2764 268710 2776 268762
rect 2828 268710 2840 268762
rect 2892 268710 5982 268762
rect 6034 268710 6046 268762
rect 6098 268710 6110 268762
rect 6162 268710 6174 268762
rect 6226 268710 8832 268762
rect 1104 268688 8832 268710
rect 1104 268218 8832 268240
rect 1104 268166 4315 268218
rect 4367 268166 4379 268218
rect 4431 268166 4443 268218
rect 4495 268166 4507 268218
rect 4559 268166 7648 268218
rect 7700 268166 7712 268218
rect 7764 268166 7776 268218
rect 7828 268166 7840 268218
rect 7892 268166 8832 268218
rect 1104 268144 8832 268166
rect 1104 267674 8832 267696
rect 1104 267622 2648 267674
rect 2700 267622 2712 267674
rect 2764 267622 2776 267674
rect 2828 267622 2840 267674
rect 2892 267622 5982 267674
rect 6034 267622 6046 267674
rect 6098 267622 6110 267674
rect 6162 267622 6174 267674
rect 6226 267622 8832 267674
rect 1104 267600 8832 267622
rect 1104 267130 8832 267152
rect 1104 267078 4315 267130
rect 4367 267078 4379 267130
rect 4431 267078 4443 267130
rect 4495 267078 4507 267130
rect 4559 267078 7648 267130
rect 7700 267078 7712 267130
rect 7764 267078 7776 267130
rect 7828 267078 7840 267130
rect 7892 267078 8832 267130
rect 1104 267056 8832 267078
rect 1104 266586 8832 266608
rect 1104 266534 2648 266586
rect 2700 266534 2712 266586
rect 2764 266534 2776 266586
rect 2828 266534 2840 266586
rect 2892 266534 5982 266586
rect 6034 266534 6046 266586
rect 6098 266534 6110 266586
rect 6162 266534 6174 266586
rect 6226 266534 8832 266586
rect 1104 266512 8832 266534
rect 1104 266042 8832 266064
rect 1104 265990 4315 266042
rect 4367 265990 4379 266042
rect 4431 265990 4443 266042
rect 4495 265990 4507 266042
rect 4559 265990 7648 266042
rect 7700 265990 7712 266042
rect 7764 265990 7776 266042
rect 7828 265990 7840 266042
rect 7892 265990 8832 266042
rect 1104 265968 8832 265990
rect 1104 265498 8832 265520
rect 1104 265446 2648 265498
rect 2700 265446 2712 265498
rect 2764 265446 2776 265498
rect 2828 265446 2840 265498
rect 2892 265446 5982 265498
rect 6034 265446 6046 265498
rect 6098 265446 6110 265498
rect 6162 265446 6174 265498
rect 6226 265446 8832 265498
rect 1104 265424 8832 265446
rect 1104 264954 8832 264976
rect 1104 264902 4315 264954
rect 4367 264902 4379 264954
rect 4431 264902 4443 264954
rect 4495 264902 4507 264954
rect 4559 264902 7648 264954
rect 7700 264902 7712 264954
rect 7764 264902 7776 264954
rect 7828 264902 7840 264954
rect 7892 264902 8832 264954
rect 1104 264880 8832 264902
rect 1104 264410 8832 264432
rect 1104 264358 2648 264410
rect 2700 264358 2712 264410
rect 2764 264358 2776 264410
rect 2828 264358 2840 264410
rect 2892 264358 5982 264410
rect 6034 264358 6046 264410
rect 6098 264358 6110 264410
rect 6162 264358 6174 264410
rect 6226 264358 8832 264410
rect 1104 264336 8832 264358
rect 1104 263866 8832 263888
rect 1104 263814 4315 263866
rect 4367 263814 4379 263866
rect 4431 263814 4443 263866
rect 4495 263814 4507 263866
rect 4559 263814 7648 263866
rect 7700 263814 7712 263866
rect 7764 263814 7776 263866
rect 7828 263814 7840 263866
rect 7892 263814 8832 263866
rect 1104 263792 8832 263814
rect 1104 263322 8832 263344
rect 1104 263270 2648 263322
rect 2700 263270 2712 263322
rect 2764 263270 2776 263322
rect 2828 263270 2840 263322
rect 2892 263270 5982 263322
rect 6034 263270 6046 263322
rect 6098 263270 6110 263322
rect 6162 263270 6174 263322
rect 6226 263270 8832 263322
rect 1104 263248 8832 263270
rect 1104 262778 8832 262800
rect 1104 262726 4315 262778
rect 4367 262726 4379 262778
rect 4431 262726 4443 262778
rect 4495 262726 4507 262778
rect 4559 262726 7648 262778
rect 7700 262726 7712 262778
rect 7764 262726 7776 262778
rect 7828 262726 7840 262778
rect 7892 262726 8832 262778
rect 1104 262704 8832 262726
rect 1104 262234 8832 262256
rect 1104 262182 2648 262234
rect 2700 262182 2712 262234
rect 2764 262182 2776 262234
rect 2828 262182 2840 262234
rect 2892 262182 5982 262234
rect 6034 262182 6046 262234
rect 6098 262182 6110 262234
rect 6162 262182 6174 262234
rect 6226 262182 8832 262234
rect 1104 262160 8832 262182
rect 1104 261690 8832 261712
rect 1104 261638 4315 261690
rect 4367 261638 4379 261690
rect 4431 261638 4443 261690
rect 4495 261638 4507 261690
rect 4559 261638 7648 261690
rect 7700 261638 7712 261690
rect 7764 261638 7776 261690
rect 7828 261638 7840 261690
rect 7892 261638 8832 261690
rect 1104 261616 8832 261638
rect 1104 261146 8832 261168
rect 1104 261094 2648 261146
rect 2700 261094 2712 261146
rect 2764 261094 2776 261146
rect 2828 261094 2840 261146
rect 2892 261094 5982 261146
rect 6034 261094 6046 261146
rect 6098 261094 6110 261146
rect 6162 261094 6174 261146
rect 6226 261094 8832 261146
rect 1104 261072 8832 261094
rect 1104 260602 8832 260624
rect 1104 260550 4315 260602
rect 4367 260550 4379 260602
rect 4431 260550 4443 260602
rect 4495 260550 4507 260602
rect 4559 260550 7648 260602
rect 7700 260550 7712 260602
rect 7764 260550 7776 260602
rect 7828 260550 7840 260602
rect 7892 260550 8832 260602
rect 1104 260528 8832 260550
rect 1104 260058 8832 260080
rect 1104 260006 2648 260058
rect 2700 260006 2712 260058
rect 2764 260006 2776 260058
rect 2828 260006 2840 260058
rect 2892 260006 5982 260058
rect 6034 260006 6046 260058
rect 6098 260006 6110 260058
rect 6162 260006 6174 260058
rect 6226 260006 8832 260058
rect 1104 259984 8832 260006
rect 1104 259514 8832 259536
rect 1104 259462 4315 259514
rect 4367 259462 4379 259514
rect 4431 259462 4443 259514
rect 4495 259462 4507 259514
rect 4559 259462 7648 259514
rect 7700 259462 7712 259514
rect 7764 259462 7776 259514
rect 7828 259462 7840 259514
rect 7892 259462 8832 259514
rect 1104 259440 8832 259462
rect 1104 258970 8832 258992
rect 1104 258918 2648 258970
rect 2700 258918 2712 258970
rect 2764 258918 2776 258970
rect 2828 258918 2840 258970
rect 2892 258918 5982 258970
rect 6034 258918 6046 258970
rect 6098 258918 6110 258970
rect 6162 258918 6174 258970
rect 6226 258918 8832 258970
rect 1104 258896 8832 258918
rect 1104 258426 8832 258448
rect 1104 258374 4315 258426
rect 4367 258374 4379 258426
rect 4431 258374 4443 258426
rect 4495 258374 4507 258426
rect 4559 258374 7648 258426
rect 7700 258374 7712 258426
rect 7764 258374 7776 258426
rect 7828 258374 7840 258426
rect 7892 258374 8832 258426
rect 1104 258352 8832 258374
rect 1104 257882 8832 257904
rect 1104 257830 2648 257882
rect 2700 257830 2712 257882
rect 2764 257830 2776 257882
rect 2828 257830 2840 257882
rect 2892 257830 5982 257882
rect 6034 257830 6046 257882
rect 6098 257830 6110 257882
rect 6162 257830 6174 257882
rect 6226 257830 8832 257882
rect 1104 257808 8832 257830
rect 1104 257338 8832 257360
rect 1104 257286 4315 257338
rect 4367 257286 4379 257338
rect 4431 257286 4443 257338
rect 4495 257286 4507 257338
rect 4559 257286 7648 257338
rect 7700 257286 7712 257338
rect 7764 257286 7776 257338
rect 7828 257286 7840 257338
rect 7892 257286 8832 257338
rect 1104 257264 8832 257286
rect 1104 256794 8832 256816
rect 1104 256742 2648 256794
rect 2700 256742 2712 256794
rect 2764 256742 2776 256794
rect 2828 256742 2840 256794
rect 2892 256742 5982 256794
rect 6034 256742 6046 256794
rect 6098 256742 6110 256794
rect 6162 256742 6174 256794
rect 6226 256742 8832 256794
rect 1104 256720 8832 256742
rect 1104 256250 8832 256272
rect 1104 256198 4315 256250
rect 4367 256198 4379 256250
rect 4431 256198 4443 256250
rect 4495 256198 4507 256250
rect 4559 256198 7648 256250
rect 7700 256198 7712 256250
rect 7764 256198 7776 256250
rect 7828 256198 7840 256250
rect 7892 256198 8832 256250
rect 1104 256176 8832 256198
rect 1104 255706 8832 255728
rect 1104 255654 2648 255706
rect 2700 255654 2712 255706
rect 2764 255654 2776 255706
rect 2828 255654 2840 255706
rect 2892 255654 5982 255706
rect 6034 255654 6046 255706
rect 6098 255654 6110 255706
rect 6162 255654 6174 255706
rect 6226 255654 8832 255706
rect 1104 255632 8832 255654
rect 1104 255162 8832 255184
rect 1104 255110 4315 255162
rect 4367 255110 4379 255162
rect 4431 255110 4443 255162
rect 4495 255110 4507 255162
rect 4559 255110 7648 255162
rect 7700 255110 7712 255162
rect 7764 255110 7776 255162
rect 7828 255110 7840 255162
rect 7892 255110 8832 255162
rect 1104 255088 8832 255110
rect 1104 254618 8832 254640
rect 1104 254566 2648 254618
rect 2700 254566 2712 254618
rect 2764 254566 2776 254618
rect 2828 254566 2840 254618
rect 2892 254566 5982 254618
rect 6034 254566 6046 254618
rect 6098 254566 6110 254618
rect 6162 254566 6174 254618
rect 6226 254566 8832 254618
rect 1104 254544 8832 254566
rect 1104 254074 8832 254096
rect 1104 254022 4315 254074
rect 4367 254022 4379 254074
rect 4431 254022 4443 254074
rect 4495 254022 4507 254074
rect 4559 254022 7648 254074
rect 7700 254022 7712 254074
rect 7764 254022 7776 254074
rect 7828 254022 7840 254074
rect 7892 254022 8832 254074
rect 1104 254000 8832 254022
rect 1104 253530 8832 253552
rect 1104 253478 2648 253530
rect 2700 253478 2712 253530
rect 2764 253478 2776 253530
rect 2828 253478 2840 253530
rect 2892 253478 5982 253530
rect 6034 253478 6046 253530
rect 6098 253478 6110 253530
rect 6162 253478 6174 253530
rect 6226 253478 8832 253530
rect 1104 253456 8832 253478
rect 1104 252986 8832 253008
rect 1104 252934 4315 252986
rect 4367 252934 4379 252986
rect 4431 252934 4443 252986
rect 4495 252934 4507 252986
rect 4559 252934 7648 252986
rect 7700 252934 7712 252986
rect 7764 252934 7776 252986
rect 7828 252934 7840 252986
rect 7892 252934 8832 252986
rect 1104 252912 8832 252934
rect 1104 252442 8832 252464
rect 1104 252390 2648 252442
rect 2700 252390 2712 252442
rect 2764 252390 2776 252442
rect 2828 252390 2840 252442
rect 2892 252390 5982 252442
rect 6034 252390 6046 252442
rect 6098 252390 6110 252442
rect 6162 252390 6174 252442
rect 6226 252390 8832 252442
rect 1104 252368 8832 252390
rect 1104 251898 8832 251920
rect 1104 251846 4315 251898
rect 4367 251846 4379 251898
rect 4431 251846 4443 251898
rect 4495 251846 4507 251898
rect 4559 251846 7648 251898
rect 7700 251846 7712 251898
rect 7764 251846 7776 251898
rect 7828 251846 7840 251898
rect 7892 251846 8832 251898
rect 1104 251824 8832 251846
rect 1104 251354 8832 251376
rect 1104 251302 2648 251354
rect 2700 251302 2712 251354
rect 2764 251302 2776 251354
rect 2828 251302 2840 251354
rect 2892 251302 5982 251354
rect 6034 251302 6046 251354
rect 6098 251302 6110 251354
rect 6162 251302 6174 251354
rect 6226 251302 8832 251354
rect 1104 251280 8832 251302
rect 1104 250810 8832 250832
rect 1104 250758 4315 250810
rect 4367 250758 4379 250810
rect 4431 250758 4443 250810
rect 4495 250758 4507 250810
rect 4559 250758 7648 250810
rect 7700 250758 7712 250810
rect 7764 250758 7776 250810
rect 7828 250758 7840 250810
rect 7892 250758 8832 250810
rect 1104 250736 8832 250758
rect 1104 250266 8832 250288
rect 1104 250214 2648 250266
rect 2700 250214 2712 250266
rect 2764 250214 2776 250266
rect 2828 250214 2840 250266
rect 2892 250214 5982 250266
rect 6034 250214 6046 250266
rect 6098 250214 6110 250266
rect 6162 250214 6174 250266
rect 6226 250214 8832 250266
rect 1104 250192 8832 250214
rect 1104 249722 8832 249744
rect 1104 249670 4315 249722
rect 4367 249670 4379 249722
rect 4431 249670 4443 249722
rect 4495 249670 4507 249722
rect 4559 249670 7648 249722
rect 7700 249670 7712 249722
rect 7764 249670 7776 249722
rect 7828 249670 7840 249722
rect 7892 249670 8832 249722
rect 1104 249648 8832 249670
rect 1104 249178 8832 249200
rect 1104 249126 2648 249178
rect 2700 249126 2712 249178
rect 2764 249126 2776 249178
rect 2828 249126 2840 249178
rect 2892 249126 5982 249178
rect 6034 249126 6046 249178
rect 6098 249126 6110 249178
rect 6162 249126 6174 249178
rect 6226 249126 8832 249178
rect 1104 249104 8832 249126
rect 1104 248634 8832 248656
rect 1104 248582 4315 248634
rect 4367 248582 4379 248634
rect 4431 248582 4443 248634
rect 4495 248582 4507 248634
rect 4559 248582 7648 248634
rect 7700 248582 7712 248634
rect 7764 248582 7776 248634
rect 7828 248582 7840 248634
rect 7892 248582 8832 248634
rect 1104 248560 8832 248582
rect 1104 248090 8832 248112
rect 1104 248038 2648 248090
rect 2700 248038 2712 248090
rect 2764 248038 2776 248090
rect 2828 248038 2840 248090
rect 2892 248038 5982 248090
rect 6034 248038 6046 248090
rect 6098 248038 6110 248090
rect 6162 248038 6174 248090
rect 6226 248038 8832 248090
rect 1104 248016 8832 248038
rect 1104 247546 8832 247568
rect 1104 247494 4315 247546
rect 4367 247494 4379 247546
rect 4431 247494 4443 247546
rect 4495 247494 4507 247546
rect 4559 247494 7648 247546
rect 7700 247494 7712 247546
rect 7764 247494 7776 247546
rect 7828 247494 7840 247546
rect 7892 247494 8832 247546
rect 1104 247472 8832 247494
rect 1104 247002 8832 247024
rect 1104 246950 2648 247002
rect 2700 246950 2712 247002
rect 2764 246950 2776 247002
rect 2828 246950 2840 247002
rect 2892 246950 5982 247002
rect 6034 246950 6046 247002
rect 6098 246950 6110 247002
rect 6162 246950 6174 247002
rect 6226 246950 8832 247002
rect 1104 246928 8832 246950
rect 1104 246458 8832 246480
rect 1104 246406 4315 246458
rect 4367 246406 4379 246458
rect 4431 246406 4443 246458
rect 4495 246406 4507 246458
rect 4559 246406 7648 246458
rect 7700 246406 7712 246458
rect 7764 246406 7776 246458
rect 7828 246406 7840 246458
rect 7892 246406 8832 246458
rect 1104 246384 8832 246406
rect 1104 245914 8832 245936
rect 1104 245862 2648 245914
rect 2700 245862 2712 245914
rect 2764 245862 2776 245914
rect 2828 245862 2840 245914
rect 2892 245862 5982 245914
rect 6034 245862 6046 245914
rect 6098 245862 6110 245914
rect 6162 245862 6174 245914
rect 6226 245862 8832 245914
rect 1104 245840 8832 245862
rect 1104 245370 8832 245392
rect 1104 245318 4315 245370
rect 4367 245318 4379 245370
rect 4431 245318 4443 245370
rect 4495 245318 4507 245370
rect 4559 245318 7648 245370
rect 7700 245318 7712 245370
rect 7764 245318 7776 245370
rect 7828 245318 7840 245370
rect 7892 245318 8832 245370
rect 1104 245296 8832 245318
rect 1104 244826 8832 244848
rect 1104 244774 2648 244826
rect 2700 244774 2712 244826
rect 2764 244774 2776 244826
rect 2828 244774 2840 244826
rect 2892 244774 5982 244826
rect 6034 244774 6046 244826
rect 6098 244774 6110 244826
rect 6162 244774 6174 244826
rect 6226 244774 8832 244826
rect 1104 244752 8832 244774
rect 2222 244712 2228 244724
rect 2183 244684 2228 244712
rect 2222 244672 2228 244684
rect 2280 244672 2286 244724
rect 2041 244511 2099 244517
rect 2041 244477 2053 244511
rect 2087 244508 2099 244511
rect 2087 244480 2728 244508
rect 2087 244477 2099 244480
rect 2041 244471 2099 244477
rect 2700 244381 2728 244480
rect 2685 244375 2743 244381
rect 2685 244341 2697 244375
rect 2731 244372 2743 244375
rect 3510 244372 3516 244384
rect 2731 244344 3516 244372
rect 2731 244341 2743 244344
rect 2685 244335 2743 244341
rect 3510 244332 3516 244344
rect 3568 244332 3574 244384
rect 1104 244282 8832 244304
rect 1104 244230 4315 244282
rect 4367 244230 4379 244282
rect 4431 244230 4443 244282
rect 4495 244230 4507 244282
rect 4559 244230 7648 244282
rect 7700 244230 7712 244282
rect 7764 244230 7776 244282
rect 7828 244230 7840 244282
rect 7892 244230 8832 244282
rect 1104 244208 8832 244230
rect 1104 243738 8832 243760
rect 1104 243686 2648 243738
rect 2700 243686 2712 243738
rect 2764 243686 2776 243738
rect 2828 243686 2840 243738
rect 2892 243686 5982 243738
rect 6034 243686 6046 243738
rect 6098 243686 6110 243738
rect 6162 243686 6174 243738
rect 6226 243686 8832 243738
rect 1104 243664 8832 243686
rect 1104 243194 8832 243216
rect 1104 243142 4315 243194
rect 4367 243142 4379 243194
rect 4431 243142 4443 243194
rect 4495 243142 4507 243194
rect 4559 243142 7648 243194
rect 7700 243142 7712 243194
rect 7764 243142 7776 243194
rect 7828 243142 7840 243194
rect 7892 243142 8832 243194
rect 1104 243120 8832 243142
rect 1104 242650 8832 242672
rect 1104 242598 2648 242650
rect 2700 242598 2712 242650
rect 2764 242598 2776 242650
rect 2828 242598 2840 242650
rect 2892 242598 5982 242650
rect 6034 242598 6046 242650
rect 6098 242598 6110 242650
rect 6162 242598 6174 242650
rect 6226 242598 8832 242650
rect 1104 242576 8832 242598
rect 1104 242106 8832 242128
rect 1104 242054 4315 242106
rect 4367 242054 4379 242106
rect 4431 242054 4443 242106
rect 4495 242054 4507 242106
rect 4559 242054 7648 242106
rect 7700 242054 7712 242106
rect 7764 242054 7776 242106
rect 7828 242054 7840 242106
rect 7892 242054 8832 242106
rect 1104 242032 8832 242054
rect 7374 241952 7380 242004
rect 7432 241992 7438 242004
rect 7653 241995 7711 242001
rect 7653 241992 7665 241995
rect 7432 241964 7665 241992
rect 7432 241952 7438 241964
rect 7653 241961 7665 241964
rect 7699 241961 7711 241995
rect 7653 241955 7711 241961
rect 7466 241856 7472 241868
rect 7427 241828 7472 241856
rect 7466 241816 7472 241828
rect 7524 241816 7530 241868
rect 1104 241562 8832 241584
rect 1104 241510 2648 241562
rect 2700 241510 2712 241562
rect 2764 241510 2776 241562
rect 2828 241510 2840 241562
rect 2892 241510 5982 241562
rect 6034 241510 6046 241562
rect 6098 241510 6110 241562
rect 6162 241510 6174 241562
rect 6226 241510 8832 241562
rect 1104 241488 8832 241510
rect 7466 241108 7472 241120
rect 7427 241080 7472 241108
rect 7466 241068 7472 241080
rect 7524 241068 7530 241120
rect 1104 241018 8832 241040
rect 1104 240966 4315 241018
rect 4367 240966 4379 241018
rect 4431 240966 4443 241018
rect 4495 240966 4507 241018
rect 4559 240966 7648 241018
rect 7700 240966 7712 241018
rect 7764 240966 7776 241018
rect 7828 240966 7840 241018
rect 7892 240966 8832 241018
rect 1104 240944 8832 240966
rect 1104 240474 8832 240496
rect 1104 240422 2648 240474
rect 2700 240422 2712 240474
rect 2764 240422 2776 240474
rect 2828 240422 2840 240474
rect 2892 240422 5982 240474
rect 6034 240422 6046 240474
rect 6098 240422 6110 240474
rect 6162 240422 6174 240474
rect 6226 240422 8832 240474
rect 1104 240400 8832 240422
rect 1104 239930 8832 239952
rect 1104 239878 4315 239930
rect 4367 239878 4379 239930
rect 4431 239878 4443 239930
rect 4495 239878 4507 239930
rect 4559 239878 7648 239930
rect 7700 239878 7712 239930
rect 7764 239878 7776 239930
rect 7828 239878 7840 239930
rect 7892 239878 8832 239930
rect 1104 239856 8832 239878
rect 1104 239386 8832 239408
rect 1104 239334 2648 239386
rect 2700 239334 2712 239386
rect 2764 239334 2776 239386
rect 2828 239334 2840 239386
rect 2892 239334 5982 239386
rect 6034 239334 6046 239386
rect 6098 239334 6110 239386
rect 6162 239334 6174 239386
rect 6226 239334 8832 239386
rect 1104 239312 8832 239334
rect 6362 239232 6368 239284
rect 6420 239272 6426 239284
rect 7009 239275 7067 239281
rect 7009 239272 7021 239275
rect 6420 239244 7021 239272
rect 6420 239232 6426 239244
rect 7009 239241 7021 239244
rect 7055 239241 7067 239275
rect 7009 239235 7067 239241
rect 6822 239068 6828 239080
rect 6783 239040 6828 239068
rect 6822 239028 6828 239040
rect 6880 239068 6886 239080
rect 7377 239071 7435 239077
rect 7377 239068 7389 239071
rect 6880 239040 7389 239068
rect 6880 239028 6886 239040
rect 7377 239037 7389 239040
rect 7423 239037 7435 239071
rect 7377 239031 7435 239037
rect 1104 238842 8832 238864
rect 1104 238790 4315 238842
rect 4367 238790 4379 238842
rect 4431 238790 4443 238842
rect 4495 238790 4507 238842
rect 4559 238790 7648 238842
rect 7700 238790 7712 238842
rect 7764 238790 7776 238842
rect 7828 238790 7840 238842
rect 7892 238790 8832 238842
rect 1104 238768 8832 238790
rect 1104 238298 8832 238320
rect 1104 238246 2648 238298
rect 2700 238246 2712 238298
rect 2764 238246 2776 238298
rect 2828 238246 2840 238298
rect 2892 238246 5982 238298
rect 6034 238246 6046 238298
rect 6098 238246 6110 238298
rect 6162 238246 6174 238298
rect 6226 238246 8832 238298
rect 1104 238224 8832 238246
rect 1104 237754 8832 237776
rect 1104 237702 4315 237754
rect 4367 237702 4379 237754
rect 4431 237702 4443 237754
rect 4495 237702 4507 237754
rect 4559 237702 7648 237754
rect 7700 237702 7712 237754
rect 7764 237702 7776 237754
rect 7828 237702 7840 237754
rect 7892 237702 8832 237754
rect 1104 237680 8832 237702
rect 2498 237504 2504 237516
rect 2459 237476 2504 237504
rect 2498 237464 2504 237476
rect 2556 237464 2562 237516
rect 2685 237439 2743 237445
rect 2685 237405 2697 237439
rect 2731 237436 2743 237439
rect 2958 237436 2964 237448
rect 2731 237408 2964 237436
rect 2731 237405 2743 237408
rect 2685 237399 2743 237405
rect 2958 237396 2964 237408
rect 3016 237396 3022 237448
rect 3145 237303 3203 237309
rect 3145 237269 3157 237303
rect 3191 237300 3203 237303
rect 3510 237300 3516 237312
rect 3191 237272 3516 237300
rect 3191 237269 3203 237272
rect 3145 237263 3203 237269
rect 3510 237260 3516 237272
rect 3568 237260 3574 237312
rect 1104 237210 8832 237232
rect 1104 237158 2648 237210
rect 2700 237158 2712 237210
rect 2764 237158 2776 237210
rect 2828 237158 2840 237210
rect 2892 237158 5982 237210
rect 6034 237158 6046 237210
rect 6098 237158 6110 237210
rect 6162 237158 6174 237210
rect 6226 237158 8832 237210
rect 1104 237136 8832 237158
rect 2498 237096 2504 237108
rect 2459 237068 2504 237096
rect 2498 237056 2504 237068
rect 2556 237056 2562 237108
rect 2958 236756 2964 236768
rect 2871 236728 2964 236756
rect 2958 236716 2964 236728
rect 3016 236756 3022 236768
rect 3786 236756 3792 236768
rect 3016 236728 3792 236756
rect 3016 236716 3022 236728
rect 3786 236716 3792 236728
rect 3844 236716 3850 236768
rect 1104 236666 8832 236688
rect 1104 236614 4315 236666
rect 4367 236614 4379 236666
rect 4431 236614 4443 236666
rect 4495 236614 4507 236666
rect 4559 236614 7648 236666
rect 7700 236614 7712 236666
rect 7764 236614 7776 236666
rect 7828 236614 7840 236666
rect 7892 236614 8832 236666
rect 1104 236592 8832 236614
rect 1104 236122 8832 236144
rect 1104 236070 2648 236122
rect 2700 236070 2712 236122
rect 2764 236070 2776 236122
rect 2828 236070 2840 236122
rect 2892 236070 5982 236122
rect 6034 236070 6046 236122
rect 6098 236070 6110 236122
rect 6162 236070 6174 236122
rect 6226 236070 8832 236122
rect 1104 236048 8832 236070
rect 1104 235578 8832 235600
rect 1104 235526 4315 235578
rect 4367 235526 4379 235578
rect 4431 235526 4443 235578
rect 4495 235526 4507 235578
rect 4559 235526 7648 235578
rect 7700 235526 7712 235578
rect 7764 235526 7776 235578
rect 7828 235526 7840 235578
rect 7892 235526 8832 235578
rect 1104 235504 8832 235526
rect 1104 235034 8832 235056
rect 1104 234982 2648 235034
rect 2700 234982 2712 235034
rect 2764 234982 2776 235034
rect 2828 234982 2840 235034
rect 2892 234982 5982 235034
rect 6034 234982 6046 235034
rect 6098 234982 6110 235034
rect 6162 234982 6174 235034
rect 6226 234982 8832 235034
rect 1104 234960 8832 234982
rect 1104 234490 8832 234512
rect 1104 234438 4315 234490
rect 4367 234438 4379 234490
rect 4431 234438 4443 234490
rect 4495 234438 4507 234490
rect 4559 234438 7648 234490
rect 7700 234438 7712 234490
rect 7764 234438 7776 234490
rect 7828 234438 7840 234490
rect 7892 234438 8832 234490
rect 1104 234416 8832 234438
rect 4154 234268 4160 234320
rect 4212 234308 4218 234320
rect 4386 234311 4444 234317
rect 4386 234308 4398 234311
rect 4212 234280 4398 234308
rect 4212 234268 4218 234280
rect 4386 234277 4398 234280
rect 4432 234277 4444 234311
rect 4386 234271 4444 234277
rect 6730 234240 6736 234252
rect 6691 234212 6736 234240
rect 6730 234200 6736 234212
rect 6788 234200 6794 234252
rect 3970 234132 3976 234184
rect 4028 234172 4034 234184
rect 4065 234175 4123 234181
rect 4065 234172 4077 234175
rect 4028 234144 4077 234172
rect 4028 234132 4034 234144
rect 4065 234141 4077 234144
rect 4111 234141 4123 234175
rect 6914 234172 6920 234184
rect 6875 234144 6920 234172
rect 4065 234135 4123 234141
rect 6914 234132 6920 234144
rect 6972 234132 6978 234184
rect 4982 234036 4988 234048
rect 4943 234008 4988 234036
rect 4982 233996 4988 234008
rect 5040 233996 5046 234048
rect 7377 234039 7435 234045
rect 7377 234005 7389 234039
rect 7423 234036 7435 234039
rect 7466 234036 7472 234048
rect 7423 234008 7472 234036
rect 7423 234005 7435 234008
rect 7377 233999 7435 234005
rect 7466 233996 7472 234008
rect 7524 234036 7530 234048
rect 8202 234036 8208 234048
rect 7524 234008 8208 234036
rect 7524 233996 7530 234008
rect 8202 233996 8208 234008
rect 8260 233996 8266 234048
rect 1104 233946 8832 233968
rect 1104 233894 2648 233946
rect 2700 233894 2712 233946
rect 2764 233894 2776 233946
rect 2828 233894 2840 233946
rect 2892 233894 5982 233946
rect 6034 233894 6046 233946
rect 6098 233894 6110 233946
rect 6162 233894 6174 233946
rect 6226 233894 8832 233946
rect 1104 233872 8832 233894
rect 6730 233792 6736 233844
rect 6788 233832 6794 233844
rect 7009 233835 7067 233841
rect 7009 233832 7021 233835
rect 6788 233804 7021 233832
rect 6788 233792 6794 233804
rect 7009 233801 7021 233804
rect 7055 233801 7067 233835
rect 7009 233795 7067 233801
rect 3694 233724 3700 233776
rect 3752 233764 3758 233776
rect 5077 233767 5135 233773
rect 5077 233764 5089 233767
rect 3752 233736 5089 233764
rect 3752 233724 3758 233736
rect 5077 233733 5089 233736
rect 5123 233764 5135 233767
rect 6822 233764 6828 233776
rect 5123 233736 6828 233764
rect 5123 233733 5135 233736
rect 5077 233727 5135 233733
rect 6822 233724 6828 233736
rect 6880 233724 6886 233776
rect 4617 233699 4675 233705
rect 4617 233665 4629 233699
rect 4663 233696 4675 233699
rect 4982 233696 4988 233708
rect 4663 233668 4988 233696
rect 4663 233665 4675 233668
rect 4617 233659 4675 233665
rect 4982 233656 4988 233668
rect 5040 233656 5046 233708
rect 4433 233631 4491 233637
rect 4433 233597 4445 233631
rect 4479 233628 4491 233631
rect 4706 233628 4712 233640
rect 4479 233600 4712 233628
rect 4479 233597 4491 233600
rect 4433 233591 4491 233597
rect 4706 233588 4712 233600
rect 4764 233628 4770 233640
rect 5534 233628 5540 233640
rect 4764 233600 5540 233628
rect 4764 233588 4770 233600
rect 5534 233588 5540 233600
rect 5592 233588 5598 233640
rect 3789 233495 3847 233501
rect 3789 233461 3801 233495
rect 3835 233492 3847 233495
rect 3970 233492 3976 233504
rect 3835 233464 3976 233492
rect 3835 233461 3847 233464
rect 3789 233455 3847 233461
rect 3970 233452 3976 233464
rect 4028 233452 4034 233504
rect 4154 233452 4160 233504
rect 4212 233492 4218 233504
rect 4212 233464 4257 233492
rect 4212 233452 4218 233464
rect 5350 233452 5356 233504
rect 5408 233492 5414 233504
rect 6914 233492 6920 233504
rect 5408 233464 6920 233492
rect 5408 233452 5414 233464
rect 6914 233452 6920 233464
rect 6972 233492 6978 233504
rect 7377 233495 7435 233501
rect 7377 233492 7389 233495
rect 6972 233464 7389 233492
rect 6972 233452 6978 233464
rect 7377 233461 7389 233464
rect 7423 233461 7435 233495
rect 7377 233455 7435 233461
rect 1104 233402 8832 233424
rect 1104 233350 4315 233402
rect 4367 233350 4379 233402
rect 4431 233350 4443 233402
rect 4495 233350 4507 233402
rect 4559 233350 7648 233402
rect 7700 233350 7712 233402
rect 7764 233350 7776 233402
rect 7828 233350 7840 233402
rect 7892 233350 8832 233402
rect 1104 233328 8832 233350
rect 4525 233291 4583 233297
rect 4525 233257 4537 233291
rect 4571 233288 4583 233291
rect 4706 233288 4712 233300
rect 4571 233260 4712 233288
rect 4571 233257 4583 233260
rect 4525 233251 4583 233257
rect 4706 233248 4712 233260
rect 4764 233248 4770 233300
rect 4893 233291 4951 233297
rect 4893 233257 4905 233291
rect 4939 233288 4951 233291
rect 4982 233288 4988 233300
rect 4939 233260 4988 233288
rect 4939 233257 4951 233260
rect 4893 233251 4951 233257
rect 4982 233248 4988 233260
rect 5040 233248 5046 233300
rect 1104 232858 8832 232880
rect 1104 232806 2648 232858
rect 2700 232806 2712 232858
rect 2764 232806 2776 232858
rect 2828 232806 2840 232858
rect 2892 232806 5982 232858
rect 6034 232806 6046 232858
rect 6098 232806 6110 232858
rect 6162 232806 6174 232858
rect 6226 232806 8832 232858
rect 1104 232784 8832 232806
rect 3786 232744 3792 232756
rect 3747 232716 3792 232744
rect 3786 232704 3792 232716
rect 3844 232704 3850 232756
rect 2869 232543 2927 232549
rect 2869 232509 2881 232543
rect 2915 232540 2927 232543
rect 2958 232540 2964 232552
rect 2915 232512 2964 232540
rect 2915 232509 2927 232512
rect 2869 232503 2927 232509
rect 2958 232500 2964 232512
rect 3016 232500 3022 232552
rect 2777 232475 2835 232481
rect 2777 232441 2789 232475
rect 2823 232472 2835 232475
rect 3231 232475 3289 232481
rect 3231 232472 3243 232475
rect 2823 232444 3243 232472
rect 2823 232441 2835 232444
rect 2777 232435 2835 232441
rect 3231 232441 3243 232444
rect 3277 232472 3289 232475
rect 4062 232472 4068 232484
rect 3277 232444 4068 232472
rect 3277 232441 3289 232444
rect 3231 232435 3289 232441
rect 4062 232432 4068 232444
rect 4120 232472 4126 232484
rect 4154 232472 4160 232484
rect 4120 232444 4160 232472
rect 4120 232432 4126 232444
rect 4154 232432 4160 232444
rect 4212 232432 4218 232484
rect 1104 232314 8832 232336
rect 1104 232262 4315 232314
rect 4367 232262 4379 232314
rect 4431 232262 4443 232314
rect 4495 232262 4507 232314
rect 4559 232262 7648 232314
rect 7700 232262 7712 232314
rect 7764 232262 7776 232314
rect 7828 232262 7840 232314
rect 7892 232262 8832 232314
rect 1104 232240 8832 232262
rect 2958 231860 2964 231872
rect 2919 231832 2964 231860
rect 2958 231820 2964 231832
rect 3016 231820 3022 231872
rect 1104 231770 8832 231792
rect 1104 231718 2648 231770
rect 2700 231718 2712 231770
rect 2764 231718 2776 231770
rect 2828 231718 2840 231770
rect 2892 231718 5982 231770
rect 6034 231718 6046 231770
rect 6098 231718 6110 231770
rect 6162 231718 6174 231770
rect 6226 231718 8832 231770
rect 1104 231696 8832 231718
rect 1104 231226 8832 231248
rect 1104 231174 4315 231226
rect 4367 231174 4379 231226
rect 4431 231174 4443 231226
rect 4495 231174 4507 231226
rect 4559 231174 7648 231226
rect 7700 231174 7712 231226
rect 7764 231174 7776 231226
rect 7828 231174 7840 231226
rect 7892 231174 8832 231226
rect 1104 231152 8832 231174
rect 4706 231072 4712 231124
rect 4764 231112 4770 231124
rect 4801 231115 4859 231121
rect 4801 231112 4813 231115
rect 4764 231084 4813 231112
rect 4764 231072 4770 231084
rect 4801 231081 4813 231084
rect 4847 231081 4859 231115
rect 5350 231112 5356 231124
rect 5311 231084 5356 231112
rect 4801 231075 4859 231081
rect 5350 231072 5356 231084
rect 5408 231072 5414 231124
rect 4062 231004 4068 231056
rect 4120 231044 4126 231056
rect 4724 231044 4752 231072
rect 4120 231016 4752 231044
rect 4120 231004 4126 231016
rect 4433 230911 4491 230917
rect 4433 230877 4445 230911
rect 4479 230908 4491 230911
rect 4982 230908 4988 230920
rect 4479 230880 4988 230908
rect 4479 230877 4491 230880
rect 4433 230871 4491 230877
rect 4982 230868 4988 230880
rect 5040 230868 5046 230920
rect 2961 230775 3019 230781
rect 2961 230741 2973 230775
rect 3007 230772 3019 230775
rect 3786 230772 3792 230784
rect 3007 230744 3792 230772
rect 3007 230741 3019 230744
rect 2961 230735 3019 230741
rect 3786 230732 3792 230744
rect 3844 230732 3850 230784
rect 1104 230682 8832 230704
rect 1104 230630 2648 230682
rect 2700 230630 2712 230682
rect 2764 230630 2776 230682
rect 2828 230630 2840 230682
rect 2892 230630 5982 230682
rect 6034 230630 6046 230682
rect 6098 230630 6110 230682
rect 6162 230630 6174 230682
rect 6226 230630 8832 230682
rect 1104 230608 8832 230630
rect 2777 230503 2835 230509
rect 2777 230469 2789 230503
rect 2823 230500 2835 230503
rect 4062 230500 4068 230512
rect 2823 230472 4068 230500
rect 2823 230469 2835 230472
rect 2777 230463 2835 230469
rect 3160 230373 3188 230472
rect 4062 230460 4068 230472
rect 4120 230460 4126 230512
rect 3145 230367 3203 230373
rect 3145 230333 3157 230367
rect 3191 230333 3203 230367
rect 3145 230327 3203 230333
rect 3329 230367 3387 230373
rect 3329 230333 3341 230367
rect 3375 230333 3387 230367
rect 3329 230327 3387 230333
rect 3344 230296 3372 230327
rect 3418 230324 3424 230376
rect 3476 230364 3482 230376
rect 3697 230367 3755 230373
rect 3697 230364 3709 230367
rect 3476 230336 3709 230364
rect 3476 230324 3482 230336
rect 3697 230333 3709 230336
rect 3743 230333 3755 230367
rect 3697 230327 3755 230333
rect 3786 230324 3792 230376
rect 3844 230364 3850 230376
rect 4065 230367 4123 230373
rect 4065 230364 4077 230367
rect 3844 230336 4077 230364
rect 3844 230324 3850 230336
rect 4065 230333 4077 230336
rect 4111 230333 4123 230367
rect 4065 230327 4123 230333
rect 2424 230268 3372 230296
rect 2424 230240 2452 230268
rect 2406 230228 2412 230240
rect 2367 230200 2412 230228
rect 2406 230188 2412 230200
rect 2464 230188 2470 230240
rect 3970 230188 3976 230240
rect 4028 230228 4034 230240
rect 4065 230231 4123 230237
rect 4065 230228 4077 230231
rect 4028 230200 4077 230228
rect 4028 230188 4034 230200
rect 4065 230197 4077 230200
rect 4111 230197 4123 230231
rect 4706 230228 4712 230240
rect 4667 230200 4712 230228
rect 4065 230191 4123 230197
rect 4706 230188 4712 230200
rect 4764 230188 4770 230240
rect 4982 230228 4988 230240
rect 4943 230200 4988 230228
rect 4982 230188 4988 230200
rect 5040 230188 5046 230240
rect 1104 230138 8832 230160
rect 1104 230086 4315 230138
rect 4367 230086 4379 230138
rect 4431 230086 4443 230138
rect 4495 230086 4507 230138
rect 4559 230086 7648 230138
rect 7700 230086 7712 230138
rect 7764 230086 7776 230138
rect 7828 230086 7840 230138
rect 7892 230086 8832 230138
rect 1104 230064 8832 230086
rect 2961 230027 3019 230033
rect 2961 229993 2973 230027
rect 3007 230024 3019 230027
rect 3418 230024 3424 230036
rect 3007 229996 3424 230024
rect 3007 229993 3019 229996
rect 2961 229987 3019 229993
rect 3418 229984 3424 229996
rect 3476 229984 3482 230036
rect 3712 229996 4568 230024
rect 1486 229916 1492 229968
rect 1544 229956 1550 229968
rect 3712 229956 3740 229996
rect 1544 229928 3740 229956
rect 1544 229916 1550 229928
rect 3786 229916 3792 229968
rect 3844 229956 3850 229968
rect 4433 229959 4491 229965
rect 4433 229956 4445 229959
rect 3844 229928 4445 229956
rect 3844 229916 3850 229928
rect 4433 229925 4445 229928
rect 4479 229925 4491 229959
rect 4433 229919 4491 229925
rect 4062 229888 4068 229900
rect 4023 229860 4068 229888
rect 4062 229848 4068 229860
rect 4120 229848 4126 229900
rect 4249 229891 4307 229897
rect 4249 229857 4261 229891
rect 4295 229857 4307 229891
rect 4249 229851 4307 229857
rect 4341 229891 4399 229897
rect 4341 229857 4353 229891
rect 4387 229888 4399 229891
rect 4540 229888 4568 229996
rect 5074 229888 5080 229900
rect 4387 229860 5080 229888
rect 4387 229857 4399 229860
rect 4341 229851 4399 229857
rect 3050 229712 3056 229764
rect 3108 229752 3114 229764
rect 4264 229752 4292 229851
rect 5074 229848 5080 229860
rect 5132 229848 5138 229900
rect 4614 229780 4620 229832
rect 4672 229820 4678 229832
rect 4801 229823 4859 229829
rect 4801 229820 4813 229823
rect 4672 229792 4813 229820
rect 4672 229780 4678 229792
rect 4801 229789 4813 229792
rect 4847 229789 4859 229823
rect 4801 229783 4859 229789
rect 5350 229752 5356 229764
rect 3108 229724 5356 229752
rect 3108 229712 3114 229724
rect 5350 229712 5356 229724
rect 5408 229712 5414 229764
rect 2498 229644 2504 229696
rect 2556 229684 2562 229696
rect 3237 229687 3295 229693
rect 3237 229684 3249 229687
rect 2556 229656 3249 229684
rect 2556 229644 2562 229656
rect 3237 229653 3249 229656
rect 3283 229684 3295 229687
rect 3786 229684 3792 229696
rect 3283 229656 3792 229684
rect 3283 229653 3295 229656
rect 3237 229647 3295 229653
rect 3786 229644 3792 229656
rect 3844 229644 3850 229696
rect 1104 229594 8832 229616
rect 1104 229542 2648 229594
rect 2700 229542 2712 229594
rect 2764 229542 2776 229594
rect 2828 229542 2840 229594
rect 2892 229542 5982 229594
rect 6034 229542 6046 229594
rect 6098 229542 6110 229594
rect 6162 229542 6174 229594
rect 6226 229542 8832 229594
rect 1104 229520 8832 229542
rect 2777 229483 2835 229489
rect 2777 229449 2789 229483
rect 2823 229480 2835 229483
rect 3418 229480 3424 229492
rect 2823 229452 3424 229480
rect 2823 229449 2835 229452
rect 2777 229443 2835 229449
rect 3418 229440 3424 229452
rect 3476 229440 3482 229492
rect 5350 229480 5356 229492
rect 5311 229452 5356 229480
rect 5350 229440 5356 229452
rect 5408 229440 5414 229492
rect 5074 229412 5080 229424
rect 5035 229384 5080 229412
rect 5074 229372 5080 229384
rect 5132 229372 5138 229424
rect 2041 229347 2099 229353
rect 2041 229313 2053 229347
rect 2087 229344 2099 229347
rect 2406 229344 2412 229356
rect 2087 229316 2412 229344
rect 2087 229313 2099 229316
rect 2041 229307 2099 229313
rect 2406 229304 2412 229316
rect 2464 229344 2470 229356
rect 4341 229347 4399 229353
rect 2464 229316 3372 229344
rect 2464 229304 2470 229316
rect 3344 229285 3372 229316
rect 4341 229313 4353 229347
rect 4387 229344 4399 229347
rect 4982 229344 4988 229356
rect 4387 229316 4988 229344
rect 4387 229313 4399 229316
rect 4341 229307 4399 229313
rect 4982 229304 4988 229316
rect 5040 229304 5046 229356
rect 2869 229279 2927 229285
rect 2869 229276 2881 229279
rect 2424 229248 2881 229276
rect 2424 229152 2452 229248
rect 2869 229245 2881 229248
rect 2915 229245 2927 229279
rect 2869 229239 2927 229245
rect 3329 229279 3387 229285
rect 3329 229245 3341 229279
rect 3375 229245 3387 229279
rect 3329 229239 3387 229245
rect 3344 229208 3372 229239
rect 3418 229236 3424 229288
rect 3476 229276 3482 229288
rect 3697 229279 3755 229285
rect 3697 229276 3709 229279
rect 3476 229248 3709 229276
rect 3476 229236 3482 229248
rect 3697 229245 3709 229248
rect 3743 229245 3755 229279
rect 3697 229239 3755 229245
rect 3786 229236 3792 229288
rect 3844 229276 3850 229288
rect 4065 229279 4123 229285
rect 4065 229276 4077 229279
rect 3844 229248 4077 229276
rect 3844 229236 3850 229248
rect 4065 229245 4077 229248
rect 4111 229276 4123 229279
rect 5721 229279 5779 229285
rect 5721 229276 5733 229279
rect 4111 229248 5733 229276
rect 4111 229245 4123 229248
rect 4065 229239 4123 229245
rect 5721 229245 5733 229248
rect 5767 229245 5779 229279
rect 5721 229239 5779 229245
rect 3602 229208 3608 229220
rect 3344 229180 3608 229208
rect 3602 229168 3608 229180
rect 3660 229168 3666 229220
rect 2406 229140 2412 229152
rect 2367 229112 2412 229140
rect 2406 229100 2412 229112
rect 2464 229100 2470 229152
rect 4062 229100 4068 229152
rect 4120 229140 4126 229152
rect 4709 229143 4767 229149
rect 4709 229140 4721 229143
rect 4120 229112 4721 229140
rect 4120 229100 4126 229112
rect 4709 229109 4721 229112
rect 4755 229140 4767 229143
rect 4798 229140 4804 229152
rect 4755 229112 4804 229140
rect 4755 229109 4767 229112
rect 4709 229103 4767 229109
rect 4798 229100 4804 229112
rect 4856 229100 4862 229152
rect 1104 229050 8832 229072
rect 1104 228998 4315 229050
rect 4367 228998 4379 229050
rect 4431 228998 4443 229050
rect 4495 228998 4507 229050
rect 4559 228998 7648 229050
rect 7700 228998 7712 229050
rect 7764 228998 7776 229050
rect 7828 228998 7840 229050
rect 7892 228998 8832 229050
rect 1104 228976 8832 228998
rect 2593 228939 2651 228945
rect 2593 228905 2605 228939
rect 2639 228936 2651 228939
rect 3050 228936 3056 228948
rect 2639 228908 3056 228936
rect 2639 228905 2651 228908
rect 2593 228899 2651 228905
rect 3050 228896 3056 228908
rect 3108 228896 3114 228948
rect 3418 228936 3424 228948
rect 3379 228908 3424 228936
rect 3418 228896 3424 228908
rect 3476 228896 3482 228948
rect 2498 228828 2504 228880
rect 2556 228868 2562 228880
rect 2777 228871 2835 228877
rect 2777 228868 2789 228871
rect 2556 228840 2789 228868
rect 2556 228828 2562 228840
rect 2777 228837 2789 228840
rect 2823 228837 2835 228871
rect 2777 228831 2835 228837
rect 1486 228760 1492 228812
rect 1544 228800 1550 228812
rect 2685 228803 2743 228809
rect 2685 228800 2697 228803
rect 1544 228772 2697 228800
rect 1544 228760 1550 228772
rect 2685 228769 2697 228772
rect 2731 228769 2743 228803
rect 4065 228803 4123 228809
rect 4065 228800 4077 228803
rect 2685 228763 2743 228769
rect 2792 228772 4077 228800
rect 1762 228692 1768 228744
rect 1820 228732 1826 228744
rect 2406 228732 2412 228744
rect 1820 228704 2412 228732
rect 1820 228692 1826 228704
rect 2406 228692 2412 228704
rect 2464 228732 2470 228744
rect 2792 228732 2820 228772
rect 4065 228769 4077 228772
rect 4111 228769 4123 228803
rect 4065 228763 4123 228769
rect 4709 228803 4767 228809
rect 4709 228769 4721 228803
rect 4755 228800 4767 228803
rect 4798 228800 4804 228812
rect 4755 228772 4804 228800
rect 4755 228769 4767 228772
rect 4709 228763 4767 228769
rect 4798 228760 4804 228772
rect 4856 228760 4862 228812
rect 3142 228732 3148 228744
rect 2464 228704 2820 228732
rect 3103 228704 3148 228732
rect 2464 228692 2470 228704
rect 3142 228692 3148 228704
rect 3200 228692 3206 228744
rect 2317 228599 2375 228605
rect 2317 228565 2329 228599
rect 2363 228596 2375 228599
rect 2406 228596 2412 228608
rect 2363 228568 2412 228596
rect 2363 228565 2375 228568
rect 2317 228559 2375 228565
rect 2406 228556 2412 228568
rect 2464 228556 2470 228608
rect 1104 228506 8832 228528
rect 1104 228454 2648 228506
rect 2700 228454 2712 228506
rect 2764 228454 2776 228506
rect 2828 228454 2840 228506
rect 2892 228454 5982 228506
rect 6034 228454 6046 228506
rect 6098 228454 6110 228506
rect 6162 228454 6174 228506
rect 6226 228454 8832 228506
rect 1104 228432 8832 228454
rect 1486 228352 1492 228404
rect 1544 228392 1550 228404
rect 2038 228392 2044 228404
rect 1544 228364 2044 228392
rect 1544 228352 1550 228364
rect 2038 228352 2044 228364
rect 2096 228352 2102 228404
rect 1210 228284 1216 228336
rect 1268 228324 1274 228336
rect 2409 228327 2467 228333
rect 2409 228324 2421 228327
rect 1268 228296 2421 228324
rect 1268 228284 1274 228296
rect 2409 228293 2421 228296
rect 2455 228293 2467 228327
rect 2409 228287 2467 228293
rect 2869 228327 2927 228333
rect 2869 228293 2881 228327
rect 2915 228324 2927 228327
rect 3234 228324 3240 228336
rect 2915 228296 3240 228324
rect 2915 228293 2927 228296
rect 2869 228287 2927 228293
rect 1762 228052 1768 228064
rect 1723 228024 1768 228052
rect 1762 228012 1768 228024
rect 1820 228012 1826 228064
rect 2314 228012 2320 228064
rect 2372 228052 2378 228064
rect 2424 228052 2452 228287
rect 3234 228284 3240 228296
rect 3292 228284 3298 228336
rect 2958 228216 2964 228268
rect 3016 228256 3022 228268
rect 3697 228259 3755 228265
rect 3697 228256 3709 228259
rect 3016 228228 3709 228256
rect 3016 228216 3022 228228
rect 3697 228225 3709 228228
rect 3743 228225 3755 228259
rect 3697 228219 3755 228225
rect 3050 228148 3056 228200
rect 3108 228188 3114 228200
rect 3313 228191 3371 228197
rect 3313 228188 3325 228191
rect 3108 228160 3325 228188
rect 3108 228148 3114 228160
rect 3313 228157 3325 228160
rect 3359 228157 3371 228191
rect 3313 228151 3371 228157
rect 2958 228120 2964 228132
rect 2919 228092 2964 228120
rect 2958 228080 2964 228092
rect 3016 228080 3022 228132
rect 3145 228055 3203 228061
rect 3145 228052 3157 228055
rect 2372 228024 3157 228052
rect 2372 228012 2378 228024
rect 3145 228021 3157 228024
rect 3191 228021 3203 228055
rect 3145 228015 3203 228021
rect 3234 228012 3240 228064
rect 3292 228052 3298 228064
rect 4157 228055 4215 228061
rect 4157 228052 4169 228055
rect 3292 228024 4169 228052
rect 3292 228012 3298 228024
rect 4157 228021 4169 228024
rect 4203 228052 4215 228055
rect 4798 228052 4804 228064
rect 4203 228024 4804 228052
rect 4203 228021 4215 228024
rect 4157 228015 4215 228021
rect 4798 228012 4804 228024
rect 4856 228012 4862 228064
rect 1104 227962 8832 227984
rect 1104 227910 4315 227962
rect 4367 227910 4379 227962
rect 4431 227910 4443 227962
rect 4495 227910 4507 227962
rect 4559 227910 7648 227962
rect 7700 227910 7712 227962
rect 7764 227910 7776 227962
rect 7828 227910 7840 227962
rect 7892 227910 8832 227962
rect 1104 227888 8832 227910
rect 2958 227808 2964 227860
rect 3016 227848 3022 227860
rect 3053 227851 3111 227857
rect 3053 227848 3065 227851
rect 3016 227820 3065 227848
rect 3016 227808 3022 227820
rect 3053 227817 3065 227820
rect 3099 227848 3111 227851
rect 3418 227848 3424 227860
rect 3099 227820 3424 227848
rect 3099 227817 3111 227820
rect 3053 227811 3111 227817
rect 3418 227808 3424 227820
rect 3476 227808 3482 227860
rect 2038 227672 2044 227724
rect 2096 227712 2102 227724
rect 2869 227715 2927 227721
rect 2869 227712 2881 227715
rect 2096 227684 2881 227712
rect 2096 227672 2102 227684
rect 2869 227681 2881 227684
rect 2915 227681 2927 227715
rect 2869 227675 2927 227681
rect 2501 227511 2559 227517
rect 2501 227477 2513 227511
rect 2547 227508 2559 227511
rect 3050 227508 3056 227520
rect 2547 227480 3056 227508
rect 2547 227477 2559 227480
rect 2501 227471 2559 227477
rect 3050 227468 3056 227480
rect 3108 227508 3114 227520
rect 3326 227508 3332 227520
rect 3108 227480 3332 227508
rect 3108 227468 3114 227480
rect 3326 227468 3332 227480
rect 3384 227468 3390 227520
rect 3602 227468 3608 227520
rect 3660 227508 3666 227520
rect 3697 227511 3755 227517
rect 3697 227508 3709 227511
rect 3660 227480 3709 227508
rect 3660 227468 3666 227480
rect 3697 227477 3709 227480
rect 3743 227477 3755 227511
rect 3697 227471 3755 227477
rect 1104 227418 8832 227440
rect 1104 227366 2648 227418
rect 2700 227366 2712 227418
rect 2764 227366 2776 227418
rect 2828 227366 2840 227418
rect 2892 227366 5982 227418
rect 6034 227366 6046 227418
rect 6098 227366 6110 227418
rect 6162 227366 6174 227418
rect 6226 227366 8832 227418
rect 1104 227344 8832 227366
rect 2038 227304 2044 227316
rect 1999 227276 2044 227304
rect 2038 227264 2044 227276
rect 2096 227264 2102 227316
rect 2314 227304 2320 227316
rect 2275 227276 2320 227304
rect 2314 227264 2320 227276
rect 2372 227264 2378 227316
rect 2314 227128 2320 227180
rect 2372 227168 2378 227180
rect 2372 227140 4108 227168
rect 2372 227128 2378 227140
rect 2777 227103 2835 227109
rect 2777 227069 2789 227103
rect 2823 227100 2835 227103
rect 3145 227103 3203 227109
rect 3145 227100 3157 227103
rect 2823 227072 3157 227100
rect 2823 227069 2835 227072
rect 2777 227063 2835 227069
rect 3145 227069 3157 227072
rect 3191 227100 3203 227103
rect 3234 227100 3240 227112
rect 3191 227072 3240 227100
rect 3191 227069 3203 227072
rect 3145 227063 3203 227069
rect 3234 227060 3240 227072
rect 3292 227060 3298 227112
rect 3329 227103 3387 227109
rect 3329 227069 3341 227103
rect 3375 227069 3387 227103
rect 3329 227063 3387 227069
rect 3344 227032 3372 227063
rect 3418 227060 3424 227112
rect 3476 227100 3482 227112
rect 4080 227109 4108 227140
rect 3697 227103 3755 227109
rect 3697 227100 3709 227103
rect 3476 227072 3709 227100
rect 3476 227060 3482 227072
rect 3697 227069 3709 227072
rect 3743 227069 3755 227103
rect 3697 227063 3755 227069
rect 4065 227103 4123 227109
rect 4065 227069 4077 227103
rect 4111 227069 4123 227103
rect 4065 227063 4123 227069
rect 3602 227032 3608 227044
rect 3344 227004 3608 227032
rect 3050 226924 3056 226976
rect 3108 226964 3114 226976
rect 3344 226964 3372 227004
rect 3602 226992 3608 227004
rect 3660 226992 3666 227044
rect 4062 226964 4068 226976
rect 3108 226936 3372 226964
rect 4023 226936 4068 226964
rect 3108 226924 3114 226936
rect 4062 226924 4068 226936
rect 4120 226924 4126 226976
rect 1104 226874 8832 226896
rect 1104 226822 4315 226874
rect 4367 226822 4379 226874
rect 4431 226822 4443 226874
rect 4495 226822 4507 226874
rect 4559 226822 7648 226874
rect 7700 226822 7712 226874
rect 7764 226822 7776 226874
rect 7828 226822 7840 226874
rect 7892 226822 8832 226874
rect 1104 226800 8832 226822
rect 3418 226760 3424 226772
rect 3379 226732 3424 226760
rect 3418 226720 3424 226732
rect 3476 226720 3482 226772
rect 4706 226720 4712 226772
rect 4764 226760 4770 226772
rect 4801 226763 4859 226769
rect 4801 226760 4813 226763
rect 4764 226732 4813 226760
rect 4764 226720 4770 226732
rect 4801 226729 4813 226732
rect 4847 226729 4859 226763
rect 4801 226723 4859 226729
rect 2406 226692 2412 226704
rect 2367 226664 2412 226692
rect 2406 226652 2412 226664
rect 2464 226652 2470 226704
rect 2314 226584 2320 226636
rect 2372 226624 2378 226636
rect 2501 226627 2559 226633
rect 2501 226624 2513 226627
rect 2372 226596 2513 226624
rect 2372 226584 2378 226596
rect 2501 226593 2513 226596
rect 2547 226593 2559 226627
rect 2501 226587 2559 226593
rect 4433 226627 4491 226633
rect 4433 226593 4445 226627
rect 4479 226624 4491 226627
rect 4614 226624 4620 226636
rect 4479 226596 4620 226624
rect 4479 226593 4491 226596
rect 4433 226587 4491 226593
rect 4614 226584 4620 226596
rect 4672 226584 4678 226636
rect 5353 226423 5411 226429
rect 5353 226389 5365 226423
rect 5399 226420 5411 226423
rect 5810 226420 5816 226432
rect 5399 226392 5816 226420
rect 5399 226389 5411 226392
rect 5353 226383 5411 226389
rect 5810 226380 5816 226392
rect 5868 226380 5874 226432
rect 1104 226330 8832 226352
rect 1104 226278 2648 226330
rect 2700 226278 2712 226330
rect 2764 226278 2776 226330
rect 2828 226278 2840 226330
rect 2892 226278 5982 226330
rect 6034 226278 6046 226330
rect 6098 226278 6110 226330
rect 6162 226278 6174 226330
rect 6226 226278 8832 226330
rect 1104 226256 8832 226278
rect 2314 226176 2320 226228
rect 2372 226216 2378 226228
rect 2409 226219 2467 226225
rect 2409 226216 2421 226219
rect 2372 226188 2421 226216
rect 2372 226176 2378 226188
rect 2409 226185 2421 226188
rect 2455 226185 2467 226219
rect 2409 226179 2467 226185
rect 3142 226176 3148 226228
rect 3200 226216 3206 226228
rect 3513 226219 3571 226225
rect 3513 226216 3525 226219
rect 3200 226188 3525 226216
rect 3200 226176 3206 226188
rect 3513 226185 3525 226188
rect 3559 226216 3571 226219
rect 3559 226188 4476 226216
rect 3559 226185 3571 226188
rect 3513 226179 3571 226185
rect 4448 226089 4476 226188
rect 4614 226176 4620 226228
rect 4672 226216 4678 226228
rect 5629 226219 5687 226225
rect 5629 226216 5641 226219
rect 4672 226188 5641 226216
rect 4672 226176 4678 226188
rect 5629 226185 5641 226188
rect 5675 226185 5687 226219
rect 5629 226179 5687 226185
rect 4433 226083 4491 226089
rect 4433 226049 4445 226083
rect 4479 226049 4491 226083
rect 4433 226043 4491 226049
rect 3973 226015 4031 226021
rect 3973 225981 3985 226015
rect 4019 226012 4031 226015
rect 4019 225984 4154 226012
rect 4019 225981 4031 225984
rect 3973 225975 4031 225981
rect 4126 225944 4154 225984
rect 4341 225947 4399 225953
rect 4341 225944 4353 225947
rect 4126 225916 4353 225944
rect 4341 225913 4353 225916
rect 4387 225944 4399 225947
rect 4706 225944 4712 225956
rect 4387 225916 4712 225944
rect 4387 225913 4399 225916
rect 4341 225907 4399 225913
rect 4706 225904 4712 225916
rect 4764 225953 4770 225956
rect 4764 225947 4812 225953
rect 4764 225913 4766 225947
rect 4800 225913 4812 225947
rect 4764 225907 4812 225913
rect 4764 225904 4770 225907
rect 5353 225879 5411 225885
rect 5353 225845 5365 225879
rect 5399 225876 5411 225879
rect 7006 225876 7012 225888
rect 5399 225848 7012 225876
rect 5399 225845 5411 225848
rect 5353 225839 5411 225845
rect 7006 225836 7012 225848
rect 7064 225836 7070 225888
rect 1104 225786 8832 225808
rect 1104 225734 4315 225786
rect 4367 225734 4379 225786
rect 4431 225734 4443 225786
rect 4495 225734 4507 225786
rect 4559 225734 7648 225786
rect 7700 225734 7712 225786
rect 7764 225734 7776 225786
rect 7828 225734 7840 225786
rect 7892 225734 8832 225786
rect 1104 225712 8832 225734
rect 4706 225632 4712 225684
rect 4764 225672 4770 225684
rect 4801 225675 4859 225681
rect 4801 225672 4813 225675
rect 4764 225644 4813 225672
rect 4764 225632 4770 225644
rect 4801 225641 4813 225644
rect 4847 225641 4859 225675
rect 4801 225635 4859 225641
rect 4062 225496 4068 225548
rect 4120 225536 4126 225548
rect 4433 225539 4491 225545
rect 4433 225536 4445 225539
rect 4120 225508 4445 225536
rect 4120 225496 4126 225508
rect 4433 225505 4445 225508
rect 4479 225505 4491 225539
rect 6270 225536 6276 225548
rect 6231 225508 6276 225536
rect 4433 225499 4491 225505
rect 6270 225496 6276 225508
rect 6328 225496 6334 225548
rect 5810 225428 5816 225480
rect 5868 225468 5874 225480
rect 6457 225471 6515 225477
rect 6457 225468 6469 225471
rect 5868 225440 6469 225468
rect 5868 225428 5874 225440
rect 6457 225437 6469 225440
rect 6503 225437 6515 225471
rect 6457 225431 6515 225437
rect 5350 225332 5356 225344
rect 5311 225304 5356 225332
rect 5350 225292 5356 225304
rect 5408 225292 5414 225344
rect 5626 225292 5632 225344
rect 5684 225332 5690 225344
rect 6641 225335 6699 225341
rect 6641 225332 6653 225335
rect 5684 225304 6653 225332
rect 5684 225292 5690 225304
rect 6641 225301 6653 225304
rect 6687 225301 6699 225335
rect 6641 225295 6699 225301
rect 1104 225242 8832 225264
rect 1104 225190 2648 225242
rect 2700 225190 2712 225242
rect 2764 225190 2776 225242
rect 2828 225190 2840 225242
rect 2892 225190 5982 225242
rect 6034 225190 6046 225242
rect 6098 225190 6110 225242
rect 6162 225190 6174 225242
rect 6226 225190 8832 225242
rect 1104 225168 8832 225190
rect 4062 225088 4068 225140
rect 4120 225128 4126 225140
rect 4801 225131 4859 225137
rect 4801 225128 4813 225131
rect 4120 225100 4813 225128
rect 4120 225088 4126 225100
rect 4801 225097 4813 225100
rect 4847 225097 4859 225131
rect 4801 225091 4859 225097
rect 5810 225088 5816 225140
rect 5868 225128 5874 225140
rect 5905 225131 5963 225137
rect 5905 225128 5917 225131
rect 5868 225100 5917 225128
rect 5868 225088 5874 225100
rect 5905 225097 5917 225100
rect 5951 225097 5963 225131
rect 6270 225128 6276 225140
rect 6231 225100 6276 225128
rect 5905 225091 5963 225097
rect 6270 225088 6276 225100
rect 6328 225088 6334 225140
rect 3970 225020 3976 225072
rect 4028 225060 4034 225072
rect 4525 225063 4583 225069
rect 4525 225060 4537 225063
rect 4028 225032 4537 225060
rect 4028 225020 4034 225032
rect 4525 225029 4537 225032
rect 4571 225060 4583 225063
rect 4706 225060 4712 225072
rect 4571 225032 4712 225060
rect 4571 225029 4583 225032
rect 4525 225023 4583 225029
rect 4706 225020 4712 225032
rect 4764 225020 4770 225072
rect 6825 224995 6883 225001
rect 6825 224961 6837 224995
rect 6871 224992 6883 224995
rect 6914 224992 6920 225004
rect 6871 224964 6920 224992
rect 6871 224961 6883 224964
rect 6825 224955 6883 224961
rect 6914 224952 6920 224964
rect 6972 224992 6978 225004
rect 8294 224992 8300 225004
rect 6972 224964 8300 224992
rect 6972 224952 6978 224964
rect 8294 224952 8300 224964
rect 8352 224952 8358 225004
rect 7006 224924 7012 224936
rect 6967 224896 7012 224924
rect 7006 224884 7012 224896
rect 7064 224884 7070 224936
rect 7469 224791 7527 224797
rect 7469 224757 7481 224791
rect 7515 224788 7527 224791
rect 8018 224788 8024 224800
rect 7515 224760 8024 224788
rect 7515 224757 7527 224760
rect 7469 224751 7527 224757
rect 8018 224748 8024 224760
rect 8076 224748 8082 224800
rect 1104 224698 8832 224720
rect 1104 224646 4315 224698
rect 4367 224646 4379 224698
rect 4431 224646 4443 224698
rect 4495 224646 4507 224698
rect 4559 224646 7648 224698
rect 7700 224646 7712 224698
rect 7764 224646 7776 224698
rect 7828 224646 7840 224698
rect 7892 224646 8832 224698
rect 1104 224624 8832 224646
rect 1762 224544 1768 224596
rect 1820 224584 1826 224596
rect 2498 224584 2504 224596
rect 1820 224556 2504 224584
rect 1820 224544 1826 224556
rect 2498 224544 2504 224556
rect 2556 224584 2562 224596
rect 2593 224587 2651 224593
rect 2593 224584 2605 224587
rect 2556 224556 2605 224584
rect 2556 224544 2562 224556
rect 2593 224553 2605 224556
rect 2639 224553 2651 224587
rect 6914 224584 6920 224596
rect 6875 224556 6920 224584
rect 2593 224547 2651 224553
rect 6914 224544 6920 224556
rect 6972 224544 6978 224596
rect 7006 224544 7012 224596
rect 7064 224584 7070 224596
rect 7193 224587 7251 224593
rect 7193 224584 7205 224587
rect 7064 224556 7205 224584
rect 7064 224544 7070 224556
rect 7193 224553 7205 224556
rect 7239 224553 7251 224587
rect 7193 224547 7251 224553
rect 5442 224408 5448 224460
rect 5500 224448 5506 224460
rect 5810 224448 5816 224460
rect 5500 224420 5816 224448
rect 5500 224408 5506 224420
rect 5810 224408 5816 224420
rect 5868 224408 5874 224460
rect 5350 224340 5356 224392
rect 5408 224380 5414 224392
rect 5997 224383 6055 224389
rect 5997 224380 6009 224383
rect 5408 224352 6009 224380
rect 5408 224340 5414 224352
rect 5997 224349 6009 224352
rect 6043 224380 6055 224383
rect 6270 224380 6276 224392
rect 6043 224352 6276 224380
rect 6043 224349 6055 224352
rect 5997 224343 6055 224349
rect 6270 224340 6276 224352
rect 6328 224340 6334 224392
rect 6457 224247 6515 224253
rect 6457 224213 6469 224247
rect 6503 224244 6515 224247
rect 6546 224244 6552 224256
rect 6503 224216 6552 224244
rect 6503 224213 6515 224216
rect 6457 224207 6515 224213
rect 6546 224204 6552 224216
rect 6604 224204 6610 224256
rect 1104 224154 8832 224176
rect 1104 224102 2648 224154
rect 2700 224102 2712 224154
rect 2764 224102 2776 224154
rect 2828 224102 2840 224154
rect 2892 224102 5982 224154
rect 6034 224102 6046 224154
rect 6098 224102 6110 224154
rect 6162 224102 6174 224154
rect 6226 224102 8832 224154
rect 1104 224080 8832 224102
rect 2314 224000 2320 224052
rect 2372 224040 2378 224052
rect 2409 224043 2467 224049
rect 2409 224040 2421 224043
rect 2372 224012 2421 224040
rect 2372 224000 2378 224012
rect 2409 224009 2421 224012
rect 2455 224009 2467 224043
rect 5810 224040 5816 224052
rect 5771 224012 5816 224040
rect 2409 224003 2467 224009
rect 2424 223904 2452 224003
rect 5810 224000 5816 224012
rect 5868 224000 5874 224052
rect 6270 224040 6276 224052
rect 6231 224012 6276 224040
rect 6270 224000 6276 224012
rect 6328 224000 6334 224052
rect 2958 223904 2964 223916
rect 2424 223876 2964 223904
rect 2958 223864 2964 223876
rect 3016 223904 3022 223916
rect 3016 223876 3832 223904
rect 3016 223864 3022 223876
rect 2498 223796 2504 223848
rect 2556 223836 2562 223848
rect 2593 223839 2651 223845
rect 2593 223836 2605 223839
rect 2556 223808 2605 223836
rect 2556 223796 2562 223808
rect 2593 223805 2605 223808
rect 2639 223805 2651 223839
rect 3234 223836 3240 223848
rect 3195 223808 3240 223836
rect 2593 223799 2651 223805
rect 3234 223796 3240 223808
rect 3292 223796 3298 223848
rect 3418 223836 3424 223848
rect 3379 223808 3424 223836
rect 3418 223796 3424 223808
rect 3476 223796 3482 223848
rect 3804 223845 3832 223876
rect 3789 223839 3847 223845
rect 3789 223805 3801 223839
rect 3835 223805 3847 223839
rect 3789 223799 3847 223805
rect 2133 223771 2191 223777
rect 2133 223737 2145 223771
rect 2179 223768 2191 223771
rect 3050 223768 3056 223780
rect 2179 223740 3056 223768
rect 2179 223737 2191 223740
rect 2133 223731 2191 223737
rect 3050 223728 3056 223740
rect 3108 223768 3114 223780
rect 3252 223768 3280 223796
rect 3108 223740 3280 223768
rect 3108 223728 3114 223740
rect 2869 223703 2927 223709
rect 2869 223669 2881 223703
rect 2915 223700 2927 223703
rect 3142 223700 3148 223712
rect 2915 223672 3148 223700
rect 2915 223669 2927 223672
rect 2869 223663 2927 223669
rect 3142 223660 3148 223672
rect 3200 223660 3206 223712
rect 1104 223610 8832 223632
rect 1104 223558 4315 223610
rect 4367 223558 4379 223610
rect 4431 223558 4443 223610
rect 4495 223558 4507 223610
rect 4559 223558 7648 223610
rect 7700 223558 7712 223610
rect 7764 223558 7776 223610
rect 7828 223558 7840 223610
rect 7892 223558 8832 223610
rect 1104 223536 8832 223558
rect 2685 223499 2743 223505
rect 2685 223465 2697 223499
rect 2731 223496 2743 223499
rect 3050 223496 3056 223508
rect 2731 223468 3056 223496
rect 2731 223465 2743 223468
rect 2685 223459 2743 223465
rect 3050 223456 3056 223468
rect 3108 223496 3114 223508
rect 3418 223496 3424 223508
rect 3108 223468 3424 223496
rect 3108 223456 3114 223468
rect 3418 223456 3424 223468
rect 3476 223456 3482 223508
rect 1104 223066 8832 223088
rect 1104 223014 2648 223066
rect 2700 223014 2712 223066
rect 2764 223014 2776 223066
rect 2828 223014 2840 223066
rect 2892 223014 5982 223066
rect 6034 223014 6046 223066
rect 6098 223014 6110 223066
rect 6162 223014 6174 223066
rect 6226 223014 8832 223066
rect 1104 222992 8832 223014
rect 1104 222522 8832 222544
rect 1104 222470 4315 222522
rect 4367 222470 4379 222522
rect 4431 222470 4443 222522
rect 4495 222470 4507 222522
rect 4559 222470 7648 222522
rect 7700 222470 7712 222522
rect 7764 222470 7776 222522
rect 7828 222470 7840 222522
rect 7892 222470 8832 222522
rect 1104 222448 8832 222470
rect 3050 222408 3056 222420
rect 3011 222380 3056 222408
rect 3050 222368 3056 222380
rect 3108 222368 3114 222420
rect 1104 221978 8832 222000
rect 1104 221926 2648 221978
rect 2700 221926 2712 221978
rect 2764 221926 2776 221978
rect 2828 221926 2840 221978
rect 2892 221926 5982 221978
rect 6034 221926 6046 221978
rect 6098 221926 6110 221978
rect 6162 221926 6174 221978
rect 6226 221926 8832 221978
rect 1104 221904 8832 221926
rect 2498 221864 2504 221876
rect 2459 221836 2504 221864
rect 2498 221824 2504 221836
rect 2556 221824 2562 221876
rect 2869 221867 2927 221873
rect 2869 221833 2881 221867
rect 2915 221864 2927 221867
rect 2958 221864 2964 221876
rect 2915 221836 2964 221864
rect 2915 221833 2927 221836
rect 2869 221827 2927 221833
rect 2958 221824 2964 221836
rect 3016 221824 3022 221876
rect 3234 221756 3240 221808
rect 3292 221796 3298 221808
rect 3292 221768 4154 221796
rect 3292 221756 3298 221768
rect 2961 221731 3019 221737
rect 2961 221697 2973 221731
rect 3007 221728 3019 221731
rect 3050 221728 3056 221740
rect 3007 221700 3056 221728
rect 3007 221697 3019 221700
rect 2961 221691 3019 221697
rect 3050 221688 3056 221700
rect 3108 221688 3114 221740
rect 4126 221728 4154 221768
rect 4525 221731 4583 221737
rect 4525 221728 4537 221731
rect 4126 221700 4537 221728
rect 4525 221697 4537 221700
rect 4571 221697 4583 221731
rect 4525 221691 4583 221697
rect 2498 221620 2504 221672
rect 2556 221660 2562 221672
rect 3237 221663 3295 221669
rect 3237 221660 3249 221663
rect 2556 221632 3249 221660
rect 2556 221620 2562 221632
rect 3237 221629 3249 221632
rect 3283 221629 3295 221663
rect 4433 221663 4491 221669
rect 4433 221660 4445 221663
rect 3237 221623 3295 221629
rect 4126 221632 4445 221660
rect 2958 221552 2964 221604
rect 3016 221592 3022 221604
rect 3145 221595 3203 221601
rect 3145 221592 3157 221595
rect 3016 221564 3157 221592
rect 3016 221552 3022 221564
rect 3145 221561 3157 221564
rect 3191 221561 3203 221595
rect 3326 221592 3332 221604
rect 3287 221564 3332 221592
rect 3145 221555 3203 221561
rect 3326 221552 3332 221564
rect 3384 221552 3390 221604
rect 3694 221592 3700 221604
rect 3655 221564 3700 221592
rect 3694 221552 3700 221564
rect 3752 221552 3758 221604
rect 3344 221524 3372 221552
rect 4126 221524 4154 221632
rect 4433 221629 4445 221632
rect 4479 221660 4491 221663
rect 4617 221663 4675 221669
rect 4617 221660 4629 221663
rect 4479 221632 4629 221660
rect 4479 221629 4491 221632
rect 4433 221623 4491 221629
rect 4617 221629 4629 221632
rect 4663 221629 4675 221663
rect 4617 221623 4675 221629
rect 3344 221496 4154 221524
rect 1104 221434 8832 221456
rect 1104 221382 4315 221434
rect 4367 221382 4379 221434
rect 4431 221382 4443 221434
rect 4495 221382 4507 221434
rect 4559 221382 7648 221434
rect 7700 221382 7712 221434
rect 7764 221382 7776 221434
rect 7828 221382 7840 221434
rect 7892 221382 8832 221434
rect 1104 221360 8832 221382
rect 1394 220940 1400 220992
rect 1452 220980 1458 220992
rect 2961 220983 3019 220989
rect 2961 220980 2973 220983
rect 1452 220952 2973 220980
rect 1452 220940 1458 220952
rect 2961 220949 2973 220952
rect 3007 220980 3019 220983
rect 3326 220980 3332 220992
rect 3007 220952 3332 220980
rect 3007 220949 3019 220952
rect 2961 220943 3019 220949
rect 3326 220940 3332 220952
rect 3384 220940 3390 220992
rect 1104 220890 8832 220912
rect 1104 220838 2648 220890
rect 2700 220838 2712 220890
rect 2764 220838 2776 220890
rect 2828 220838 2840 220890
rect 2892 220838 5982 220890
rect 6034 220838 6046 220890
rect 6098 220838 6110 220890
rect 6162 220838 6174 220890
rect 6226 220838 8832 220890
rect 1104 220816 8832 220838
rect 1104 220346 8832 220368
rect 1104 220294 4315 220346
rect 4367 220294 4379 220346
rect 4431 220294 4443 220346
rect 4495 220294 4507 220346
rect 4559 220294 7648 220346
rect 7700 220294 7712 220346
rect 7764 220294 7776 220346
rect 7828 220294 7840 220346
rect 7892 220294 8832 220346
rect 1104 220272 8832 220294
rect 1104 219802 8832 219824
rect 1104 219750 2648 219802
rect 2700 219750 2712 219802
rect 2764 219750 2776 219802
rect 2828 219750 2840 219802
rect 2892 219750 5982 219802
rect 6034 219750 6046 219802
rect 6098 219750 6110 219802
rect 6162 219750 6174 219802
rect 6226 219750 8832 219802
rect 1104 219728 8832 219750
rect 1104 219258 8832 219280
rect 1104 219206 4315 219258
rect 4367 219206 4379 219258
rect 4431 219206 4443 219258
rect 4495 219206 4507 219258
rect 4559 219206 7648 219258
rect 7700 219206 7712 219258
rect 7764 219206 7776 219258
rect 7828 219206 7840 219258
rect 7892 219206 8832 219258
rect 1104 219184 8832 219206
rect 1104 218714 8832 218736
rect 1104 218662 2648 218714
rect 2700 218662 2712 218714
rect 2764 218662 2776 218714
rect 2828 218662 2840 218714
rect 2892 218662 5982 218714
rect 6034 218662 6046 218714
rect 6098 218662 6110 218714
rect 6162 218662 6174 218714
rect 6226 218662 8832 218714
rect 1104 218640 8832 218662
rect 1104 218170 8832 218192
rect 1104 218118 4315 218170
rect 4367 218118 4379 218170
rect 4431 218118 4443 218170
rect 4495 218118 4507 218170
rect 4559 218118 7648 218170
rect 7700 218118 7712 218170
rect 7764 218118 7776 218170
rect 7828 218118 7840 218170
rect 7892 218118 8832 218170
rect 1104 218096 8832 218118
rect 1104 217626 8832 217648
rect 1104 217574 2648 217626
rect 2700 217574 2712 217626
rect 2764 217574 2776 217626
rect 2828 217574 2840 217626
rect 2892 217574 5982 217626
rect 6034 217574 6046 217626
rect 6098 217574 6110 217626
rect 6162 217574 6174 217626
rect 6226 217574 8832 217626
rect 1104 217552 8832 217574
rect 1104 217082 8832 217104
rect 1104 217030 4315 217082
rect 4367 217030 4379 217082
rect 4431 217030 4443 217082
rect 4495 217030 4507 217082
rect 4559 217030 7648 217082
rect 7700 217030 7712 217082
rect 7764 217030 7776 217082
rect 7828 217030 7840 217082
rect 7892 217030 8832 217082
rect 1104 217008 8832 217030
rect 1104 216538 8832 216560
rect 1104 216486 2648 216538
rect 2700 216486 2712 216538
rect 2764 216486 2776 216538
rect 2828 216486 2840 216538
rect 2892 216486 5982 216538
rect 6034 216486 6046 216538
rect 6098 216486 6110 216538
rect 6162 216486 6174 216538
rect 6226 216486 8832 216538
rect 1104 216464 8832 216486
rect 1104 215994 8832 216016
rect 1104 215942 4315 215994
rect 4367 215942 4379 215994
rect 4431 215942 4443 215994
rect 4495 215942 4507 215994
rect 4559 215942 7648 215994
rect 7700 215942 7712 215994
rect 7764 215942 7776 215994
rect 7828 215942 7840 215994
rect 7892 215942 8832 215994
rect 1104 215920 8832 215942
rect 1104 215450 8832 215472
rect 1104 215398 2648 215450
rect 2700 215398 2712 215450
rect 2764 215398 2776 215450
rect 2828 215398 2840 215450
rect 2892 215398 5982 215450
rect 6034 215398 6046 215450
rect 6098 215398 6110 215450
rect 6162 215398 6174 215450
rect 6226 215398 8832 215450
rect 1104 215376 8832 215398
rect 3605 215203 3663 215209
rect 3605 215169 3617 215203
rect 3651 215200 3663 215203
rect 3694 215200 3700 215212
rect 3651 215172 3700 215200
rect 3651 215169 3663 215172
rect 3605 215163 3663 215169
rect 3694 215160 3700 215172
rect 3752 215160 3758 215212
rect 3326 214956 3332 215008
rect 3384 214996 3390 215008
rect 3513 214999 3571 215005
rect 3513 214996 3525 214999
rect 3384 214968 3525 214996
rect 3384 214956 3390 214968
rect 3513 214965 3525 214968
rect 3559 214996 3571 214999
rect 3970 214996 3976 215008
rect 3559 214968 3976 214996
rect 3559 214965 3571 214968
rect 3513 214959 3571 214965
rect 3970 214956 3976 214968
rect 4028 214956 4034 215008
rect 4525 214999 4583 215005
rect 4525 214965 4537 214999
rect 4571 214996 4583 214999
rect 4614 214996 4620 215008
rect 4571 214968 4620 214996
rect 4571 214965 4583 214968
rect 4525 214959 4583 214965
rect 4614 214956 4620 214968
rect 4672 214956 4678 215008
rect 1104 214906 8832 214928
rect 1104 214854 4315 214906
rect 4367 214854 4379 214906
rect 4431 214854 4443 214906
rect 4495 214854 4507 214906
rect 4559 214854 7648 214906
rect 7700 214854 7712 214906
rect 7764 214854 7776 214906
rect 7828 214854 7840 214906
rect 7892 214854 8832 214906
rect 1104 214832 8832 214854
rect 3694 214792 3700 214804
rect 3655 214764 3700 214792
rect 3694 214752 3700 214764
rect 3752 214752 3758 214804
rect 1104 214362 8832 214384
rect 1104 214310 2648 214362
rect 2700 214310 2712 214362
rect 2764 214310 2776 214362
rect 2828 214310 2840 214362
rect 2892 214310 5982 214362
rect 6034 214310 6046 214362
rect 6098 214310 6110 214362
rect 6162 214310 6174 214362
rect 6226 214310 8832 214362
rect 1104 214288 8832 214310
rect 7282 214208 7288 214260
rect 7340 214248 7346 214260
rect 7653 214251 7711 214257
rect 7653 214248 7665 214251
rect 7340 214220 7665 214248
rect 7340 214208 7346 214220
rect 7653 214217 7665 214220
rect 7699 214217 7711 214251
rect 7653 214211 7711 214217
rect 6730 214004 6736 214056
rect 6788 214044 6794 214056
rect 7469 214047 7527 214053
rect 7469 214044 7481 214047
rect 6788 214016 7481 214044
rect 6788 214004 6794 214016
rect 7469 214013 7481 214016
rect 7515 214044 7527 214047
rect 8021 214047 8079 214053
rect 8021 214044 8033 214047
rect 7515 214016 8033 214044
rect 7515 214013 7527 214016
rect 7469 214007 7527 214013
rect 8021 214013 8033 214016
rect 8067 214013 8079 214047
rect 8021 214007 8079 214013
rect 1104 213818 8832 213840
rect 1104 213766 4315 213818
rect 4367 213766 4379 213818
rect 4431 213766 4443 213818
rect 4495 213766 4507 213818
rect 4559 213766 7648 213818
rect 7700 213766 7712 213818
rect 7764 213766 7776 213818
rect 7828 213766 7840 213818
rect 7892 213766 8832 213818
rect 1104 213744 8832 213766
rect 1104 213274 8832 213296
rect 1104 213222 2648 213274
rect 2700 213222 2712 213274
rect 2764 213222 2776 213274
rect 2828 213222 2840 213274
rect 2892 213222 5982 213274
rect 6034 213222 6046 213274
rect 6098 213222 6110 213274
rect 6162 213222 6174 213274
rect 6226 213222 8832 213274
rect 1104 213200 8832 213222
rect 1104 212730 8832 212752
rect 1104 212678 4315 212730
rect 4367 212678 4379 212730
rect 4431 212678 4443 212730
rect 4495 212678 4507 212730
rect 4559 212678 7648 212730
rect 7700 212678 7712 212730
rect 7764 212678 7776 212730
rect 7828 212678 7840 212730
rect 7892 212678 8832 212730
rect 1104 212656 8832 212678
rect 1104 212186 8832 212208
rect 1104 212134 2648 212186
rect 2700 212134 2712 212186
rect 2764 212134 2776 212186
rect 2828 212134 2840 212186
rect 2892 212134 5982 212186
rect 6034 212134 6046 212186
rect 6098 212134 6110 212186
rect 6162 212134 6174 212186
rect 6226 212134 8832 212186
rect 1104 212112 8832 212134
rect 106 212032 112 212084
rect 164 212072 170 212084
rect 4249 212075 4307 212081
rect 4249 212072 4261 212075
rect 164 212044 4261 212072
rect 164 212032 170 212044
rect 4249 212041 4261 212044
rect 4295 212072 4307 212075
rect 4295 212044 4476 212072
rect 4295 212041 4307 212044
rect 4249 212035 4307 212041
rect 4448 211945 4476 212044
rect 4433 211939 4491 211945
rect 4433 211905 4445 211939
rect 4479 211905 4491 211939
rect 4614 211936 4620 211948
rect 4575 211908 4620 211936
rect 4433 211899 4491 211905
rect 4614 211896 4620 211908
rect 4672 211896 4678 211948
rect 5077 211735 5135 211741
rect 5077 211701 5089 211735
rect 5123 211732 5135 211735
rect 6730 211732 6736 211744
rect 5123 211704 6736 211732
rect 5123 211701 5135 211704
rect 5077 211695 5135 211701
rect 6730 211692 6736 211704
rect 6788 211692 6794 211744
rect 1104 211642 8832 211664
rect 1104 211590 4315 211642
rect 4367 211590 4379 211642
rect 4431 211590 4443 211642
rect 4495 211590 4507 211642
rect 4559 211590 7648 211642
rect 7700 211590 7712 211642
rect 7764 211590 7776 211642
rect 7828 211590 7840 211642
rect 7892 211590 8832 211642
rect 1104 211568 8832 211590
rect 4525 211531 4583 211537
rect 4525 211497 4537 211531
rect 4571 211528 4583 211531
rect 4614 211528 4620 211540
rect 4571 211500 4620 211528
rect 4571 211497 4583 211500
rect 4525 211491 4583 211497
rect 4614 211488 4620 211500
rect 4672 211488 4678 211540
rect 1104 211098 8832 211120
rect 1104 211046 2648 211098
rect 2700 211046 2712 211098
rect 2764 211046 2776 211098
rect 2828 211046 2840 211098
rect 2892 211046 5982 211098
rect 6034 211046 6046 211098
rect 6098 211046 6110 211098
rect 6162 211046 6174 211098
rect 6226 211046 8832 211098
rect 1104 211024 8832 211046
rect 7006 210984 7012 210996
rect 6967 210956 7012 210984
rect 7006 210944 7012 210956
rect 7064 210944 7070 210996
rect 3878 210740 3884 210792
rect 3936 210780 3942 210792
rect 6825 210783 6883 210789
rect 6825 210780 6837 210783
rect 3936 210752 6837 210780
rect 3936 210740 3942 210752
rect 6825 210749 6837 210752
rect 6871 210780 6883 210783
rect 7377 210783 7435 210789
rect 7377 210780 7389 210783
rect 6871 210752 7389 210780
rect 6871 210749 6883 210752
rect 6825 210743 6883 210749
rect 7377 210749 7389 210752
rect 7423 210749 7435 210783
rect 7377 210743 7435 210749
rect 1104 210554 8832 210576
rect 1104 210502 4315 210554
rect 4367 210502 4379 210554
rect 4431 210502 4443 210554
rect 4495 210502 4507 210554
rect 4559 210502 7648 210554
rect 7700 210502 7712 210554
rect 7764 210502 7776 210554
rect 7828 210502 7840 210554
rect 7892 210502 8832 210554
rect 1104 210480 8832 210502
rect 1104 210010 8832 210032
rect 1104 209958 2648 210010
rect 2700 209958 2712 210010
rect 2764 209958 2776 210010
rect 2828 209958 2840 210010
rect 2892 209958 5982 210010
rect 6034 209958 6046 210010
rect 6098 209958 6110 210010
rect 6162 209958 6174 210010
rect 6226 209958 8832 210010
rect 1104 209936 8832 209958
rect 3329 209899 3387 209905
rect 3329 209865 3341 209899
rect 3375 209896 3387 209899
rect 3878 209896 3884 209908
rect 3375 209868 3884 209896
rect 3375 209865 3387 209868
rect 3329 209859 3387 209865
rect 3878 209856 3884 209868
rect 3936 209856 3942 209908
rect 2685 209695 2743 209701
rect 2685 209692 2697 209695
rect 2516 209664 2697 209692
rect 14 209516 20 209568
rect 72 209556 78 209568
rect 2516 209565 2544 209664
rect 2685 209661 2697 209664
rect 2731 209661 2743 209695
rect 2685 209655 2743 209661
rect 2869 209695 2927 209701
rect 2869 209661 2881 209695
rect 2915 209692 2927 209695
rect 2958 209692 2964 209704
rect 2915 209664 2964 209692
rect 2915 209661 2927 209664
rect 2869 209655 2927 209661
rect 2958 209652 2964 209664
rect 3016 209652 3022 209704
rect 2501 209559 2559 209565
rect 2501 209556 2513 209559
rect 72 209528 2513 209556
rect 72 209516 78 209528
rect 2501 209525 2513 209528
rect 2547 209525 2559 209559
rect 2501 209519 2559 209525
rect 1104 209466 8832 209488
rect 1104 209414 4315 209466
rect 4367 209414 4379 209466
rect 4431 209414 4443 209466
rect 4495 209414 4507 209466
rect 4559 209414 7648 209466
rect 7700 209414 7712 209466
rect 7764 209414 7776 209466
rect 7828 209414 7840 209466
rect 7892 209414 8832 209466
rect 1104 209392 8832 209414
rect 2777 209015 2835 209021
rect 2777 208981 2789 209015
rect 2823 209012 2835 209015
rect 2958 209012 2964 209024
rect 2823 208984 2964 209012
rect 2823 208981 2835 208984
rect 2777 208975 2835 208981
rect 2958 208972 2964 208984
rect 3016 209012 3022 209024
rect 3694 209012 3700 209024
rect 3016 208984 3700 209012
rect 3016 208972 3022 208984
rect 3694 208972 3700 208984
rect 3752 208972 3758 209024
rect 1104 208922 8832 208944
rect 1104 208870 2648 208922
rect 2700 208870 2712 208922
rect 2764 208870 2776 208922
rect 2828 208870 2840 208922
rect 2892 208870 5982 208922
rect 6034 208870 6046 208922
rect 6098 208870 6110 208922
rect 6162 208870 6174 208922
rect 6226 208870 8832 208922
rect 1104 208848 8832 208870
rect 3694 208808 3700 208820
rect 3655 208780 3700 208808
rect 3694 208768 3700 208780
rect 3752 208768 3758 208820
rect 2777 208675 2835 208681
rect 2777 208641 2789 208675
rect 2823 208672 2835 208675
rect 3142 208672 3148 208684
rect 2823 208644 3148 208672
rect 2823 208641 2835 208644
rect 2777 208635 2835 208641
rect 3142 208632 3148 208644
rect 3200 208632 3206 208684
rect 2685 208539 2743 208545
rect 2685 208505 2697 208539
rect 2731 208536 2743 208539
rect 2958 208536 2964 208548
rect 2731 208508 2964 208536
rect 2731 208505 2743 208508
rect 2685 208499 2743 208505
rect 2958 208496 2964 208508
rect 3016 208536 3022 208548
rect 3139 208539 3197 208545
rect 3139 208536 3151 208539
rect 3016 208508 3151 208536
rect 3016 208496 3022 208508
rect 3139 208505 3151 208508
rect 3185 208536 3197 208539
rect 3326 208536 3332 208548
rect 3185 208508 3332 208536
rect 3185 208505 3197 208508
rect 3139 208499 3197 208505
rect 3326 208496 3332 208508
rect 3384 208496 3390 208548
rect 1104 208378 8832 208400
rect 1104 208326 4315 208378
rect 4367 208326 4379 208378
rect 4431 208326 4443 208378
rect 4495 208326 4507 208378
rect 4559 208326 7648 208378
rect 7700 208326 7712 208378
rect 7764 208326 7776 208378
rect 7828 208326 7840 208378
rect 7892 208326 8832 208378
rect 1104 208304 8832 208326
rect 2869 208267 2927 208273
rect 2869 208233 2881 208267
rect 2915 208264 2927 208267
rect 3142 208264 3148 208276
rect 2915 208236 3148 208264
rect 2915 208233 2927 208236
rect 2869 208227 2927 208233
rect 3142 208224 3148 208236
rect 3200 208224 3206 208276
rect 1104 207834 8832 207856
rect 1104 207782 2648 207834
rect 2700 207782 2712 207834
rect 2764 207782 2776 207834
rect 2828 207782 2840 207834
rect 2892 207782 5982 207834
rect 6034 207782 6046 207834
rect 6098 207782 6110 207834
rect 6162 207782 6174 207834
rect 6226 207782 8832 207834
rect 1104 207760 8832 207782
rect 1104 207290 8832 207312
rect 1104 207238 4315 207290
rect 4367 207238 4379 207290
rect 4431 207238 4443 207290
rect 4495 207238 4507 207290
rect 4559 207238 7648 207290
rect 7700 207238 7712 207290
rect 7764 207238 7776 207290
rect 7828 207238 7840 207290
rect 7892 207238 8832 207290
rect 1104 207216 8832 207238
rect 1104 206746 8832 206768
rect 1104 206694 2648 206746
rect 2700 206694 2712 206746
rect 2764 206694 2776 206746
rect 2828 206694 2840 206746
rect 2892 206694 5982 206746
rect 6034 206694 6046 206746
rect 6098 206694 6110 206746
rect 6162 206694 6174 206746
rect 6226 206694 8832 206746
rect 1104 206672 8832 206694
rect 1104 206202 8832 206224
rect 1104 206150 4315 206202
rect 4367 206150 4379 206202
rect 4431 206150 4443 206202
rect 4495 206150 4507 206202
rect 4559 206150 7648 206202
rect 7700 206150 7712 206202
rect 7764 206150 7776 206202
rect 7828 206150 7840 206202
rect 7892 206150 8832 206202
rect 1104 206128 8832 206150
rect 1104 205658 8832 205680
rect 1104 205606 2648 205658
rect 2700 205606 2712 205658
rect 2764 205606 2776 205658
rect 2828 205606 2840 205658
rect 2892 205606 5982 205658
rect 6034 205606 6046 205658
rect 6098 205606 6110 205658
rect 6162 205606 6174 205658
rect 6226 205606 8832 205658
rect 1104 205584 8832 205606
rect 1104 205114 8832 205136
rect 1104 205062 4315 205114
rect 4367 205062 4379 205114
rect 4431 205062 4443 205114
rect 4495 205062 4507 205114
rect 4559 205062 7648 205114
rect 7700 205062 7712 205114
rect 7764 205062 7776 205114
rect 7828 205062 7840 205114
rect 7892 205062 8832 205114
rect 1104 205040 8832 205062
rect 1104 204570 8832 204592
rect 1104 204518 2648 204570
rect 2700 204518 2712 204570
rect 2764 204518 2776 204570
rect 2828 204518 2840 204570
rect 2892 204518 5982 204570
rect 6034 204518 6046 204570
rect 6098 204518 6110 204570
rect 6162 204518 6174 204570
rect 6226 204518 8832 204570
rect 1104 204496 8832 204518
rect 1104 204026 8832 204048
rect 1104 203974 4315 204026
rect 4367 203974 4379 204026
rect 4431 203974 4443 204026
rect 4495 203974 4507 204026
rect 4559 203974 7648 204026
rect 7700 203974 7712 204026
rect 7764 203974 7776 204026
rect 7828 203974 7840 204026
rect 7892 203974 8832 204026
rect 1104 203952 8832 203974
rect 1104 203482 8832 203504
rect 1104 203430 2648 203482
rect 2700 203430 2712 203482
rect 2764 203430 2776 203482
rect 2828 203430 2840 203482
rect 2892 203430 5982 203482
rect 6034 203430 6046 203482
rect 6098 203430 6110 203482
rect 6162 203430 6174 203482
rect 6226 203430 8832 203482
rect 1104 203408 8832 203430
rect 1104 202938 8832 202960
rect 1104 202886 4315 202938
rect 4367 202886 4379 202938
rect 4431 202886 4443 202938
rect 4495 202886 4507 202938
rect 4559 202886 7648 202938
rect 7700 202886 7712 202938
rect 7764 202886 7776 202938
rect 7828 202886 7840 202938
rect 7892 202886 8832 202938
rect 1104 202864 8832 202886
rect 1104 202394 8832 202416
rect 1104 202342 2648 202394
rect 2700 202342 2712 202394
rect 2764 202342 2776 202394
rect 2828 202342 2840 202394
rect 2892 202342 5982 202394
rect 6034 202342 6046 202394
rect 6098 202342 6110 202394
rect 6162 202342 6174 202394
rect 6226 202342 8832 202394
rect 1104 202320 8832 202342
rect 1104 201850 8832 201872
rect 1104 201798 4315 201850
rect 4367 201798 4379 201850
rect 4431 201798 4443 201850
rect 4495 201798 4507 201850
rect 4559 201798 7648 201850
rect 7700 201798 7712 201850
rect 7764 201798 7776 201850
rect 7828 201798 7840 201850
rect 7892 201798 8832 201850
rect 1104 201776 8832 201798
rect 1104 201306 8832 201328
rect 1104 201254 2648 201306
rect 2700 201254 2712 201306
rect 2764 201254 2776 201306
rect 2828 201254 2840 201306
rect 2892 201254 5982 201306
rect 6034 201254 6046 201306
rect 6098 201254 6110 201306
rect 6162 201254 6174 201306
rect 6226 201254 8832 201306
rect 1104 201232 8832 201254
rect 1104 200762 8832 200784
rect 1104 200710 4315 200762
rect 4367 200710 4379 200762
rect 4431 200710 4443 200762
rect 4495 200710 4507 200762
rect 4559 200710 7648 200762
rect 7700 200710 7712 200762
rect 7764 200710 7776 200762
rect 7828 200710 7840 200762
rect 7892 200710 8832 200762
rect 1104 200688 8832 200710
rect 1104 200218 8832 200240
rect 1104 200166 2648 200218
rect 2700 200166 2712 200218
rect 2764 200166 2776 200218
rect 2828 200166 2840 200218
rect 2892 200166 5982 200218
rect 6034 200166 6046 200218
rect 6098 200166 6110 200218
rect 6162 200166 6174 200218
rect 6226 200166 8832 200218
rect 1104 200144 8832 200166
rect 1104 199674 8832 199696
rect 1104 199622 4315 199674
rect 4367 199622 4379 199674
rect 4431 199622 4443 199674
rect 4495 199622 4507 199674
rect 4559 199622 7648 199674
rect 7700 199622 7712 199674
rect 7764 199622 7776 199674
rect 7828 199622 7840 199674
rect 7892 199622 8832 199674
rect 1104 199600 8832 199622
rect 1104 199130 8832 199152
rect 1104 199078 2648 199130
rect 2700 199078 2712 199130
rect 2764 199078 2776 199130
rect 2828 199078 2840 199130
rect 2892 199078 5982 199130
rect 6034 199078 6046 199130
rect 6098 199078 6110 199130
rect 6162 199078 6174 199130
rect 6226 199078 8832 199130
rect 1104 199056 8832 199078
rect 1104 198586 8832 198608
rect 1104 198534 4315 198586
rect 4367 198534 4379 198586
rect 4431 198534 4443 198586
rect 4495 198534 4507 198586
rect 4559 198534 7648 198586
rect 7700 198534 7712 198586
rect 7764 198534 7776 198586
rect 7828 198534 7840 198586
rect 7892 198534 8832 198586
rect 1104 198512 8832 198534
rect 1104 198042 8832 198064
rect 1104 197990 2648 198042
rect 2700 197990 2712 198042
rect 2764 197990 2776 198042
rect 2828 197990 2840 198042
rect 2892 197990 5982 198042
rect 6034 197990 6046 198042
rect 6098 197990 6110 198042
rect 6162 197990 6174 198042
rect 6226 197990 8832 198042
rect 1104 197968 8832 197990
rect 1104 197498 8832 197520
rect 1104 197446 4315 197498
rect 4367 197446 4379 197498
rect 4431 197446 4443 197498
rect 4495 197446 4507 197498
rect 4559 197446 7648 197498
rect 7700 197446 7712 197498
rect 7764 197446 7776 197498
rect 7828 197446 7840 197498
rect 7892 197446 8832 197498
rect 1104 197424 8832 197446
rect 1104 196954 8832 196976
rect 1104 196902 2648 196954
rect 2700 196902 2712 196954
rect 2764 196902 2776 196954
rect 2828 196902 2840 196954
rect 2892 196902 5982 196954
rect 6034 196902 6046 196954
rect 6098 196902 6110 196954
rect 6162 196902 6174 196954
rect 6226 196902 8832 196954
rect 1104 196880 8832 196902
rect 1104 196410 8832 196432
rect 1104 196358 4315 196410
rect 4367 196358 4379 196410
rect 4431 196358 4443 196410
rect 4495 196358 4507 196410
rect 4559 196358 7648 196410
rect 7700 196358 7712 196410
rect 7764 196358 7776 196410
rect 7828 196358 7840 196410
rect 7892 196358 8832 196410
rect 1104 196336 8832 196358
rect 1104 195866 8832 195888
rect 1104 195814 2648 195866
rect 2700 195814 2712 195866
rect 2764 195814 2776 195866
rect 2828 195814 2840 195866
rect 2892 195814 5982 195866
rect 6034 195814 6046 195866
rect 6098 195814 6110 195866
rect 6162 195814 6174 195866
rect 6226 195814 8832 195866
rect 1104 195792 8832 195814
rect 1104 195322 8832 195344
rect 1104 195270 4315 195322
rect 4367 195270 4379 195322
rect 4431 195270 4443 195322
rect 4495 195270 4507 195322
rect 4559 195270 7648 195322
rect 7700 195270 7712 195322
rect 7764 195270 7776 195322
rect 7828 195270 7840 195322
rect 7892 195270 8832 195322
rect 1104 195248 8832 195270
rect 1104 194778 8832 194800
rect 1104 194726 2648 194778
rect 2700 194726 2712 194778
rect 2764 194726 2776 194778
rect 2828 194726 2840 194778
rect 2892 194726 5982 194778
rect 6034 194726 6046 194778
rect 6098 194726 6110 194778
rect 6162 194726 6174 194778
rect 6226 194726 8832 194778
rect 1104 194704 8832 194726
rect 1104 194234 8832 194256
rect 1104 194182 4315 194234
rect 4367 194182 4379 194234
rect 4431 194182 4443 194234
rect 4495 194182 4507 194234
rect 4559 194182 7648 194234
rect 7700 194182 7712 194234
rect 7764 194182 7776 194234
rect 7828 194182 7840 194234
rect 7892 194182 8832 194234
rect 1104 194160 8832 194182
rect 1104 193690 8832 193712
rect 1104 193638 2648 193690
rect 2700 193638 2712 193690
rect 2764 193638 2776 193690
rect 2828 193638 2840 193690
rect 2892 193638 5982 193690
rect 6034 193638 6046 193690
rect 6098 193638 6110 193690
rect 6162 193638 6174 193690
rect 6226 193638 8832 193690
rect 1104 193616 8832 193638
rect 1104 193146 8832 193168
rect 1104 193094 4315 193146
rect 4367 193094 4379 193146
rect 4431 193094 4443 193146
rect 4495 193094 4507 193146
rect 4559 193094 7648 193146
rect 7700 193094 7712 193146
rect 7764 193094 7776 193146
rect 7828 193094 7840 193146
rect 7892 193094 8832 193146
rect 1104 193072 8832 193094
rect 1104 192602 8832 192624
rect 1104 192550 2648 192602
rect 2700 192550 2712 192602
rect 2764 192550 2776 192602
rect 2828 192550 2840 192602
rect 2892 192550 5982 192602
rect 6034 192550 6046 192602
rect 6098 192550 6110 192602
rect 6162 192550 6174 192602
rect 6226 192550 8832 192602
rect 1104 192528 8832 192550
rect 1104 192058 8832 192080
rect 1104 192006 4315 192058
rect 4367 192006 4379 192058
rect 4431 192006 4443 192058
rect 4495 192006 4507 192058
rect 4559 192006 7648 192058
rect 7700 192006 7712 192058
rect 7764 192006 7776 192058
rect 7828 192006 7840 192058
rect 7892 192006 8832 192058
rect 1104 191984 8832 192006
rect 1104 191514 8832 191536
rect 1104 191462 2648 191514
rect 2700 191462 2712 191514
rect 2764 191462 2776 191514
rect 2828 191462 2840 191514
rect 2892 191462 5982 191514
rect 6034 191462 6046 191514
rect 6098 191462 6110 191514
rect 6162 191462 6174 191514
rect 6226 191462 8832 191514
rect 1104 191440 8832 191462
rect 1104 190970 8832 190992
rect 1104 190918 4315 190970
rect 4367 190918 4379 190970
rect 4431 190918 4443 190970
rect 4495 190918 4507 190970
rect 4559 190918 7648 190970
rect 7700 190918 7712 190970
rect 7764 190918 7776 190970
rect 7828 190918 7840 190970
rect 7892 190918 8832 190970
rect 1104 190896 8832 190918
rect 1104 190426 8832 190448
rect 1104 190374 2648 190426
rect 2700 190374 2712 190426
rect 2764 190374 2776 190426
rect 2828 190374 2840 190426
rect 2892 190374 5982 190426
rect 6034 190374 6046 190426
rect 6098 190374 6110 190426
rect 6162 190374 6174 190426
rect 6226 190374 8832 190426
rect 1104 190352 8832 190374
rect 1104 189882 8832 189904
rect 1104 189830 4315 189882
rect 4367 189830 4379 189882
rect 4431 189830 4443 189882
rect 4495 189830 4507 189882
rect 4559 189830 7648 189882
rect 7700 189830 7712 189882
rect 7764 189830 7776 189882
rect 7828 189830 7840 189882
rect 7892 189830 8832 189882
rect 1104 189808 8832 189830
rect 1104 189338 8832 189360
rect 1104 189286 2648 189338
rect 2700 189286 2712 189338
rect 2764 189286 2776 189338
rect 2828 189286 2840 189338
rect 2892 189286 5982 189338
rect 6034 189286 6046 189338
rect 6098 189286 6110 189338
rect 6162 189286 6174 189338
rect 6226 189286 8832 189338
rect 1104 189264 8832 189286
rect 1104 188794 8832 188816
rect 1104 188742 4315 188794
rect 4367 188742 4379 188794
rect 4431 188742 4443 188794
rect 4495 188742 4507 188794
rect 4559 188742 7648 188794
rect 7700 188742 7712 188794
rect 7764 188742 7776 188794
rect 7828 188742 7840 188794
rect 7892 188742 8832 188794
rect 1104 188720 8832 188742
rect 1104 188250 8832 188272
rect 1104 188198 2648 188250
rect 2700 188198 2712 188250
rect 2764 188198 2776 188250
rect 2828 188198 2840 188250
rect 2892 188198 5982 188250
rect 6034 188198 6046 188250
rect 6098 188198 6110 188250
rect 6162 188198 6174 188250
rect 6226 188198 8832 188250
rect 1104 188176 8832 188198
rect 1104 187706 8832 187728
rect 1104 187654 4315 187706
rect 4367 187654 4379 187706
rect 4431 187654 4443 187706
rect 4495 187654 4507 187706
rect 4559 187654 7648 187706
rect 7700 187654 7712 187706
rect 7764 187654 7776 187706
rect 7828 187654 7840 187706
rect 7892 187654 8832 187706
rect 1104 187632 8832 187654
rect 1104 187162 8832 187184
rect 1104 187110 2648 187162
rect 2700 187110 2712 187162
rect 2764 187110 2776 187162
rect 2828 187110 2840 187162
rect 2892 187110 5982 187162
rect 6034 187110 6046 187162
rect 6098 187110 6110 187162
rect 6162 187110 6174 187162
rect 6226 187110 8832 187162
rect 1104 187088 8832 187110
rect 1104 186618 8832 186640
rect 1104 186566 4315 186618
rect 4367 186566 4379 186618
rect 4431 186566 4443 186618
rect 4495 186566 4507 186618
rect 4559 186566 7648 186618
rect 7700 186566 7712 186618
rect 7764 186566 7776 186618
rect 7828 186566 7840 186618
rect 7892 186566 8832 186618
rect 1104 186544 8832 186566
rect 1104 186074 8832 186096
rect 1104 186022 2648 186074
rect 2700 186022 2712 186074
rect 2764 186022 2776 186074
rect 2828 186022 2840 186074
rect 2892 186022 5982 186074
rect 6034 186022 6046 186074
rect 6098 186022 6110 186074
rect 6162 186022 6174 186074
rect 6226 186022 8832 186074
rect 1104 186000 8832 186022
rect 1104 185530 8832 185552
rect 1104 185478 4315 185530
rect 4367 185478 4379 185530
rect 4431 185478 4443 185530
rect 4495 185478 4507 185530
rect 4559 185478 7648 185530
rect 7700 185478 7712 185530
rect 7764 185478 7776 185530
rect 7828 185478 7840 185530
rect 7892 185478 8832 185530
rect 1104 185456 8832 185478
rect 1104 184986 8832 185008
rect 1104 184934 2648 184986
rect 2700 184934 2712 184986
rect 2764 184934 2776 184986
rect 2828 184934 2840 184986
rect 2892 184934 5982 184986
rect 6034 184934 6046 184986
rect 6098 184934 6110 184986
rect 6162 184934 6174 184986
rect 6226 184934 8832 184986
rect 1104 184912 8832 184934
rect 1104 184442 8832 184464
rect 1104 184390 4315 184442
rect 4367 184390 4379 184442
rect 4431 184390 4443 184442
rect 4495 184390 4507 184442
rect 4559 184390 7648 184442
rect 7700 184390 7712 184442
rect 7764 184390 7776 184442
rect 7828 184390 7840 184442
rect 7892 184390 8832 184442
rect 1104 184368 8832 184390
rect 1104 183898 8832 183920
rect 1104 183846 2648 183898
rect 2700 183846 2712 183898
rect 2764 183846 2776 183898
rect 2828 183846 2840 183898
rect 2892 183846 5982 183898
rect 6034 183846 6046 183898
rect 6098 183846 6110 183898
rect 6162 183846 6174 183898
rect 6226 183846 8832 183898
rect 1104 183824 8832 183846
rect 1104 183354 8832 183376
rect 1104 183302 4315 183354
rect 4367 183302 4379 183354
rect 4431 183302 4443 183354
rect 4495 183302 4507 183354
rect 4559 183302 7648 183354
rect 7700 183302 7712 183354
rect 7764 183302 7776 183354
rect 7828 183302 7840 183354
rect 7892 183302 8832 183354
rect 1104 183280 8832 183302
rect 1104 182810 8832 182832
rect 1104 182758 2648 182810
rect 2700 182758 2712 182810
rect 2764 182758 2776 182810
rect 2828 182758 2840 182810
rect 2892 182758 5982 182810
rect 6034 182758 6046 182810
rect 6098 182758 6110 182810
rect 6162 182758 6174 182810
rect 6226 182758 8832 182810
rect 1104 182736 8832 182758
rect 1104 182266 8832 182288
rect 1104 182214 4315 182266
rect 4367 182214 4379 182266
rect 4431 182214 4443 182266
rect 4495 182214 4507 182266
rect 4559 182214 7648 182266
rect 7700 182214 7712 182266
rect 7764 182214 7776 182266
rect 7828 182214 7840 182266
rect 7892 182214 8832 182266
rect 1104 182192 8832 182214
rect 1104 181722 8832 181744
rect 1104 181670 2648 181722
rect 2700 181670 2712 181722
rect 2764 181670 2776 181722
rect 2828 181670 2840 181722
rect 2892 181670 5982 181722
rect 6034 181670 6046 181722
rect 6098 181670 6110 181722
rect 6162 181670 6174 181722
rect 6226 181670 8832 181722
rect 1104 181648 8832 181670
rect 1104 181178 8832 181200
rect 1104 181126 4315 181178
rect 4367 181126 4379 181178
rect 4431 181126 4443 181178
rect 4495 181126 4507 181178
rect 4559 181126 7648 181178
rect 7700 181126 7712 181178
rect 7764 181126 7776 181178
rect 7828 181126 7840 181178
rect 7892 181126 8832 181178
rect 1104 181104 8832 181126
rect 1104 180634 8832 180656
rect 1104 180582 2648 180634
rect 2700 180582 2712 180634
rect 2764 180582 2776 180634
rect 2828 180582 2840 180634
rect 2892 180582 5982 180634
rect 6034 180582 6046 180634
rect 6098 180582 6110 180634
rect 6162 180582 6174 180634
rect 6226 180582 8832 180634
rect 1104 180560 8832 180582
rect 1104 180090 8832 180112
rect 1104 180038 4315 180090
rect 4367 180038 4379 180090
rect 4431 180038 4443 180090
rect 4495 180038 4507 180090
rect 4559 180038 7648 180090
rect 7700 180038 7712 180090
rect 7764 180038 7776 180090
rect 7828 180038 7840 180090
rect 7892 180038 8832 180090
rect 1104 180016 8832 180038
rect 1104 179546 8832 179568
rect 1104 179494 2648 179546
rect 2700 179494 2712 179546
rect 2764 179494 2776 179546
rect 2828 179494 2840 179546
rect 2892 179494 5982 179546
rect 6034 179494 6046 179546
rect 6098 179494 6110 179546
rect 6162 179494 6174 179546
rect 6226 179494 8832 179546
rect 1104 179472 8832 179494
rect 1104 179002 8832 179024
rect 1104 178950 4315 179002
rect 4367 178950 4379 179002
rect 4431 178950 4443 179002
rect 4495 178950 4507 179002
rect 4559 178950 7648 179002
rect 7700 178950 7712 179002
rect 7764 178950 7776 179002
rect 7828 178950 7840 179002
rect 7892 178950 8832 179002
rect 1104 178928 8832 178950
rect 1104 178458 8832 178480
rect 1104 178406 2648 178458
rect 2700 178406 2712 178458
rect 2764 178406 2776 178458
rect 2828 178406 2840 178458
rect 2892 178406 5982 178458
rect 6034 178406 6046 178458
rect 6098 178406 6110 178458
rect 6162 178406 6174 178458
rect 6226 178406 8832 178458
rect 1104 178384 8832 178406
rect 1104 177914 8832 177936
rect 1104 177862 4315 177914
rect 4367 177862 4379 177914
rect 4431 177862 4443 177914
rect 4495 177862 4507 177914
rect 4559 177862 7648 177914
rect 7700 177862 7712 177914
rect 7764 177862 7776 177914
rect 7828 177862 7840 177914
rect 7892 177862 8832 177914
rect 1104 177840 8832 177862
rect 1104 177370 8832 177392
rect 1104 177318 2648 177370
rect 2700 177318 2712 177370
rect 2764 177318 2776 177370
rect 2828 177318 2840 177370
rect 2892 177318 5982 177370
rect 6034 177318 6046 177370
rect 6098 177318 6110 177370
rect 6162 177318 6174 177370
rect 6226 177318 8832 177370
rect 1104 177296 8832 177318
rect 1104 176826 8832 176848
rect 1104 176774 4315 176826
rect 4367 176774 4379 176826
rect 4431 176774 4443 176826
rect 4495 176774 4507 176826
rect 4559 176774 7648 176826
rect 7700 176774 7712 176826
rect 7764 176774 7776 176826
rect 7828 176774 7840 176826
rect 7892 176774 8832 176826
rect 1104 176752 8832 176774
rect 1104 176282 8832 176304
rect 1104 176230 2648 176282
rect 2700 176230 2712 176282
rect 2764 176230 2776 176282
rect 2828 176230 2840 176282
rect 2892 176230 5982 176282
rect 6034 176230 6046 176282
rect 6098 176230 6110 176282
rect 6162 176230 6174 176282
rect 6226 176230 8832 176282
rect 1104 176208 8832 176230
rect 1104 175738 8832 175760
rect 1104 175686 4315 175738
rect 4367 175686 4379 175738
rect 4431 175686 4443 175738
rect 4495 175686 4507 175738
rect 4559 175686 7648 175738
rect 7700 175686 7712 175738
rect 7764 175686 7776 175738
rect 7828 175686 7840 175738
rect 7892 175686 8832 175738
rect 1104 175664 8832 175686
rect 1104 175194 8832 175216
rect 1104 175142 2648 175194
rect 2700 175142 2712 175194
rect 2764 175142 2776 175194
rect 2828 175142 2840 175194
rect 2892 175142 5982 175194
rect 6034 175142 6046 175194
rect 6098 175142 6110 175194
rect 6162 175142 6174 175194
rect 6226 175142 8832 175194
rect 1104 175120 8832 175142
rect 1104 174650 8832 174672
rect 1104 174598 4315 174650
rect 4367 174598 4379 174650
rect 4431 174598 4443 174650
rect 4495 174598 4507 174650
rect 4559 174598 7648 174650
rect 7700 174598 7712 174650
rect 7764 174598 7776 174650
rect 7828 174598 7840 174650
rect 7892 174598 8832 174650
rect 1104 174576 8832 174598
rect 1104 174106 8832 174128
rect 1104 174054 2648 174106
rect 2700 174054 2712 174106
rect 2764 174054 2776 174106
rect 2828 174054 2840 174106
rect 2892 174054 5982 174106
rect 6034 174054 6046 174106
rect 6098 174054 6110 174106
rect 6162 174054 6174 174106
rect 6226 174054 8832 174106
rect 1104 174032 8832 174054
rect 1104 173562 8832 173584
rect 1104 173510 4315 173562
rect 4367 173510 4379 173562
rect 4431 173510 4443 173562
rect 4495 173510 4507 173562
rect 4559 173510 7648 173562
rect 7700 173510 7712 173562
rect 7764 173510 7776 173562
rect 7828 173510 7840 173562
rect 7892 173510 8832 173562
rect 1104 173488 8832 173510
rect 1104 173018 8832 173040
rect 1104 172966 2648 173018
rect 2700 172966 2712 173018
rect 2764 172966 2776 173018
rect 2828 172966 2840 173018
rect 2892 172966 5982 173018
rect 6034 172966 6046 173018
rect 6098 172966 6110 173018
rect 6162 172966 6174 173018
rect 6226 172966 8832 173018
rect 1104 172944 8832 172966
rect 1104 172474 8832 172496
rect 1104 172422 4315 172474
rect 4367 172422 4379 172474
rect 4431 172422 4443 172474
rect 4495 172422 4507 172474
rect 4559 172422 7648 172474
rect 7700 172422 7712 172474
rect 7764 172422 7776 172474
rect 7828 172422 7840 172474
rect 7892 172422 8832 172474
rect 1104 172400 8832 172422
rect 6638 172320 6644 172372
rect 6696 172360 6702 172372
rect 7653 172363 7711 172369
rect 7653 172360 7665 172363
rect 6696 172332 7665 172360
rect 6696 172320 6702 172332
rect 7653 172329 7665 172332
rect 7699 172329 7711 172363
rect 7653 172323 7711 172329
rect 6546 172184 6552 172236
rect 6604 172224 6610 172236
rect 6822 172224 6828 172236
rect 6604 172196 6828 172224
rect 6604 172184 6610 172196
rect 6822 172184 6828 172196
rect 6880 172224 6886 172236
rect 7466 172224 7472 172236
rect 6880 172196 7472 172224
rect 6880 172184 6886 172196
rect 7466 172184 7472 172196
rect 7524 172184 7530 172236
rect 1104 171930 8832 171952
rect 1104 171878 2648 171930
rect 2700 171878 2712 171930
rect 2764 171878 2776 171930
rect 2828 171878 2840 171930
rect 2892 171878 5982 171930
rect 6034 171878 6046 171930
rect 6098 171878 6110 171930
rect 6162 171878 6174 171930
rect 6226 171878 8832 171930
rect 1104 171856 8832 171878
rect 7466 171816 7472 171828
rect 7427 171788 7472 171816
rect 7466 171776 7472 171788
rect 7524 171776 7530 171828
rect 1104 171386 8832 171408
rect 1104 171334 4315 171386
rect 4367 171334 4379 171386
rect 4431 171334 4443 171386
rect 4495 171334 4507 171386
rect 4559 171334 7648 171386
rect 7700 171334 7712 171386
rect 7764 171334 7776 171386
rect 7828 171334 7840 171386
rect 7892 171334 8832 171386
rect 1104 171312 8832 171334
rect 1104 170842 8832 170864
rect 1104 170790 2648 170842
rect 2700 170790 2712 170842
rect 2764 170790 2776 170842
rect 2828 170790 2840 170842
rect 2892 170790 5982 170842
rect 6034 170790 6046 170842
rect 6098 170790 6110 170842
rect 6162 170790 6174 170842
rect 6226 170790 8832 170842
rect 1104 170768 8832 170790
rect 1104 170298 8832 170320
rect 1104 170246 4315 170298
rect 4367 170246 4379 170298
rect 4431 170246 4443 170298
rect 4495 170246 4507 170298
rect 4559 170246 7648 170298
rect 7700 170246 7712 170298
rect 7764 170246 7776 170298
rect 7828 170246 7840 170298
rect 7892 170246 8832 170298
rect 1104 170224 8832 170246
rect 1104 169754 8832 169776
rect 1104 169702 2648 169754
rect 2700 169702 2712 169754
rect 2764 169702 2776 169754
rect 2828 169702 2840 169754
rect 2892 169702 5982 169754
rect 6034 169702 6046 169754
rect 6098 169702 6110 169754
rect 6162 169702 6174 169754
rect 6226 169702 8832 169754
rect 1104 169680 8832 169702
rect 1104 169210 8832 169232
rect 1104 169158 4315 169210
rect 4367 169158 4379 169210
rect 4431 169158 4443 169210
rect 4495 169158 4507 169210
rect 4559 169158 7648 169210
rect 7700 169158 7712 169210
rect 7764 169158 7776 169210
rect 7828 169158 7840 169210
rect 7892 169158 8832 169210
rect 1104 169136 8832 169158
rect 1104 168666 8832 168688
rect 1104 168614 2648 168666
rect 2700 168614 2712 168666
rect 2764 168614 2776 168666
rect 2828 168614 2840 168666
rect 2892 168614 5982 168666
rect 6034 168614 6046 168666
rect 6098 168614 6110 168666
rect 6162 168614 6174 168666
rect 6226 168614 8832 168666
rect 1104 168592 8832 168614
rect 1104 168122 8832 168144
rect 1104 168070 4315 168122
rect 4367 168070 4379 168122
rect 4431 168070 4443 168122
rect 4495 168070 4507 168122
rect 4559 168070 7648 168122
rect 7700 168070 7712 168122
rect 7764 168070 7776 168122
rect 7828 168070 7840 168122
rect 7892 168070 8832 168122
rect 1104 168048 8832 168070
rect 1104 167578 8832 167600
rect 1104 167526 2648 167578
rect 2700 167526 2712 167578
rect 2764 167526 2776 167578
rect 2828 167526 2840 167578
rect 2892 167526 5982 167578
rect 6034 167526 6046 167578
rect 6098 167526 6110 167578
rect 6162 167526 6174 167578
rect 6226 167526 8832 167578
rect 1104 167504 8832 167526
rect 1104 167034 8832 167056
rect 1104 166982 4315 167034
rect 4367 166982 4379 167034
rect 4431 166982 4443 167034
rect 4495 166982 4507 167034
rect 4559 166982 7648 167034
rect 7700 166982 7712 167034
rect 7764 166982 7776 167034
rect 7828 166982 7840 167034
rect 7892 166982 8832 167034
rect 1104 166960 8832 166982
rect 1104 166490 8832 166512
rect 1104 166438 2648 166490
rect 2700 166438 2712 166490
rect 2764 166438 2776 166490
rect 2828 166438 2840 166490
rect 2892 166438 5982 166490
rect 6034 166438 6046 166490
rect 6098 166438 6110 166490
rect 6162 166438 6174 166490
rect 6226 166438 8832 166490
rect 1104 166416 8832 166438
rect 1104 165946 8832 165968
rect 1104 165894 4315 165946
rect 4367 165894 4379 165946
rect 4431 165894 4443 165946
rect 4495 165894 4507 165946
rect 4559 165894 7648 165946
rect 7700 165894 7712 165946
rect 7764 165894 7776 165946
rect 7828 165894 7840 165946
rect 7892 165894 8832 165946
rect 1104 165872 8832 165894
rect 1104 165402 8832 165424
rect 1104 165350 2648 165402
rect 2700 165350 2712 165402
rect 2764 165350 2776 165402
rect 2828 165350 2840 165402
rect 2892 165350 5982 165402
rect 6034 165350 6046 165402
rect 6098 165350 6110 165402
rect 6162 165350 6174 165402
rect 6226 165350 8832 165402
rect 1104 165328 8832 165350
rect 1104 164858 8832 164880
rect 1104 164806 4315 164858
rect 4367 164806 4379 164858
rect 4431 164806 4443 164858
rect 4495 164806 4507 164858
rect 4559 164806 7648 164858
rect 7700 164806 7712 164858
rect 7764 164806 7776 164858
rect 7828 164806 7840 164858
rect 7892 164806 8832 164858
rect 1104 164784 8832 164806
rect 1104 164314 8832 164336
rect 1104 164262 2648 164314
rect 2700 164262 2712 164314
rect 2764 164262 2776 164314
rect 2828 164262 2840 164314
rect 2892 164262 5982 164314
rect 6034 164262 6046 164314
rect 6098 164262 6110 164314
rect 6162 164262 6174 164314
rect 6226 164262 8832 164314
rect 1104 164240 8832 164262
rect 1104 163770 8832 163792
rect 1104 163718 4315 163770
rect 4367 163718 4379 163770
rect 4431 163718 4443 163770
rect 4495 163718 4507 163770
rect 4559 163718 7648 163770
rect 7700 163718 7712 163770
rect 7764 163718 7776 163770
rect 7828 163718 7840 163770
rect 7892 163718 8832 163770
rect 1104 163696 8832 163718
rect 1104 163226 8832 163248
rect 1104 163174 2648 163226
rect 2700 163174 2712 163226
rect 2764 163174 2776 163226
rect 2828 163174 2840 163226
rect 2892 163174 5982 163226
rect 6034 163174 6046 163226
rect 6098 163174 6110 163226
rect 6162 163174 6174 163226
rect 6226 163174 8832 163226
rect 1104 163152 8832 163174
rect 1104 162682 8832 162704
rect 1104 162630 4315 162682
rect 4367 162630 4379 162682
rect 4431 162630 4443 162682
rect 4495 162630 4507 162682
rect 4559 162630 7648 162682
rect 7700 162630 7712 162682
rect 7764 162630 7776 162682
rect 7828 162630 7840 162682
rect 7892 162630 8832 162682
rect 1104 162608 8832 162630
rect 1104 162138 8832 162160
rect 1104 162086 2648 162138
rect 2700 162086 2712 162138
rect 2764 162086 2776 162138
rect 2828 162086 2840 162138
rect 2892 162086 5982 162138
rect 6034 162086 6046 162138
rect 6098 162086 6110 162138
rect 6162 162086 6174 162138
rect 6226 162086 8832 162138
rect 1104 162064 8832 162086
rect 1104 161594 8832 161616
rect 1104 161542 4315 161594
rect 4367 161542 4379 161594
rect 4431 161542 4443 161594
rect 4495 161542 4507 161594
rect 4559 161542 7648 161594
rect 7700 161542 7712 161594
rect 7764 161542 7776 161594
rect 7828 161542 7840 161594
rect 7892 161542 8832 161594
rect 1104 161520 8832 161542
rect 1104 161050 8832 161072
rect 1104 160998 2648 161050
rect 2700 160998 2712 161050
rect 2764 160998 2776 161050
rect 2828 160998 2840 161050
rect 2892 160998 5982 161050
rect 6034 160998 6046 161050
rect 6098 160998 6110 161050
rect 6162 160998 6174 161050
rect 6226 160998 8832 161050
rect 1104 160976 8832 160998
rect 1104 160506 8832 160528
rect 1104 160454 4315 160506
rect 4367 160454 4379 160506
rect 4431 160454 4443 160506
rect 4495 160454 4507 160506
rect 4559 160454 7648 160506
rect 7700 160454 7712 160506
rect 7764 160454 7776 160506
rect 7828 160454 7840 160506
rect 7892 160454 8832 160506
rect 1104 160432 8832 160454
rect 1104 159962 8832 159984
rect 1104 159910 2648 159962
rect 2700 159910 2712 159962
rect 2764 159910 2776 159962
rect 2828 159910 2840 159962
rect 2892 159910 5982 159962
rect 6034 159910 6046 159962
rect 6098 159910 6110 159962
rect 6162 159910 6174 159962
rect 6226 159910 8832 159962
rect 1104 159888 8832 159910
rect 1104 159418 8832 159440
rect 1104 159366 4315 159418
rect 4367 159366 4379 159418
rect 4431 159366 4443 159418
rect 4495 159366 4507 159418
rect 4559 159366 7648 159418
rect 7700 159366 7712 159418
rect 7764 159366 7776 159418
rect 7828 159366 7840 159418
rect 7892 159366 8832 159418
rect 1104 159344 8832 159366
rect 1104 158874 8832 158896
rect 1104 158822 2648 158874
rect 2700 158822 2712 158874
rect 2764 158822 2776 158874
rect 2828 158822 2840 158874
rect 2892 158822 5982 158874
rect 6034 158822 6046 158874
rect 6098 158822 6110 158874
rect 6162 158822 6174 158874
rect 6226 158822 8832 158874
rect 1104 158800 8832 158822
rect 1104 158330 8832 158352
rect 1104 158278 4315 158330
rect 4367 158278 4379 158330
rect 4431 158278 4443 158330
rect 4495 158278 4507 158330
rect 4559 158278 7648 158330
rect 7700 158278 7712 158330
rect 7764 158278 7776 158330
rect 7828 158278 7840 158330
rect 7892 158278 8832 158330
rect 1104 158256 8832 158278
rect 3418 158176 3424 158228
rect 3476 158216 3482 158228
rect 4249 158219 4307 158225
rect 4249 158216 4261 158219
rect 3476 158188 4261 158216
rect 3476 158176 3482 158188
rect 4249 158185 4261 158188
rect 4295 158185 4307 158219
rect 4249 158179 4307 158185
rect 6914 158148 6920 158160
rect 4080 158120 6920 158148
rect 4080 158092 4108 158120
rect 6914 158108 6920 158120
rect 6972 158148 6978 158160
rect 8018 158148 8024 158160
rect 6972 158120 8024 158148
rect 6972 158108 6978 158120
rect 8018 158108 8024 158120
rect 8076 158108 8082 158160
rect 4062 158089 4068 158092
rect 4053 158083 4068 158089
rect 4053 158080 4065 158083
rect 3975 158052 4065 158080
rect 4053 158049 4065 158052
rect 4053 158043 4068 158049
rect 4062 158040 4068 158043
rect 4120 158040 4126 158092
rect 1104 157786 8832 157808
rect 1104 157734 2648 157786
rect 2700 157734 2712 157786
rect 2764 157734 2776 157786
rect 2828 157734 2840 157786
rect 2892 157734 5982 157786
rect 6034 157734 6046 157786
rect 6098 157734 6110 157786
rect 6162 157734 6174 157786
rect 6226 157734 8832 157786
rect 1104 157712 8832 157734
rect 4062 157672 4068 157684
rect 4023 157644 4068 157672
rect 4062 157632 4068 157644
rect 4120 157632 4126 157684
rect 1104 157242 8832 157264
rect 1104 157190 4315 157242
rect 4367 157190 4379 157242
rect 4431 157190 4443 157242
rect 4495 157190 4507 157242
rect 4559 157190 7648 157242
rect 7700 157190 7712 157242
rect 7764 157190 7776 157242
rect 7828 157190 7840 157242
rect 7892 157190 8832 157242
rect 1104 157168 8832 157190
rect 1104 156698 8832 156720
rect 1104 156646 2648 156698
rect 2700 156646 2712 156698
rect 2764 156646 2776 156698
rect 2828 156646 2840 156698
rect 2892 156646 5982 156698
rect 6034 156646 6046 156698
rect 6098 156646 6110 156698
rect 6162 156646 6174 156698
rect 6226 156646 8832 156698
rect 1104 156624 8832 156646
rect 1104 156154 8832 156176
rect 1104 156102 4315 156154
rect 4367 156102 4379 156154
rect 4431 156102 4443 156154
rect 4495 156102 4507 156154
rect 4559 156102 7648 156154
rect 7700 156102 7712 156154
rect 7764 156102 7776 156154
rect 7828 156102 7840 156154
rect 7892 156102 8832 156154
rect 1104 156080 8832 156102
rect 1104 155610 8832 155632
rect 1104 155558 2648 155610
rect 2700 155558 2712 155610
rect 2764 155558 2776 155610
rect 2828 155558 2840 155610
rect 2892 155558 5982 155610
rect 6034 155558 6046 155610
rect 6098 155558 6110 155610
rect 6162 155558 6174 155610
rect 6226 155558 8832 155610
rect 1104 155536 8832 155558
rect 1104 155066 8832 155088
rect 1104 155014 4315 155066
rect 4367 155014 4379 155066
rect 4431 155014 4443 155066
rect 4495 155014 4507 155066
rect 4559 155014 7648 155066
rect 7700 155014 7712 155066
rect 7764 155014 7776 155066
rect 7828 155014 7840 155066
rect 7892 155014 8832 155066
rect 1104 154992 8832 155014
rect 1104 154522 8832 154544
rect 1104 154470 2648 154522
rect 2700 154470 2712 154522
rect 2764 154470 2776 154522
rect 2828 154470 2840 154522
rect 2892 154470 5982 154522
rect 6034 154470 6046 154522
rect 6098 154470 6110 154522
rect 6162 154470 6174 154522
rect 6226 154470 8832 154522
rect 1104 154448 8832 154470
rect 1104 153978 8832 154000
rect 1104 153926 4315 153978
rect 4367 153926 4379 153978
rect 4431 153926 4443 153978
rect 4495 153926 4507 153978
rect 4559 153926 7648 153978
rect 7700 153926 7712 153978
rect 7764 153926 7776 153978
rect 7828 153926 7840 153978
rect 7892 153926 8832 153978
rect 1104 153904 8832 153926
rect 1104 153434 8832 153456
rect 1104 153382 2648 153434
rect 2700 153382 2712 153434
rect 2764 153382 2776 153434
rect 2828 153382 2840 153434
rect 2892 153382 5982 153434
rect 6034 153382 6046 153434
rect 6098 153382 6110 153434
rect 6162 153382 6174 153434
rect 6226 153382 8832 153434
rect 1104 153360 8832 153382
rect 1104 152890 8832 152912
rect 1104 152838 4315 152890
rect 4367 152838 4379 152890
rect 4431 152838 4443 152890
rect 4495 152838 4507 152890
rect 4559 152838 7648 152890
rect 7700 152838 7712 152890
rect 7764 152838 7776 152890
rect 7828 152838 7840 152890
rect 7892 152838 8832 152890
rect 1104 152816 8832 152838
rect 1104 152346 8832 152368
rect 1104 152294 2648 152346
rect 2700 152294 2712 152346
rect 2764 152294 2776 152346
rect 2828 152294 2840 152346
rect 2892 152294 5982 152346
rect 6034 152294 6046 152346
rect 6098 152294 6110 152346
rect 6162 152294 6174 152346
rect 6226 152294 8832 152346
rect 1104 152272 8832 152294
rect 1104 151802 8832 151824
rect 1104 151750 4315 151802
rect 4367 151750 4379 151802
rect 4431 151750 4443 151802
rect 4495 151750 4507 151802
rect 4559 151750 7648 151802
rect 7700 151750 7712 151802
rect 7764 151750 7776 151802
rect 7828 151750 7840 151802
rect 7892 151750 8832 151802
rect 1104 151728 8832 151750
rect 1104 151258 8832 151280
rect 1104 151206 2648 151258
rect 2700 151206 2712 151258
rect 2764 151206 2776 151258
rect 2828 151206 2840 151258
rect 2892 151206 5982 151258
rect 6034 151206 6046 151258
rect 6098 151206 6110 151258
rect 6162 151206 6174 151258
rect 6226 151206 8832 151258
rect 1104 151184 8832 151206
rect 1104 150714 8832 150736
rect 1104 150662 4315 150714
rect 4367 150662 4379 150714
rect 4431 150662 4443 150714
rect 4495 150662 4507 150714
rect 4559 150662 7648 150714
rect 7700 150662 7712 150714
rect 7764 150662 7776 150714
rect 7828 150662 7840 150714
rect 7892 150662 8832 150714
rect 1104 150640 8832 150662
rect 1104 150170 8832 150192
rect 1104 150118 2648 150170
rect 2700 150118 2712 150170
rect 2764 150118 2776 150170
rect 2828 150118 2840 150170
rect 2892 150118 5982 150170
rect 6034 150118 6046 150170
rect 6098 150118 6110 150170
rect 6162 150118 6174 150170
rect 6226 150118 8832 150170
rect 1104 150096 8832 150118
rect 1104 149626 8832 149648
rect 1104 149574 4315 149626
rect 4367 149574 4379 149626
rect 4431 149574 4443 149626
rect 4495 149574 4507 149626
rect 4559 149574 7648 149626
rect 7700 149574 7712 149626
rect 7764 149574 7776 149626
rect 7828 149574 7840 149626
rect 7892 149574 8832 149626
rect 1104 149552 8832 149574
rect 1104 149082 8832 149104
rect 1104 149030 2648 149082
rect 2700 149030 2712 149082
rect 2764 149030 2776 149082
rect 2828 149030 2840 149082
rect 2892 149030 5982 149082
rect 6034 149030 6046 149082
rect 6098 149030 6110 149082
rect 6162 149030 6174 149082
rect 6226 149030 8832 149082
rect 1104 149008 8832 149030
rect 1104 148538 8832 148560
rect 1104 148486 4315 148538
rect 4367 148486 4379 148538
rect 4431 148486 4443 148538
rect 4495 148486 4507 148538
rect 4559 148486 7648 148538
rect 7700 148486 7712 148538
rect 7764 148486 7776 148538
rect 7828 148486 7840 148538
rect 7892 148486 8832 148538
rect 1104 148464 8832 148486
rect 1104 147994 8832 148016
rect 1104 147942 2648 147994
rect 2700 147942 2712 147994
rect 2764 147942 2776 147994
rect 2828 147942 2840 147994
rect 2892 147942 5982 147994
rect 6034 147942 6046 147994
rect 6098 147942 6110 147994
rect 6162 147942 6174 147994
rect 6226 147942 8832 147994
rect 1104 147920 8832 147942
rect 1104 147450 8832 147472
rect 1104 147398 4315 147450
rect 4367 147398 4379 147450
rect 4431 147398 4443 147450
rect 4495 147398 4507 147450
rect 4559 147398 7648 147450
rect 7700 147398 7712 147450
rect 7764 147398 7776 147450
rect 7828 147398 7840 147450
rect 7892 147398 8832 147450
rect 1104 147376 8832 147398
rect 1104 146906 8832 146928
rect 1104 146854 2648 146906
rect 2700 146854 2712 146906
rect 2764 146854 2776 146906
rect 2828 146854 2840 146906
rect 2892 146854 5982 146906
rect 6034 146854 6046 146906
rect 6098 146854 6110 146906
rect 6162 146854 6174 146906
rect 6226 146854 8832 146906
rect 1104 146832 8832 146854
rect 1104 146362 8832 146384
rect 1104 146310 4315 146362
rect 4367 146310 4379 146362
rect 4431 146310 4443 146362
rect 4495 146310 4507 146362
rect 4559 146310 7648 146362
rect 7700 146310 7712 146362
rect 7764 146310 7776 146362
rect 7828 146310 7840 146362
rect 7892 146310 8832 146362
rect 1104 146288 8832 146310
rect 1104 145818 8832 145840
rect 1104 145766 2648 145818
rect 2700 145766 2712 145818
rect 2764 145766 2776 145818
rect 2828 145766 2840 145818
rect 2892 145766 5982 145818
rect 6034 145766 6046 145818
rect 6098 145766 6110 145818
rect 6162 145766 6174 145818
rect 6226 145766 8832 145818
rect 1104 145744 8832 145766
rect 1104 145274 8832 145296
rect 1104 145222 4315 145274
rect 4367 145222 4379 145274
rect 4431 145222 4443 145274
rect 4495 145222 4507 145274
rect 4559 145222 7648 145274
rect 7700 145222 7712 145274
rect 7764 145222 7776 145274
rect 7828 145222 7840 145274
rect 7892 145222 8832 145274
rect 1104 145200 8832 145222
rect 1104 144730 8832 144752
rect 1104 144678 2648 144730
rect 2700 144678 2712 144730
rect 2764 144678 2776 144730
rect 2828 144678 2840 144730
rect 2892 144678 5982 144730
rect 6034 144678 6046 144730
rect 6098 144678 6110 144730
rect 6162 144678 6174 144730
rect 6226 144678 8832 144730
rect 1104 144656 8832 144678
rect 1104 144186 8832 144208
rect 1104 144134 4315 144186
rect 4367 144134 4379 144186
rect 4431 144134 4443 144186
rect 4495 144134 4507 144186
rect 4559 144134 7648 144186
rect 7700 144134 7712 144186
rect 7764 144134 7776 144186
rect 7828 144134 7840 144186
rect 7892 144134 8832 144186
rect 1104 144112 8832 144134
rect 1104 143642 8832 143664
rect 1104 143590 2648 143642
rect 2700 143590 2712 143642
rect 2764 143590 2776 143642
rect 2828 143590 2840 143642
rect 2892 143590 5982 143642
rect 6034 143590 6046 143642
rect 6098 143590 6110 143642
rect 6162 143590 6174 143642
rect 6226 143590 8832 143642
rect 1104 143568 8832 143590
rect 1104 143098 8832 143120
rect 1104 143046 4315 143098
rect 4367 143046 4379 143098
rect 4431 143046 4443 143098
rect 4495 143046 4507 143098
rect 4559 143046 7648 143098
rect 7700 143046 7712 143098
rect 7764 143046 7776 143098
rect 7828 143046 7840 143098
rect 7892 143046 8832 143098
rect 1104 143024 8832 143046
rect 1104 142554 8832 142576
rect 1104 142502 2648 142554
rect 2700 142502 2712 142554
rect 2764 142502 2776 142554
rect 2828 142502 2840 142554
rect 2892 142502 5982 142554
rect 6034 142502 6046 142554
rect 6098 142502 6110 142554
rect 6162 142502 6174 142554
rect 6226 142502 8832 142554
rect 1104 142480 8832 142502
rect 1104 142010 8832 142032
rect 1104 141958 4315 142010
rect 4367 141958 4379 142010
rect 4431 141958 4443 142010
rect 4495 141958 4507 142010
rect 4559 141958 7648 142010
rect 7700 141958 7712 142010
rect 7764 141958 7776 142010
rect 7828 141958 7840 142010
rect 7892 141958 8832 142010
rect 1104 141936 8832 141958
rect 1104 141466 8832 141488
rect 1104 141414 2648 141466
rect 2700 141414 2712 141466
rect 2764 141414 2776 141466
rect 2828 141414 2840 141466
rect 2892 141414 5982 141466
rect 6034 141414 6046 141466
rect 6098 141414 6110 141466
rect 6162 141414 6174 141466
rect 6226 141414 8832 141466
rect 1104 141392 8832 141414
rect 1104 140922 8832 140944
rect 1104 140870 4315 140922
rect 4367 140870 4379 140922
rect 4431 140870 4443 140922
rect 4495 140870 4507 140922
rect 4559 140870 7648 140922
rect 7700 140870 7712 140922
rect 7764 140870 7776 140922
rect 7828 140870 7840 140922
rect 7892 140870 8832 140922
rect 1104 140848 8832 140870
rect 1104 140378 8832 140400
rect 1104 140326 2648 140378
rect 2700 140326 2712 140378
rect 2764 140326 2776 140378
rect 2828 140326 2840 140378
rect 2892 140326 5982 140378
rect 6034 140326 6046 140378
rect 6098 140326 6110 140378
rect 6162 140326 6174 140378
rect 6226 140326 8832 140378
rect 1104 140304 8832 140326
rect 1104 139834 8832 139856
rect 1104 139782 4315 139834
rect 4367 139782 4379 139834
rect 4431 139782 4443 139834
rect 4495 139782 4507 139834
rect 4559 139782 7648 139834
rect 7700 139782 7712 139834
rect 7764 139782 7776 139834
rect 7828 139782 7840 139834
rect 7892 139782 8832 139834
rect 1104 139760 8832 139782
rect 1104 139290 8832 139312
rect 1104 139238 2648 139290
rect 2700 139238 2712 139290
rect 2764 139238 2776 139290
rect 2828 139238 2840 139290
rect 2892 139238 5982 139290
rect 6034 139238 6046 139290
rect 6098 139238 6110 139290
rect 6162 139238 6174 139290
rect 6226 139238 8832 139290
rect 1104 139216 8832 139238
rect 1104 138746 8832 138768
rect 1104 138694 4315 138746
rect 4367 138694 4379 138746
rect 4431 138694 4443 138746
rect 4495 138694 4507 138746
rect 4559 138694 7648 138746
rect 7700 138694 7712 138746
rect 7764 138694 7776 138746
rect 7828 138694 7840 138746
rect 7892 138694 8832 138746
rect 1104 138672 8832 138694
rect 1104 138202 8832 138224
rect 1104 138150 2648 138202
rect 2700 138150 2712 138202
rect 2764 138150 2776 138202
rect 2828 138150 2840 138202
rect 2892 138150 5982 138202
rect 6034 138150 6046 138202
rect 6098 138150 6110 138202
rect 6162 138150 6174 138202
rect 6226 138150 8832 138202
rect 1104 138128 8832 138150
rect 1104 137658 8832 137680
rect 1104 137606 4315 137658
rect 4367 137606 4379 137658
rect 4431 137606 4443 137658
rect 4495 137606 4507 137658
rect 4559 137606 7648 137658
rect 7700 137606 7712 137658
rect 7764 137606 7776 137658
rect 7828 137606 7840 137658
rect 7892 137606 8832 137658
rect 1104 137584 8832 137606
rect 1104 137114 8832 137136
rect 1104 137062 2648 137114
rect 2700 137062 2712 137114
rect 2764 137062 2776 137114
rect 2828 137062 2840 137114
rect 2892 137062 5982 137114
rect 6034 137062 6046 137114
rect 6098 137062 6110 137114
rect 6162 137062 6174 137114
rect 6226 137062 8832 137114
rect 1104 137040 8832 137062
rect 1104 136570 8832 136592
rect 1104 136518 4315 136570
rect 4367 136518 4379 136570
rect 4431 136518 4443 136570
rect 4495 136518 4507 136570
rect 4559 136518 7648 136570
rect 7700 136518 7712 136570
rect 7764 136518 7776 136570
rect 7828 136518 7840 136570
rect 7892 136518 8832 136570
rect 1104 136496 8832 136518
rect 1104 136026 8832 136048
rect 1104 135974 2648 136026
rect 2700 135974 2712 136026
rect 2764 135974 2776 136026
rect 2828 135974 2840 136026
rect 2892 135974 5982 136026
rect 6034 135974 6046 136026
rect 6098 135974 6110 136026
rect 6162 135974 6174 136026
rect 6226 135974 8832 136026
rect 1104 135952 8832 135974
rect 1104 135482 8832 135504
rect 1104 135430 4315 135482
rect 4367 135430 4379 135482
rect 4431 135430 4443 135482
rect 4495 135430 4507 135482
rect 4559 135430 7648 135482
rect 7700 135430 7712 135482
rect 7764 135430 7776 135482
rect 7828 135430 7840 135482
rect 7892 135430 8832 135482
rect 1104 135408 8832 135430
rect 1104 134938 8832 134960
rect 1104 134886 2648 134938
rect 2700 134886 2712 134938
rect 2764 134886 2776 134938
rect 2828 134886 2840 134938
rect 2892 134886 5982 134938
rect 6034 134886 6046 134938
rect 6098 134886 6110 134938
rect 6162 134886 6174 134938
rect 6226 134886 8832 134938
rect 1104 134864 8832 134886
rect 1104 134394 8832 134416
rect 1104 134342 4315 134394
rect 4367 134342 4379 134394
rect 4431 134342 4443 134394
rect 4495 134342 4507 134394
rect 4559 134342 7648 134394
rect 7700 134342 7712 134394
rect 7764 134342 7776 134394
rect 7828 134342 7840 134394
rect 7892 134342 8832 134394
rect 1104 134320 8832 134342
rect 1104 133850 8832 133872
rect 1104 133798 2648 133850
rect 2700 133798 2712 133850
rect 2764 133798 2776 133850
rect 2828 133798 2840 133850
rect 2892 133798 5982 133850
rect 6034 133798 6046 133850
rect 6098 133798 6110 133850
rect 6162 133798 6174 133850
rect 6226 133798 8832 133850
rect 1104 133776 8832 133798
rect 1104 133306 8832 133328
rect 1104 133254 4315 133306
rect 4367 133254 4379 133306
rect 4431 133254 4443 133306
rect 4495 133254 4507 133306
rect 4559 133254 7648 133306
rect 7700 133254 7712 133306
rect 7764 133254 7776 133306
rect 7828 133254 7840 133306
rect 7892 133254 8832 133306
rect 1104 133232 8832 133254
rect 1104 132762 8832 132784
rect 1104 132710 2648 132762
rect 2700 132710 2712 132762
rect 2764 132710 2776 132762
rect 2828 132710 2840 132762
rect 2892 132710 5982 132762
rect 6034 132710 6046 132762
rect 6098 132710 6110 132762
rect 6162 132710 6174 132762
rect 6226 132710 8832 132762
rect 1104 132688 8832 132710
rect 1104 132218 8832 132240
rect 1104 132166 4315 132218
rect 4367 132166 4379 132218
rect 4431 132166 4443 132218
rect 4495 132166 4507 132218
rect 4559 132166 7648 132218
rect 7700 132166 7712 132218
rect 7764 132166 7776 132218
rect 7828 132166 7840 132218
rect 7892 132166 8832 132218
rect 1104 132144 8832 132166
rect 1104 131674 8832 131696
rect 1104 131622 2648 131674
rect 2700 131622 2712 131674
rect 2764 131622 2776 131674
rect 2828 131622 2840 131674
rect 2892 131622 5982 131674
rect 6034 131622 6046 131674
rect 6098 131622 6110 131674
rect 6162 131622 6174 131674
rect 6226 131622 8832 131674
rect 1104 131600 8832 131622
rect 1104 131130 8832 131152
rect 1104 131078 4315 131130
rect 4367 131078 4379 131130
rect 4431 131078 4443 131130
rect 4495 131078 4507 131130
rect 4559 131078 7648 131130
rect 7700 131078 7712 131130
rect 7764 131078 7776 131130
rect 7828 131078 7840 131130
rect 7892 131078 8832 131130
rect 1104 131056 8832 131078
rect 1104 130586 8832 130608
rect 1104 130534 2648 130586
rect 2700 130534 2712 130586
rect 2764 130534 2776 130586
rect 2828 130534 2840 130586
rect 2892 130534 5982 130586
rect 6034 130534 6046 130586
rect 6098 130534 6110 130586
rect 6162 130534 6174 130586
rect 6226 130534 8832 130586
rect 1104 130512 8832 130534
rect 1104 130042 8832 130064
rect 1104 129990 4315 130042
rect 4367 129990 4379 130042
rect 4431 129990 4443 130042
rect 4495 129990 4507 130042
rect 4559 129990 7648 130042
rect 7700 129990 7712 130042
rect 7764 129990 7776 130042
rect 7828 129990 7840 130042
rect 7892 129990 8832 130042
rect 1104 129968 8832 129990
rect 1104 129498 8832 129520
rect 1104 129446 2648 129498
rect 2700 129446 2712 129498
rect 2764 129446 2776 129498
rect 2828 129446 2840 129498
rect 2892 129446 5982 129498
rect 6034 129446 6046 129498
rect 6098 129446 6110 129498
rect 6162 129446 6174 129498
rect 6226 129446 8832 129498
rect 1104 129424 8832 129446
rect 1104 128954 8832 128976
rect 1104 128902 4315 128954
rect 4367 128902 4379 128954
rect 4431 128902 4443 128954
rect 4495 128902 4507 128954
rect 4559 128902 7648 128954
rect 7700 128902 7712 128954
rect 7764 128902 7776 128954
rect 7828 128902 7840 128954
rect 7892 128902 8832 128954
rect 1104 128880 8832 128902
rect 1104 128410 8832 128432
rect 1104 128358 2648 128410
rect 2700 128358 2712 128410
rect 2764 128358 2776 128410
rect 2828 128358 2840 128410
rect 2892 128358 5982 128410
rect 6034 128358 6046 128410
rect 6098 128358 6110 128410
rect 6162 128358 6174 128410
rect 6226 128358 8832 128410
rect 1104 128336 8832 128358
rect 1104 127866 8832 127888
rect 1104 127814 4315 127866
rect 4367 127814 4379 127866
rect 4431 127814 4443 127866
rect 4495 127814 4507 127866
rect 4559 127814 7648 127866
rect 7700 127814 7712 127866
rect 7764 127814 7776 127866
rect 7828 127814 7840 127866
rect 7892 127814 8832 127866
rect 1104 127792 8832 127814
rect 1104 127322 8832 127344
rect 1104 127270 2648 127322
rect 2700 127270 2712 127322
rect 2764 127270 2776 127322
rect 2828 127270 2840 127322
rect 2892 127270 5982 127322
rect 6034 127270 6046 127322
rect 6098 127270 6110 127322
rect 6162 127270 6174 127322
rect 6226 127270 8832 127322
rect 1104 127248 8832 127270
rect 1104 126778 8832 126800
rect 1104 126726 4315 126778
rect 4367 126726 4379 126778
rect 4431 126726 4443 126778
rect 4495 126726 4507 126778
rect 4559 126726 7648 126778
rect 7700 126726 7712 126778
rect 7764 126726 7776 126778
rect 7828 126726 7840 126778
rect 7892 126726 8832 126778
rect 1104 126704 8832 126726
rect 1104 126234 8832 126256
rect 1104 126182 2648 126234
rect 2700 126182 2712 126234
rect 2764 126182 2776 126234
rect 2828 126182 2840 126234
rect 2892 126182 5982 126234
rect 6034 126182 6046 126234
rect 6098 126182 6110 126234
rect 6162 126182 6174 126234
rect 6226 126182 8832 126234
rect 1104 126160 8832 126182
rect 1104 125690 8832 125712
rect 1104 125638 4315 125690
rect 4367 125638 4379 125690
rect 4431 125638 4443 125690
rect 4495 125638 4507 125690
rect 4559 125638 7648 125690
rect 7700 125638 7712 125690
rect 7764 125638 7776 125690
rect 7828 125638 7840 125690
rect 7892 125638 8832 125690
rect 1104 125616 8832 125638
rect 1104 125146 8832 125168
rect 1104 125094 2648 125146
rect 2700 125094 2712 125146
rect 2764 125094 2776 125146
rect 2828 125094 2840 125146
rect 2892 125094 5982 125146
rect 6034 125094 6046 125146
rect 6098 125094 6110 125146
rect 6162 125094 6174 125146
rect 6226 125094 8832 125146
rect 1104 125072 8832 125094
rect 1104 124602 8832 124624
rect 1104 124550 4315 124602
rect 4367 124550 4379 124602
rect 4431 124550 4443 124602
rect 4495 124550 4507 124602
rect 4559 124550 7648 124602
rect 7700 124550 7712 124602
rect 7764 124550 7776 124602
rect 7828 124550 7840 124602
rect 7892 124550 8832 124602
rect 1104 124528 8832 124550
rect 1104 124058 8832 124080
rect 1104 124006 2648 124058
rect 2700 124006 2712 124058
rect 2764 124006 2776 124058
rect 2828 124006 2840 124058
rect 2892 124006 5982 124058
rect 6034 124006 6046 124058
rect 6098 124006 6110 124058
rect 6162 124006 6174 124058
rect 6226 124006 8832 124058
rect 1104 123984 8832 124006
rect 1104 123514 8832 123536
rect 1104 123462 4315 123514
rect 4367 123462 4379 123514
rect 4431 123462 4443 123514
rect 4495 123462 4507 123514
rect 4559 123462 7648 123514
rect 7700 123462 7712 123514
rect 7764 123462 7776 123514
rect 7828 123462 7840 123514
rect 7892 123462 8832 123514
rect 1104 123440 8832 123462
rect 1104 122970 8832 122992
rect 1104 122918 2648 122970
rect 2700 122918 2712 122970
rect 2764 122918 2776 122970
rect 2828 122918 2840 122970
rect 2892 122918 5982 122970
rect 6034 122918 6046 122970
rect 6098 122918 6110 122970
rect 6162 122918 6174 122970
rect 6226 122918 8832 122970
rect 1104 122896 8832 122918
rect 1104 122426 8832 122448
rect 1104 122374 4315 122426
rect 4367 122374 4379 122426
rect 4431 122374 4443 122426
rect 4495 122374 4507 122426
rect 4559 122374 7648 122426
rect 7700 122374 7712 122426
rect 7764 122374 7776 122426
rect 7828 122374 7840 122426
rect 7892 122374 8832 122426
rect 1104 122352 8832 122374
rect 1104 121882 8832 121904
rect 1104 121830 2648 121882
rect 2700 121830 2712 121882
rect 2764 121830 2776 121882
rect 2828 121830 2840 121882
rect 2892 121830 5982 121882
rect 6034 121830 6046 121882
rect 6098 121830 6110 121882
rect 6162 121830 6174 121882
rect 6226 121830 8832 121882
rect 1104 121808 8832 121830
rect 1104 121338 8832 121360
rect 1104 121286 4315 121338
rect 4367 121286 4379 121338
rect 4431 121286 4443 121338
rect 4495 121286 4507 121338
rect 4559 121286 7648 121338
rect 7700 121286 7712 121338
rect 7764 121286 7776 121338
rect 7828 121286 7840 121338
rect 7892 121286 8832 121338
rect 1104 121264 8832 121286
rect 1104 120794 8832 120816
rect 1104 120742 2648 120794
rect 2700 120742 2712 120794
rect 2764 120742 2776 120794
rect 2828 120742 2840 120794
rect 2892 120742 5982 120794
rect 6034 120742 6046 120794
rect 6098 120742 6110 120794
rect 6162 120742 6174 120794
rect 6226 120742 8832 120794
rect 1104 120720 8832 120742
rect 1104 120250 8832 120272
rect 1104 120198 4315 120250
rect 4367 120198 4379 120250
rect 4431 120198 4443 120250
rect 4495 120198 4507 120250
rect 4559 120198 7648 120250
rect 7700 120198 7712 120250
rect 7764 120198 7776 120250
rect 7828 120198 7840 120250
rect 7892 120198 8832 120250
rect 1104 120176 8832 120198
rect 1104 119706 8832 119728
rect 1104 119654 2648 119706
rect 2700 119654 2712 119706
rect 2764 119654 2776 119706
rect 2828 119654 2840 119706
rect 2892 119654 5982 119706
rect 6034 119654 6046 119706
rect 6098 119654 6110 119706
rect 6162 119654 6174 119706
rect 6226 119654 8832 119706
rect 1104 119632 8832 119654
rect 1104 119162 8832 119184
rect 1104 119110 4315 119162
rect 4367 119110 4379 119162
rect 4431 119110 4443 119162
rect 4495 119110 4507 119162
rect 4559 119110 7648 119162
rect 7700 119110 7712 119162
rect 7764 119110 7776 119162
rect 7828 119110 7840 119162
rect 7892 119110 8832 119162
rect 1104 119088 8832 119110
rect 1104 118618 8832 118640
rect 1104 118566 2648 118618
rect 2700 118566 2712 118618
rect 2764 118566 2776 118618
rect 2828 118566 2840 118618
rect 2892 118566 5982 118618
rect 6034 118566 6046 118618
rect 6098 118566 6110 118618
rect 6162 118566 6174 118618
rect 6226 118566 8832 118618
rect 1104 118544 8832 118566
rect 1104 118074 8832 118096
rect 1104 118022 4315 118074
rect 4367 118022 4379 118074
rect 4431 118022 4443 118074
rect 4495 118022 4507 118074
rect 4559 118022 7648 118074
rect 7700 118022 7712 118074
rect 7764 118022 7776 118074
rect 7828 118022 7840 118074
rect 7892 118022 8832 118074
rect 1104 118000 8832 118022
rect 1104 117530 8832 117552
rect 1104 117478 2648 117530
rect 2700 117478 2712 117530
rect 2764 117478 2776 117530
rect 2828 117478 2840 117530
rect 2892 117478 5982 117530
rect 6034 117478 6046 117530
rect 6098 117478 6110 117530
rect 6162 117478 6174 117530
rect 6226 117478 8832 117530
rect 1104 117456 8832 117478
rect 1104 116986 8832 117008
rect 1104 116934 4315 116986
rect 4367 116934 4379 116986
rect 4431 116934 4443 116986
rect 4495 116934 4507 116986
rect 4559 116934 7648 116986
rect 7700 116934 7712 116986
rect 7764 116934 7776 116986
rect 7828 116934 7840 116986
rect 7892 116934 8832 116986
rect 1104 116912 8832 116934
rect 1104 116442 8832 116464
rect 1104 116390 2648 116442
rect 2700 116390 2712 116442
rect 2764 116390 2776 116442
rect 2828 116390 2840 116442
rect 2892 116390 5982 116442
rect 6034 116390 6046 116442
rect 6098 116390 6110 116442
rect 6162 116390 6174 116442
rect 6226 116390 8832 116442
rect 1104 116368 8832 116390
rect 1104 115898 8832 115920
rect 1104 115846 4315 115898
rect 4367 115846 4379 115898
rect 4431 115846 4443 115898
rect 4495 115846 4507 115898
rect 4559 115846 7648 115898
rect 7700 115846 7712 115898
rect 7764 115846 7776 115898
rect 7828 115846 7840 115898
rect 7892 115846 8832 115898
rect 1104 115824 8832 115846
rect 1104 115354 8832 115376
rect 1104 115302 2648 115354
rect 2700 115302 2712 115354
rect 2764 115302 2776 115354
rect 2828 115302 2840 115354
rect 2892 115302 5982 115354
rect 6034 115302 6046 115354
rect 6098 115302 6110 115354
rect 6162 115302 6174 115354
rect 6226 115302 8832 115354
rect 1104 115280 8832 115302
rect 1104 114810 8832 114832
rect 1104 114758 4315 114810
rect 4367 114758 4379 114810
rect 4431 114758 4443 114810
rect 4495 114758 4507 114810
rect 4559 114758 7648 114810
rect 7700 114758 7712 114810
rect 7764 114758 7776 114810
rect 7828 114758 7840 114810
rect 7892 114758 8832 114810
rect 1104 114736 8832 114758
rect 1104 114266 8832 114288
rect 1104 114214 2648 114266
rect 2700 114214 2712 114266
rect 2764 114214 2776 114266
rect 2828 114214 2840 114266
rect 2892 114214 5982 114266
rect 6034 114214 6046 114266
rect 6098 114214 6110 114266
rect 6162 114214 6174 114266
rect 6226 114214 8832 114266
rect 1104 114192 8832 114214
rect 1104 113722 8832 113744
rect 1104 113670 4315 113722
rect 4367 113670 4379 113722
rect 4431 113670 4443 113722
rect 4495 113670 4507 113722
rect 4559 113670 7648 113722
rect 7700 113670 7712 113722
rect 7764 113670 7776 113722
rect 7828 113670 7840 113722
rect 7892 113670 8832 113722
rect 1104 113648 8832 113670
rect 1104 113178 8832 113200
rect 1104 113126 2648 113178
rect 2700 113126 2712 113178
rect 2764 113126 2776 113178
rect 2828 113126 2840 113178
rect 2892 113126 5982 113178
rect 6034 113126 6046 113178
rect 6098 113126 6110 113178
rect 6162 113126 6174 113178
rect 6226 113126 8832 113178
rect 1104 113104 8832 113126
rect 1104 112634 8832 112656
rect 1104 112582 4315 112634
rect 4367 112582 4379 112634
rect 4431 112582 4443 112634
rect 4495 112582 4507 112634
rect 4559 112582 7648 112634
rect 7700 112582 7712 112634
rect 7764 112582 7776 112634
rect 7828 112582 7840 112634
rect 7892 112582 8832 112634
rect 1104 112560 8832 112582
rect 1104 112090 8832 112112
rect 1104 112038 2648 112090
rect 2700 112038 2712 112090
rect 2764 112038 2776 112090
rect 2828 112038 2840 112090
rect 2892 112038 5982 112090
rect 6034 112038 6046 112090
rect 6098 112038 6110 112090
rect 6162 112038 6174 112090
rect 6226 112038 8832 112090
rect 1104 112016 8832 112038
rect 1104 111546 8832 111568
rect 1104 111494 4315 111546
rect 4367 111494 4379 111546
rect 4431 111494 4443 111546
rect 4495 111494 4507 111546
rect 4559 111494 7648 111546
rect 7700 111494 7712 111546
rect 7764 111494 7776 111546
rect 7828 111494 7840 111546
rect 7892 111494 8832 111546
rect 1104 111472 8832 111494
rect 1104 111002 8832 111024
rect 1104 110950 2648 111002
rect 2700 110950 2712 111002
rect 2764 110950 2776 111002
rect 2828 110950 2840 111002
rect 2892 110950 5982 111002
rect 6034 110950 6046 111002
rect 6098 110950 6110 111002
rect 6162 110950 6174 111002
rect 6226 110950 8832 111002
rect 1104 110928 8832 110950
rect 1104 110458 8832 110480
rect 1104 110406 4315 110458
rect 4367 110406 4379 110458
rect 4431 110406 4443 110458
rect 4495 110406 4507 110458
rect 4559 110406 7648 110458
rect 7700 110406 7712 110458
rect 7764 110406 7776 110458
rect 7828 110406 7840 110458
rect 7892 110406 8832 110458
rect 1104 110384 8832 110406
rect 1104 109914 8832 109936
rect 1104 109862 2648 109914
rect 2700 109862 2712 109914
rect 2764 109862 2776 109914
rect 2828 109862 2840 109914
rect 2892 109862 5982 109914
rect 6034 109862 6046 109914
rect 6098 109862 6110 109914
rect 6162 109862 6174 109914
rect 6226 109862 8832 109914
rect 1104 109840 8832 109862
rect 1104 109370 8832 109392
rect 1104 109318 4315 109370
rect 4367 109318 4379 109370
rect 4431 109318 4443 109370
rect 4495 109318 4507 109370
rect 4559 109318 7648 109370
rect 7700 109318 7712 109370
rect 7764 109318 7776 109370
rect 7828 109318 7840 109370
rect 7892 109318 8832 109370
rect 1104 109296 8832 109318
rect 1104 108826 8832 108848
rect 1104 108774 2648 108826
rect 2700 108774 2712 108826
rect 2764 108774 2776 108826
rect 2828 108774 2840 108826
rect 2892 108774 5982 108826
rect 6034 108774 6046 108826
rect 6098 108774 6110 108826
rect 6162 108774 6174 108826
rect 6226 108774 8832 108826
rect 1104 108752 8832 108774
rect 1104 108282 8832 108304
rect 1104 108230 4315 108282
rect 4367 108230 4379 108282
rect 4431 108230 4443 108282
rect 4495 108230 4507 108282
rect 4559 108230 7648 108282
rect 7700 108230 7712 108282
rect 7764 108230 7776 108282
rect 7828 108230 7840 108282
rect 7892 108230 8832 108282
rect 1104 108208 8832 108230
rect 1104 107738 8832 107760
rect 1104 107686 2648 107738
rect 2700 107686 2712 107738
rect 2764 107686 2776 107738
rect 2828 107686 2840 107738
rect 2892 107686 5982 107738
rect 6034 107686 6046 107738
rect 6098 107686 6110 107738
rect 6162 107686 6174 107738
rect 6226 107686 8832 107738
rect 1104 107664 8832 107686
rect 1104 107194 8832 107216
rect 1104 107142 4315 107194
rect 4367 107142 4379 107194
rect 4431 107142 4443 107194
rect 4495 107142 4507 107194
rect 4559 107142 7648 107194
rect 7700 107142 7712 107194
rect 7764 107142 7776 107194
rect 7828 107142 7840 107194
rect 7892 107142 8832 107194
rect 1104 107120 8832 107142
rect 1104 106650 8832 106672
rect 1104 106598 2648 106650
rect 2700 106598 2712 106650
rect 2764 106598 2776 106650
rect 2828 106598 2840 106650
rect 2892 106598 5982 106650
rect 6034 106598 6046 106650
rect 6098 106598 6110 106650
rect 6162 106598 6174 106650
rect 6226 106598 8832 106650
rect 1104 106576 8832 106598
rect 1104 106106 8832 106128
rect 1104 106054 4315 106106
rect 4367 106054 4379 106106
rect 4431 106054 4443 106106
rect 4495 106054 4507 106106
rect 4559 106054 7648 106106
rect 7700 106054 7712 106106
rect 7764 106054 7776 106106
rect 7828 106054 7840 106106
rect 7892 106054 8832 106106
rect 1104 106032 8832 106054
rect 1104 105562 8832 105584
rect 1104 105510 2648 105562
rect 2700 105510 2712 105562
rect 2764 105510 2776 105562
rect 2828 105510 2840 105562
rect 2892 105510 5982 105562
rect 6034 105510 6046 105562
rect 6098 105510 6110 105562
rect 6162 105510 6174 105562
rect 6226 105510 8832 105562
rect 1104 105488 8832 105510
rect 1104 105018 8832 105040
rect 1104 104966 4315 105018
rect 4367 104966 4379 105018
rect 4431 104966 4443 105018
rect 4495 104966 4507 105018
rect 4559 104966 7648 105018
rect 7700 104966 7712 105018
rect 7764 104966 7776 105018
rect 7828 104966 7840 105018
rect 7892 104966 8832 105018
rect 1104 104944 8832 104966
rect 1104 104474 8832 104496
rect 1104 104422 2648 104474
rect 2700 104422 2712 104474
rect 2764 104422 2776 104474
rect 2828 104422 2840 104474
rect 2892 104422 5982 104474
rect 6034 104422 6046 104474
rect 6098 104422 6110 104474
rect 6162 104422 6174 104474
rect 6226 104422 8832 104474
rect 1104 104400 8832 104422
rect 1104 103930 8832 103952
rect 1104 103878 4315 103930
rect 4367 103878 4379 103930
rect 4431 103878 4443 103930
rect 4495 103878 4507 103930
rect 4559 103878 7648 103930
rect 7700 103878 7712 103930
rect 7764 103878 7776 103930
rect 7828 103878 7840 103930
rect 7892 103878 8832 103930
rect 1104 103856 8832 103878
rect 1104 103386 8832 103408
rect 1104 103334 2648 103386
rect 2700 103334 2712 103386
rect 2764 103334 2776 103386
rect 2828 103334 2840 103386
rect 2892 103334 5982 103386
rect 6034 103334 6046 103386
rect 6098 103334 6110 103386
rect 6162 103334 6174 103386
rect 6226 103334 8832 103386
rect 1104 103312 8832 103334
rect 1104 102842 8832 102864
rect 1104 102790 4315 102842
rect 4367 102790 4379 102842
rect 4431 102790 4443 102842
rect 4495 102790 4507 102842
rect 4559 102790 7648 102842
rect 7700 102790 7712 102842
rect 7764 102790 7776 102842
rect 7828 102790 7840 102842
rect 7892 102790 8832 102842
rect 1104 102768 8832 102790
rect 1104 102298 8832 102320
rect 1104 102246 2648 102298
rect 2700 102246 2712 102298
rect 2764 102246 2776 102298
rect 2828 102246 2840 102298
rect 2892 102246 5982 102298
rect 6034 102246 6046 102298
rect 6098 102246 6110 102298
rect 6162 102246 6174 102298
rect 6226 102246 8832 102298
rect 1104 102224 8832 102246
rect 1104 101754 8832 101776
rect 1104 101702 4315 101754
rect 4367 101702 4379 101754
rect 4431 101702 4443 101754
rect 4495 101702 4507 101754
rect 4559 101702 7648 101754
rect 7700 101702 7712 101754
rect 7764 101702 7776 101754
rect 7828 101702 7840 101754
rect 7892 101702 8832 101754
rect 1104 101680 8832 101702
rect 1104 101210 8832 101232
rect 1104 101158 2648 101210
rect 2700 101158 2712 101210
rect 2764 101158 2776 101210
rect 2828 101158 2840 101210
rect 2892 101158 5982 101210
rect 6034 101158 6046 101210
rect 6098 101158 6110 101210
rect 6162 101158 6174 101210
rect 6226 101158 8832 101210
rect 1104 101136 8832 101158
rect 1104 100666 8832 100688
rect 1104 100614 4315 100666
rect 4367 100614 4379 100666
rect 4431 100614 4443 100666
rect 4495 100614 4507 100666
rect 4559 100614 7648 100666
rect 7700 100614 7712 100666
rect 7764 100614 7776 100666
rect 7828 100614 7840 100666
rect 7892 100614 8832 100666
rect 1104 100592 8832 100614
rect 1104 100122 8832 100144
rect 1104 100070 2648 100122
rect 2700 100070 2712 100122
rect 2764 100070 2776 100122
rect 2828 100070 2840 100122
rect 2892 100070 5982 100122
rect 6034 100070 6046 100122
rect 6098 100070 6110 100122
rect 6162 100070 6174 100122
rect 6226 100070 8832 100122
rect 1104 100048 8832 100070
rect 1104 99578 8832 99600
rect 1104 99526 4315 99578
rect 4367 99526 4379 99578
rect 4431 99526 4443 99578
rect 4495 99526 4507 99578
rect 4559 99526 7648 99578
rect 7700 99526 7712 99578
rect 7764 99526 7776 99578
rect 7828 99526 7840 99578
rect 7892 99526 8832 99578
rect 1104 99504 8832 99526
rect 1104 99034 8832 99056
rect 1104 98982 2648 99034
rect 2700 98982 2712 99034
rect 2764 98982 2776 99034
rect 2828 98982 2840 99034
rect 2892 98982 5982 99034
rect 6034 98982 6046 99034
rect 6098 98982 6110 99034
rect 6162 98982 6174 99034
rect 6226 98982 8832 99034
rect 1104 98960 8832 98982
rect 1104 98490 8832 98512
rect 1104 98438 4315 98490
rect 4367 98438 4379 98490
rect 4431 98438 4443 98490
rect 4495 98438 4507 98490
rect 4559 98438 7648 98490
rect 7700 98438 7712 98490
rect 7764 98438 7776 98490
rect 7828 98438 7840 98490
rect 7892 98438 8832 98490
rect 1104 98416 8832 98438
rect 1104 97946 8832 97968
rect 1104 97894 2648 97946
rect 2700 97894 2712 97946
rect 2764 97894 2776 97946
rect 2828 97894 2840 97946
rect 2892 97894 5982 97946
rect 6034 97894 6046 97946
rect 6098 97894 6110 97946
rect 6162 97894 6174 97946
rect 6226 97894 8832 97946
rect 1104 97872 8832 97894
rect 1104 97402 8832 97424
rect 1104 97350 4315 97402
rect 4367 97350 4379 97402
rect 4431 97350 4443 97402
rect 4495 97350 4507 97402
rect 4559 97350 7648 97402
rect 7700 97350 7712 97402
rect 7764 97350 7776 97402
rect 7828 97350 7840 97402
rect 7892 97350 8832 97402
rect 1104 97328 8832 97350
rect 1104 96858 8832 96880
rect 1104 96806 2648 96858
rect 2700 96806 2712 96858
rect 2764 96806 2776 96858
rect 2828 96806 2840 96858
rect 2892 96806 5982 96858
rect 6034 96806 6046 96858
rect 6098 96806 6110 96858
rect 6162 96806 6174 96858
rect 6226 96806 8832 96858
rect 1104 96784 8832 96806
rect 1104 96314 8832 96336
rect 1104 96262 4315 96314
rect 4367 96262 4379 96314
rect 4431 96262 4443 96314
rect 4495 96262 4507 96314
rect 4559 96262 7648 96314
rect 7700 96262 7712 96314
rect 7764 96262 7776 96314
rect 7828 96262 7840 96314
rect 7892 96262 8832 96314
rect 1104 96240 8832 96262
rect 1104 95770 8832 95792
rect 1104 95718 2648 95770
rect 2700 95718 2712 95770
rect 2764 95718 2776 95770
rect 2828 95718 2840 95770
rect 2892 95718 5982 95770
rect 6034 95718 6046 95770
rect 6098 95718 6110 95770
rect 6162 95718 6174 95770
rect 6226 95718 8832 95770
rect 1104 95696 8832 95718
rect 1104 95226 8832 95248
rect 1104 95174 4315 95226
rect 4367 95174 4379 95226
rect 4431 95174 4443 95226
rect 4495 95174 4507 95226
rect 4559 95174 7648 95226
rect 7700 95174 7712 95226
rect 7764 95174 7776 95226
rect 7828 95174 7840 95226
rect 7892 95174 8832 95226
rect 1104 95152 8832 95174
rect 1104 94682 8832 94704
rect 1104 94630 2648 94682
rect 2700 94630 2712 94682
rect 2764 94630 2776 94682
rect 2828 94630 2840 94682
rect 2892 94630 5982 94682
rect 6034 94630 6046 94682
rect 6098 94630 6110 94682
rect 6162 94630 6174 94682
rect 6226 94630 8832 94682
rect 1104 94608 8832 94630
rect 1104 94138 8832 94160
rect 1104 94086 4315 94138
rect 4367 94086 4379 94138
rect 4431 94086 4443 94138
rect 4495 94086 4507 94138
rect 4559 94086 7648 94138
rect 7700 94086 7712 94138
rect 7764 94086 7776 94138
rect 7828 94086 7840 94138
rect 7892 94086 8832 94138
rect 1104 94064 8832 94086
rect 1104 93594 8832 93616
rect 1104 93542 2648 93594
rect 2700 93542 2712 93594
rect 2764 93542 2776 93594
rect 2828 93542 2840 93594
rect 2892 93542 5982 93594
rect 6034 93542 6046 93594
rect 6098 93542 6110 93594
rect 6162 93542 6174 93594
rect 6226 93542 8832 93594
rect 1104 93520 8832 93542
rect 1104 93050 8832 93072
rect 1104 92998 4315 93050
rect 4367 92998 4379 93050
rect 4431 92998 4443 93050
rect 4495 92998 4507 93050
rect 4559 92998 7648 93050
rect 7700 92998 7712 93050
rect 7764 92998 7776 93050
rect 7828 92998 7840 93050
rect 7892 92998 8832 93050
rect 1104 92976 8832 92998
rect 1104 92506 8832 92528
rect 1104 92454 2648 92506
rect 2700 92454 2712 92506
rect 2764 92454 2776 92506
rect 2828 92454 2840 92506
rect 2892 92454 5982 92506
rect 6034 92454 6046 92506
rect 6098 92454 6110 92506
rect 6162 92454 6174 92506
rect 6226 92454 8832 92506
rect 1104 92432 8832 92454
rect 1104 91962 8832 91984
rect 1104 91910 4315 91962
rect 4367 91910 4379 91962
rect 4431 91910 4443 91962
rect 4495 91910 4507 91962
rect 4559 91910 7648 91962
rect 7700 91910 7712 91962
rect 7764 91910 7776 91962
rect 7828 91910 7840 91962
rect 7892 91910 8832 91962
rect 1104 91888 8832 91910
rect 1104 91418 8832 91440
rect 1104 91366 2648 91418
rect 2700 91366 2712 91418
rect 2764 91366 2776 91418
rect 2828 91366 2840 91418
rect 2892 91366 5982 91418
rect 6034 91366 6046 91418
rect 6098 91366 6110 91418
rect 6162 91366 6174 91418
rect 6226 91366 8832 91418
rect 1104 91344 8832 91366
rect 1104 90874 8832 90896
rect 1104 90822 4315 90874
rect 4367 90822 4379 90874
rect 4431 90822 4443 90874
rect 4495 90822 4507 90874
rect 4559 90822 7648 90874
rect 7700 90822 7712 90874
rect 7764 90822 7776 90874
rect 7828 90822 7840 90874
rect 7892 90822 8832 90874
rect 1104 90800 8832 90822
rect 1104 90330 8832 90352
rect 1104 90278 2648 90330
rect 2700 90278 2712 90330
rect 2764 90278 2776 90330
rect 2828 90278 2840 90330
rect 2892 90278 5982 90330
rect 6034 90278 6046 90330
rect 6098 90278 6110 90330
rect 6162 90278 6174 90330
rect 6226 90278 8832 90330
rect 1104 90256 8832 90278
rect 1104 89786 8832 89808
rect 1104 89734 4315 89786
rect 4367 89734 4379 89786
rect 4431 89734 4443 89786
rect 4495 89734 4507 89786
rect 4559 89734 7648 89786
rect 7700 89734 7712 89786
rect 7764 89734 7776 89786
rect 7828 89734 7840 89786
rect 7892 89734 8832 89786
rect 1104 89712 8832 89734
rect 1104 89242 8832 89264
rect 1104 89190 2648 89242
rect 2700 89190 2712 89242
rect 2764 89190 2776 89242
rect 2828 89190 2840 89242
rect 2892 89190 5982 89242
rect 6034 89190 6046 89242
rect 6098 89190 6110 89242
rect 6162 89190 6174 89242
rect 6226 89190 8832 89242
rect 1104 89168 8832 89190
rect 1104 88698 8832 88720
rect 1104 88646 4315 88698
rect 4367 88646 4379 88698
rect 4431 88646 4443 88698
rect 4495 88646 4507 88698
rect 4559 88646 7648 88698
rect 7700 88646 7712 88698
rect 7764 88646 7776 88698
rect 7828 88646 7840 88698
rect 7892 88646 8832 88698
rect 1104 88624 8832 88646
rect 1104 88154 8832 88176
rect 1104 88102 2648 88154
rect 2700 88102 2712 88154
rect 2764 88102 2776 88154
rect 2828 88102 2840 88154
rect 2892 88102 5982 88154
rect 6034 88102 6046 88154
rect 6098 88102 6110 88154
rect 6162 88102 6174 88154
rect 6226 88102 8832 88154
rect 1104 88080 8832 88102
rect 1104 87610 8832 87632
rect 1104 87558 4315 87610
rect 4367 87558 4379 87610
rect 4431 87558 4443 87610
rect 4495 87558 4507 87610
rect 4559 87558 7648 87610
rect 7700 87558 7712 87610
rect 7764 87558 7776 87610
rect 7828 87558 7840 87610
rect 7892 87558 8832 87610
rect 1104 87536 8832 87558
rect 1104 87066 8832 87088
rect 1104 87014 2648 87066
rect 2700 87014 2712 87066
rect 2764 87014 2776 87066
rect 2828 87014 2840 87066
rect 2892 87014 5982 87066
rect 6034 87014 6046 87066
rect 6098 87014 6110 87066
rect 6162 87014 6174 87066
rect 6226 87014 8832 87066
rect 1104 86992 8832 87014
rect 1104 86522 8832 86544
rect 1104 86470 4315 86522
rect 4367 86470 4379 86522
rect 4431 86470 4443 86522
rect 4495 86470 4507 86522
rect 4559 86470 7648 86522
rect 7700 86470 7712 86522
rect 7764 86470 7776 86522
rect 7828 86470 7840 86522
rect 7892 86470 8832 86522
rect 1104 86448 8832 86470
rect 1104 85978 8832 86000
rect 1104 85926 2648 85978
rect 2700 85926 2712 85978
rect 2764 85926 2776 85978
rect 2828 85926 2840 85978
rect 2892 85926 5982 85978
rect 6034 85926 6046 85978
rect 6098 85926 6110 85978
rect 6162 85926 6174 85978
rect 6226 85926 8832 85978
rect 1104 85904 8832 85926
rect 1104 85434 8832 85456
rect 1104 85382 4315 85434
rect 4367 85382 4379 85434
rect 4431 85382 4443 85434
rect 4495 85382 4507 85434
rect 4559 85382 7648 85434
rect 7700 85382 7712 85434
rect 7764 85382 7776 85434
rect 7828 85382 7840 85434
rect 7892 85382 8832 85434
rect 1104 85360 8832 85382
rect 1104 84890 8832 84912
rect 1104 84838 2648 84890
rect 2700 84838 2712 84890
rect 2764 84838 2776 84890
rect 2828 84838 2840 84890
rect 2892 84838 5982 84890
rect 6034 84838 6046 84890
rect 6098 84838 6110 84890
rect 6162 84838 6174 84890
rect 6226 84838 8832 84890
rect 1104 84816 8832 84838
rect 1104 84346 8832 84368
rect 1104 84294 4315 84346
rect 4367 84294 4379 84346
rect 4431 84294 4443 84346
rect 4495 84294 4507 84346
rect 4559 84294 7648 84346
rect 7700 84294 7712 84346
rect 7764 84294 7776 84346
rect 7828 84294 7840 84346
rect 7892 84294 8832 84346
rect 1104 84272 8832 84294
rect 1104 83802 8832 83824
rect 1104 83750 2648 83802
rect 2700 83750 2712 83802
rect 2764 83750 2776 83802
rect 2828 83750 2840 83802
rect 2892 83750 5982 83802
rect 6034 83750 6046 83802
rect 6098 83750 6110 83802
rect 6162 83750 6174 83802
rect 6226 83750 8832 83802
rect 1104 83728 8832 83750
rect 1104 83258 8832 83280
rect 1104 83206 4315 83258
rect 4367 83206 4379 83258
rect 4431 83206 4443 83258
rect 4495 83206 4507 83258
rect 4559 83206 7648 83258
rect 7700 83206 7712 83258
rect 7764 83206 7776 83258
rect 7828 83206 7840 83258
rect 7892 83206 8832 83258
rect 1104 83184 8832 83206
rect 1104 82714 8832 82736
rect 1104 82662 2648 82714
rect 2700 82662 2712 82714
rect 2764 82662 2776 82714
rect 2828 82662 2840 82714
rect 2892 82662 5982 82714
rect 6034 82662 6046 82714
rect 6098 82662 6110 82714
rect 6162 82662 6174 82714
rect 6226 82662 8832 82714
rect 1104 82640 8832 82662
rect 1104 82170 8832 82192
rect 1104 82118 4315 82170
rect 4367 82118 4379 82170
rect 4431 82118 4443 82170
rect 4495 82118 4507 82170
rect 4559 82118 7648 82170
rect 7700 82118 7712 82170
rect 7764 82118 7776 82170
rect 7828 82118 7840 82170
rect 7892 82118 8832 82170
rect 1104 82096 8832 82118
rect 1104 81626 8832 81648
rect 1104 81574 2648 81626
rect 2700 81574 2712 81626
rect 2764 81574 2776 81626
rect 2828 81574 2840 81626
rect 2892 81574 5982 81626
rect 6034 81574 6046 81626
rect 6098 81574 6110 81626
rect 6162 81574 6174 81626
rect 6226 81574 8832 81626
rect 1104 81552 8832 81574
rect 1104 81082 8832 81104
rect 1104 81030 4315 81082
rect 4367 81030 4379 81082
rect 4431 81030 4443 81082
rect 4495 81030 4507 81082
rect 4559 81030 7648 81082
rect 7700 81030 7712 81082
rect 7764 81030 7776 81082
rect 7828 81030 7840 81082
rect 7892 81030 8832 81082
rect 1104 81008 8832 81030
rect 1104 80538 8832 80560
rect 1104 80486 2648 80538
rect 2700 80486 2712 80538
rect 2764 80486 2776 80538
rect 2828 80486 2840 80538
rect 2892 80486 5982 80538
rect 6034 80486 6046 80538
rect 6098 80486 6110 80538
rect 6162 80486 6174 80538
rect 6226 80486 8832 80538
rect 1104 80464 8832 80486
rect 1104 79994 8832 80016
rect 1104 79942 4315 79994
rect 4367 79942 4379 79994
rect 4431 79942 4443 79994
rect 4495 79942 4507 79994
rect 4559 79942 7648 79994
rect 7700 79942 7712 79994
rect 7764 79942 7776 79994
rect 7828 79942 7840 79994
rect 7892 79942 8832 79994
rect 1104 79920 8832 79942
rect 1104 79450 8832 79472
rect 1104 79398 2648 79450
rect 2700 79398 2712 79450
rect 2764 79398 2776 79450
rect 2828 79398 2840 79450
rect 2892 79398 5982 79450
rect 6034 79398 6046 79450
rect 6098 79398 6110 79450
rect 6162 79398 6174 79450
rect 6226 79398 8832 79450
rect 1104 79376 8832 79398
rect 1104 78906 8832 78928
rect 1104 78854 4315 78906
rect 4367 78854 4379 78906
rect 4431 78854 4443 78906
rect 4495 78854 4507 78906
rect 4559 78854 7648 78906
rect 7700 78854 7712 78906
rect 7764 78854 7776 78906
rect 7828 78854 7840 78906
rect 7892 78854 8832 78906
rect 1104 78832 8832 78854
rect 1104 78362 8832 78384
rect 1104 78310 2648 78362
rect 2700 78310 2712 78362
rect 2764 78310 2776 78362
rect 2828 78310 2840 78362
rect 2892 78310 5982 78362
rect 6034 78310 6046 78362
rect 6098 78310 6110 78362
rect 6162 78310 6174 78362
rect 6226 78310 8832 78362
rect 1104 78288 8832 78310
rect 1104 77818 8832 77840
rect 1104 77766 4315 77818
rect 4367 77766 4379 77818
rect 4431 77766 4443 77818
rect 4495 77766 4507 77818
rect 4559 77766 7648 77818
rect 7700 77766 7712 77818
rect 7764 77766 7776 77818
rect 7828 77766 7840 77818
rect 7892 77766 8832 77818
rect 1104 77744 8832 77766
rect 1104 77274 8832 77296
rect 1104 77222 2648 77274
rect 2700 77222 2712 77274
rect 2764 77222 2776 77274
rect 2828 77222 2840 77274
rect 2892 77222 5982 77274
rect 6034 77222 6046 77274
rect 6098 77222 6110 77274
rect 6162 77222 6174 77274
rect 6226 77222 8832 77274
rect 1104 77200 8832 77222
rect 1104 76730 8832 76752
rect 1104 76678 4315 76730
rect 4367 76678 4379 76730
rect 4431 76678 4443 76730
rect 4495 76678 4507 76730
rect 4559 76678 7648 76730
rect 7700 76678 7712 76730
rect 7764 76678 7776 76730
rect 7828 76678 7840 76730
rect 7892 76678 8832 76730
rect 1104 76656 8832 76678
rect 1104 76186 8832 76208
rect 1104 76134 2648 76186
rect 2700 76134 2712 76186
rect 2764 76134 2776 76186
rect 2828 76134 2840 76186
rect 2892 76134 5982 76186
rect 6034 76134 6046 76186
rect 6098 76134 6110 76186
rect 6162 76134 6174 76186
rect 6226 76134 8832 76186
rect 1104 76112 8832 76134
rect 1104 75642 8832 75664
rect 1104 75590 4315 75642
rect 4367 75590 4379 75642
rect 4431 75590 4443 75642
rect 4495 75590 4507 75642
rect 4559 75590 7648 75642
rect 7700 75590 7712 75642
rect 7764 75590 7776 75642
rect 7828 75590 7840 75642
rect 7892 75590 8832 75642
rect 1104 75568 8832 75590
rect 1104 75098 8832 75120
rect 1104 75046 2648 75098
rect 2700 75046 2712 75098
rect 2764 75046 2776 75098
rect 2828 75046 2840 75098
rect 2892 75046 5982 75098
rect 6034 75046 6046 75098
rect 6098 75046 6110 75098
rect 6162 75046 6174 75098
rect 6226 75046 8832 75098
rect 1104 75024 8832 75046
rect 1104 74554 8832 74576
rect 1104 74502 4315 74554
rect 4367 74502 4379 74554
rect 4431 74502 4443 74554
rect 4495 74502 4507 74554
rect 4559 74502 7648 74554
rect 7700 74502 7712 74554
rect 7764 74502 7776 74554
rect 7828 74502 7840 74554
rect 7892 74502 8832 74554
rect 1104 74480 8832 74502
rect 1104 74010 8832 74032
rect 1104 73958 2648 74010
rect 2700 73958 2712 74010
rect 2764 73958 2776 74010
rect 2828 73958 2840 74010
rect 2892 73958 5982 74010
rect 6034 73958 6046 74010
rect 6098 73958 6110 74010
rect 6162 73958 6174 74010
rect 6226 73958 8832 74010
rect 1104 73936 8832 73958
rect 1104 73466 8832 73488
rect 1104 73414 4315 73466
rect 4367 73414 4379 73466
rect 4431 73414 4443 73466
rect 4495 73414 4507 73466
rect 4559 73414 7648 73466
rect 7700 73414 7712 73466
rect 7764 73414 7776 73466
rect 7828 73414 7840 73466
rect 7892 73414 8832 73466
rect 1104 73392 8832 73414
rect 1104 72922 8832 72944
rect 1104 72870 2648 72922
rect 2700 72870 2712 72922
rect 2764 72870 2776 72922
rect 2828 72870 2840 72922
rect 2892 72870 5982 72922
rect 6034 72870 6046 72922
rect 6098 72870 6110 72922
rect 6162 72870 6174 72922
rect 6226 72870 8832 72922
rect 1104 72848 8832 72870
rect 1104 72378 8832 72400
rect 1104 72326 4315 72378
rect 4367 72326 4379 72378
rect 4431 72326 4443 72378
rect 4495 72326 4507 72378
rect 4559 72326 7648 72378
rect 7700 72326 7712 72378
rect 7764 72326 7776 72378
rect 7828 72326 7840 72378
rect 7892 72326 8832 72378
rect 1104 72304 8832 72326
rect 106 72020 112 72072
rect 164 72060 170 72072
rect 5626 72060 5632 72072
rect 164 72032 5632 72060
rect 164 72020 170 72032
rect 5626 72020 5632 72032
rect 5684 72020 5690 72072
rect 5626 71884 5632 71936
rect 5684 71924 5690 71936
rect 6730 71924 6736 71936
rect 5684 71896 6736 71924
rect 5684 71884 5690 71896
rect 6730 71884 6736 71896
rect 6788 71884 6794 71936
rect 1104 71834 8832 71856
rect 1104 71782 2648 71834
rect 2700 71782 2712 71834
rect 2764 71782 2776 71834
rect 2828 71782 2840 71834
rect 2892 71782 5982 71834
rect 6034 71782 6046 71834
rect 6098 71782 6110 71834
rect 6162 71782 6174 71834
rect 6226 71782 8832 71834
rect 1104 71760 8832 71782
rect 1104 71290 8832 71312
rect 1104 71238 4315 71290
rect 4367 71238 4379 71290
rect 4431 71238 4443 71290
rect 4495 71238 4507 71290
rect 4559 71238 7648 71290
rect 7700 71238 7712 71290
rect 7764 71238 7776 71290
rect 7828 71238 7840 71290
rect 7892 71238 8832 71290
rect 1104 71216 8832 71238
rect 1104 70746 8832 70768
rect 1104 70694 2648 70746
rect 2700 70694 2712 70746
rect 2764 70694 2776 70746
rect 2828 70694 2840 70746
rect 2892 70694 5982 70746
rect 6034 70694 6046 70746
rect 6098 70694 6110 70746
rect 6162 70694 6174 70746
rect 6226 70694 8832 70746
rect 1104 70672 8832 70694
rect 1104 70202 8832 70224
rect 1104 70150 4315 70202
rect 4367 70150 4379 70202
rect 4431 70150 4443 70202
rect 4495 70150 4507 70202
rect 4559 70150 7648 70202
rect 7700 70150 7712 70202
rect 7764 70150 7776 70202
rect 7828 70150 7840 70202
rect 7892 70150 8832 70202
rect 1104 70128 8832 70150
rect 1104 69658 8832 69680
rect 1104 69606 2648 69658
rect 2700 69606 2712 69658
rect 2764 69606 2776 69658
rect 2828 69606 2840 69658
rect 2892 69606 5982 69658
rect 6034 69606 6046 69658
rect 6098 69606 6110 69658
rect 6162 69606 6174 69658
rect 6226 69606 8832 69658
rect 1104 69584 8832 69606
rect 1104 69114 8832 69136
rect 1104 69062 4315 69114
rect 4367 69062 4379 69114
rect 4431 69062 4443 69114
rect 4495 69062 4507 69114
rect 4559 69062 7648 69114
rect 7700 69062 7712 69114
rect 7764 69062 7776 69114
rect 7828 69062 7840 69114
rect 7892 69062 8832 69114
rect 1104 69040 8832 69062
rect 1104 68570 8832 68592
rect 1104 68518 2648 68570
rect 2700 68518 2712 68570
rect 2764 68518 2776 68570
rect 2828 68518 2840 68570
rect 2892 68518 5982 68570
rect 6034 68518 6046 68570
rect 6098 68518 6110 68570
rect 6162 68518 6174 68570
rect 6226 68518 8832 68570
rect 1104 68496 8832 68518
rect 1104 68026 8832 68048
rect 1104 67974 4315 68026
rect 4367 67974 4379 68026
rect 4431 67974 4443 68026
rect 4495 67974 4507 68026
rect 4559 67974 7648 68026
rect 7700 67974 7712 68026
rect 7764 67974 7776 68026
rect 7828 67974 7840 68026
rect 7892 67974 8832 68026
rect 1104 67952 8832 67974
rect 1104 67482 8832 67504
rect 1104 67430 2648 67482
rect 2700 67430 2712 67482
rect 2764 67430 2776 67482
rect 2828 67430 2840 67482
rect 2892 67430 5982 67482
rect 6034 67430 6046 67482
rect 6098 67430 6110 67482
rect 6162 67430 6174 67482
rect 6226 67430 8832 67482
rect 1104 67408 8832 67430
rect 1104 66938 8832 66960
rect 1104 66886 4315 66938
rect 4367 66886 4379 66938
rect 4431 66886 4443 66938
rect 4495 66886 4507 66938
rect 4559 66886 7648 66938
rect 7700 66886 7712 66938
rect 7764 66886 7776 66938
rect 7828 66886 7840 66938
rect 7892 66886 8832 66938
rect 1104 66864 8832 66886
rect 1104 66394 8832 66416
rect 1104 66342 2648 66394
rect 2700 66342 2712 66394
rect 2764 66342 2776 66394
rect 2828 66342 2840 66394
rect 2892 66342 5982 66394
rect 6034 66342 6046 66394
rect 6098 66342 6110 66394
rect 6162 66342 6174 66394
rect 6226 66342 8832 66394
rect 1104 66320 8832 66342
rect 1104 65850 8832 65872
rect 1104 65798 4315 65850
rect 4367 65798 4379 65850
rect 4431 65798 4443 65850
rect 4495 65798 4507 65850
rect 4559 65798 7648 65850
rect 7700 65798 7712 65850
rect 7764 65798 7776 65850
rect 7828 65798 7840 65850
rect 7892 65798 8832 65850
rect 1104 65776 8832 65798
rect 1104 65306 8832 65328
rect 1104 65254 2648 65306
rect 2700 65254 2712 65306
rect 2764 65254 2776 65306
rect 2828 65254 2840 65306
rect 2892 65254 5982 65306
rect 6034 65254 6046 65306
rect 6098 65254 6110 65306
rect 6162 65254 6174 65306
rect 6226 65254 8832 65306
rect 1104 65232 8832 65254
rect 1104 64762 8832 64784
rect 1104 64710 4315 64762
rect 4367 64710 4379 64762
rect 4431 64710 4443 64762
rect 4495 64710 4507 64762
rect 4559 64710 7648 64762
rect 7700 64710 7712 64762
rect 7764 64710 7776 64762
rect 7828 64710 7840 64762
rect 7892 64710 8832 64762
rect 1104 64688 8832 64710
rect 1104 64218 8832 64240
rect 1104 64166 2648 64218
rect 2700 64166 2712 64218
rect 2764 64166 2776 64218
rect 2828 64166 2840 64218
rect 2892 64166 5982 64218
rect 6034 64166 6046 64218
rect 6098 64166 6110 64218
rect 6162 64166 6174 64218
rect 6226 64166 8832 64218
rect 1104 64144 8832 64166
rect 1104 63674 8832 63696
rect 1104 63622 4315 63674
rect 4367 63622 4379 63674
rect 4431 63622 4443 63674
rect 4495 63622 4507 63674
rect 4559 63622 7648 63674
rect 7700 63622 7712 63674
rect 7764 63622 7776 63674
rect 7828 63622 7840 63674
rect 7892 63622 8832 63674
rect 1104 63600 8832 63622
rect 1104 63130 8832 63152
rect 1104 63078 2648 63130
rect 2700 63078 2712 63130
rect 2764 63078 2776 63130
rect 2828 63078 2840 63130
rect 2892 63078 5982 63130
rect 6034 63078 6046 63130
rect 6098 63078 6110 63130
rect 6162 63078 6174 63130
rect 6226 63078 8832 63130
rect 1104 63056 8832 63078
rect 1104 62586 8832 62608
rect 1104 62534 4315 62586
rect 4367 62534 4379 62586
rect 4431 62534 4443 62586
rect 4495 62534 4507 62586
rect 4559 62534 7648 62586
rect 7700 62534 7712 62586
rect 7764 62534 7776 62586
rect 7828 62534 7840 62586
rect 7892 62534 8832 62586
rect 1104 62512 8832 62534
rect 1104 62042 8832 62064
rect 1104 61990 2648 62042
rect 2700 61990 2712 62042
rect 2764 61990 2776 62042
rect 2828 61990 2840 62042
rect 2892 61990 5982 62042
rect 6034 61990 6046 62042
rect 6098 61990 6110 62042
rect 6162 61990 6174 62042
rect 6226 61990 8832 62042
rect 1104 61968 8832 61990
rect 1104 61498 8832 61520
rect 1104 61446 4315 61498
rect 4367 61446 4379 61498
rect 4431 61446 4443 61498
rect 4495 61446 4507 61498
rect 4559 61446 7648 61498
rect 7700 61446 7712 61498
rect 7764 61446 7776 61498
rect 7828 61446 7840 61498
rect 7892 61446 8832 61498
rect 1104 61424 8832 61446
rect 1104 60954 8832 60976
rect 1104 60902 2648 60954
rect 2700 60902 2712 60954
rect 2764 60902 2776 60954
rect 2828 60902 2840 60954
rect 2892 60902 5982 60954
rect 6034 60902 6046 60954
rect 6098 60902 6110 60954
rect 6162 60902 6174 60954
rect 6226 60902 8832 60954
rect 1104 60880 8832 60902
rect 1104 60410 8832 60432
rect 1104 60358 4315 60410
rect 4367 60358 4379 60410
rect 4431 60358 4443 60410
rect 4495 60358 4507 60410
rect 4559 60358 7648 60410
rect 7700 60358 7712 60410
rect 7764 60358 7776 60410
rect 7828 60358 7840 60410
rect 7892 60358 8832 60410
rect 1104 60336 8832 60358
rect 1104 59866 8832 59888
rect 1104 59814 2648 59866
rect 2700 59814 2712 59866
rect 2764 59814 2776 59866
rect 2828 59814 2840 59866
rect 2892 59814 5982 59866
rect 6034 59814 6046 59866
rect 6098 59814 6110 59866
rect 6162 59814 6174 59866
rect 6226 59814 8832 59866
rect 1104 59792 8832 59814
rect 1104 59322 8832 59344
rect 1104 59270 4315 59322
rect 4367 59270 4379 59322
rect 4431 59270 4443 59322
rect 4495 59270 4507 59322
rect 4559 59270 7648 59322
rect 7700 59270 7712 59322
rect 7764 59270 7776 59322
rect 7828 59270 7840 59322
rect 7892 59270 8832 59322
rect 1104 59248 8832 59270
rect 1104 58778 8832 58800
rect 1104 58726 2648 58778
rect 2700 58726 2712 58778
rect 2764 58726 2776 58778
rect 2828 58726 2840 58778
rect 2892 58726 5982 58778
rect 6034 58726 6046 58778
rect 6098 58726 6110 58778
rect 6162 58726 6174 58778
rect 6226 58726 8832 58778
rect 1104 58704 8832 58726
rect 1104 58234 8832 58256
rect 1104 58182 4315 58234
rect 4367 58182 4379 58234
rect 4431 58182 4443 58234
rect 4495 58182 4507 58234
rect 4559 58182 7648 58234
rect 7700 58182 7712 58234
rect 7764 58182 7776 58234
rect 7828 58182 7840 58234
rect 7892 58182 8832 58234
rect 1104 58160 8832 58182
rect 1104 57690 8832 57712
rect 1104 57638 2648 57690
rect 2700 57638 2712 57690
rect 2764 57638 2776 57690
rect 2828 57638 2840 57690
rect 2892 57638 5982 57690
rect 6034 57638 6046 57690
rect 6098 57638 6110 57690
rect 6162 57638 6174 57690
rect 6226 57638 8832 57690
rect 1104 57616 8832 57638
rect 1104 57146 8832 57168
rect 1104 57094 4315 57146
rect 4367 57094 4379 57146
rect 4431 57094 4443 57146
rect 4495 57094 4507 57146
rect 4559 57094 7648 57146
rect 7700 57094 7712 57146
rect 7764 57094 7776 57146
rect 7828 57094 7840 57146
rect 7892 57094 8832 57146
rect 1104 57072 8832 57094
rect 1104 56602 8832 56624
rect 1104 56550 2648 56602
rect 2700 56550 2712 56602
rect 2764 56550 2776 56602
rect 2828 56550 2840 56602
rect 2892 56550 5982 56602
rect 6034 56550 6046 56602
rect 6098 56550 6110 56602
rect 6162 56550 6174 56602
rect 6226 56550 8832 56602
rect 1104 56528 8832 56550
rect 1104 56058 8832 56080
rect 1104 56006 4315 56058
rect 4367 56006 4379 56058
rect 4431 56006 4443 56058
rect 4495 56006 4507 56058
rect 4559 56006 7648 56058
rect 7700 56006 7712 56058
rect 7764 56006 7776 56058
rect 7828 56006 7840 56058
rect 7892 56006 8832 56058
rect 1104 55984 8832 56006
rect 1104 55514 8832 55536
rect 1104 55462 2648 55514
rect 2700 55462 2712 55514
rect 2764 55462 2776 55514
rect 2828 55462 2840 55514
rect 2892 55462 5982 55514
rect 6034 55462 6046 55514
rect 6098 55462 6110 55514
rect 6162 55462 6174 55514
rect 6226 55462 8832 55514
rect 1104 55440 8832 55462
rect 1104 54970 8832 54992
rect 1104 54918 4315 54970
rect 4367 54918 4379 54970
rect 4431 54918 4443 54970
rect 4495 54918 4507 54970
rect 4559 54918 7648 54970
rect 7700 54918 7712 54970
rect 7764 54918 7776 54970
rect 7828 54918 7840 54970
rect 7892 54918 8832 54970
rect 1104 54896 8832 54918
rect 1104 54426 8832 54448
rect 1104 54374 2648 54426
rect 2700 54374 2712 54426
rect 2764 54374 2776 54426
rect 2828 54374 2840 54426
rect 2892 54374 5982 54426
rect 6034 54374 6046 54426
rect 6098 54374 6110 54426
rect 6162 54374 6174 54426
rect 6226 54374 8832 54426
rect 1104 54352 8832 54374
rect 1104 53882 8832 53904
rect 1104 53830 4315 53882
rect 4367 53830 4379 53882
rect 4431 53830 4443 53882
rect 4495 53830 4507 53882
rect 4559 53830 7648 53882
rect 7700 53830 7712 53882
rect 7764 53830 7776 53882
rect 7828 53830 7840 53882
rect 7892 53830 8832 53882
rect 1104 53808 8832 53830
rect 1104 53338 8832 53360
rect 1104 53286 2648 53338
rect 2700 53286 2712 53338
rect 2764 53286 2776 53338
rect 2828 53286 2840 53338
rect 2892 53286 5982 53338
rect 6034 53286 6046 53338
rect 6098 53286 6110 53338
rect 6162 53286 6174 53338
rect 6226 53286 8832 53338
rect 1104 53264 8832 53286
rect 1104 52794 8832 52816
rect 1104 52742 4315 52794
rect 4367 52742 4379 52794
rect 4431 52742 4443 52794
rect 4495 52742 4507 52794
rect 4559 52742 7648 52794
rect 7700 52742 7712 52794
rect 7764 52742 7776 52794
rect 7828 52742 7840 52794
rect 7892 52742 8832 52794
rect 1104 52720 8832 52742
rect 1104 52250 8832 52272
rect 1104 52198 2648 52250
rect 2700 52198 2712 52250
rect 2764 52198 2776 52250
rect 2828 52198 2840 52250
rect 2892 52198 5982 52250
rect 6034 52198 6046 52250
rect 6098 52198 6110 52250
rect 6162 52198 6174 52250
rect 6226 52198 8832 52250
rect 1104 52176 8832 52198
rect 1104 51706 8832 51728
rect 1104 51654 4315 51706
rect 4367 51654 4379 51706
rect 4431 51654 4443 51706
rect 4495 51654 4507 51706
rect 4559 51654 7648 51706
rect 7700 51654 7712 51706
rect 7764 51654 7776 51706
rect 7828 51654 7840 51706
rect 7892 51654 8832 51706
rect 1104 51632 8832 51654
rect 1104 51162 8832 51184
rect 1104 51110 2648 51162
rect 2700 51110 2712 51162
rect 2764 51110 2776 51162
rect 2828 51110 2840 51162
rect 2892 51110 5982 51162
rect 6034 51110 6046 51162
rect 6098 51110 6110 51162
rect 6162 51110 6174 51162
rect 6226 51110 8832 51162
rect 1104 51088 8832 51110
rect 7009 50983 7067 50989
rect 7009 50949 7021 50983
rect 7055 50980 7067 50983
rect 8202 50980 8208 50992
rect 7055 50952 8208 50980
rect 7055 50949 7067 50952
rect 7009 50943 7067 50949
rect 8202 50940 8208 50952
rect 8260 50940 8266 50992
rect 6730 50804 6736 50856
rect 6788 50844 6794 50856
rect 6825 50847 6883 50853
rect 6825 50844 6837 50847
rect 6788 50816 6837 50844
rect 6788 50804 6794 50816
rect 6825 50813 6837 50816
rect 6871 50844 6883 50847
rect 7377 50847 7435 50853
rect 7377 50844 7389 50847
rect 6871 50816 7389 50844
rect 6871 50813 6883 50816
rect 6825 50807 6883 50813
rect 7377 50813 7389 50816
rect 7423 50813 7435 50847
rect 7377 50807 7435 50813
rect 1104 50618 8832 50640
rect 1104 50566 4315 50618
rect 4367 50566 4379 50618
rect 4431 50566 4443 50618
rect 4495 50566 4507 50618
rect 4559 50566 7648 50618
rect 7700 50566 7712 50618
rect 7764 50566 7776 50618
rect 7828 50566 7840 50618
rect 7892 50566 8832 50618
rect 1104 50544 8832 50566
rect 1104 50074 8832 50096
rect 1104 50022 2648 50074
rect 2700 50022 2712 50074
rect 2764 50022 2776 50074
rect 2828 50022 2840 50074
rect 2892 50022 5982 50074
rect 6034 50022 6046 50074
rect 6098 50022 6110 50074
rect 6162 50022 6174 50074
rect 6226 50022 8832 50074
rect 1104 50000 8832 50022
rect 1104 49530 8832 49552
rect 1104 49478 4315 49530
rect 4367 49478 4379 49530
rect 4431 49478 4443 49530
rect 4495 49478 4507 49530
rect 4559 49478 7648 49530
rect 7700 49478 7712 49530
rect 7764 49478 7776 49530
rect 7828 49478 7840 49530
rect 7892 49478 8832 49530
rect 1104 49456 8832 49478
rect 1104 48986 8832 49008
rect 1104 48934 2648 48986
rect 2700 48934 2712 48986
rect 2764 48934 2776 48986
rect 2828 48934 2840 48986
rect 2892 48934 5982 48986
rect 6034 48934 6046 48986
rect 6098 48934 6110 48986
rect 6162 48934 6174 48986
rect 6226 48934 8832 48986
rect 1104 48912 8832 48934
rect 1104 48442 8832 48464
rect 1104 48390 4315 48442
rect 4367 48390 4379 48442
rect 4431 48390 4443 48442
rect 4495 48390 4507 48442
rect 4559 48390 7648 48442
rect 7700 48390 7712 48442
rect 7764 48390 7776 48442
rect 7828 48390 7840 48442
rect 7892 48390 8832 48442
rect 1104 48368 8832 48390
rect 1104 47898 8832 47920
rect 1104 47846 2648 47898
rect 2700 47846 2712 47898
rect 2764 47846 2776 47898
rect 2828 47846 2840 47898
rect 2892 47846 5982 47898
rect 6034 47846 6046 47898
rect 6098 47846 6110 47898
rect 6162 47846 6174 47898
rect 6226 47846 8832 47898
rect 1104 47824 8832 47846
rect 1104 47354 8832 47376
rect 1104 47302 4315 47354
rect 4367 47302 4379 47354
rect 4431 47302 4443 47354
rect 4495 47302 4507 47354
rect 4559 47302 7648 47354
rect 7700 47302 7712 47354
rect 7764 47302 7776 47354
rect 7828 47302 7840 47354
rect 7892 47302 8832 47354
rect 1104 47280 8832 47302
rect 1104 46810 8832 46832
rect 1104 46758 2648 46810
rect 2700 46758 2712 46810
rect 2764 46758 2776 46810
rect 2828 46758 2840 46810
rect 2892 46758 5982 46810
rect 6034 46758 6046 46810
rect 6098 46758 6110 46810
rect 6162 46758 6174 46810
rect 6226 46758 8832 46810
rect 1104 46736 8832 46758
rect 1104 46266 8832 46288
rect 1104 46214 4315 46266
rect 4367 46214 4379 46266
rect 4431 46214 4443 46266
rect 4495 46214 4507 46266
rect 4559 46214 7648 46266
rect 7700 46214 7712 46266
rect 7764 46214 7776 46266
rect 7828 46214 7840 46266
rect 7892 46214 8832 46266
rect 1104 46192 8832 46214
rect 1104 45722 8832 45744
rect 1104 45670 2648 45722
rect 2700 45670 2712 45722
rect 2764 45670 2776 45722
rect 2828 45670 2840 45722
rect 2892 45670 5982 45722
rect 6034 45670 6046 45722
rect 6098 45670 6110 45722
rect 6162 45670 6174 45722
rect 6226 45670 8832 45722
rect 1104 45648 8832 45670
rect 1104 45178 8832 45200
rect 1104 45126 4315 45178
rect 4367 45126 4379 45178
rect 4431 45126 4443 45178
rect 4495 45126 4507 45178
rect 4559 45126 7648 45178
rect 7700 45126 7712 45178
rect 7764 45126 7776 45178
rect 7828 45126 7840 45178
rect 7892 45126 8832 45178
rect 1104 45104 8832 45126
rect 1104 44634 8832 44656
rect 1104 44582 2648 44634
rect 2700 44582 2712 44634
rect 2764 44582 2776 44634
rect 2828 44582 2840 44634
rect 2892 44582 5982 44634
rect 6034 44582 6046 44634
rect 6098 44582 6110 44634
rect 6162 44582 6174 44634
rect 6226 44582 8832 44634
rect 1104 44560 8832 44582
rect 1104 44090 8832 44112
rect 1104 44038 4315 44090
rect 4367 44038 4379 44090
rect 4431 44038 4443 44090
rect 4495 44038 4507 44090
rect 4559 44038 7648 44090
rect 7700 44038 7712 44090
rect 7764 44038 7776 44090
rect 7828 44038 7840 44090
rect 7892 44038 8832 44090
rect 1104 44016 8832 44038
rect 1104 43546 8832 43568
rect 1104 43494 2648 43546
rect 2700 43494 2712 43546
rect 2764 43494 2776 43546
rect 2828 43494 2840 43546
rect 2892 43494 5982 43546
rect 6034 43494 6046 43546
rect 6098 43494 6110 43546
rect 6162 43494 6174 43546
rect 6226 43494 8832 43546
rect 1104 43472 8832 43494
rect 1104 43002 8832 43024
rect 1104 42950 4315 43002
rect 4367 42950 4379 43002
rect 4431 42950 4443 43002
rect 4495 42950 4507 43002
rect 4559 42950 7648 43002
rect 7700 42950 7712 43002
rect 7764 42950 7776 43002
rect 7828 42950 7840 43002
rect 7892 42950 8832 43002
rect 1104 42928 8832 42950
rect 1104 42458 8832 42480
rect 1104 42406 2648 42458
rect 2700 42406 2712 42458
rect 2764 42406 2776 42458
rect 2828 42406 2840 42458
rect 2892 42406 5982 42458
rect 6034 42406 6046 42458
rect 6098 42406 6110 42458
rect 6162 42406 6174 42458
rect 6226 42406 8832 42458
rect 1104 42384 8832 42406
rect 1104 41914 8832 41936
rect 1104 41862 4315 41914
rect 4367 41862 4379 41914
rect 4431 41862 4443 41914
rect 4495 41862 4507 41914
rect 4559 41862 7648 41914
rect 7700 41862 7712 41914
rect 7764 41862 7776 41914
rect 7828 41862 7840 41914
rect 7892 41862 8832 41914
rect 1104 41840 8832 41862
rect 1104 41370 8832 41392
rect 1104 41318 2648 41370
rect 2700 41318 2712 41370
rect 2764 41318 2776 41370
rect 2828 41318 2840 41370
rect 2892 41318 5982 41370
rect 6034 41318 6046 41370
rect 6098 41318 6110 41370
rect 6162 41318 6174 41370
rect 6226 41318 8832 41370
rect 1104 41296 8832 41318
rect 1104 40826 8832 40848
rect 1104 40774 4315 40826
rect 4367 40774 4379 40826
rect 4431 40774 4443 40826
rect 4495 40774 4507 40826
rect 4559 40774 7648 40826
rect 7700 40774 7712 40826
rect 7764 40774 7776 40826
rect 7828 40774 7840 40826
rect 7892 40774 8832 40826
rect 1104 40752 8832 40774
rect 1104 40282 8832 40304
rect 1104 40230 2648 40282
rect 2700 40230 2712 40282
rect 2764 40230 2776 40282
rect 2828 40230 2840 40282
rect 2892 40230 5982 40282
rect 6034 40230 6046 40282
rect 6098 40230 6110 40282
rect 6162 40230 6174 40282
rect 6226 40230 8832 40282
rect 1104 40208 8832 40230
rect 1104 39738 8832 39760
rect 1104 39686 4315 39738
rect 4367 39686 4379 39738
rect 4431 39686 4443 39738
rect 4495 39686 4507 39738
rect 4559 39686 7648 39738
rect 7700 39686 7712 39738
rect 7764 39686 7776 39738
rect 7828 39686 7840 39738
rect 7892 39686 8832 39738
rect 1104 39664 8832 39686
rect 1104 39194 8832 39216
rect 1104 39142 2648 39194
rect 2700 39142 2712 39194
rect 2764 39142 2776 39194
rect 2828 39142 2840 39194
rect 2892 39142 5982 39194
rect 6034 39142 6046 39194
rect 6098 39142 6110 39194
rect 6162 39142 6174 39194
rect 6226 39142 8832 39194
rect 1104 39120 8832 39142
rect 1104 38650 8832 38672
rect 1104 38598 4315 38650
rect 4367 38598 4379 38650
rect 4431 38598 4443 38650
rect 4495 38598 4507 38650
rect 4559 38598 7648 38650
rect 7700 38598 7712 38650
rect 7764 38598 7776 38650
rect 7828 38598 7840 38650
rect 7892 38598 8832 38650
rect 1104 38576 8832 38598
rect 1104 38106 8832 38128
rect 1104 38054 2648 38106
rect 2700 38054 2712 38106
rect 2764 38054 2776 38106
rect 2828 38054 2840 38106
rect 2892 38054 5982 38106
rect 6034 38054 6046 38106
rect 6098 38054 6110 38106
rect 6162 38054 6174 38106
rect 6226 38054 8832 38106
rect 1104 38032 8832 38054
rect 1104 37562 8832 37584
rect 1104 37510 4315 37562
rect 4367 37510 4379 37562
rect 4431 37510 4443 37562
rect 4495 37510 4507 37562
rect 4559 37510 7648 37562
rect 7700 37510 7712 37562
rect 7764 37510 7776 37562
rect 7828 37510 7840 37562
rect 7892 37510 8832 37562
rect 1104 37488 8832 37510
rect 1104 37018 8832 37040
rect 1104 36966 2648 37018
rect 2700 36966 2712 37018
rect 2764 36966 2776 37018
rect 2828 36966 2840 37018
rect 2892 36966 5982 37018
rect 6034 36966 6046 37018
rect 6098 36966 6110 37018
rect 6162 36966 6174 37018
rect 6226 36966 8832 37018
rect 1104 36944 8832 36966
rect 1104 36474 8832 36496
rect 1104 36422 4315 36474
rect 4367 36422 4379 36474
rect 4431 36422 4443 36474
rect 4495 36422 4507 36474
rect 4559 36422 7648 36474
rect 7700 36422 7712 36474
rect 7764 36422 7776 36474
rect 7828 36422 7840 36474
rect 7892 36422 8832 36474
rect 1104 36400 8832 36422
rect 1104 35930 8832 35952
rect 1104 35878 2648 35930
rect 2700 35878 2712 35930
rect 2764 35878 2776 35930
rect 2828 35878 2840 35930
rect 2892 35878 5982 35930
rect 6034 35878 6046 35930
rect 6098 35878 6110 35930
rect 6162 35878 6174 35930
rect 6226 35878 8832 35930
rect 1104 35856 8832 35878
rect 1104 35386 8832 35408
rect 1104 35334 4315 35386
rect 4367 35334 4379 35386
rect 4431 35334 4443 35386
rect 4495 35334 4507 35386
rect 4559 35334 7648 35386
rect 7700 35334 7712 35386
rect 7764 35334 7776 35386
rect 7828 35334 7840 35386
rect 7892 35334 8832 35386
rect 1104 35312 8832 35334
rect 1104 34842 8832 34864
rect 1104 34790 2648 34842
rect 2700 34790 2712 34842
rect 2764 34790 2776 34842
rect 2828 34790 2840 34842
rect 2892 34790 5982 34842
rect 6034 34790 6046 34842
rect 6098 34790 6110 34842
rect 6162 34790 6174 34842
rect 6226 34790 8832 34842
rect 1104 34768 8832 34790
rect 1104 34298 8832 34320
rect 1104 34246 4315 34298
rect 4367 34246 4379 34298
rect 4431 34246 4443 34298
rect 4495 34246 4507 34298
rect 4559 34246 7648 34298
rect 7700 34246 7712 34298
rect 7764 34246 7776 34298
rect 7828 34246 7840 34298
rect 7892 34246 8832 34298
rect 1104 34224 8832 34246
rect 1104 33754 8832 33776
rect 1104 33702 2648 33754
rect 2700 33702 2712 33754
rect 2764 33702 2776 33754
rect 2828 33702 2840 33754
rect 2892 33702 5982 33754
rect 6034 33702 6046 33754
rect 6098 33702 6110 33754
rect 6162 33702 6174 33754
rect 6226 33702 8832 33754
rect 1104 33680 8832 33702
rect 1104 33210 8832 33232
rect 1104 33158 4315 33210
rect 4367 33158 4379 33210
rect 4431 33158 4443 33210
rect 4495 33158 4507 33210
rect 4559 33158 7648 33210
rect 7700 33158 7712 33210
rect 7764 33158 7776 33210
rect 7828 33158 7840 33210
rect 7892 33158 8832 33210
rect 1104 33136 8832 33158
rect 1104 32666 8832 32688
rect 1104 32614 2648 32666
rect 2700 32614 2712 32666
rect 2764 32614 2776 32666
rect 2828 32614 2840 32666
rect 2892 32614 5982 32666
rect 6034 32614 6046 32666
rect 6098 32614 6110 32666
rect 6162 32614 6174 32666
rect 6226 32614 8832 32666
rect 1104 32592 8832 32614
rect 1104 32122 8832 32144
rect 1104 32070 4315 32122
rect 4367 32070 4379 32122
rect 4431 32070 4443 32122
rect 4495 32070 4507 32122
rect 4559 32070 7648 32122
rect 7700 32070 7712 32122
rect 7764 32070 7776 32122
rect 7828 32070 7840 32122
rect 7892 32070 8832 32122
rect 1104 32048 8832 32070
rect 1104 31578 8832 31600
rect 1104 31526 2648 31578
rect 2700 31526 2712 31578
rect 2764 31526 2776 31578
rect 2828 31526 2840 31578
rect 2892 31526 5982 31578
rect 6034 31526 6046 31578
rect 6098 31526 6110 31578
rect 6162 31526 6174 31578
rect 6226 31526 8832 31578
rect 1104 31504 8832 31526
rect 1104 31034 8832 31056
rect 1104 30982 4315 31034
rect 4367 30982 4379 31034
rect 4431 30982 4443 31034
rect 4495 30982 4507 31034
rect 4559 30982 7648 31034
rect 7700 30982 7712 31034
rect 7764 30982 7776 31034
rect 7828 30982 7840 31034
rect 7892 30982 8832 31034
rect 1104 30960 8832 30982
rect 1104 30490 8832 30512
rect 1104 30438 2648 30490
rect 2700 30438 2712 30490
rect 2764 30438 2776 30490
rect 2828 30438 2840 30490
rect 2892 30438 5982 30490
rect 6034 30438 6046 30490
rect 6098 30438 6110 30490
rect 6162 30438 6174 30490
rect 6226 30438 8832 30490
rect 1104 30416 8832 30438
rect 1104 29946 8832 29968
rect 1104 29894 4315 29946
rect 4367 29894 4379 29946
rect 4431 29894 4443 29946
rect 4495 29894 4507 29946
rect 4559 29894 7648 29946
rect 7700 29894 7712 29946
rect 7764 29894 7776 29946
rect 7828 29894 7840 29946
rect 7892 29894 8832 29946
rect 1104 29872 8832 29894
rect 1104 29402 8832 29424
rect 1104 29350 2648 29402
rect 2700 29350 2712 29402
rect 2764 29350 2776 29402
rect 2828 29350 2840 29402
rect 2892 29350 5982 29402
rect 6034 29350 6046 29402
rect 6098 29350 6110 29402
rect 6162 29350 6174 29402
rect 6226 29350 8832 29402
rect 1104 29328 8832 29350
rect 1104 28858 8832 28880
rect 1104 28806 4315 28858
rect 4367 28806 4379 28858
rect 4431 28806 4443 28858
rect 4495 28806 4507 28858
rect 4559 28806 7648 28858
rect 7700 28806 7712 28858
rect 7764 28806 7776 28858
rect 7828 28806 7840 28858
rect 7892 28806 8832 28858
rect 1104 28784 8832 28806
rect 1104 28314 8832 28336
rect 1104 28262 2648 28314
rect 2700 28262 2712 28314
rect 2764 28262 2776 28314
rect 2828 28262 2840 28314
rect 2892 28262 5982 28314
rect 6034 28262 6046 28314
rect 6098 28262 6110 28314
rect 6162 28262 6174 28314
rect 6226 28262 8832 28314
rect 1104 28240 8832 28262
rect 1104 27770 8832 27792
rect 1104 27718 4315 27770
rect 4367 27718 4379 27770
rect 4431 27718 4443 27770
rect 4495 27718 4507 27770
rect 4559 27718 7648 27770
rect 7700 27718 7712 27770
rect 7764 27718 7776 27770
rect 7828 27718 7840 27770
rect 7892 27718 8832 27770
rect 1104 27696 8832 27718
rect 1104 27226 8832 27248
rect 1104 27174 2648 27226
rect 2700 27174 2712 27226
rect 2764 27174 2776 27226
rect 2828 27174 2840 27226
rect 2892 27174 5982 27226
rect 6034 27174 6046 27226
rect 6098 27174 6110 27226
rect 6162 27174 6174 27226
rect 6226 27174 8832 27226
rect 1104 27152 8832 27174
rect 1104 26682 8832 26704
rect 1104 26630 4315 26682
rect 4367 26630 4379 26682
rect 4431 26630 4443 26682
rect 4495 26630 4507 26682
rect 4559 26630 7648 26682
rect 7700 26630 7712 26682
rect 7764 26630 7776 26682
rect 7828 26630 7840 26682
rect 7892 26630 8832 26682
rect 1104 26608 8832 26630
rect 1104 26138 8832 26160
rect 1104 26086 2648 26138
rect 2700 26086 2712 26138
rect 2764 26086 2776 26138
rect 2828 26086 2840 26138
rect 2892 26086 5982 26138
rect 6034 26086 6046 26138
rect 6098 26086 6110 26138
rect 6162 26086 6174 26138
rect 6226 26086 8832 26138
rect 1104 26064 8832 26086
rect 1104 25594 8832 25616
rect 1104 25542 4315 25594
rect 4367 25542 4379 25594
rect 4431 25542 4443 25594
rect 4495 25542 4507 25594
rect 4559 25542 7648 25594
rect 7700 25542 7712 25594
rect 7764 25542 7776 25594
rect 7828 25542 7840 25594
rect 7892 25542 8832 25594
rect 1104 25520 8832 25542
rect 1104 25050 8832 25072
rect 1104 24998 2648 25050
rect 2700 24998 2712 25050
rect 2764 24998 2776 25050
rect 2828 24998 2840 25050
rect 2892 24998 5982 25050
rect 6034 24998 6046 25050
rect 6098 24998 6110 25050
rect 6162 24998 6174 25050
rect 6226 24998 8832 25050
rect 1104 24976 8832 24998
rect 1104 24506 8832 24528
rect 1104 24454 4315 24506
rect 4367 24454 4379 24506
rect 4431 24454 4443 24506
rect 4495 24454 4507 24506
rect 4559 24454 7648 24506
rect 7700 24454 7712 24506
rect 7764 24454 7776 24506
rect 7828 24454 7840 24506
rect 7892 24454 8832 24506
rect 1104 24432 8832 24454
rect 1104 23962 8832 23984
rect 1104 23910 2648 23962
rect 2700 23910 2712 23962
rect 2764 23910 2776 23962
rect 2828 23910 2840 23962
rect 2892 23910 5982 23962
rect 6034 23910 6046 23962
rect 6098 23910 6110 23962
rect 6162 23910 6174 23962
rect 6226 23910 8832 23962
rect 1104 23888 8832 23910
rect 1104 23418 8832 23440
rect 1104 23366 4315 23418
rect 4367 23366 4379 23418
rect 4431 23366 4443 23418
rect 4495 23366 4507 23418
rect 4559 23366 7648 23418
rect 7700 23366 7712 23418
rect 7764 23366 7776 23418
rect 7828 23366 7840 23418
rect 7892 23366 8832 23418
rect 1104 23344 8832 23366
rect 1104 22874 8832 22896
rect 1104 22822 2648 22874
rect 2700 22822 2712 22874
rect 2764 22822 2776 22874
rect 2828 22822 2840 22874
rect 2892 22822 5982 22874
rect 6034 22822 6046 22874
rect 6098 22822 6110 22874
rect 6162 22822 6174 22874
rect 6226 22822 8832 22874
rect 1104 22800 8832 22822
rect 1104 22330 8832 22352
rect 1104 22278 4315 22330
rect 4367 22278 4379 22330
rect 4431 22278 4443 22330
rect 4495 22278 4507 22330
rect 4559 22278 7648 22330
rect 7700 22278 7712 22330
rect 7764 22278 7776 22330
rect 7828 22278 7840 22330
rect 7892 22278 8832 22330
rect 1104 22256 8832 22278
rect 1104 21786 8832 21808
rect 1104 21734 2648 21786
rect 2700 21734 2712 21786
rect 2764 21734 2776 21786
rect 2828 21734 2840 21786
rect 2892 21734 5982 21786
rect 6034 21734 6046 21786
rect 6098 21734 6110 21786
rect 6162 21734 6174 21786
rect 6226 21734 8832 21786
rect 1104 21712 8832 21734
rect 1104 21242 8832 21264
rect 1104 21190 4315 21242
rect 4367 21190 4379 21242
rect 4431 21190 4443 21242
rect 4495 21190 4507 21242
rect 4559 21190 7648 21242
rect 7700 21190 7712 21242
rect 7764 21190 7776 21242
rect 7828 21190 7840 21242
rect 7892 21190 8832 21242
rect 1104 21168 8832 21190
rect 1104 20698 8832 20720
rect 1104 20646 2648 20698
rect 2700 20646 2712 20698
rect 2764 20646 2776 20698
rect 2828 20646 2840 20698
rect 2892 20646 5982 20698
rect 6034 20646 6046 20698
rect 6098 20646 6110 20698
rect 6162 20646 6174 20698
rect 6226 20646 8832 20698
rect 1104 20624 8832 20646
rect 1104 20154 8832 20176
rect 1104 20102 4315 20154
rect 4367 20102 4379 20154
rect 4431 20102 4443 20154
rect 4495 20102 4507 20154
rect 4559 20102 7648 20154
rect 7700 20102 7712 20154
rect 7764 20102 7776 20154
rect 7828 20102 7840 20154
rect 7892 20102 8832 20154
rect 1104 20080 8832 20102
rect 1104 19610 8832 19632
rect 1104 19558 2648 19610
rect 2700 19558 2712 19610
rect 2764 19558 2776 19610
rect 2828 19558 2840 19610
rect 2892 19558 5982 19610
rect 6034 19558 6046 19610
rect 6098 19558 6110 19610
rect 6162 19558 6174 19610
rect 6226 19558 8832 19610
rect 1104 19536 8832 19558
rect 1104 19066 8832 19088
rect 1104 19014 4315 19066
rect 4367 19014 4379 19066
rect 4431 19014 4443 19066
rect 4495 19014 4507 19066
rect 4559 19014 7648 19066
rect 7700 19014 7712 19066
rect 7764 19014 7776 19066
rect 7828 19014 7840 19066
rect 7892 19014 8832 19066
rect 1104 18992 8832 19014
rect 1104 18522 8832 18544
rect 1104 18470 2648 18522
rect 2700 18470 2712 18522
rect 2764 18470 2776 18522
rect 2828 18470 2840 18522
rect 2892 18470 5982 18522
rect 6034 18470 6046 18522
rect 6098 18470 6110 18522
rect 6162 18470 6174 18522
rect 6226 18470 8832 18522
rect 1104 18448 8832 18470
rect 1104 17978 8832 18000
rect 1104 17926 4315 17978
rect 4367 17926 4379 17978
rect 4431 17926 4443 17978
rect 4495 17926 4507 17978
rect 4559 17926 7648 17978
rect 7700 17926 7712 17978
rect 7764 17926 7776 17978
rect 7828 17926 7840 17978
rect 7892 17926 8832 17978
rect 1104 17904 8832 17926
rect 1104 17434 8832 17456
rect 1104 17382 2648 17434
rect 2700 17382 2712 17434
rect 2764 17382 2776 17434
rect 2828 17382 2840 17434
rect 2892 17382 5982 17434
rect 6034 17382 6046 17434
rect 6098 17382 6110 17434
rect 6162 17382 6174 17434
rect 6226 17382 8832 17434
rect 1104 17360 8832 17382
rect 1104 16890 8832 16912
rect 1104 16838 4315 16890
rect 4367 16838 4379 16890
rect 4431 16838 4443 16890
rect 4495 16838 4507 16890
rect 4559 16838 7648 16890
rect 7700 16838 7712 16890
rect 7764 16838 7776 16890
rect 7828 16838 7840 16890
rect 7892 16838 8832 16890
rect 1104 16816 8832 16838
rect 1104 16346 8832 16368
rect 1104 16294 2648 16346
rect 2700 16294 2712 16346
rect 2764 16294 2776 16346
rect 2828 16294 2840 16346
rect 2892 16294 5982 16346
rect 6034 16294 6046 16346
rect 6098 16294 6110 16346
rect 6162 16294 6174 16346
rect 6226 16294 8832 16346
rect 1104 16272 8832 16294
rect 1104 15802 8832 15824
rect 1104 15750 4315 15802
rect 4367 15750 4379 15802
rect 4431 15750 4443 15802
rect 4495 15750 4507 15802
rect 4559 15750 7648 15802
rect 7700 15750 7712 15802
rect 7764 15750 7776 15802
rect 7828 15750 7840 15802
rect 7892 15750 8832 15802
rect 1104 15728 8832 15750
rect 1104 15258 8832 15280
rect 1104 15206 2648 15258
rect 2700 15206 2712 15258
rect 2764 15206 2776 15258
rect 2828 15206 2840 15258
rect 2892 15206 5982 15258
rect 6034 15206 6046 15258
rect 6098 15206 6110 15258
rect 6162 15206 6174 15258
rect 6226 15206 8832 15258
rect 1104 15184 8832 15206
rect 1104 14714 8832 14736
rect 1104 14662 4315 14714
rect 4367 14662 4379 14714
rect 4431 14662 4443 14714
rect 4495 14662 4507 14714
rect 4559 14662 7648 14714
rect 7700 14662 7712 14714
rect 7764 14662 7776 14714
rect 7828 14662 7840 14714
rect 7892 14662 8832 14714
rect 1104 14640 8832 14662
rect 1104 14170 8832 14192
rect 1104 14118 2648 14170
rect 2700 14118 2712 14170
rect 2764 14118 2776 14170
rect 2828 14118 2840 14170
rect 2892 14118 5982 14170
rect 6034 14118 6046 14170
rect 6098 14118 6110 14170
rect 6162 14118 6174 14170
rect 6226 14118 8832 14170
rect 1104 14096 8832 14118
rect 1104 13626 8832 13648
rect 1104 13574 4315 13626
rect 4367 13574 4379 13626
rect 4431 13574 4443 13626
rect 4495 13574 4507 13626
rect 4559 13574 7648 13626
rect 7700 13574 7712 13626
rect 7764 13574 7776 13626
rect 7828 13574 7840 13626
rect 7892 13574 8832 13626
rect 1104 13552 8832 13574
rect 1104 13082 8832 13104
rect 1104 13030 2648 13082
rect 2700 13030 2712 13082
rect 2764 13030 2776 13082
rect 2828 13030 2840 13082
rect 2892 13030 5982 13082
rect 6034 13030 6046 13082
rect 6098 13030 6110 13082
rect 6162 13030 6174 13082
rect 6226 13030 8832 13082
rect 1104 13008 8832 13030
rect 1104 12538 8832 12560
rect 1104 12486 4315 12538
rect 4367 12486 4379 12538
rect 4431 12486 4443 12538
rect 4495 12486 4507 12538
rect 4559 12486 7648 12538
rect 7700 12486 7712 12538
rect 7764 12486 7776 12538
rect 7828 12486 7840 12538
rect 7892 12486 8832 12538
rect 1104 12464 8832 12486
rect 1104 11994 8832 12016
rect 1104 11942 2648 11994
rect 2700 11942 2712 11994
rect 2764 11942 2776 11994
rect 2828 11942 2840 11994
rect 2892 11942 5982 11994
rect 6034 11942 6046 11994
rect 6098 11942 6110 11994
rect 6162 11942 6174 11994
rect 6226 11942 8832 11994
rect 1104 11920 8832 11942
rect 1104 11450 8832 11472
rect 1104 11398 4315 11450
rect 4367 11398 4379 11450
rect 4431 11398 4443 11450
rect 4495 11398 4507 11450
rect 4559 11398 7648 11450
rect 7700 11398 7712 11450
rect 7764 11398 7776 11450
rect 7828 11398 7840 11450
rect 7892 11398 8832 11450
rect 1104 11376 8832 11398
rect 1104 10906 8832 10928
rect 1104 10854 2648 10906
rect 2700 10854 2712 10906
rect 2764 10854 2776 10906
rect 2828 10854 2840 10906
rect 2892 10854 5982 10906
rect 6034 10854 6046 10906
rect 6098 10854 6110 10906
rect 6162 10854 6174 10906
rect 6226 10854 8832 10906
rect 1104 10832 8832 10854
rect 1104 10362 8832 10384
rect 1104 10310 4315 10362
rect 4367 10310 4379 10362
rect 4431 10310 4443 10362
rect 4495 10310 4507 10362
rect 4559 10310 7648 10362
rect 7700 10310 7712 10362
rect 7764 10310 7776 10362
rect 7828 10310 7840 10362
rect 7892 10310 8832 10362
rect 1104 10288 8832 10310
rect 1104 9818 8832 9840
rect 1104 9766 2648 9818
rect 2700 9766 2712 9818
rect 2764 9766 2776 9818
rect 2828 9766 2840 9818
rect 2892 9766 5982 9818
rect 6034 9766 6046 9818
rect 6098 9766 6110 9818
rect 6162 9766 6174 9818
rect 6226 9766 8832 9818
rect 1104 9744 8832 9766
rect 1104 9274 8832 9296
rect 1104 9222 4315 9274
rect 4367 9222 4379 9274
rect 4431 9222 4443 9274
rect 4495 9222 4507 9274
rect 4559 9222 7648 9274
rect 7700 9222 7712 9274
rect 7764 9222 7776 9274
rect 7828 9222 7840 9274
rect 7892 9222 8832 9274
rect 1104 9200 8832 9222
rect 1104 8730 8832 8752
rect 1104 8678 2648 8730
rect 2700 8678 2712 8730
rect 2764 8678 2776 8730
rect 2828 8678 2840 8730
rect 2892 8678 5982 8730
rect 6034 8678 6046 8730
rect 6098 8678 6110 8730
rect 6162 8678 6174 8730
rect 6226 8678 8832 8730
rect 1104 8656 8832 8678
rect 1104 8186 8832 8208
rect 1104 8134 4315 8186
rect 4367 8134 4379 8186
rect 4431 8134 4443 8186
rect 4495 8134 4507 8186
rect 4559 8134 7648 8186
rect 7700 8134 7712 8186
rect 7764 8134 7776 8186
rect 7828 8134 7840 8186
rect 7892 8134 8832 8186
rect 1104 8112 8832 8134
rect 1104 7642 8832 7664
rect 1104 7590 2648 7642
rect 2700 7590 2712 7642
rect 2764 7590 2776 7642
rect 2828 7590 2840 7642
rect 2892 7590 5982 7642
rect 6034 7590 6046 7642
rect 6098 7590 6110 7642
rect 6162 7590 6174 7642
rect 6226 7590 8832 7642
rect 1104 7568 8832 7590
rect 1104 7098 8832 7120
rect 1104 7046 4315 7098
rect 4367 7046 4379 7098
rect 4431 7046 4443 7098
rect 4495 7046 4507 7098
rect 4559 7046 7648 7098
rect 7700 7046 7712 7098
rect 7764 7046 7776 7098
rect 7828 7046 7840 7098
rect 7892 7046 8832 7098
rect 1104 7024 8832 7046
rect 1104 6554 8832 6576
rect 1104 6502 2648 6554
rect 2700 6502 2712 6554
rect 2764 6502 2776 6554
rect 2828 6502 2840 6554
rect 2892 6502 5982 6554
rect 6034 6502 6046 6554
rect 6098 6502 6110 6554
rect 6162 6502 6174 6554
rect 6226 6502 8832 6554
rect 1104 6480 8832 6502
rect 1104 6010 8832 6032
rect 1104 5958 4315 6010
rect 4367 5958 4379 6010
rect 4431 5958 4443 6010
rect 4495 5958 4507 6010
rect 4559 5958 7648 6010
rect 7700 5958 7712 6010
rect 7764 5958 7776 6010
rect 7828 5958 7840 6010
rect 7892 5958 8832 6010
rect 1104 5936 8832 5958
rect 1104 5466 8832 5488
rect 1104 5414 2648 5466
rect 2700 5414 2712 5466
rect 2764 5414 2776 5466
rect 2828 5414 2840 5466
rect 2892 5414 5982 5466
rect 6034 5414 6046 5466
rect 6098 5414 6110 5466
rect 6162 5414 6174 5466
rect 6226 5414 8832 5466
rect 1104 5392 8832 5414
rect 1104 4922 8832 4944
rect 1104 4870 4315 4922
rect 4367 4870 4379 4922
rect 4431 4870 4443 4922
rect 4495 4870 4507 4922
rect 4559 4870 7648 4922
rect 7700 4870 7712 4922
rect 7764 4870 7776 4922
rect 7828 4870 7840 4922
rect 7892 4870 8832 4922
rect 1104 4848 8832 4870
rect 1104 4378 8832 4400
rect 1104 4326 2648 4378
rect 2700 4326 2712 4378
rect 2764 4326 2776 4378
rect 2828 4326 2840 4378
rect 2892 4326 5982 4378
rect 6034 4326 6046 4378
rect 6098 4326 6110 4378
rect 6162 4326 6174 4378
rect 6226 4326 8832 4378
rect 1104 4304 8832 4326
rect 1104 3834 8832 3856
rect 1104 3782 4315 3834
rect 4367 3782 4379 3834
rect 4431 3782 4443 3834
rect 4495 3782 4507 3834
rect 4559 3782 7648 3834
rect 7700 3782 7712 3834
rect 7764 3782 7776 3834
rect 7828 3782 7840 3834
rect 7892 3782 8832 3834
rect 1104 3760 8832 3782
rect 1104 3290 8832 3312
rect 1104 3238 2648 3290
rect 2700 3238 2712 3290
rect 2764 3238 2776 3290
rect 2828 3238 2840 3290
rect 2892 3238 5982 3290
rect 6034 3238 6046 3290
rect 6098 3238 6110 3290
rect 6162 3238 6174 3290
rect 6226 3238 8832 3290
rect 1104 3216 8832 3238
rect 1104 2746 8832 2768
rect 1104 2694 4315 2746
rect 4367 2694 4379 2746
rect 4431 2694 4443 2746
rect 4495 2694 4507 2746
rect 4559 2694 7648 2746
rect 7700 2694 7712 2746
rect 7764 2694 7776 2746
rect 7828 2694 7840 2746
rect 7892 2694 8832 2746
rect 1104 2672 8832 2694
rect 1104 2202 8832 2224
rect 1104 2150 2648 2202
rect 2700 2150 2712 2202
rect 2764 2150 2776 2202
rect 2828 2150 2840 2202
rect 2892 2150 5982 2202
rect 6034 2150 6046 2202
rect 6098 2150 6110 2202
rect 6162 2150 6174 2202
rect 6226 2150 8832 2202
rect 1104 2128 8832 2150
rect 8202 76 8208 128
rect 8260 116 8266 128
rect 8938 116 8944 128
rect 8260 88 8944 116
rect 8260 76 8266 88
rect 8938 76 8944 88
rect 8996 76 9002 128
<< via1 >>
rect 572 332528 624 332580
rect 1216 332528 1268 332580
rect 3056 332528 3108 332580
rect 3884 332528 3936 332580
rect 4252 332528 4304 332580
rect 5448 332528 5500 332580
rect 8300 332528 8352 332580
rect 9312 332528 9364 332580
rect 2648 330726 2700 330778
rect 2712 330726 2764 330778
rect 2776 330726 2828 330778
rect 2840 330726 2892 330778
rect 5982 330726 6034 330778
rect 6046 330726 6098 330778
rect 6110 330726 6162 330778
rect 6174 330726 6226 330778
rect 4315 330182 4367 330234
rect 4379 330182 4431 330234
rect 4443 330182 4495 330234
rect 4507 330182 4559 330234
rect 7648 330182 7700 330234
rect 7712 330182 7764 330234
rect 7776 330182 7828 330234
rect 7840 330182 7892 330234
rect 2648 329638 2700 329690
rect 2712 329638 2764 329690
rect 2776 329638 2828 329690
rect 2840 329638 2892 329690
rect 5982 329638 6034 329690
rect 6046 329638 6098 329690
rect 6110 329638 6162 329690
rect 6174 329638 6226 329690
rect 4315 329094 4367 329146
rect 4379 329094 4431 329146
rect 4443 329094 4495 329146
rect 4507 329094 4559 329146
rect 7648 329094 7700 329146
rect 7712 329094 7764 329146
rect 7776 329094 7828 329146
rect 7840 329094 7892 329146
rect 2648 328550 2700 328602
rect 2712 328550 2764 328602
rect 2776 328550 2828 328602
rect 2840 328550 2892 328602
rect 5982 328550 6034 328602
rect 6046 328550 6098 328602
rect 6110 328550 6162 328602
rect 6174 328550 6226 328602
rect 4315 328006 4367 328058
rect 4379 328006 4431 328058
rect 4443 328006 4495 328058
rect 4507 328006 4559 328058
rect 7648 328006 7700 328058
rect 7712 328006 7764 328058
rect 7776 328006 7828 328058
rect 7840 328006 7892 328058
rect 2648 327462 2700 327514
rect 2712 327462 2764 327514
rect 2776 327462 2828 327514
rect 2840 327462 2892 327514
rect 5982 327462 6034 327514
rect 6046 327462 6098 327514
rect 6110 327462 6162 327514
rect 6174 327462 6226 327514
rect 4315 326918 4367 326970
rect 4379 326918 4431 326970
rect 4443 326918 4495 326970
rect 4507 326918 4559 326970
rect 7648 326918 7700 326970
rect 7712 326918 7764 326970
rect 7776 326918 7828 326970
rect 7840 326918 7892 326970
rect 2648 326374 2700 326426
rect 2712 326374 2764 326426
rect 2776 326374 2828 326426
rect 2840 326374 2892 326426
rect 5982 326374 6034 326426
rect 6046 326374 6098 326426
rect 6110 326374 6162 326426
rect 6174 326374 6226 326426
rect 4315 325830 4367 325882
rect 4379 325830 4431 325882
rect 4443 325830 4495 325882
rect 4507 325830 4559 325882
rect 7648 325830 7700 325882
rect 7712 325830 7764 325882
rect 7776 325830 7828 325882
rect 7840 325830 7892 325882
rect 2648 325286 2700 325338
rect 2712 325286 2764 325338
rect 2776 325286 2828 325338
rect 2840 325286 2892 325338
rect 5982 325286 6034 325338
rect 6046 325286 6098 325338
rect 6110 325286 6162 325338
rect 6174 325286 6226 325338
rect 4315 324742 4367 324794
rect 4379 324742 4431 324794
rect 4443 324742 4495 324794
rect 4507 324742 4559 324794
rect 7648 324742 7700 324794
rect 7712 324742 7764 324794
rect 7776 324742 7828 324794
rect 7840 324742 7892 324794
rect 2648 324198 2700 324250
rect 2712 324198 2764 324250
rect 2776 324198 2828 324250
rect 2840 324198 2892 324250
rect 5982 324198 6034 324250
rect 6046 324198 6098 324250
rect 6110 324198 6162 324250
rect 6174 324198 6226 324250
rect 4315 323654 4367 323706
rect 4379 323654 4431 323706
rect 4443 323654 4495 323706
rect 4507 323654 4559 323706
rect 7648 323654 7700 323706
rect 7712 323654 7764 323706
rect 7776 323654 7828 323706
rect 7840 323654 7892 323706
rect 2648 323110 2700 323162
rect 2712 323110 2764 323162
rect 2776 323110 2828 323162
rect 2840 323110 2892 323162
rect 5982 323110 6034 323162
rect 6046 323110 6098 323162
rect 6110 323110 6162 323162
rect 6174 323110 6226 323162
rect 4315 322566 4367 322618
rect 4379 322566 4431 322618
rect 4443 322566 4495 322618
rect 4507 322566 4559 322618
rect 7648 322566 7700 322618
rect 7712 322566 7764 322618
rect 7776 322566 7828 322618
rect 7840 322566 7892 322618
rect 2648 322022 2700 322074
rect 2712 322022 2764 322074
rect 2776 322022 2828 322074
rect 2840 322022 2892 322074
rect 5982 322022 6034 322074
rect 6046 322022 6098 322074
rect 6110 322022 6162 322074
rect 6174 322022 6226 322074
rect 4315 321478 4367 321530
rect 4379 321478 4431 321530
rect 4443 321478 4495 321530
rect 4507 321478 4559 321530
rect 7648 321478 7700 321530
rect 7712 321478 7764 321530
rect 7776 321478 7828 321530
rect 7840 321478 7892 321530
rect 2648 320934 2700 320986
rect 2712 320934 2764 320986
rect 2776 320934 2828 320986
rect 2840 320934 2892 320986
rect 5982 320934 6034 320986
rect 6046 320934 6098 320986
rect 6110 320934 6162 320986
rect 6174 320934 6226 320986
rect 4315 320390 4367 320442
rect 4379 320390 4431 320442
rect 4443 320390 4495 320442
rect 4507 320390 4559 320442
rect 7648 320390 7700 320442
rect 7712 320390 7764 320442
rect 7776 320390 7828 320442
rect 7840 320390 7892 320442
rect 2648 319846 2700 319898
rect 2712 319846 2764 319898
rect 2776 319846 2828 319898
rect 2840 319846 2892 319898
rect 5982 319846 6034 319898
rect 6046 319846 6098 319898
rect 6110 319846 6162 319898
rect 6174 319846 6226 319898
rect 4315 319302 4367 319354
rect 4379 319302 4431 319354
rect 4443 319302 4495 319354
rect 4507 319302 4559 319354
rect 7648 319302 7700 319354
rect 7712 319302 7764 319354
rect 7776 319302 7828 319354
rect 7840 319302 7892 319354
rect 2648 318758 2700 318810
rect 2712 318758 2764 318810
rect 2776 318758 2828 318810
rect 2840 318758 2892 318810
rect 5982 318758 6034 318810
rect 6046 318758 6098 318810
rect 6110 318758 6162 318810
rect 6174 318758 6226 318810
rect 4315 318214 4367 318266
rect 4379 318214 4431 318266
rect 4443 318214 4495 318266
rect 4507 318214 4559 318266
rect 7648 318214 7700 318266
rect 7712 318214 7764 318266
rect 7776 318214 7828 318266
rect 7840 318214 7892 318266
rect 2648 317670 2700 317722
rect 2712 317670 2764 317722
rect 2776 317670 2828 317722
rect 2840 317670 2892 317722
rect 5982 317670 6034 317722
rect 6046 317670 6098 317722
rect 6110 317670 6162 317722
rect 6174 317670 6226 317722
rect 4315 317126 4367 317178
rect 4379 317126 4431 317178
rect 4443 317126 4495 317178
rect 4507 317126 4559 317178
rect 7648 317126 7700 317178
rect 7712 317126 7764 317178
rect 7776 317126 7828 317178
rect 7840 317126 7892 317178
rect 2648 316582 2700 316634
rect 2712 316582 2764 316634
rect 2776 316582 2828 316634
rect 2840 316582 2892 316634
rect 5982 316582 6034 316634
rect 6046 316582 6098 316634
rect 6110 316582 6162 316634
rect 6174 316582 6226 316634
rect 4315 316038 4367 316090
rect 4379 316038 4431 316090
rect 4443 316038 4495 316090
rect 4507 316038 4559 316090
rect 7648 316038 7700 316090
rect 7712 316038 7764 316090
rect 7776 316038 7828 316090
rect 7840 316038 7892 316090
rect 2648 315494 2700 315546
rect 2712 315494 2764 315546
rect 2776 315494 2828 315546
rect 2840 315494 2892 315546
rect 5982 315494 6034 315546
rect 6046 315494 6098 315546
rect 6110 315494 6162 315546
rect 6174 315494 6226 315546
rect 7380 315120 7432 315172
rect 8024 315120 8076 315172
rect 4315 314950 4367 315002
rect 4379 314950 4431 315002
rect 4443 314950 4495 315002
rect 4507 314950 4559 315002
rect 7648 314950 7700 315002
rect 7712 314950 7764 315002
rect 7776 314950 7828 315002
rect 7840 314950 7892 315002
rect 2648 314406 2700 314458
rect 2712 314406 2764 314458
rect 2776 314406 2828 314458
rect 2840 314406 2892 314458
rect 5982 314406 6034 314458
rect 6046 314406 6098 314458
rect 6110 314406 6162 314458
rect 6174 314406 6226 314458
rect 4315 313862 4367 313914
rect 4379 313862 4431 313914
rect 4443 313862 4495 313914
rect 4507 313862 4559 313914
rect 7648 313862 7700 313914
rect 7712 313862 7764 313914
rect 7776 313862 7828 313914
rect 7840 313862 7892 313914
rect 2648 313318 2700 313370
rect 2712 313318 2764 313370
rect 2776 313318 2828 313370
rect 2840 313318 2892 313370
rect 5982 313318 6034 313370
rect 6046 313318 6098 313370
rect 6110 313318 6162 313370
rect 6174 313318 6226 313370
rect 4315 312774 4367 312826
rect 4379 312774 4431 312826
rect 4443 312774 4495 312826
rect 4507 312774 4559 312826
rect 7648 312774 7700 312826
rect 7712 312774 7764 312826
rect 7776 312774 7828 312826
rect 7840 312774 7892 312826
rect 2648 312230 2700 312282
rect 2712 312230 2764 312282
rect 2776 312230 2828 312282
rect 2840 312230 2892 312282
rect 5982 312230 6034 312282
rect 6046 312230 6098 312282
rect 6110 312230 6162 312282
rect 6174 312230 6226 312282
rect 4315 311686 4367 311738
rect 4379 311686 4431 311738
rect 4443 311686 4495 311738
rect 4507 311686 4559 311738
rect 7648 311686 7700 311738
rect 7712 311686 7764 311738
rect 7776 311686 7828 311738
rect 7840 311686 7892 311738
rect 2648 311142 2700 311194
rect 2712 311142 2764 311194
rect 2776 311142 2828 311194
rect 2840 311142 2892 311194
rect 5982 311142 6034 311194
rect 6046 311142 6098 311194
rect 6110 311142 6162 311194
rect 6174 311142 6226 311194
rect 4315 310598 4367 310650
rect 4379 310598 4431 310650
rect 4443 310598 4495 310650
rect 4507 310598 4559 310650
rect 7648 310598 7700 310650
rect 7712 310598 7764 310650
rect 7776 310598 7828 310650
rect 7840 310598 7892 310650
rect 2648 310054 2700 310106
rect 2712 310054 2764 310106
rect 2776 310054 2828 310106
rect 2840 310054 2892 310106
rect 5982 310054 6034 310106
rect 6046 310054 6098 310106
rect 6110 310054 6162 310106
rect 6174 310054 6226 310106
rect 4315 309510 4367 309562
rect 4379 309510 4431 309562
rect 4443 309510 4495 309562
rect 4507 309510 4559 309562
rect 7648 309510 7700 309562
rect 7712 309510 7764 309562
rect 7776 309510 7828 309562
rect 7840 309510 7892 309562
rect 2648 308966 2700 309018
rect 2712 308966 2764 309018
rect 2776 308966 2828 309018
rect 2840 308966 2892 309018
rect 5982 308966 6034 309018
rect 6046 308966 6098 309018
rect 6110 308966 6162 309018
rect 6174 308966 6226 309018
rect 4315 308422 4367 308474
rect 4379 308422 4431 308474
rect 4443 308422 4495 308474
rect 4507 308422 4559 308474
rect 7648 308422 7700 308474
rect 7712 308422 7764 308474
rect 7776 308422 7828 308474
rect 7840 308422 7892 308474
rect 2648 307878 2700 307930
rect 2712 307878 2764 307930
rect 2776 307878 2828 307930
rect 2840 307878 2892 307930
rect 5982 307878 6034 307930
rect 6046 307878 6098 307930
rect 6110 307878 6162 307930
rect 6174 307878 6226 307930
rect 4315 307334 4367 307386
rect 4379 307334 4431 307386
rect 4443 307334 4495 307386
rect 4507 307334 4559 307386
rect 7648 307334 7700 307386
rect 7712 307334 7764 307386
rect 7776 307334 7828 307386
rect 7840 307334 7892 307386
rect 2648 306790 2700 306842
rect 2712 306790 2764 306842
rect 2776 306790 2828 306842
rect 2840 306790 2892 306842
rect 5982 306790 6034 306842
rect 6046 306790 6098 306842
rect 6110 306790 6162 306842
rect 6174 306790 6226 306842
rect 4315 306246 4367 306298
rect 4379 306246 4431 306298
rect 4443 306246 4495 306298
rect 4507 306246 4559 306298
rect 7648 306246 7700 306298
rect 7712 306246 7764 306298
rect 7776 306246 7828 306298
rect 7840 306246 7892 306298
rect 2648 305702 2700 305754
rect 2712 305702 2764 305754
rect 2776 305702 2828 305754
rect 2840 305702 2892 305754
rect 5982 305702 6034 305754
rect 6046 305702 6098 305754
rect 6110 305702 6162 305754
rect 6174 305702 6226 305754
rect 4315 305158 4367 305210
rect 4379 305158 4431 305210
rect 4443 305158 4495 305210
rect 4507 305158 4559 305210
rect 7648 305158 7700 305210
rect 7712 305158 7764 305210
rect 7776 305158 7828 305210
rect 7840 305158 7892 305210
rect 2648 304614 2700 304666
rect 2712 304614 2764 304666
rect 2776 304614 2828 304666
rect 2840 304614 2892 304666
rect 5982 304614 6034 304666
rect 6046 304614 6098 304666
rect 6110 304614 6162 304666
rect 6174 304614 6226 304666
rect 4315 304070 4367 304122
rect 4379 304070 4431 304122
rect 4443 304070 4495 304122
rect 4507 304070 4559 304122
rect 7648 304070 7700 304122
rect 7712 304070 7764 304122
rect 7776 304070 7828 304122
rect 7840 304070 7892 304122
rect 2648 303526 2700 303578
rect 2712 303526 2764 303578
rect 2776 303526 2828 303578
rect 2840 303526 2892 303578
rect 5982 303526 6034 303578
rect 6046 303526 6098 303578
rect 6110 303526 6162 303578
rect 6174 303526 6226 303578
rect 4315 302982 4367 303034
rect 4379 302982 4431 303034
rect 4443 302982 4495 303034
rect 4507 302982 4559 303034
rect 7648 302982 7700 303034
rect 7712 302982 7764 303034
rect 7776 302982 7828 303034
rect 7840 302982 7892 303034
rect 2648 302438 2700 302490
rect 2712 302438 2764 302490
rect 2776 302438 2828 302490
rect 2840 302438 2892 302490
rect 5982 302438 6034 302490
rect 6046 302438 6098 302490
rect 6110 302438 6162 302490
rect 6174 302438 6226 302490
rect 4315 301894 4367 301946
rect 4379 301894 4431 301946
rect 4443 301894 4495 301946
rect 4507 301894 4559 301946
rect 7648 301894 7700 301946
rect 7712 301894 7764 301946
rect 7776 301894 7828 301946
rect 7840 301894 7892 301946
rect 2648 301350 2700 301402
rect 2712 301350 2764 301402
rect 2776 301350 2828 301402
rect 2840 301350 2892 301402
rect 5982 301350 6034 301402
rect 6046 301350 6098 301402
rect 6110 301350 6162 301402
rect 6174 301350 6226 301402
rect 4315 300806 4367 300858
rect 4379 300806 4431 300858
rect 4443 300806 4495 300858
rect 4507 300806 4559 300858
rect 7648 300806 7700 300858
rect 7712 300806 7764 300858
rect 7776 300806 7828 300858
rect 7840 300806 7892 300858
rect 2648 300262 2700 300314
rect 2712 300262 2764 300314
rect 2776 300262 2828 300314
rect 2840 300262 2892 300314
rect 5982 300262 6034 300314
rect 6046 300262 6098 300314
rect 6110 300262 6162 300314
rect 6174 300262 6226 300314
rect 4315 299718 4367 299770
rect 4379 299718 4431 299770
rect 4443 299718 4495 299770
rect 4507 299718 4559 299770
rect 7648 299718 7700 299770
rect 7712 299718 7764 299770
rect 7776 299718 7828 299770
rect 7840 299718 7892 299770
rect 2648 299174 2700 299226
rect 2712 299174 2764 299226
rect 2776 299174 2828 299226
rect 2840 299174 2892 299226
rect 5982 299174 6034 299226
rect 6046 299174 6098 299226
rect 6110 299174 6162 299226
rect 6174 299174 6226 299226
rect 4315 298630 4367 298682
rect 4379 298630 4431 298682
rect 4443 298630 4495 298682
rect 4507 298630 4559 298682
rect 7648 298630 7700 298682
rect 7712 298630 7764 298682
rect 7776 298630 7828 298682
rect 7840 298630 7892 298682
rect 2648 298086 2700 298138
rect 2712 298086 2764 298138
rect 2776 298086 2828 298138
rect 2840 298086 2892 298138
rect 5982 298086 6034 298138
rect 6046 298086 6098 298138
rect 6110 298086 6162 298138
rect 6174 298086 6226 298138
rect 4315 297542 4367 297594
rect 4379 297542 4431 297594
rect 4443 297542 4495 297594
rect 4507 297542 4559 297594
rect 7648 297542 7700 297594
rect 7712 297542 7764 297594
rect 7776 297542 7828 297594
rect 7840 297542 7892 297594
rect 2648 296998 2700 297050
rect 2712 296998 2764 297050
rect 2776 296998 2828 297050
rect 2840 296998 2892 297050
rect 5982 296998 6034 297050
rect 6046 296998 6098 297050
rect 6110 296998 6162 297050
rect 6174 296998 6226 297050
rect 4315 296454 4367 296506
rect 4379 296454 4431 296506
rect 4443 296454 4495 296506
rect 4507 296454 4559 296506
rect 7648 296454 7700 296506
rect 7712 296454 7764 296506
rect 7776 296454 7828 296506
rect 7840 296454 7892 296506
rect 2648 295910 2700 295962
rect 2712 295910 2764 295962
rect 2776 295910 2828 295962
rect 2840 295910 2892 295962
rect 5982 295910 6034 295962
rect 6046 295910 6098 295962
rect 6110 295910 6162 295962
rect 6174 295910 6226 295962
rect 4315 295366 4367 295418
rect 4379 295366 4431 295418
rect 4443 295366 4495 295418
rect 4507 295366 4559 295418
rect 7648 295366 7700 295418
rect 7712 295366 7764 295418
rect 7776 295366 7828 295418
rect 7840 295366 7892 295418
rect 2648 294822 2700 294874
rect 2712 294822 2764 294874
rect 2776 294822 2828 294874
rect 2840 294822 2892 294874
rect 5982 294822 6034 294874
rect 6046 294822 6098 294874
rect 6110 294822 6162 294874
rect 6174 294822 6226 294874
rect 4315 294278 4367 294330
rect 4379 294278 4431 294330
rect 4443 294278 4495 294330
rect 4507 294278 4559 294330
rect 7648 294278 7700 294330
rect 7712 294278 7764 294330
rect 7776 294278 7828 294330
rect 7840 294278 7892 294330
rect 2648 293734 2700 293786
rect 2712 293734 2764 293786
rect 2776 293734 2828 293786
rect 2840 293734 2892 293786
rect 5982 293734 6034 293786
rect 6046 293734 6098 293786
rect 6110 293734 6162 293786
rect 6174 293734 6226 293786
rect 4315 293190 4367 293242
rect 4379 293190 4431 293242
rect 4443 293190 4495 293242
rect 4507 293190 4559 293242
rect 7648 293190 7700 293242
rect 7712 293190 7764 293242
rect 7776 293190 7828 293242
rect 7840 293190 7892 293242
rect 2648 292646 2700 292698
rect 2712 292646 2764 292698
rect 2776 292646 2828 292698
rect 2840 292646 2892 292698
rect 5982 292646 6034 292698
rect 6046 292646 6098 292698
rect 6110 292646 6162 292698
rect 6174 292646 6226 292698
rect 4315 292102 4367 292154
rect 4379 292102 4431 292154
rect 4443 292102 4495 292154
rect 4507 292102 4559 292154
rect 7648 292102 7700 292154
rect 7712 292102 7764 292154
rect 7776 292102 7828 292154
rect 7840 292102 7892 292154
rect 2648 291558 2700 291610
rect 2712 291558 2764 291610
rect 2776 291558 2828 291610
rect 2840 291558 2892 291610
rect 5982 291558 6034 291610
rect 6046 291558 6098 291610
rect 6110 291558 6162 291610
rect 6174 291558 6226 291610
rect 4315 291014 4367 291066
rect 4379 291014 4431 291066
rect 4443 291014 4495 291066
rect 4507 291014 4559 291066
rect 7648 291014 7700 291066
rect 7712 291014 7764 291066
rect 7776 291014 7828 291066
rect 7840 291014 7892 291066
rect 2648 290470 2700 290522
rect 2712 290470 2764 290522
rect 2776 290470 2828 290522
rect 2840 290470 2892 290522
rect 5982 290470 6034 290522
rect 6046 290470 6098 290522
rect 6110 290470 6162 290522
rect 6174 290470 6226 290522
rect 4315 289926 4367 289978
rect 4379 289926 4431 289978
rect 4443 289926 4495 289978
rect 4507 289926 4559 289978
rect 7648 289926 7700 289978
rect 7712 289926 7764 289978
rect 7776 289926 7828 289978
rect 7840 289926 7892 289978
rect 2648 289382 2700 289434
rect 2712 289382 2764 289434
rect 2776 289382 2828 289434
rect 2840 289382 2892 289434
rect 5982 289382 6034 289434
rect 6046 289382 6098 289434
rect 6110 289382 6162 289434
rect 6174 289382 6226 289434
rect 4315 288838 4367 288890
rect 4379 288838 4431 288890
rect 4443 288838 4495 288890
rect 4507 288838 4559 288890
rect 7648 288838 7700 288890
rect 7712 288838 7764 288890
rect 7776 288838 7828 288890
rect 7840 288838 7892 288890
rect 2648 288294 2700 288346
rect 2712 288294 2764 288346
rect 2776 288294 2828 288346
rect 2840 288294 2892 288346
rect 5982 288294 6034 288346
rect 6046 288294 6098 288346
rect 6110 288294 6162 288346
rect 6174 288294 6226 288346
rect 4315 287750 4367 287802
rect 4379 287750 4431 287802
rect 4443 287750 4495 287802
rect 4507 287750 4559 287802
rect 7648 287750 7700 287802
rect 7712 287750 7764 287802
rect 7776 287750 7828 287802
rect 7840 287750 7892 287802
rect 2648 287206 2700 287258
rect 2712 287206 2764 287258
rect 2776 287206 2828 287258
rect 2840 287206 2892 287258
rect 5982 287206 6034 287258
rect 6046 287206 6098 287258
rect 6110 287206 6162 287258
rect 6174 287206 6226 287258
rect 4315 286662 4367 286714
rect 4379 286662 4431 286714
rect 4443 286662 4495 286714
rect 4507 286662 4559 286714
rect 7648 286662 7700 286714
rect 7712 286662 7764 286714
rect 7776 286662 7828 286714
rect 7840 286662 7892 286714
rect 2648 286118 2700 286170
rect 2712 286118 2764 286170
rect 2776 286118 2828 286170
rect 2840 286118 2892 286170
rect 5982 286118 6034 286170
rect 6046 286118 6098 286170
rect 6110 286118 6162 286170
rect 6174 286118 6226 286170
rect 4315 285574 4367 285626
rect 4379 285574 4431 285626
rect 4443 285574 4495 285626
rect 4507 285574 4559 285626
rect 7648 285574 7700 285626
rect 7712 285574 7764 285626
rect 7776 285574 7828 285626
rect 7840 285574 7892 285626
rect 2648 285030 2700 285082
rect 2712 285030 2764 285082
rect 2776 285030 2828 285082
rect 2840 285030 2892 285082
rect 5982 285030 6034 285082
rect 6046 285030 6098 285082
rect 6110 285030 6162 285082
rect 6174 285030 6226 285082
rect 4315 284486 4367 284538
rect 4379 284486 4431 284538
rect 4443 284486 4495 284538
rect 4507 284486 4559 284538
rect 7648 284486 7700 284538
rect 7712 284486 7764 284538
rect 7776 284486 7828 284538
rect 7840 284486 7892 284538
rect 2648 283942 2700 283994
rect 2712 283942 2764 283994
rect 2776 283942 2828 283994
rect 2840 283942 2892 283994
rect 5982 283942 6034 283994
rect 6046 283942 6098 283994
rect 6110 283942 6162 283994
rect 6174 283942 6226 283994
rect 4315 283398 4367 283450
rect 4379 283398 4431 283450
rect 4443 283398 4495 283450
rect 4507 283398 4559 283450
rect 7648 283398 7700 283450
rect 7712 283398 7764 283450
rect 7776 283398 7828 283450
rect 7840 283398 7892 283450
rect 2648 282854 2700 282906
rect 2712 282854 2764 282906
rect 2776 282854 2828 282906
rect 2840 282854 2892 282906
rect 5982 282854 6034 282906
rect 6046 282854 6098 282906
rect 6110 282854 6162 282906
rect 6174 282854 6226 282906
rect 4315 282310 4367 282362
rect 4379 282310 4431 282362
rect 4443 282310 4495 282362
rect 4507 282310 4559 282362
rect 7648 282310 7700 282362
rect 7712 282310 7764 282362
rect 7776 282310 7828 282362
rect 7840 282310 7892 282362
rect 2648 281766 2700 281818
rect 2712 281766 2764 281818
rect 2776 281766 2828 281818
rect 2840 281766 2892 281818
rect 5982 281766 6034 281818
rect 6046 281766 6098 281818
rect 6110 281766 6162 281818
rect 6174 281766 6226 281818
rect 4315 281222 4367 281274
rect 4379 281222 4431 281274
rect 4443 281222 4495 281274
rect 4507 281222 4559 281274
rect 7648 281222 7700 281274
rect 7712 281222 7764 281274
rect 7776 281222 7828 281274
rect 7840 281222 7892 281274
rect 2648 280678 2700 280730
rect 2712 280678 2764 280730
rect 2776 280678 2828 280730
rect 2840 280678 2892 280730
rect 5982 280678 6034 280730
rect 6046 280678 6098 280730
rect 6110 280678 6162 280730
rect 6174 280678 6226 280730
rect 4315 280134 4367 280186
rect 4379 280134 4431 280186
rect 4443 280134 4495 280186
rect 4507 280134 4559 280186
rect 7648 280134 7700 280186
rect 7712 280134 7764 280186
rect 7776 280134 7828 280186
rect 7840 280134 7892 280186
rect 2648 279590 2700 279642
rect 2712 279590 2764 279642
rect 2776 279590 2828 279642
rect 2840 279590 2892 279642
rect 5982 279590 6034 279642
rect 6046 279590 6098 279642
rect 6110 279590 6162 279642
rect 6174 279590 6226 279642
rect 4315 279046 4367 279098
rect 4379 279046 4431 279098
rect 4443 279046 4495 279098
rect 4507 279046 4559 279098
rect 7648 279046 7700 279098
rect 7712 279046 7764 279098
rect 7776 279046 7828 279098
rect 7840 279046 7892 279098
rect 2648 278502 2700 278554
rect 2712 278502 2764 278554
rect 2776 278502 2828 278554
rect 2840 278502 2892 278554
rect 5982 278502 6034 278554
rect 6046 278502 6098 278554
rect 6110 278502 6162 278554
rect 6174 278502 6226 278554
rect 4315 277958 4367 278010
rect 4379 277958 4431 278010
rect 4443 277958 4495 278010
rect 4507 277958 4559 278010
rect 7648 277958 7700 278010
rect 7712 277958 7764 278010
rect 7776 277958 7828 278010
rect 7840 277958 7892 278010
rect 2648 277414 2700 277466
rect 2712 277414 2764 277466
rect 2776 277414 2828 277466
rect 2840 277414 2892 277466
rect 5982 277414 6034 277466
rect 6046 277414 6098 277466
rect 6110 277414 6162 277466
rect 6174 277414 6226 277466
rect 4315 276870 4367 276922
rect 4379 276870 4431 276922
rect 4443 276870 4495 276922
rect 4507 276870 4559 276922
rect 7648 276870 7700 276922
rect 7712 276870 7764 276922
rect 7776 276870 7828 276922
rect 7840 276870 7892 276922
rect 2648 276326 2700 276378
rect 2712 276326 2764 276378
rect 2776 276326 2828 276378
rect 2840 276326 2892 276378
rect 5982 276326 6034 276378
rect 6046 276326 6098 276378
rect 6110 276326 6162 276378
rect 6174 276326 6226 276378
rect 4315 275782 4367 275834
rect 4379 275782 4431 275834
rect 4443 275782 4495 275834
rect 4507 275782 4559 275834
rect 7648 275782 7700 275834
rect 7712 275782 7764 275834
rect 7776 275782 7828 275834
rect 7840 275782 7892 275834
rect 2648 275238 2700 275290
rect 2712 275238 2764 275290
rect 2776 275238 2828 275290
rect 2840 275238 2892 275290
rect 5982 275238 6034 275290
rect 6046 275238 6098 275290
rect 6110 275238 6162 275290
rect 6174 275238 6226 275290
rect 4315 274694 4367 274746
rect 4379 274694 4431 274746
rect 4443 274694 4495 274746
rect 4507 274694 4559 274746
rect 7648 274694 7700 274746
rect 7712 274694 7764 274746
rect 7776 274694 7828 274746
rect 7840 274694 7892 274746
rect 2648 274150 2700 274202
rect 2712 274150 2764 274202
rect 2776 274150 2828 274202
rect 2840 274150 2892 274202
rect 5982 274150 6034 274202
rect 6046 274150 6098 274202
rect 6110 274150 6162 274202
rect 6174 274150 6226 274202
rect 4315 273606 4367 273658
rect 4379 273606 4431 273658
rect 4443 273606 4495 273658
rect 4507 273606 4559 273658
rect 7648 273606 7700 273658
rect 7712 273606 7764 273658
rect 7776 273606 7828 273658
rect 7840 273606 7892 273658
rect 2648 273062 2700 273114
rect 2712 273062 2764 273114
rect 2776 273062 2828 273114
rect 2840 273062 2892 273114
rect 5982 273062 6034 273114
rect 6046 273062 6098 273114
rect 6110 273062 6162 273114
rect 6174 273062 6226 273114
rect 4315 272518 4367 272570
rect 4379 272518 4431 272570
rect 4443 272518 4495 272570
rect 4507 272518 4559 272570
rect 7648 272518 7700 272570
rect 7712 272518 7764 272570
rect 7776 272518 7828 272570
rect 7840 272518 7892 272570
rect 2648 271974 2700 272026
rect 2712 271974 2764 272026
rect 2776 271974 2828 272026
rect 2840 271974 2892 272026
rect 5982 271974 6034 272026
rect 6046 271974 6098 272026
rect 6110 271974 6162 272026
rect 6174 271974 6226 272026
rect 4315 271430 4367 271482
rect 4379 271430 4431 271482
rect 4443 271430 4495 271482
rect 4507 271430 4559 271482
rect 7648 271430 7700 271482
rect 7712 271430 7764 271482
rect 7776 271430 7828 271482
rect 7840 271430 7892 271482
rect 2648 270886 2700 270938
rect 2712 270886 2764 270938
rect 2776 270886 2828 270938
rect 2840 270886 2892 270938
rect 5982 270886 6034 270938
rect 6046 270886 6098 270938
rect 6110 270886 6162 270938
rect 6174 270886 6226 270938
rect 4315 270342 4367 270394
rect 4379 270342 4431 270394
rect 4443 270342 4495 270394
rect 4507 270342 4559 270394
rect 7648 270342 7700 270394
rect 7712 270342 7764 270394
rect 7776 270342 7828 270394
rect 7840 270342 7892 270394
rect 2648 269798 2700 269850
rect 2712 269798 2764 269850
rect 2776 269798 2828 269850
rect 2840 269798 2892 269850
rect 5982 269798 6034 269850
rect 6046 269798 6098 269850
rect 6110 269798 6162 269850
rect 6174 269798 6226 269850
rect 4315 269254 4367 269306
rect 4379 269254 4431 269306
rect 4443 269254 4495 269306
rect 4507 269254 4559 269306
rect 7648 269254 7700 269306
rect 7712 269254 7764 269306
rect 7776 269254 7828 269306
rect 7840 269254 7892 269306
rect 2648 268710 2700 268762
rect 2712 268710 2764 268762
rect 2776 268710 2828 268762
rect 2840 268710 2892 268762
rect 5982 268710 6034 268762
rect 6046 268710 6098 268762
rect 6110 268710 6162 268762
rect 6174 268710 6226 268762
rect 4315 268166 4367 268218
rect 4379 268166 4431 268218
rect 4443 268166 4495 268218
rect 4507 268166 4559 268218
rect 7648 268166 7700 268218
rect 7712 268166 7764 268218
rect 7776 268166 7828 268218
rect 7840 268166 7892 268218
rect 2648 267622 2700 267674
rect 2712 267622 2764 267674
rect 2776 267622 2828 267674
rect 2840 267622 2892 267674
rect 5982 267622 6034 267674
rect 6046 267622 6098 267674
rect 6110 267622 6162 267674
rect 6174 267622 6226 267674
rect 4315 267078 4367 267130
rect 4379 267078 4431 267130
rect 4443 267078 4495 267130
rect 4507 267078 4559 267130
rect 7648 267078 7700 267130
rect 7712 267078 7764 267130
rect 7776 267078 7828 267130
rect 7840 267078 7892 267130
rect 2648 266534 2700 266586
rect 2712 266534 2764 266586
rect 2776 266534 2828 266586
rect 2840 266534 2892 266586
rect 5982 266534 6034 266586
rect 6046 266534 6098 266586
rect 6110 266534 6162 266586
rect 6174 266534 6226 266586
rect 4315 265990 4367 266042
rect 4379 265990 4431 266042
rect 4443 265990 4495 266042
rect 4507 265990 4559 266042
rect 7648 265990 7700 266042
rect 7712 265990 7764 266042
rect 7776 265990 7828 266042
rect 7840 265990 7892 266042
rect 2648 265446 2700 265498
rect 2712 265446 2764 265498
rect 2776 265446 2828 265498
rect 2840 265446 2892 265498
rect 5982 265446 6034 265498
rect 6046 265446 6098 265498
rect 6110 265446 6162 265498
rect 6174 265446 6226 265498
rect 4315 264902 4367 264954
rect 4379 264902 4431 264954
rect 4443 264902 4495 264954
rect 4507 264902 4559 264954
rect 7648 264902 7700 264954
rect 7712 264902 7764 264954
rect 7776 264902 7828 264954
rect 7840 264902 7892 264954
rect 2648 264358 2700 264410
rect 2712 264358 2764 264410
rect 2776 264358 2828 264410
rect 2840 264358 2892 264410
rect 5982 264358 6034 264410
rect 6046 264358 6098 264410
rect 6110 264358 6162 264410
rect 6174 264358 6226 264410
rect 4315 263814 4367 263866
rect 4379 263814 4431 263866
rect 4443 263814 4495 263866
rect 4507 263814 4559 263866
rect 7648 263814 7700 263866
rect 7712 263814 7764 263866
rect 7776 263814 7828 263866
rect 7840 263814 7892 263866
rect 2648 263270 2700 263322
rect 2712 263270 2764 263322
rect 2776 263270 2828 263322
rect 2840 263270 2892 263322
rect 5982 263270 6034 263322
rect 6046 263270 6098 263322
rect 6110 263270 6162 263322
rect 6174 263270 6226 263322
rect 4315 262726 4367 262778
rect 4379 262726 4431 262778
rect 4443 262726 4495 262778
rect 4507 262726 4559 262778
rect 7648 262726 7700 262778
rect 7712 262726 7764 262778
rect 7776 262726 7828 262778
rect 7840 262726 7892 262778
rect 2648 262182 2700 262234
rect 2712 262182 2764 262234
rect 2776 262182 2828 262234
rect 2840 262182 2892 262234
rect 5982 262182 6034 262234
rect 6046 262182 6098 262234
rect 6110 262182 6162 262234
rect 6174 262182 6226 262234
rect 4315 261638 4367 261690
rect 4379 261638 4431 261690
rect 4443 261638 4495 261690
rect 4507 261638 4559 261690
rect 7648 261638 7700 261690
rect 7712 261638 7764 261690
rect 7776 261638 7828 261690
rect 7840 261638 7892 261690
rect 2648 261094 2700 261146
rect 2712 261094 2764 261146
rect 2776 261094 2828 261146
rect 2840 261094 2892 261146
rect 5982 261094 6034 261146
rect 6046 261094 6098 261146
rect 6110 261094 6162 261146
rect 6174 261094 6226 261146
rect 4315 260550 4367 260602
rect 4379 260550 4431 260602
rect 4443 260550 4495 260602
rect 4507 260550 4559 260602
rect 7648 260550 7700 260602
rect 7712 260550 7764 260602
rect 7776 260550 7828 260602
rect 7840 260550 7892 260602
rect 2648 260006 2700 260058
rect 2712 260006 2764 260058
rect 2776 260006 2828 260058
rect 2840 260006 2892 260058
rect 5982 260006 6034 260058
rect 6046 260006 6098 260058
rect 6110 260006 6162 260058
rect 6174 260006 6226 260058
rect 4315 259462 4367 259514
rect 4379 259462 4431 259514
rect 4443 259462 4495 259514
rect 4507 259462 4559 259514
rect 7648 259462 7700 259514
rect 7712 259462 7764 259514
rect 7776 259462 7828 259514
rect 7840 259462 7892 259514
rect 2648 258918 2700 258970
rect 2712 258918 2764 258970
rect 2776 258918 2828 258970
rect 2840 258918 2892 258970
rect 5982 258918 6034 258970
rect 6046 258918 6098 258970
rect 6110 258918 6162 258970
rect 6174 258918 6226 258970
rect 4315 258374 4367 258426
rect 4379 258374 4431 258426
rect 4443 258374 4495 258426
rect 4507 258374 4559 258426
rect 7648 258374 7700 258426
rect 7712 258374 7764 258426
rect 7776 258374 7828 258426
rect 7840 258374 7892 258426
rect 2648 257830 2700 257882
rect 2712 257830 2764 257882
rect 2776 257830 2828 257882
rect 2840 257830 2892 257882
rect 5982 257830 6034 257882
rect 6046 257830 6098 257882
rect 6110 257830 6162 257882
rect 6174 257830 6226 257882
rect 4315 257286 4367 257338
rect 4379 257286 4431 257338
rect 4443 257286 4495 257338
rect 4507 257286 4559 257338
rect 7648 257286 7700 257338
rect 7712 257286 7764 257338
rect 7776 257286 7828 257338
rect 7840 257286 7892 257338
rect 2648 256742 2700 256794
rect 2712 256742 2764 256794
rect 2776 256742 2828 256794
rect 2840 256742 2892 256794
rect 5982 256742 6034 256794
rect 6046 256742 6098 256794
rect 6110 256742 6162 256794
rect 6174 256742 6226 256794
rect 4315 256198 4367 256250
rect 4379 256198 4431 256250
rect 4443 256198 4495 256250
rect 4507 256198 4559 256250
rect 7648 256198 7700 256250
rect 7712 256198 7764 256250
rect 7776 256198 7828 256250
rect 7840 256198 7892 256250
rect 2648 255654 2700 255706
rect 2712 255654 2764 255706
rect 2776 255654 2828 255706
rect 2840 255654 2892 255706
rect 5982 255654 6034 255706
rect 6046 255654 6098 255706
rect 6110 255654 6162 255706
rect 6174 255654 6226 255706
rect 4315 255110 4367 255162
rect 4379 255110 4431 255162
rect 4443 255110 4495 255162
rect 4507 255110 4559 255162
rect 7648 255110 7700 255162
rect 7712 255110 7764 255162
rect 7776 255110 7828 255162
rect 7840 255110 7892 255162
rect 2648 254566 2700 254618
rect 2712 254566 2764 254618
rect 2776 254566 2828 254618
rect 2840 254566 2892 254618
rect 5982 254566 6034 254618
rect 6046 254566 6098 254618
rect 6110 254566 6162 254618
rect 6174 254566 6226 254618
rect 4315 254022 4367 254074
rect 4379 254022 4431 254074
rect 4443 254022 4495 254074
rect 4507 254022 4559 254074
rect 7648 254022 7700 254074
rect 7712 254022 7764 254074
rect 7776 254022 7828 254074
rect 7840 254022 7892 254074
rect 2648 253478 2700 253530
rect 2712 253478 2764 253530
rect 2776 253478 2828 253530
rect 2840 253478 2892 253530
rect 5982 253478 6034 253530
rect 6046 253478 6098 253530
rect 6110 253478 6162 253530
rect 6174 253478 6226 253530
rect 4315 252934 4367 252986
rect 4379 252934 4431 252986
rect 4443 252934 4495 252986
rect 4507 252934 4559 252986
rect 7648 252934 7700 252986
rect 7712 252934 7764 252986
rect 7776 252934 7828 252986
rect 7840 252934 7892 252986
rect 2648 252390 2700 252442
rect 2712 252390 2764 252442
rect 2776 252390 2828 252442
rect 2840 252390 2892 252442
rect 5982 252390 6034 252442
rect 6046 252390 6098 252442
rect 6110 252390 6162 252442
rect 6174 252390 6226 252442
rect 4315 251846 4367 251898
rect 4379 251846 4431 251898
rect 4443 251846 4495 251898
rect 4507 251846 4559 251898
rect 7648 251846 7700 251898
rect 7712 251846 7764 251898
rect 7776 251846 7828 251898
rect 7840 251846 7892 251898
rect 2648 251302 2700 251354
rect 2712 251302 2764 251354
rect 2776 251302 2828 251354
rect 2840 251302 2892 251354
rect 5982 251302 6034 251354
rect 6046 251302 6098 251354
rect 6110 251302 6162 251354
rect 6174 251302 6226 251354
rect 4315 250758 4367 250810
rect 4379 250758 4431 250810
rect 4443 250758 4495 250810
rect 4507 250758 4559 250810
rect 7648 250758 7700 250810
rect 7712 250758 7764 250810
rect 7776 250758 7828 250810
rect 7840 250758 7892 250810
rect 2648 250214 2700 250266
rect 2712 250214 2764 250266
rect 2776 250214 2828 250266
rect 2840 250214 2892 250266
rect 5982 250214 6034 250266
rect 6046 250214 6098 250266
rect 6110 250214 6162 250266
rect 6174 250214 6226 250266
rect 4315 249670 4367 249722
rect 4379 249670 4431 249722
rect 4443 249670 4495 249722
rect 4507 249670 4559 249722
rect 7648 249670 7700 249722
rect 7712 249670 7764 249722
rect 7776 249670 7828 249722
rect 7840 249670 7892 249722
rect 2648 249126 2700 249178
rect 2712 249126 2764 249178
rect 2776 249126 2828 249178
rect 2840 249126 2892 249178
rect 5982 249126 6034 249178
rect 6046 249126 6098 249178
rect 6110 249126 6162 249178
rect 6174 249126 6226 249178
rect 4315 248582 4367 248634
rect 4379 248582 4431 248634
rect 4443 248582 4495 248634
rect 4507 248582 4559 248634
rect 7648 248582 7700 248634
rect 7712 248582 7764 248634
rect 7776 248582 7828 248634
rect 7840 248582 7892 248634
rect 2648 248038 2700 248090
rect 2712 248038 2764 248090
rect 2776 248038 2828 248090
rect 2840 248038 2892 248090
rect 5982 248038 6034 248090
rect 6046 248038 6098 248090
rect 6110 248038 6162 248090
rect 6174 248038 6226 248090
rect 4315 247494 4367 247546
rect 4379 247494 4431 247546
rect 4443 247494 4495 247546
rect 4507 247494 4559 247546
rect 7648 247494 7700 247546
rect 7712 247494 7764 247546
rect 7776 247494 7828 247546
rect 7840 247494 7892 247546
rect 2648 246950 2700 247002
rect 2712 246950 2764 247002
rect 2776 246950 2828 247002
rect 2840 246950 2892 247002
rect 5982 246950 6034 247002
rect 6046 246950 6098 247002
rect 6110 246950 6162 247002
rect 6174 246950 6226 247002
rect 4315 246406 4367 246458
rect 4379 246406 4431 246458
rect 4443 246406 4495 246458
rect 4507 246406 4559 246458
rect 7648 246406 7700 246458
rect 7712 246406 7764 246458
rect 7776 246406 7828 246458
rect 7840 246406 7892 246458
rect 2648 245862 2700 245914
rect 2712 245862 2764 245914
rect 2776 245862 2828 245914
rect 2840 245862 2892 245914
rect 5982 245862 6034 245914
rect 6046 245862 6098 245914
rect 6110 245862 6162 245914
rect 6174 245862 6226 245914
rect 4315 245318 4367 245370
rect 4379 245318 4431 245370
rect 4443 245318 4495 245370
rect 4507 245318 4559 245370
rect 7648 245318 7700 245370
rect 7712 245318 7764 245370
rect 7776 245318 7828 245370
rect 7840 245318 7892 245370
rect 2648 244774 2700 244826
rect 2712 244774 2764 244826
rect 2776 244774 2828 244826
rect 2840 244774 2892 244826
rect 5982 244774 6034 244826
rect 6046 244774 6098 244826
rect 6110 244774 6162 244826
rect 6174 244774 6226 244826
rect 2228 244715 2280 244724
rect 2228 244681 2237 244715
rect 2237 244681 2271 244715
rect 2271 244681 2280 244715
rect 2228 244672 2280 244681
rect 3516 244332 3568 244384
rect 4315 244230 4367 244282
rect 4379 244230 4431 244282
rect 4443 244230 4495 244282
rect 4507 244230 4559 244282
rect 7648 244230 7700 244282
rect 7712 244230 7764 244282
rect 7776 244230 7828 244282
rect 7840 244230 7892 244282
rect 2648 243686 2700 243738
rect 2712 243686 2764 243738
rect 2776 243686 2828 243738
rect 2840 243686 2892 243738
rect 5982 243686 6034 243738
rect 6046 243686 6098 243738
rect 6110 243686 6162 243738
rect 6174 243686 6226 243738
rect 4315 243142 4367 243194
rect 4379 243142 4431 243194
rect 4443 243142 4495 243194
rect 4507 243142 4559 243194
rect 7648 243142 7700 243194
rect 7712 243142 7764 243194
rect 7776 243142 7828 243194
rect 7840 243142 7892 243194
rect 2648 242598 2700 242650
rect 2712 242598 2764 242650
rect 2776 242598 2828 242650
rect 2840 242598 2892 242650
rect 5982 242598 6034 242650
rect 6046 242598 6098 242650
rect 6110 242598 6162 242650
rect 6174 242598 6226 242650
rect 4315 242054 4367 242106
rect 4379 242054 4431 242106
rect 4443 242054 4495 242106
rect 4507 242054 4559 242106
rect 7648 242054 7700 242106
rect 7712 242054 7764 242106
rect 7776 242054 7828 242106
rect 7840 242054 7892 242106
rect 7380 241952 7432 242004
rect 7472 241859 7524 241868
rect 7472 241825 7481 241859
rect 7481 241825 7515 241859
rect 7515 241825 7524 241859
rect 7472 241816 7524 241825
rect 2648 241510 2700 241562
rect 2712 241510 2764 241562
rect 2776 241510 2828 241562
rect 2840 241510 2892 241562
rect 5982 241510 6034 241562
rect 6046 241510 6098 241562
rect 6110 241510 6162 241562
rect 6174 241510 6226 241562
rect 7472 241111 7524 241120
rect 7472 241077 7481 241111
rect 7481 241077 7515 241111
rect 7515 241077 7524 241111
rect 7472 241068 7524 241077
rect 4315 240966 4367 241018
rect 4379 240966 4431 241018
rect 4443 240966 4495 241018
rect 4507 240966 4559 241018
rect 7648 240966 7700 241018
rect 7712 240966 7764 241018
rect 7776 240966 7828 241018
rect 7840 240966 7892 241018
rect 2648 240422 2700 240474
rect 2712 240422 2764 240474
rect 2776 240422 2828 240474
rect 2840 240422 2892 240474
rect 5982 240422 6034 240474
rect 6046 240422 6098 240474
rect 6110 240422 6162 240474
rect 6174 240422 6226 240474
rect 4315 239878 4367 239930
rect 4379 239878 4431 239930
rect 4443 239878 4495 239930
rect 4507 239878 4559 239930
rect 7648 239878 7700 239930
rect 7712 239878 7764 239930
rect 7776 239878 7828 239930
rect 7840 239878 7892 239930
rect 2648 239334 2700 239386
rect 2712 239334 2764 239386
rect 2776 239334 2828 239386
rect 2840 239334 2892 239386
rect 5982 239334 6034 239386
rect 6046 239334 6098 239386
rect 6110 239334 6162 239386
rect 6174 239334 6226 239386
rect 6368 239232 6420 239284
rect 6828 239071 6880 239080
rect 6828 239037 6837 239071
rect 6837 239037 6871 239071
rect 6871 239037 6880 239071
rect 6828 239028 6880 239037
rect 4315 238790 4367 238842
rect 4379 238790 4431 238842
rect 4443 238790 4495 238842
rect 4507 238790 4559 238842
rect 7648 238790 7700 238842
rect 7712 238790 7764 238842
rect 7776 238790 7828 238842
rect 7840 238790 7892 238842
rect 2648 238246 2700 238298
rect 2712 238246 2764 238298
rect 2776 238246 2828 238298
rect 2840 238246 2892 238298
rect 5982 238246 6034 238298
rect 6046 238246 6098 238298
rect 6110 238246 6162 238298
rect 6174 238246 6226 238298
rect 4315 237702 4367 237754
rect 4379 237702 4431 237754
rect 4443 237702 4495 237754
rect 4507 237702 4559 237754
rect 7648 237702 7700 237754
rect 7712 237702 7764 237754
rect 7776 237702 7828 237754
rect 7840 237702 7892 237754
rect 2504 237507 2556 237516
rect 2504 237473 2513 237507
rect 2513 237473 2547 237507
rect 2547 237473 2556 237507
rect 2504 237464 2556 237473
rect 2964 237396 3016 237448
rect 3516 237260 3568 237312
rect 2648 237158 2700 237210
rect 2712 237158 2764 237210
rect 2776 237158 2828 237210
rect 2840 237158 2892 237210
rect 5982 237158 6034 237210
rect 6046 237158 6098 237210
rect 6110 237158 6162 237210
rect 6174 237158 6226 237210
rect 2504 237099 2556 237108
rect 2504 237065 2513 237099
rect 2513 237065 2547 237099
rect 2547 237065 2556 237099
rect 2504 237056 2556 237065
rect 2964 236759 3016 236768
rect 2964 236725 2973 236759
rect 2973 236725 3007 236759
rect 3007 236725 3016 236759
rect 2964 236716 3016 236725
rect 3792 236716 3844 236768
rect 4315 236614 4367 236666
rect 4379 236614 4431 236666
rect 4443 236614 4495 236666
rect 4507 236614 4559 236666
rect 7648 236614 7700 236666
rect 7712 236614 7764 236666
rect 7776 236614 7828 236666
rect 7840 236614 7892 236666
rect 2648 236070 2700 236122
rect 2712 236070 2764 236122
rect 2776 236070 2828 236122
rect 2840 236070 2892 236122
rect 5982 236070 6034 236122
rect 6046 236070 6098 236122
rect 6110 236070 6162 236122
rect 6174 236070 6226 236122
rect 4315 235526 4367 235578
rect 4379 235526 4431 235578
rect 4443 235526 4495 235578
rect 4507 235526 4559 235578
rect 7648 235526 7700 235578
rect 7712 235526 7764 235578
rect 7776 235526 7828 235578
rect 7840 235526 7892 235578
rect 2648 234982 2700 235034
rect 2712 234982 2764 235034
rect 2776 234982 2828 235034
rect 2840 234982 2892 235034
rect 5982 234982 6034 235034
rect 6046 234982 6098 235034
rect 6110 234982 6162 235034
rect 6174 234982 6226 235034
rect 4315 234438 4367 234490
rect 4379 234438 4431 234490
rect 4443 234438 4495 234490
rect 4507 234438 4559 234490
rect 7648 234438 7700 234490
rect 7712 234438 7764 234490
rect 7776 234438 7828 234490
rect 7840 234438 7892 234490
rect 4160 234268 4212 234320
rect 6736 234243 6788 234252
rect 6736 234209 6745 234243
rect 6745 234209 6779 234243
rect 6779 234209 6788 234243
rect 6736 234200 6788 234209
rect 3976 234132 4028 234184
rect 6920 234175 6972 234184
rect 6920 234141 6929 234175
rect 6929 234141 6963 234175
rect 6963 234141 6972 234175
rect 6920 234132 6972 234141
rect 4988 234039 5040 234048
rect 4988 234005 4997 234039
rect 4997 234005 5031 234039
rect 5031 234005 5040 234039
rect 4988 233996 5040 234005
rect 7472 233996 7524 234048
rect 8208 233996 8260 234048
rect 2648 233894 2700 233946
rect 2712 233894 2764 233946
rect 2776 233894 2828 233946
rect 2840 233894 2892 233946
rect 5982 233894 6034 233946
rect 6046 233894 6098 233946
rect 6110 233894 6162 233946
rect 6174 233894 6226 233946
rect 6736 233792 6788 233844
rect 3700 233724 3752 233776
rect 6828 233724 6880 233776
rect 4988 233656 5040 233708
rect 4712 233588 4764 233640
rect 5540 233588 5592 233640
rect 3976 233452 4028 233504
rect 4160 233495 4212 233504
rect 4160 233461 4169 233495
rect 4169 233461 4203 233495
rect 4203 233461 4212 233495
rect 4160 233452 4212 233461
rect 5356 233452 5408 233504
rect 6920 233452 6972 233504
rect 4315 233350 4367 233402
rect 4379 233350 4431 233402
rect 4443 233350 4495 233402
rect 4507 233350 4559 233402
rect 7648 233350 7700 233402
rect 7712 233350 7764 233402
rect 7776 233350 7828 233402
rect 7840 233350 7892 233402
rect 4712 233248 4764 233300
rect 4988 233248 5040 233300
rect 2648 232806 2700 232858
rect 2712 232806 2764 232858
rect 2776 232806 2828 232858
rect 2840 232806 2892 232858
rect 5982 232806 6034 232858
rect 6046 232806 6098 232858
rect 6110 232806 6162 232858
rect 6174 232806 6226 232858
rect 3792 232747 3844 232756
rect 3792 232713 3801 232747
rect 3801 232713 3835 232747
rect 3835 232713 3844 232747
rect 3792 232704 3844 232713
rect 2964 232500 3016 232552
rect 4068 232432 4120 232484
rect 4160 232432 4212 232484
rect 4315 232262 4367 232314
rect 4379 232262 4431 232314
rect 4443 232262 4495 232314
rect 4507 232262 4559 232314
rect 7648 232262 7700 232314
rect 7712 232262 7764 232314
rect 7776 232262 7828 232314
rect 7840 232262 7892 232314
rect 2964 231863 3016 231872
rect 2964 231829 2973 231863
rect 2973 231829 3007 231863
rect 3007 231829 3016 231863
rect 2964 231820 3016 231829
rect 2648 231718 2700 231770
rect 2712 231718 2764 231770
rect 2776 231718 2828 231770
rect 2840 231718 2892 231770
rect 5982 231718 6034 231770
rect 6046 231718 6098 231770
rect 6110 231718 6162 231770
rect 6174 231718 6226 231770
rect 4315 231174 4367 231226
rect 4379 231174 4431 231226
rect 4443 231174 4495 231226
rect 4507 231174 4559 231226
rect 7648 231174 7700 231226
rect 7712 231174 7764 231226
rect 7776 231174 7828 231226
rect 7840 231174 7892 231226
rect 4712 231072 4764 231124
rect 5356 231115 5408 231124
rect 5356 231081 5365 231115
rect 5365 231081 5399 231115
rect 5399 231081 5408 231115
rect 5356 231072 5408 231081
rect 4068 231004 4120 231056
rect 4988 230868 5040 230920
rect 3792 230732 3844 230784
rect 2648 230630 2700 230682
rect 2712 230630 2764 230682
rect 2776 230630 2828 230682
rect 2840 230630 2892 230682
rect 5982 230630 6034 230682
rect 6046 230630 6098 230682
rect 6110 230630 6162 230682
rect 6174 230630 6226 230682
rect 4068 230460 4120 230512
rect 3424 230324 3476 230376
rect 3792 230324 3844 230376
rect 2412 230231 2464 230240
rect 2412 230197 2421 230231
rect 2421 230197 2455 230231
rect 2455 230197 2464 230231
rect 2412 230188 2464 230197
rect 3976 230188 4028 230240
rect 4712 230231 4764 230240
rect 4712 230197 4721 230231
rect 4721 230197 4755 230231
rect 4755 230197 4764 230231
rect 4712 230188 4764 230197
rect 4988 230231 5040 230240
rect 4988 230197 4997 230231
rect 4997 230197 5031 230231
rect 5031 230197 5040 230231
rect 4988 230188 5040 230197
rect 4315 230086 4367 230138
rect 4379 230086 4431 230138
rect 4443 230086 4495 230138
rect 4507 230086 4559 230138
rect 7648 230086 7700 230138
rect 7712 230086 7764 230138
rect 7776 230086 7828 230138
rect 7840 230086 7892 230138
rect 3424 229984 3476 230036
rect 1492 229916 1544 229968
rect 3792 229916 3844 229968
rect 4068 229891 4120 229900
rect 4068 229857 4077 229891
rect 4077 229857 4111 229891
rect 4111 229857 4120 229891
rect 4068 229848 4120 229857
rect 3056 229712 3108 229764
rect 5080 229848 5132 229900
rect 4620 229780 4672 229832
rect 5356 229712 5408 229764
rect 2504 229644 2556 229696
rect 3792 229644 3844 229696
rect 2648 229542 2700 229594
rect 2712 229542 2764 229594
rect 2776 229542 2828 229594
rect 2840 229542 2892 229594
rect 5982 229542 6034 229594
rect 6046 229542 6098 229594
rect 6110 229542 6162 229594
rect 6174 229542 6226 229594
rect 3424 229440 3476 229492
rect 5356 229483 5408 229492
rect 5356 229449 5365 229483
rect 5365 229449 5399 229483
rect 5399 229449 5408 229483
rect 5356 229440 5408 229449
rect 5080 229415 5132 229424
rect 5080 229381 5089 229415
rect 5089 229381 5123 229415
rect 5123 229381 5132 229415
rect 5080 229372 5132 229381
rect 2412 229304 2464 229356
rect 4988 229304 5040 229356
rect 3424 229236 3476 229288
rect 3792 229236 3844 229288
rect 3608 229168 3660 229220
rect 2412 229143 2464 229152
rect 2412 229109 2421 229143
rect 2421 229109 2455 229143
rect 2455 229109 2464 229143
rect 2412 229100 2464 229109
rect 4068 229100 4120 229152
rect 4804 229100 4856 229152
rect 4315 228998 4367 229050
rect 4379 228998 4431 229050
rect 4443 228998 4495 229050
rect 4507 228998 4559 229050
rect 7648 228998 7700 229050
rect 7712 228998 7764 229050
rect 7776 228998 7828 229050
rect 7840 228998 7892 229050
rect 3056 228896 3108 228948
rect 3424 228939 3476 228948
rect 3424 228905 3433 228939
rect 3433 228905 3467 228939
rect 3467 228905 3476 228939
rect 3424 228896 3476 228905
rect 2504 228828 2556 228880
rect 1492 228760 1544 228812
rect 1768 228692 1820 228744
rect 2412 228735 2464 228744
rect 2412 228701 2421 228735
rect 2421 228701 2455 228735
rect 2455 228701 2464 228735
rect 4804 228760 4856 228812
rect 3148 228735 3200 228744
rect 2412 228692 2464 228701
rect 3148 228701 3157 228735
rect 3157 228701 3191 228735
rect 3191 228701 3200 228735
rect 3148 228692 3200 228701
rect 2412 228556 2464 228608
rect 2648 228454 2700 228506
rect 2712 228454 2764 228506
rect 2776 228454 2828 228506
rect 2840 228454 2892 228506
rect 5982 228454 6034 228506
rect 6046 228454 6098 228506
rect 6110 228454 6162 228506
rect 6174 228454 6226 228506
rect 1492 228352 1544 228404
rect 2044 228395 2096 228404
rect 2044 228361 2053 228395
rect 2053 228361 2087 228395
rect 2087 228361 2096 228395
rect 2044 228352 2096 228361
rect 1216 228284 1268 228336
rect 1768 228055 1820 228064
rect 1768 228021 1777 228055
rect 1777 228021 1811 228055
rect 1811 228021 1820 228055
rect 1768 228012 1820 228021
rect 2320 228012 2372 228064
rect 3240 228284 3292 228336
rect 2964 228216 3016 228268
rect 3056 228148 3108 228200
rect 2964 228123 3016 228132
rect 2964 228089 2973 228123
rect 2973 228089 3007 228123
rect 3007 228089 3016 228123
rect 2964 228080 3016 228089
rect 3240 228055 3292 228064
rect 3240 228021 3249 228055
rect 3249 228021 3283 228055
rect 3283 228021 3292 228055
rect 3240 228012 3292 228021
rect 4804 228012 4856 228064
rect 4315 227910 4367 227962
rect 4379 227910 4431 227962
rect 4443 227910 4495 227962
rect 4507 227910 4559 227962
rect 7648 227910 7700 227962
rect 7712 227910 7764 227962
rect 7776 227910 7828 227962
rect 7840 227910 7892 227962
rect 2964 227808 3016 227860
rect 3424 227808 3476 227860
rect 2044 227672 2096 227724
rect 3056 227468 3108 227520
rect 3332 227511 3384 227520
rect 3332 227477 3341 227511
rect 3341 227477 3375 227511
rect 3375 227477 3384 227511
rect 3332 227468 3384 227477
rect 3608 227468 3660 227520
rect 2648 227366 2700 227418
rect 2712 227366 2764 227418
rect 2776 227366 2828 227418
rect 2840 227366 2892 227418
rect 5982 227366 6034 227418
rect 6046 227366 6098 227418
rect 6110 227366 6162 227418
rect 6174 227366 6226 227418
rect 2044 227307 2096 227316
rect 2044 227273 2053 227307
rect 2053 227273 2087 227307
rect 2087 227273 2096 227307
rect 2044 227264 2096 227273
rect 2320 227307 2372 227316
rect 2320 227273 2329 227307
rect 2329 227273 2363 227307
rect 2363 227273 2372 227307
rect 2320 227264 2372 227273
rect 2320 227128 2372 227180
rect 3240 227060 3292 227112
rect 3424 227060 3476 227112
rect 3056 226924 3108 226976
rect 3608 226992 3660 227044
rect 4068 226967 4120 226976
rect 4068 226933 4077 226967
rect 4077 226933 4111 226967
rect 4111 226933 4120 226967
rect 4068 226924 4120 226933
rect 4315 226822 4367 226874
rect 4379 226822 4431 226874
rect 4443 226822 4495 226874
rect 4507 226822 4559 226874
rect 7648 226822 7700 226874
rect 7712 226822 7764 226874
rect 7776 226822 7828 226874
rect 7840 226822 7892 226874
rect 3424 226763 3476 226772
rect 3424 226729 3433 226763
rect 3433 226729 3467 226763
rect 3467 226729 3476 226763
rect 3424 226720 3476 226729
rect 4712 226720 4764 226772
rect 2412 226695 2464 226704
rect 2412 226661 2421 226695
rect 2421 226661 2455 226695
rect 2455 226661 2464 226695
rect 2412 226652 2464 226661
rect 2320 226584 2372 226636
rect 4620 226584 4672 226636
rect 5816 226380 5868 226432
rect 2648 226278 2700 226330
rect 2712 226278 2764 226330
rect 2776 226278 2828 226330
rect 2840 226278 2892 226330
rect 5982 226278 6034 226330
rect 6046 226278 6098 226330
rect 6110 226278 6162 226330
rect 6174 226278 6226 226330
rect 2320 226176 2372 226228
rect 3148 226176 3200 226228
rect 4620 226176 4672 226228
rect 4712 225904 4764 225956
rect 7012 225836 7064 225888
rect 4315 225734 4367 225786
rect 4379 225734 4431 225786
rect 4443 225734 4495 225786
rect 4507 225734 4559 225786
rect 7648 225734 7700 225786
rect 7712 225734 7764 225786
rect 7776 225734 7828 225786
rect 7840 225734 7892 225786
rect 4712 225632 4764 225684
rect 4068 225496 4120 225548
rect 6276 225539 6328 225548
rect 6276 225505 6285 225539
rect 6285 225505 6319 225539
rect 6319 225505 6328 225539
rect 6276 225496 6328 225505
rect 5816 225428 5868 225480
rect 5356 225335 5408 225344
rect 5356 225301 5365 225335
rect 5365 225301 5399 225335
rect 5399 225301 5408 225335
rect 5356 225292 5408 225301
rect 5632 225292 5684 225344
rect 2648 225190 2700 225242
rect 2712 225190 2764 225242
rect 2776 225190 2828 225242
rect 2840 225190 2892 225242
rect 5982 225190 6034 225242
rect 6046 225190 6098 225242
rect 6110 225190 6162 225242
rect 6174 225190 6226 225242
rect 4068 225088 4120 225140
rect 5816 225088 5868 225140
rect 6276 225131 6328 225140
rect 6276 225097 6285 225131
rect 6285 225097 6319 225131
rect 6319 225097 6328 225131
rect 6276 225088 6328 225097
rect 3976 225020 4028 225072
rect 4712 225020 4764 225072
rect 6920 224952 6972 225004
rect 8300 224952 8352 225004
rect 7012 224927 7064 224936
rect 7012 224893 7021 224927
rect 7021 224893 7055 224927
rect 7055 224893 7064 224927
rect 7012 224884 7064 224893
rect 8024 224748 8076 224800
rect 4315 224646 4367 224698
rect 4379 224646 4431 224698
rect 4443 224646 4495 224698
rect 4507 224646 4559 224698
rect 7648 224646 7700 224698
rect 7712 224646 7764 224698
rect 7776 224646 7828 224698
rect 7840 224646 7892 224698
rect 1768 224544 1820 224596
rect 2504 224544 2556 224596
rect 6920 224587 6972 224596
rect 6920 224553 6929 224587
rect 6929 224553 6963 224587
rect 6963 224553 6972 224587
rect 6920 224544 6972 224553
rect 7012 224544 7064 224596
rect 5448 224408 5500 224460
rect 5816 224451 5868 224460
rect 5816 224417 5825 224451
rect 5825 224417 5859 224451
rect 5859 224417 5868 224451
rect 5816 224408 5868 224417
rect 5356 224340 5408 224392
rect 6276 224340 6328 224392
rect 6552 224204 6604 224256
rect 2648 224102 2700 224154
rect 2712 224102 2764 224154
rect 2776 224102 2828 224154
rect 2840 224102 2892 224154
rect 5982 224102 6034 224154
rect 6046 224102 6098 224154
rect 6110 224102 6162 224154
rect 6174 224102 6226 224154
rect 2320 224000 2372 224052
rect 5816 224043 5868 224052
rect 5816 224009 5825 224043
rect 5825 224009 5859 224043
rect 5859 224009 5868 224043
rect 5816 224000 5868 224009
rect 6276 224043 6328 224052
rect 6276 224009 6285 224043
rect 6285 224009 6319 224043
rect 6319 224009 6328 224043
rect 6276 224000 6328 224009
rect 2964 223864 3016 223916
rect 2504 223796 2556 223848
rect 3240 223839 3292 223848
rect 3240 223805 3249 223839
rect 3249 223805 3283 223839
rect 3283 223805 3292 223839
rect 3240 223796 3292 223805
rect 3424 223839 3476 223848
rect 3424 223805 3433 223839
rect 3433 223805 3467 223839
rect 3467 223805 3476 223839
rect 3424 223796 3476 223805
rect 3056 223728 3108 223780
rect 3148 223660 3200 223712
rect 4315 223558 4367 223610
rect 4379 223558 4431 223610
rect 4443 223558 4495 223610
rect 4507 223558 4559 223610
rect 7648 223558 7700 223610
rect 7712 223558 7764 223610
rect 7776 223558 7828 223610
rect 7840 223558 7892 223610
rect 3056 223456 3108 223508
rect 3424 223456 3476 223508
rect 2648 223014 2700 223066
rect 2712 223014 2764 223066
rect 2776 223014 2828 223066
rect 2840 223014 2892 223066
rect 5982 223014 6034 223066
rect 6046 223014 6098 223066
rect 6110 223014 6162 223066
rect 6174 223014 6226 223066
rect 4315 222470 4367 222522
rect 4379 222470 4431 222522
rect 4443 222470 4495 222522
rect 4507 222470 4559 222522
rect 7648 222470 7700 222522
rect 7712 222470 7764 222522
rect 7776 222470 7828 222522
rect 7840 222470 7892 222522
rect 3056 222411 3108 222420
rect 3056 222377 3065 222411
rect 3065 222377 3099 222411
rect 3099 222377 3108 222411
rect 3056 222368 3108 222377
rect 2648 221926 2700 221978
rect 2712 221926 2764 221978
rect 2776 221926 2828 221978
rect 2840 221926 2892 221978
rect 5982 221926 6034 221978
rect 6046 221926 6098 221978
rect 6110 221926 6162 221978
rect 6174 221926 6226 221978
rect 2504 221867 2556 221876
rect 2504 221833 2513 221867
rect 2513 221833 2547 221867
rect 2547 221833 2556 221867
rect 2504 221824 2556 221833
rect 2964 221824 3016 221876
rect 3240 221756 3292 221808
rect 3056 221688 3108 221740
rect 2504 221620 2556 221672
rect 2964 221552 3016 221604
rect 3332 221595 3384 221604
rect 3332 221561 3341 221595
rect 3341 221561 3375 221595
rect 3375 221561 3384 221595
rect 3332 221552 3384 221561
rect 3700 221595 3752 221604
rect 3700 221561 3709 221595
rect 3709 221561 3743 221595
rect 3743 221561 3752 221595
rect 3700 221552 3752 221561
rect 4315 221382 4367 221434
rect 4379 221382 4431 221434
rect 4443 221382 4495 221434
rect 4507 221382 4559 221434
rect 7648 221382 7700 221434
rect 7712 221382 7764 221434
rect 7776 221382 7828 221434
rect 7840 221382 7892 221434
rect 1400 220940 1452 220992
rect 3332 220940 3384 220992
rect 2648 220838 2700 220890
rect 2712 220838 2764 220890
rect 2776 220838 2828 220890
rect 2840 220838 2892 220890
rect 5982 220838 6034 220890
rect 6046 220838 6098 220890
rect 6110 220838 6162 220890
rect 6174 220838 6226 220890
rect 4315 220294 4367 220346
rect 4379 220294 4431 220346
rect 4443 220294 4495 220346
rect 4507 220294 4559 220346
rect 7648 220294 7700 220346
rect 7712 220294 7764 220346
rect 7776 220294 7828 220346
rect 7840 220294 7892 220346
rect 2648 219750 2700 219802
rect 2712 219750 2764 219802
rect 2776 219750 2828 219802
rect 2840 219750 2892 219802
rect 5982 219750 6034 219802
rect 6046 219750 6098 219802
rect 6110 219750 6162 219802
rect 6174 219750 6226 219802
rect 4315 219206 4367 219258
rect 4379 219206 4431 219258
rect 4443 219206 4495 219258
rect 4507 219206 4559 219258
rect 7648 219206 7700 219258
rect 7712 219206 7764 219258
rect 7776 219206 7828 219258
rect 7840 219206 7892 219258
rect 2648 218662 2700 218714
rect 2712 218662 2764 218714
rect 2776 218662 2828 218714
rect 2840 218662 2892 218714
rect 5982 218662 6034 218714
rect 6046 218662 6098 218714
rect 6110 218662 6162 218714
rect 6174 218662 6226 218714
rect 4315 218118 4367 218170
rect 4379 218118 4431 218170
rect 4443 218118 4495 218170
rect 4507 218118 4559 218170
rect 7648 218118 7700 218170
rect 7712 218118 7764 218170
rect 7776 218118 7828 218170
rect 7840 218118 7892 218170
rect 2648 217574 2700 217626
rect 2712 217574 2764 217626
rect 2776 217574 2828 217626
rect 2840 217574 2892 217626
rect 5982 217574 6034 217626
rect 6046 217574 6098 217626
rect 6110 217574 6162 217626
rect 6174 217574 6226 217626
rect 4315 217030 4367 217082
rect 4379 217030 4431 217082
rect 4443 217030 4495 217082
rect 4507 217030 4559 217082
rect 7648 217030 7700 217082
rect 7712 217030 7764 217082
rect 7776 217030 7828 217082
rect 7840 217030 7892 217082
rect 2648 216486 2700 216538
rect 2712 216486 2764 216538
rect 2776 216486 2828 216538
rect 2840 216486 2892 216538
rect 5982 216486 6034 216538
rect 6046 216486 6098 216538
rect 6110 216486 6162 216538
rect 6174 216486 6226 216538
rect 4315 215942 4367 215994
rect 4379 215942 4431 215994
rect 4443 215942 4495 215994
rect 4507 215942 4559 215994
rect 7648 215942 7700 215994
rect 7712 215942 7764 215994
rect 7776 215942 7828 215994
rect 7840 215942 7892 215994
rect 2648 215398 2700 215450
rect 2712 215398 2764 215450
rect 2776 215398 2828 215450
rect 2840 215398 2892 215450
rect 5982 215398 6034 215450
rect 6046 215398 6098 215450
rect 6110 215398 6162 215450
rect 6174 215398 6226 215450
rect 3700 215160 3752 215212
rect 3332 214956 3384 215008
rect 3976 214999 4028 215008
rect 3976 214965 3985 214999
rect 3985 214965 4019 214999
rect 4019 214965 4028 214999
rect 3976 214956 4028 214965
rect 4620 214956 4672 215008
rect 4315 214854 4367 214906
rect 4379 214854 4431 214906
rect 4443 214854 4495 214906
rect 4507 214854 4559 214906
rect 7648 214854 7700 214906
rect 7712 214854 7764 214906
rect 7776 214854 7828 214906
rect 7840 214854 7892 214906
rect 3700 214795 3752 214804
rect 3700 214761 3709 214795
rect 3709 214761 3743 214795
rect 3743 214761 3752 214795
rect 3700 214752 3752 214761
rect 2648 214310 2700 214362
rect 2712 214310 2764 214362
rect 2776 214310 2828 214362
rect 2840 214310 2892 214362
rect 5982 214310 6034 214362
rect 6046 214310 6098 214362
rect 6110 214310 6162 214362
rect 6174 214310 6226 214362
rect 7288 214208 7340 214260
rect 6736 214004 6788 214056
rect 4315 213766 4367 213818
rect 4379 213766 4431 213818
rect 4443 213766 4495 213818
rect 4507 213766 4559 213818
rect 7648 213766 7700 213818
rect 7712 213766 7764 213818
rect 7776 213766 7828 213818
rect 7840 213766 7892 213818
rect 2648 213222 2700 213274
rect 2712 213222 2764 213274
rect 2776 213222 2828 213274
rect 2840 213222 2892 213274
rect 5982 213222 6034 213274
rect 6046 213222 6098 213274
rect 6110 213222 6162 213274
rect 6174 213222 6226 213274
rect 4315 212678 4367 212730
rect 4379 212678 4431 212730
rect 4443 212678 4495 212730
rect 4507 212678 4559 212730
rect 7648 212678 7700 212730
rect 7712 212678 7764 212730
rect 7776 212678 7828 212730
rect 7840 212678 7892 212730
rect 2648 212134 2700 212186
rect 2712 212134 2764 212186
rect 2776 212134 2828 212186
rect 2840 212134 2892 212186
rect 5982 212134 6034 212186
rect 6046 212134 6098 212186
rect 6110 212134 6162 212186
rect 6174 212134 6226 212186
rect 112 212032 164 212084
rect 4620 211939 4672 211948
rect 4620 211905 4629 211939
rect 4629 211905 4663 211939
rect 4663 211905 4672 211939
rect 4620 211896 4672 211905
rect 6736 211692 6788 211744
rect 4315 211590 4367 211642
rect 4379 211590 4431 211642
rect 4443 211590 4495 211642
rect 4507 211590 4559 211642
rect 7648 211590 7700 211642
rect 7712 211590 7764 211642
rect 7776 211590 7828 211642
rect 7840 211590 7892 211642
rect 4620 211488 4672 211540
rect 2648 211046 2700 211098
rect 2712 211046 2764 211098
rect 2776 211046 2828 211098
rect 2840 211046 2892 211098
rect 5982 211046 6034 211098
rect 6046 211046 6098 211098
rect 6110 211046 6162 211098
rect 6174 211046 6226 211098
rect 7012 210987 7064 210996
rect 7012 210953 7021 210987
rect 7021 210953 7055 210987
rect 7055 210953 7064 210987
rect 7012 210944 7064 210953
rect 3884 210740 3936 210792
rect 4315 210502 4367 210554
rect 4379 210502 4431 210554
rect 4443 210502 4495 210554
rect 4507 210502 4559 210554
rect 7648 210502 7700 210554
rect 7712 210502 7764 210554
rect 7776 210502 7828 210554
rect 7840 210502 7892 210554
rect 2648 209958 2700 210010
rect 2712 209958 2764 210010
rect 2776 209958 2828 210010
rect 2840 209958 2892 210010
rect 5982 209958 6034 210010
rect 6046 209958 6098 210010
rect 6110 209958 6162 210010
rect 6174 209958 6226 210010
rect 3884 209856 3936 209908
rect 20 209516 72 209568
rect 2964 209652 3016 209704
rect 4315 209414 4367 209466
rect 4379 209414 4431 209466
rect 4443 209414 4495 209466
rect 4507 209414 4559 209466
rect 7648 209414 7700 209466
rect 7712 209414 7764 209466
rect 7776 209414 7828 209466
rect 7840 209414 7892 209466
rect 2964 208972 3016 209024
rect 3700 208972 3752 209024
rect 2648 208870 2700 208922
rect 2712 208870 2764 208922
rect 2776 208870 2828 208922
rect 2840 208870 2892 208922
rect 5982 208870 6034 208922
rect 6046 208870 6098 208922
rect 6110 208870 6162 208922
rect 6174 208870 6226 208922
rect 3700 208811 3752 208820
rect 3700 208777 3709 208811
rect 3709 208777 3743 208811
rect 3743 208777 3752 208811
rect 3700 208768 3752 208777
rect 3148 208632 3200 208684
rect 2964 208496 3016 208548
rect 3332 208496 3384 208548
rect 4315 208326 4367 208378
rect 4379 208326 4431 208378
rect 4443 208326 4495 208378
rect 4507 208326 4559 208378
rect 7648 208326 7700 208378
rect 7712 208326 7764 208378
rect 7776 208326 7828 208378
rect 7840 208326 7892 208378
rect 3148 208224 3200 208276
rect 2648 207782 2700 207834
rect 2712 207782 2764 207834
rect 2776 207782 2828 207834
rect 2840 207782 2892 207834
rect 5982 207782 6034 207834
rect 6046 207782 6098 207834
rect 6110 207782 6162 207834
rect 6174 207782 6226 207834
rect 4315 207238 4367 207290
rect 4379 207238 4431 207290
rect 4443 207238 4495 207290
rect 4507 207238 4559 207290
rect 7648 207238 7700 207290
rect 7712 207238 7764 207290
rect 7776 207238 7828 207290
rect 7840 207238 7892 207290
rect 2648 206694 2700 206746
rect 2712 206694 2764 206746
rect 2776 206694 2828 206746
rect 2840 206694 2892 206746
rect 5982 206694 6034 206746
rect 6046 206694 6098 206746
rect 6110 206694 6162 206746
rect 6174 206694 6226 206746
rect 4315 206150 4367 206202
rect 4379 206150 4431 206202
rect 4443 206150 4495 206202
rect 4507 206150 4559 206202
rect 7648 206150 7700 206202
rect 7712 206150 7764 206202
rect 7776 206150 7828 206202
rect 7840 206150 7892 206202
rect 2648 205606 2700 205658
rect 2712 205606 2764 205658
rect 2776 205606 2828 205658
rect 2840 205606 2892 205658
rect 5982 205606 6034 205658
rect 6046 205606 6098 205658
rect 6110 205606 6162 205658
rect 6174 205606 6226 205658
rect 4315 205062 4367 205114
rect 4379 205062 4431 205114
rect 4443 205062 4495 205114
rect 4507 205062 4559 205114
rect 7648 205062 7700 205114
rect 7712 205062 7764 205114
rect 7776 205062 7828 205114
rect 7840 205062 7892 205114
rect 2648 204518 2700 204570
rect 2712 204518 2764 204570
rect 2776 204518 2828 204570
rect 2840 204518 2892 204570
rect 5982 204518 6034 204570
rect 6046 204518 6098 204570
rect 6110 204518 6162 204570
rect 6174 204518 6226 204570
rect 4315 203974 4367 204026
rect 4379 203974 4431 204026
rect 4443 203974 4495 204026
rect 4507 203974 4559 204026
rect 7648 203974 7700 204026
rect 7712 203974 7764 204026
rect 7776 203974 7828 204026
rect 7840 203974 7892 204026
rect 2648 203430 2700 203482
rect 2712 203430 2764 203482
rect 2776 203430 2828 203482
rect 2840 203430 2892 203482
rect 5982 203430 6034 203482
rect 6046 203430 6098 203482
rect 6110 203430 6162 203482
rect 6174 203430 6226 203482
rect 4315 202886 4367 202938
rect 4379 202886 4431 202938
rect 4443 202886 4495 202938
rect 4507 202886 4559 202938
rect 7648 202886 7700 202938
rect 7712 202886 7764 202938
rect 7776 202886 7828 202938
rect 7840 202886 7892 202938
rect 2648 202342 2700 202394
rect 2712 202342 2764 202394
rect 2776 202342 2828 202394
rect 2840 202342 2892 202394
rect 5982 202342 6034 202394
rect 6046 202342 6098 202394
rect 6110 202342 6162 202394
rect 6174 202342 6226 202394
rect 4315 201798 4367 201850
rect 4379 201798 4431 201850
rect 4443 201798 4495 201850
rect 4507 201798 4559 201850
rect 7648 201798 7700 201850
rect 7712 201798 7764 201850
rect 7776 201798 7828 201850
rect 7840 201798 7892 201850
rect 2648 201254 2700 201306
rect 2712 201254 2764 201306
rect 2776 201254 2828 201306
rect 2840 201254 2892 201306
rect 5982 201254 6034 201306
rect 6046 201254 6098 201306
rect 6110 201254 6162 201306
rect 6174 201254 6226 201306
rect 4315 200710 4367 200762
rect 4379 200710 4431 200762
rect 4443 200710 4495 200762
rect 4507 200710 4559 200762
rect 7648 200710 7700 200762
rect 7712 200710 7764 200762
rect 7776 200710 7828 200762
rect 7840 200710 7892 200762
rect 2648 200166 2700 200218
rect 2712 200166 2764 200218
rect 2776 200166 2828 200218
rect 2840 200166 2892 200218
rect 5982 200166 6034 200218
rect 6046 200166 6098 200218
rect 6110 200166 6162 200218
rect 6174 200166 6226 200218
rect 4315 199622 4367 199674
rect 4379 199622 4431 199674
rect 4443 199622 4495 199674
rect 4507 199622 4559 199674
rect 7648 199622 7700 199674
rect 7712 199622 7764 199674
rect 7776 199622 7828 199674
rect 7840 199622 7892 199674
rect 2648 199078 2700 199130
rect 2712 199078 2764 199130
rect 2776 199078 2828 199130
rect 2840 199078 2892 199130
rect 5982 199078 6034 199130
rect 6046 199078 6098 199130
rect 6110 199078 6162 199130
rect 6174 199078 6226 199130
rect 4315 198534 4367 198586
rect 4379 198534 4431 198586
rect 4443 198534 4495 198586
rect 4507 198534 4559 198586
rect 7648 198534 7700 198586
rect 7712 198534 7764 198586
rect 7776 198534 7828 198586
rect 7840 198534 7892 198586
rect 2648 197990 2700 198042
rect 2712 197990 2764 198042
rect 2776 197990 2828 198042
rect 2840 197990 2892 198042
rect 5982 197990 6034 198042
rect 6046 197990 6098 198042
rect 6110 197990 6162 198042
rect 6174 197990 6226 198042
rect 4315 197446 4367 197498
rect 4379 197446 4431 197498
rect 4443 197446 4495 197498
rect 4507 197446 4559 197498
rect 7648 197446 7700 197498
rect 7712 197446 7764 197498
rect 7776 197446 7828 197498
rect 7840 197446 7892 197498
rect 2648 196902 2700 196954
rect 2712 196902 2764 196954
rect 2776 196902 2828 196954
rect 2840 196902 2892 196954
rect 5982 196902 6034 196954
rect 6046 196902 6098 196954
rect 6110 196902 6162 196954
rect 6174 196902 6226 196954
rect 4315 196358 4367 196410
rect 4379 196358 4431 196410
rect 4443 196358 4495 196410
rect 4507 196358 4559 196410
rect 7648 196358 7700 196410
rect 7712 196358 7764 196410
rect 7776 196358 7828 196410
rect 7840 196358 7892 196410
rect 2648 195814 2700 195866
rect 2712 195814 2764 195866
rect 2776 195814 2828 195866
rect 2840 195814 2892 195866
rect 5982 195814 6034 195866
rect 6046 195814 6098 195866
rect 6110 195814 6162 195866
rect 6174 195814 6226 195866
rect 4315 195270 4367 195322
rect 4379 195270 4431 195322
rect 4443 195270 4495 195322
rect 4507 195270 4559 195322
rect 7648 195270 7700 195322
rect 7712 195270 7764 195322
rect 7776 195270 7828 195322
rect 7840 195270 7892 195322
rect 2648 194726 2700 194778
rect 2712 194726 2764 194778
rect 2776 194726 2828 194778
rect 2840 194726 2892 194778
rect 5982 194726 6034 194778
rect 6046 194726 6098 194778
rect 6110 194726 6162 194778
rect 6174 194726 6226 194778
rect 4315 194182 4367 194234
rect 4379 194182 4431 194234
rect 4443 194182 4495 194234
rect 4507 194182 4559 194234
rect 7648 194182 7700 194234
rect 7712 194182 7764 194234
rect 7776 194182 7828 194234
rect 7840 194182 7892 194234
rect 2648 193638 2700 193690
rect 2712 193638 2764 193690
rect 2776 193638 2828 193690
rect 2840 193638 2892 193690
rect 5982 193638 6034 193690
rect 6046 193638 6098 193690
rect 6110 193638 6162 193690
rect 6174 193638 6226 193690
rect 4315 193094 4367 193146
rect 4379 193094 4431 193146
rect 4443 193094 4495 193146
rect 4507 193094 4559 193146
rect 7648 193094 7700 193146
rect 7712 193094 7764 193146
rect 7776 193094 7828 193146
rect 7840 193094 7892 193146
rect 2648 192550 2700 192602
rect 2712 192550 2764 192602
rect 2776 192550 2828 192602
rect 2840 192550 2892 192602
rect 5982 192550 6034 192602
rect 6046 192550 6098 192602
rect 6110 192550 6162 192602
rect 6174 192550 6226 192602
rect 4315 192006 4367 192058
rect 4379 192006 4431 192058
rect 4443 192006 4495 192058
rect 4507 192006 4559 192058
rect 7648 192006 7700 192058
rect 7712 192006 7764 192058
rect 7776 192006 7828 192058
rect 7840 192006 7892 192058
rect 2648 191462 2700 191514
rect 2712 191462 2764 191514
rect 2776 191462 2828 191514
rect 2840 191462 2892 191514
rect 5982 191462 6034 191514
rect 6046 191462 6098 191514
rect 6110 191462 6162 191514
rect 6174 191462 6226 191514
rect 4315 190918 4367 190970
rect 4379 190918 4431 190970
rect 4443 190918 4495 190970
rect 4507 190918 4559 190970
rect 7648 190918 7700 190970
rect 7712 190918 7764 190970
rect 7776 190918 7828 190970
rect 7840 190918 7892 190970
rect 2648 190374 2700 190426
rect 2712 190374 2764 190426
rect 2776 190374 2828 190426
rect 2840 190374 2892 190426
rect 5982 190374 6034 190426
rect 6046 190374 6098 190426
rect 6110 190374 6162 190426
rect 6174 190374 6226 190426
rect 4315 189830 4367 189882
rect 4379 189830 4431 189882
rect 4443 189830 4495 189882
rect 4507 189830 4559 189882
rect 7648 189830 7700 189882
rect 7712 189830 7764 189882
rect 7776 189830 7828 189882
rect 7840 189830 7892 189882
rect 2648 189286 2700 189338
rect 2712 189286 2764 189338
rect 2776 189286 2828 189338
rect 2840 189286 2892 189338
rect 5982 189286 6034 189338
rect 6046 189286 6098 189338
rect 6110 189286 6162 189338
rect 6174 189286 6226 189338
rect 4315 188742 4367 188794
rect 4379 188742 4431 188794
rect 4443 188742 4495 188794
rect 4507 188742 4559 188794
rect 7648 188742 7700 188794
rect 7712 188742 7764 188794
rect 7776 188742 7828 188794
rect 7840 188742 7892 188794
rect 2648 188198 2700 188250
rect 2712 188198 2764 188250
rect 2776 188198 2828 188250
rect 2840 188198 2892 188250
rect 5982 188198 6034 188250
rect 6046 188198 6098 188250
rect 6110 188198 6162 188250
rect 6174 188198 6226 188250
rect 4315 187654 4367 187706
rect 4379 187654 4431 187706
rect 4443 187654 4495 187706
rect 4507 187654 4559 187706
rect 7648 187654 7700 187706
rect 7712 187654 7764 187706
rect 7776 187654 7828 187706
rect 7840 187654 7892 187706
rect 2648 187110 2700 187162
rect 2712 187110 2764 187162
rect 2776 187110 2828 187162
rect 2840 187110 2892 187162
rect 5982 187110 6034 187162
rect 6046 187110 6098 187162
rect 6110 187110 6162 187162
rect 6174 187110 6226 187162
rect 4315 186566 4367 186618
rect 4379 186566 4431 186618
rect 4443 186566 4495 186618
rect 4507 186566 4559 186618
rect 7648 186566 7700 186618
rect 7712 186566 7764 186618
rect 7776 186566 7828 186618
rect 7840 186566 7892 186618
rect 2648 186022 2700 186074
rect 2712 186022 2764 186074
rect 2776 186022 2828 186074
rect 2840 186022 2892 186074
rect 5982 186022 6034 186074
rect 6046 186022 6098 186074
rect 6110 186022 6162 186074
rect 6174 186022 6226 186074
rect 4315 185478 4367 185530
rect 4379 185478 4431 185530
rect 4443 185478 4495 185530
rect 4507 185478 4559 185530
rect 7648 185478 7700 185530
rect 7712 185478 7764 185530
rect 7776 185478 7828 185530
rect 7840 185478 7892 185530
rect 2648 184934 2700 184986
rect 2712 184934 2764 184986
rect 2776 184934 2828 184986
rect 2840 184934 2892 184986
rect 5982 184934 6034 184986
rect 6046 184934 6098 184986
rect 6110 184934 6162 184986
rect 6174 184934 6226 184986
rect 4315 184390 4367 184442
rect 4379 184390 4431 184442
rect 4443 184390 4495 184442
rect 4507 184390 4559 184442
rect 7648 184390 7700 184442
rect 7712 184390 7764 184442
rect 7776 184390 7828 184442
rect 7840 184390 7892 184442
rect 2648 183846 2700 183898
rect 2712 183846 2764 183898
rect 2776 183846 2828 183898
rect 2840 183846 2892 183898
rect 5982 183846 6034 183898
rect 6046 183846 6098 183898
rect 6110 183846 6162 183898
rect 6174 183846 6226 183898
rect 4315 183302 4367 183354
rect 4379 183302 4431 183354
rect 4443 183302 4495 183354
rect 4507 183302 4559 183354
rect 7648 183302 7700 183354
rect 7712 183302 7764 183354
rect 7776 183302 7828 183354
rect 7840 183302 7892 183354
rect 2648 182758 2700 182810
rect 2712 182758 2764 182810
rect 2776 182758 2828 182810
rect 2840 182758 2892 182810
rect 5982 182758 6034 182810
rect 6046 182758 6098 182810
rect 6110 182758 6162 182810
rect 6174 182758 6226 182810
rect 4315 182214 4367 182266
rect 4379 182214 4431 182266
rect 4443 182214 4495 182266
rect 4507 182214 4559 182266
rect 7648 182214 7700 182266
rect 7712 182214 7764 182266
rect 7776 182214 7828 182266
rect 7840 182214 7892 182266
rect 2648 181670 2700 181722
rect 2712 181670 2764 181722
rect 2776 181670 2828 181722
rect 2840 181670 2892 181722
rect 5982 181670 6034 181722
rect 6046 181670 6098 181722
rect 6110 181670 6162 181722
rect 6174 181670 6226 181722
rect 4315 181126 4367 181178
rect 4379 181126 4431 181178
rect 4443 181126 4495 181178
rect 4507 181126 4559 181178
rect 7648 181126 7700 181178
rect 7712 181126 7764 181178
rect 7776 181126 7828 181178
rect 7840 181126 7892 181178
rect 2648 180582 2700 180634
rect 2712 180582 2764 180634
rect 2776 180582 2828 180634
rect 2840 180582 2892 180634
rect 5982 180582 6034 180634
rect 6046 180582 6098 180634
rect 6110 180582 6162 180634
rect 6174 180582 6226 180634
rect 4315 180038 4367 180090
rect 4379 180038 4431 180090
rect 4443 180038 4495 180090
rect 4507 180038 4559 180090
rect 7648 180038 7700 180090
rect 7712 180038 7764 180090
rect 7776 180038 7828 180090
rect 7840 180038 7892 180090
rect 2648 179494 2700 179546
rect 2712 179494 2764 179546
rect 2776 179494 2828 179546
rect 2840 179494 2892 179546
rect 5982 179494 6034 179546
rect 6046 179494 6098 179546
rect 6110 179494 6162 179546
rect 6174 179494 6226 179546
rect 4315 178950 4367 179002
rect 4379 178950 4431 179002
rect 4443 178950 4495 179002
rect 4507 178950 4559 179002
rect 7648 178950 7700 179002
rect 7712 178950 7764 179002
rect 7776 178950 7828 179002
rect 7840 178950 7892 179002
rect 2648 178406 2700 178458
rect 2712 178406 2764 178458
rect 2776 178406 2828 178458
rect 2840 178406 2892 178458
rect 5982 178406 6034 178458
rect 6046 178406 6098 178458
rect 6110 178406 6162 178458
rect 6174 178406 6226 178458
rect 4315 177862 4367 177914
rect 4379 177862 4431 177914
rect 4443 177862 4495 177914
rect 4507 177862 4559 177914
rect 7648 177862 7700 177914
rect 7712 177862 7764 177914
rect 7776 177862 7828 177914
rect 7840 177862 7892 177914
rect 2648 177318 2700 177370
rect 2712 177318 2764 177370
rect 2776 177318 2828 177370
rect 2840 177318 2892 177370
rect 5982 177318 6034 177370
rect 6046 177318 6098 177370
rect 6110 177318 6162 177370
rect 6174 177318 6226 177370
rect 4315 176774 4367 176826
rect 4379 176774 4431 176826
rect 4443 176774 4495 176826
rect 4507 176774 4559 176826
rect 7648 176774 7700 176826
rect 7712 176774 7764 176826
rect 7776 176774 7828 176826
rect 7840 176774 7892 176826
rect 2648 176230 2700 176282
rect 2712 176230 2764 176282
rect 2776 176230 2828 176282
rect 2840 176230 2892 176282
rect 5982 176230 6034 176282
rect 6046 176230 6098 176282
rect 6110 176230 6162 176282
rect 6174 176230 6226 176282
rect 4315 175686 4367 175738
rect 4379 175686 4431 175738
rect 4443 175686 4495 175738
rect 4507 175686 4559 175738
rect 7648 175686 7700 175738
rect 7712 175686 7764 175738
rect 7776 175686 7828 175738
rect 7840 175686 7892 175738
rect 2648 175142 2700 175194
rect 2712 175142 2764 175194
rect 2776 175142 2828 175194
rect 2840 175142 2892 175194
rect 5982 175142 6034 175194
rect 6046 175142 6098 175194
rect 6110 175142 6162 175194
rect 6174 175142 6226 175194
rect 4315 174598 4367 174650
rect 4379 174598 4431 174650
rect 4443 174598 4495 174650
rect 4507 174598 4559 174650
rect 7648 174598 7700 174650
rect 7712 174598 7764 174650
rect 7776 174598 7828 174650
rect 7840 174598 7892 174650
rect 2648 174054 2700 174106
rect 2712 174054 2764 174106
rect 2776 174054 2828 174106
rect 2840 174054 2892 174106
rect 5982 174054 6034 174106
rect 6046 174054 6098 174106
rect 6110 174054 6162 174106
rect 6174 174054 6226 174106
rect 4315 173510 4367 173562
rect 4379 173510 4431 173562
rect 4443 173510 4495 173562
rect 4507 173510 4559 173562
rect 7648 173510 7700 173562
rect 7712 173510 7764 173562
rect 7776 173510 7828 173562
rect 7840 173510 7892 173562
rect 2648 172966 2700 173018
rect 2712 172966 2764 173018
rect 2776 172966 2828 173018
rect 2840 172966 2892 173018
rect 5982 172966 6034 173018
rect 6046 172966 6098 173018
rect 6110 172966 6162 173018
rect 6174 172966 6226 173018
rect 4315 172422 4367 172474
rect 4379 172422 4431 172474
rect 4443 172422 4495 172474
rect 4507 172422 4559 172474
rect 7648 172422 7700 172474
rect 7712 172422 7764 172474
rect 7776 172422 7828 172474
rect 7840 172422 7892 172474
rect 6644 172320 6696 172372
rect 6552 172184 6604 172236
rect 6828 172184 6880 172236
rect 7472 172227 7524 172236
rect 7472 172193 7481 172227
rect 7481 172193 7515 172227
rect 7515 172193 7524 172227
rect 7472 172184 7524 172193
rect 2648 171878 2700 171930
rect 2712 171878 2764 171930
rect 2776 171878 2828 171930
rect 2840 171878 2892 171930
rect 5982 171878 6034 171930
rect 6046 171878 6098 171930
rect 6110 171878 6162 171930
rect 6174 171878 6226 171930
rect 7472 171819 7524 171828
rect 7472 171785 7481 171819
rect 7481 171785 7515 171819
rect 7515 171785 7524 171819
rect 7472 171776 7524 171785
rect 4315 171334 4367 171386
rect 4379 171334 4431 171386
rect 4443 171334 4495 171386
rect 4507 171334 4559 171386
rect 7648 171334 7700 171386
rect 7712 171334 7764 171386
rect 7776 171334 7828 171386
rect 7840 171334 7892 171386
rect 2648 170790 2700 170842
rect 2712 170790 2764 170842
rect 2776 170790 2828 170842
rect 2840 170790 2892 170842
rect 5982 170790 6034 170842
rect 6046 170790 6098 170842
rect 6110 170790 6162 170842
rect 6174 170790 6226 170842
rect 4315 170246 4367 170298
rect 4379 170246 4431 170298
rect 4443 170246 4495 170298
rect 4507 170246 4559 170298
rect 7648 170246 7700 170298
rect 7712 170246 7764 170298
rect 7776 170246 7828 170298
rect 7840 170246 7892 170298
rect 2648 169702 2700 169754
rect 2712 169702 2764 169754
rect 2776 169702 2828 169754
rect 2840 169702 2892 169754
rect 5982 169702 6034 169754
rect 6046 169702 6098 169754
rect 6110 169702 6162 169754
rect 6174 169702 6226 169754
rect 4315 169158 4367 169210
rect 4379 169158 4431 169210
rect 4443 169158 4495 169210
rect 4507 169158 4559 169210
rect 7648 169158 7700 169210
rect 7712 169158 7764 169210
rect 7776 169158 7828 169210
rect 7840 169158 7892 169210
rect 2648 168614 2700 168666
rect 2712 168614 2764 168666
rect 2776 168614 2828 168666
rect 2840 168614 2892 168666
rect 5982 168614 6034 168666
rect 6046 168614 6098 168666
rect 6110 168614 6162 168666
rect 6174 168614 6226 168666
rect 4315 168070 4367 168122
rect 4379 168070 4431 168122
rect 4443 168070 4495 168122
rect 4507 168070 4559 168122
rect 7648 168070 7700 168122
rect 7712 168070 7764 168122
rect 7776 168070 7828 168122
rect 7840 168070 7892 168122
rect 2648 167526 2700 167578
rect 2712 167526 2764 167578
rect 2776 167526 2828 167578
rect 2840 167526 2892 167578
rect 5982 167526 6034 167578
rect 6046 167526 6098 167578
rect 6110 167526 6162 167578
rect 6174 167526 6226 167578
rect 4315 166982 4367 167034
rect 4379 166982 4431 167034
rect 4443 166982 4495 167034
rect 4507 166982 4559 167034
rect 7648 166982 7700 167034
rect 7712 166982 7764 167034
rect 7776 166982 7828 167034
rect 7840 166982 7892 167034
rect 2648 166438 2700 166490
rect 2712 166438 2764 166490
rect 2776 166438 2828 166490
rect 2840 166438 2892 166490
rect 5982 166438 6034 166490
rect 6046 166438 6098 166490
rect 6110 166438 6162 166490
rect 6174 166438 6226 166490
rect 4315 165894 4367 165946
rect 4379 165894 4431 165946
rect 4443 165894 4495 165946
rect 4507 165894 4559 165946
rect 7648 165894 7700 165946
rect 7712 165894 7764 165946
rect 7776 165894 7828 165946
rect 7840 165894 7892 165946
rect 2648 165350 2700 165402
rect 2712 165350 2764 165402
rect 2776 165350 2828 165402
rect 2840 165350 2892 165402
rect 5982 165350 6034 165402
rect 6046 165350 6098 165402
rect 6110 165350 6162 165402
rect 6174 165350 6226 165402
rect 4315 164806 4367 164858
rect 4379 164806 4431 164858
rect 4443 164806 4495 164858
rect 4507 164806 4559 164858
rect 7648 164806 7700 164858
rect 7712 164806 7764 164858
rect 7776 164806 7828 164858
rect 7840 164806 7892 164858
rect 2648 164262 2700 164314
rect 2712 164262 2764 164314
rect 2776 164262 2828 164314
rect 2840 164262 2892 164314
rect 5982 164262 6034 164314
rect 6046 164262 6098 164314
rect 6110 164262 6162 164314
rect 6174 164262 6226 164314
rect 4315 163718 4367 163770
rect 4379 163718 4431 163770
rect 4443 163718 4495 163770
rect 4507 163718 4559 163770
rect 7648 163718 7700 163770
rect 7712 163718 7764 163770
rect 7776 163718 7828 163770
rect 7840 163718 7892 163770
rect 2648 163174 2700 163226
rect 2712 163174 2764 163226
rect 2776 163174 2828 163226
rect 2840 163174 2892 163226
rect 5982 163174 6034 163226
rect 6046 163174 6098 163226
rect 6110 163174 6162 163226
rect 6174 163174 6226 163226
rect 4315 162630 4367 162682
rect 4379 162630 4431 162682
rect 4443 162630 4495 162682
rect 4507 162630 4559 162682
rect 7648 162630 7700 162682
rect 7712 162630 7764 162682
rect 7776 162630 7828 162682
rect 7840 162630 7892 162682
rect 2648 162086 2700 162138
rect 2712 162086 2764 162138
rect 2776 162086 2828 162138
rect 2840 162086 2892 162138
rect 5982 162086 6034 162138
rect 6046 162086 6098 162138
rect 6110 162086 6162 162138
rect 6174 162086 6226 162138
rect 4315 161542 4367 161594
rect 4379 161542 4431 161594
rect 4443 161542 4495 161594
rect 4507 161542 4559 161594
rect 7648 161542 7700 161594
rect 7712 161542 7764 161594
rect 7776 161542 7828 161594
rect 7840 161542 7892 161594
rect 2648 160998 2700 161050
rect 2712 160998 2764 161050
rect 2776 160998 2828 161050
rect 2840 160998 2892 161050
rect 5982 160998 6034 161050
rect 6046 160998 6098 161050
rect 6110 160998 6162 161050
rect 6174 160998 6226 161050
rect 4315 160454 4367 160506
rect 4379 160454 4431 160506
rect 4443 160454 4495 160506
rect 4507 160454 4559 160506
rect 7648 160454 7700 160506
rect 7712 160454 7764 160506
rect 7776 160454 7828 160506
rect 7840 160454 7892 160506
rect 2648 159910 2700 159962
rect 2712 159910 2764 159962
rect 2776 159910 2828 159962
rect 2840 159910 2892 159962
rect 5982 159910 6034 159962
rect 6046 159910 6098 159962
rect 6110 159910 6162 159962
rect 6174 159910 6226 159962
rect 4315 159366 4367 159418
rect 4379 159366 4431 159418
rect 4443 159366 4495 159418
rect 4507 159366 4559 159418
rect 7648 159366 7700 159418
rect 7712 159366 7764 159418
rect 7776 159366 7828 159418
rect 7840 159366 7892 159418
rect 2648 158822 2700 158874
rect 2712 158822 2764 158874
rect 2776 158822 2828 158874
rect 2840 158822 2892 158874
rect 5982 158822 6034 158874
rect 6046 158822 6098 158874
rect 6110 158822 6162 158874
rect 6174 158822 6226 158874
rect 4315 158278 4367 158330
rect 4379 158278 4431 158330
rect 4443 158278 4495 158330
rect 4507 158278 4559 158330
rect 7648 158278 7700 158330
rect 7712 158278 7764 158330
rect 7776 158278 7828 158330
rect 7840 158278 7892 158330
rect 3424 158176 3476 158228
rect 6920 158108 6972 158160
rect 8024 158108 8076 158160
rect 4068 158083 4120 158092
rect 4068 158049 4099 158083
rect 4099 158049 4120 158083
rect 4068 158040 4120 158049
rect 2648 157734 2700 157786
rect 2712 157734 2764 157786
rect 2776 157734 2828 157786
rect 2840 157734 2892 157786
rect 5982 157734 6034 157786
rect 6046 157734 6098 157786
rect 6110 157734 6162 157786
rect 6174 157734 6226 157786
rect 4068 157675 4120 157684
rect 4068 157641 4077 157675
rect 4077 157641 4111 157675
rect 4111 157641 4120 157675
rect 4068 157632 4120 157641
rect 4315 157190 4367 157242
rect 4379 157190 4431 157242
rect 4443 157190 4495 157242
rect 4507 157190 4559 157242
rect 7648 157190 7700 157242
rect 7712 157190 7764 157242
rect 7776 157190 7828 157242
rect 7840 157190 7892 157242
rect 2648 156646 2700 156698
rect 2712 156646 2764 156698
rect 2776 156646 2828 156698
rect 2840 156646 2892 156698
rect 5982 156646 6034 156698
rect 6046 156646 6098 156698
rect 6110 156646 6162 156698
rect 6174 156646 6226 156698
rect 4315 156102 4367 156154
rect 4379 156102 4431 156154
rect 4443 156102 4495 156154
rect 4507 156102 4559 156154
rect 7648 156102 7700 156154
rect 7712 156102 7764 156154
rect 7776 156102 7828 156154
rect 7840 156102 7892 156154
rect 2648 155558 2700 155610
rect 2712 155558 2764 155610
rect 2776 155558 2828 155610
rect 2840 155558 2892 155610
rect 5982 155558 6034 155610
rect 6046 155558 6098 155610
rect 6110 155558 6162 155610
rect 6174 155558 6226 155610
rect 4315 155014 4367 155066
rect 4379 155014 4431 155066
rect 4443 155014 4495 155066
rect 4507 155014 4559 155066
rect 7648 155014 7700 155066
rect 7712 155014 7764 155066
rect 7776 155014 7828 155066
rect 7840 155014 7892 155066
rect 2648 154470 2700 154522
rect 2712 154470 2764 154522
rect 2776 154470 2828 154522
rect 2840 154470 2892 154522
rect 5982 154470 6034 154522
rect 6046 154470 6098 154522
rect 6110 154470 6162 154522
rect 6174 154470 6226 154522
rect 4315 153926 4367 153978
rect 4379 153926 4431 153978
rect 4443 153926 4495 153978
rect 4507 153926 4559 153978
rect 7648 153926 7700 153978
rect 7712 153926 7764 153978
rect 7776 153926 7828 153978
rect 7840 153926 7892 153978
rect 2648 153382 2700 153434
rect 2712 153382 2764 153434
rect 2776 153382 2828 153434
rect 2840 153382 2892 153434
rect 5982 153382 6034 153434
rect 6046 153382 6098 153434
rect 6110 153382 6162 153434
rect 6174 153382 6226 153434
rect 4315 152838 4367 152890
rect 4379 152838 4431 152890
rect 4443 152838 4495 152890
rect 4507 152838 4559 152890
rect 7648 152838 7700 152890
rect 7712 152838 7764 152890
rect 7776 152838 7828 152890
rect 7840 152838 7892 152890
rect 2648 152294 2700 152346
rect 2712 152294 2764 152346
rect 2776 152294 2828 152346
rect 2840 152294 2892 152346
rect 5982 152294 6034 152346
rect 6046 152294 6098 152346
rect 6110 152294 6162 152346
rect 6174 152294 6226 152346
rect 4315 151750 4367 151802
rect 4379 151750 4431 151802
rect 4443 151750 4495 151802
rect 4507 151750 4559 151802
rect 7648 151750 7700 151802
rect 7712 151750 7764 151802
rect 7776 151750 7828 151802
rect 7840 151750 7892 151802
rect 2648 151206 2700 151258
rect 2712 151206 2764 151258
rect 2776 151206 2828 151258
rect 2840 151206 2892 151258
rect 5982 151206 6034 151258
rect 6046 151206 6098 151258
rect 6110 151206 6162 151258
rect 6174 151206 6226 151258
rect 4315 150662 4367 150714
rect 4379 150662 4431 150714
rect 4443 150662 4495 150714
rect 4507 150662 4559 150714
rect 7648 150662 7700 150714
rect 7712 150662 7764 150714
rect 7776 150662 7828 150714
rect 7840 150662 7892 150714
rect 2648 150118 2700 150170
rect 2712 150118 2764 150170
rect 2776 150118 2828 150170
rect 2840 150118 2892 150170
rect 5982 150118 6034 150170
rect 6046 150118 6098 150170
rect 6110 150118 6162 150170
rect 6174 150118 6226 150170
rect 4315 149574 4367 149626
rect 4379 149574 4431 149626
rect 4443 149574 4495 149626
rect 4507 149574 4559 149626
rect 7648 149574 7700 149626
rect 7712 149574 7764 149626
rect 7776 149574 7828 149626
rect 7840 149574 7892 149626
rect 2648 149030 2700 149082
rect 2712 149030 2764 149082
rect 2776 149030 2828 149082
rect 2840 149030 2892 149082
rect 5982 149030 6034 149082
rect 6046 149030 6098 149082
rect 6110 149030 6162 149082
rect 6174 149030 6226 149082
rect 4315 148486 4367 148538
rect 4379 148486 4431 148538
rect 4443 148486 4495 148538
rect 4507 148486 4559 148538
rect 7648 148486 7700 148538
rect 7712 148486 7764 148538
rect 7776 148486 7828 148538
rect 7840 148486 7892 148538
rect 2648 147942 2700 147994
rect 2712 147942 2764 147994
rect 2776 147942 2828 147994
rect 2840 147942 2892 147994
rect 5982 147942 6034 147994
rect 6046 147942 6098 147994
rect 6110 147942 6162 147994
rect 6174 147942 6226 147994
rect 4315 147398 4367 147450
rect 4379 147398 4431 147450
rect 4443 147398 4495 147450
rect 4507 147398 4559 147450
rect 7648 147398 7700 147450
rect 7712 147398 7764 147450
rect 7776 147398 7828 147450
rect 7840 147398 7892 147450
rect 2648 146854 2700 146906
rect 2712 146854 2764 146906
rect 2776 146854 2828 146906
rect 2840 146854 2892 146906
rect 5982 146854 6034 146906
rect 6046 146854 6098 146906
rect 6110 146854 6162 146906
rect 6174 146854 6226 146906
rect 4315 146310 4367 146362
rect 4379 146310 4431 146362
rect 4443 146310 4495 146362
rect 4507 146310 4559 146362
rect 7648 146310 7700 146362
rect 7712 146310 7764 146362
rect 7776 146310 7828 146362
rect 7840 146310 7892 146362
rect 2648 145766 2700 145818
rect 2712 145766 2764 145818
rect 2776 145766 2828 145818
rect 2840 145766 2892 145818
rect 5982 145766 6034 145818
rect 6046 145766 6098 145818
rect 6110 145766 6162 145818
rect 6174 145766 6226 145818
rect 4315 145222 4367 145274
rect 4379 145222 4431 145274
rect 4443 145222 4495 145274
rect 4507 145222 4559 145274
rect 7648 145222 7700 145274
rect 7712 145222 7764 145274
rect 7776 145222 7828 145274
rect 7840 145222 7892 145274
rect 2648 144678 2700 144730
rect 2712 144678 2764 144730
rect 2776 144678 2828 144730
rect 2840 144678 2892 144730
rect 5982 144678 6034 144730
rect 6046 144678 6098 144730
rect 6110 144678 6162 144730
rect 6174 144678 6226 144730
rect 4315 144134 4367 144186
rect 4379 144134 4431 144186
rect 4443 144134 4495 144186
rect 4507 144134 4559 144186
rect 7648 144134 7700 144186
rect 7712 144134 7764 144186
rect 7776 144134 7828 144186
rect 7840 144134 7892 144186
rect 2648 143590 2700 143642
rect 2712 143590 2764 143642
rect 2776 143590 2828 143642
rect 2840 143590 2892 143642
rect 5982 143590 6034 143642
rect 6046 143590 6098 143642
rect 6110 143590 6162 143642
rect 6174 143590 6226 143642
rect 4315 143046 4367 143098
rect 4379 143046 4431 143098
rect 4443 143046 4495 143098
rect 4507 143046 4559 143098
rect 7648 143046 7700 143098
rect 7712 143046 7764 143098
rect 7776 143046 7828 143098
rect 7840 143046 7892 143098
rect 2648 142502 2700 142554
rect 2712 142502 2764 142554
rect 2776 142502 2828 142554
rect 2840 142502 2892 142554
rect 5982 142502 6034 142554
rect 6046 142502 6098 142554
rect 6110 142502 6162 142554
rect 6174 142502 6226 142554
rect 4315 141958 4367 142010
rect 4379 141958 4431 142010
rect 4443 141958 4495 142010
rect 4507 141958 4559 142010
rect 7648 141958 7700 142010
rect 7712 141958 7764 142010
rect 7776 141958 7828 142010
rect 7840 141958 7892 142010
rect 2648 141414 2700 141466
rect 2712 141414 2764 141466
rect 2776 141414 2828 141466
rect 2840 141414 2892 141466
rect 5982 141414 6034 141466
rect 6046 141414 6098 141466
rect 6110 141414 6162 141466
rect 6174 141414 6226 141466
rect 4315 140870 4367 140922
rect 4379 140870 4431 140922
rect 4443 140870 4495 140922
rect 4507 140870 4559 140922
rect 7648 140870 7700 140922
rect 7712 140870 7764 140922
rect 7776 140870 7828 140922
rect 7840 140870 7892 140922
rect 2648 140326 2700 140378
rect 2712 140326 2764 140378
rect 2776 140326 2828 140378
rect 2840 140326 2892 140378
rect 5982 140326 6034 140378
rect 6046 140326 6098 140378
rect 6110 140326 6162 140378
rect 6174 140326 6226 140378
rect 4315 139782 4367 139834
rect 4379 139782 4431 139834
rect 4443 139782 4495 139834
rect 4507 139782 4559 139834
rect 7648 139782 7700 139834
rect 7712 139782 7764 139834
rect 7776 139782 7828 139834
rect 7840 139782 7892 139834
rect 2648 139238 2700 139290
rect 2712 139238 2764 139290
rect 2776 139238 2828 139290
rect 2840 139238 2892 139290
rect 5982 139238 6034 139290
rect 6046 139238 6098 139290
rect 6110 139238 6162 139290
rect 6174 139238 6226 139290
rect 4315 138694 4367 138746
rect 4379 138694 4431 138746
rect 4443 138694 4495 138746
rect 4507 138694 4559 138746
rect 7648 138694 7700 138746
rect 7712 138694 7764 138746
rect 7776 138694 7828 138746
rect 7840 138694 7892 138746
rect 2648 138150 2700 138202
rect 2712 138150 2764 138202
rect 2776 138150 2828 138202
rect 2840 138150 2892 138202
rect 5982 138150 6034 138202
rect 6046 138150 6098 138202
rect 6110 138150 6162 138202
rect 6174 138150 6226 138202
rect 4315 137606 4367 137658
rect 4379 137606 4431 137658
rect 4443 137606 4495 137658
rect 4507 137606 4559 137658
rect 7648 137606 7700 137658
rect 7712 137606 7764 137658
rect 7776 137606 7828 137658
rect 7840 137606 7892 137658
rect 2648 137062 2700 137114
rect 2712 137062 2764 137114
rect 2776 137062 2828 137114
rect 2840 137062 2892 137114
rect 5982 137062 6034 137114
rect 6046 137062 6098 137114
rect 6110 137062 6162 137114
rect 6174 137062 6226 137114
rect 4315 136518 4367 136570
rect 4379 136518 4431 136570
rect 4443 136518 4495 136570
rect 4507 136518 4559 136570
rect 7648 136518 7700 136570
rect 7712 136518 7764 136570
rect 7776 136518 7828 136570
rect 7840 136518 7892 136570
rect 2648 135974 2700 136026
rect 2712 135974 2764 136026
rect 2776 135974 2828 136026
rect 2840 135974 2892 136026
rect 5982 135974 6034 136026
rect 6046 135974 6098 136026
rect 6110 135974 6162 136026
rect 6174 135974 6226 136026
rect 4315 135430 4367 135482
rect 4379 135430 4431 135482
rect 4443 135430 4495 135482
rect 4507 135430 4559 135482
rect 7648 135430 7700 135482
rect 7712 135430 7764 135482
rect 7776 135430 7828 135482
rect 7840 135430 7892 135482
rect 2648 134886 2700 134938
rect 2712 134886 2764 134938
rect 2776 134886 2828 134938
rect 2840 134886 2892 134938
rect 5982 134886 6034 134938
rect 6046 134886 6098 134938
rect 6110 134886 6162 134938
rect 6174 134886 6226 134938
rect 4315 134342 4367 134394
rect 4379 134342 4431 134394
rect 4443 134342 4495 134394
rect 4507 134342 4559 134394
rect 7648 134342 7700 134394
rect 7712 134342 7764 134394
rect 7776 134342 7828 134394
rect 7840 134342 7892 134394
rect 2648 133798 2700 133850
rect 2712 133798 2764 133850
rect 2776 133798 2828 133850
rect 2840 133798 2892 133850
rect 5982 133798 6034 133850
rect 6046 133798 6098 133850
rect 6110 133798 6162 133850
rect 6174 133798 6226 133850
rect 4315 133254 4367 133306
rect 4379 133254 4431 133306
rect 4443 133254 4495 133306
rect 4507 133254 4559 133306
rect 7648 133254 7700 133306
rect 7712 133254 7764 133306
rect 7776 133254 7828 133306
rect 7840 133254 7892 133306
rect 2648 132710 2700 132762
rect 2712 132710 2764 132762
rect 2776 132710 2828 132762
rect 2840 132710 2892 132762
rect 5982 132710 6034 132762
rect 6046 132710 6098 132762
rect 6110 132710 6162 132762
rect 6174 132710 6226 132762
rect 4315 132166 4367 132218
rect 4379 132166 4431 132218
rect 4443 132166 4495 132218
rect 4507 132166 4559 132218
rect 7648 132166 7700 132218
rect 7712 132166 7764 132218
rect 7776 132166 7828 132218
rect 7840 132166 7892 132218
rect 2648 131622 2700 131674
rect 2712 131622 2764 131674
rect 2776 131622 2828 131674
rect 2840 131622 2892 131674
rect 5982 131622 6034 131674
rect 6046 131622 6098 131674
rect 6110 131622 6162 131674
rect 6174 131622 6226 131674
rect 4315 131078 4367 131130
rect 4379 131078 4431 131130
rect 4443 131078 4495 131130
rect 4507 131078 4559 131130
rect 7648 131078 7700 131130
rect 7712 131078 7764 131130
rect 7776 131078 7828 131130
rect 7840 131078 7892 131130
rect 2648 130534 2700 130586
rect 2712 130534 2764 130586
rect 2776 130534 2828 130586
rect 2840 130534 2892 130586
rect 5982 130534 6034 130586
rect 6046 130534 6098 130586
rect 6110 130534 6162 130586
rect 6174 130534 6226 130586
rect 4315 129990 4367 130042
rect 4379 129990 4431 130042
rect 4443 129990 4495 130042
rect 4507 129990 4559 130042
rect 7648 129990 7700 130042
rect 7712 129990 7764 130042
rect 7776 129990 7828 130042
rect 7840 129990 7892 130042
rect 2648 129446 2700 129498
rect 2712 129446 2764 129498
rect 2776 129446 2828 129498
rect 2840 129446 2892 129498
rect 5982 129446 6034 129498
rect 6046 129446 6098 129498
rect 6110 129446 6162 129498
rect 6174 129446 6226 129498
rect 4315 128902 4367 128954
rect 4379 128902 4431 128954
rect 4443 128902 4495 128954
rect 4507 128902 4559 128954
rect 7648 128902 7700 128954
rect 7712 128902 7764 128954
rect 7776 128902 7828 128954
rect 7840 128902 7892 128954
rect 2648 128358 2700 128410
rect 2712 128358 2764 128410
rect 2776 128358 2828 128410
rect 2840 128358 2892 128410
rect 5982 128358 6034 128410
rect 6046 128358 6098 128410
rect 6110 128358 6162 128410
rect 6174 128358 6226 128410
rect 4315 127814 4367 127866
rect 4379 127814 4431 127866
rect 4443 127814 4495 127866
rect 4507 127814 4559 127866
rect 7648 127814 7700 127866
rect 7712 127814 7764 127866
rect 7776 127814 7828 127866
rect 7840 127814 7892 127866
rect 2648 127270 2700 127322
rect 2712 127270 2764 127322
rect 2776 127270 2828 127322
rect 2840 127270 2892 127322
rect 5982 127270 6034 127322
rect 6046 127270 6098 127322
rect 6110 127270 6162 127322
rect 6174 127270 6226 127322
rect 4315 126726 4367 126778
rect 4379 126726 4431 126778
rect 4443 126726 4495 126778
rect 4507 126726 4559 126778
rect 7648 126726 7700 126778
rect 7712 126726 7764 126778
rect 7776 126726 7828 126778
rect 7840 126726 7892 126778
rect 2648 126182 2700 126234
rect 2712 126182 2764 126234
rect 2776 126182 2828 126234
rect 2840 126182 2892 126234
rect 5982 126182 6034 126234
rect 6046 126182 6098 126234
rect 6110 126182 6162 126234
rect 6174 126182 6226 126234
rect 4315 125638 4367 125690
rect 4379 125638 4431 125690
rect 4443 125638 4495 125690
rect 4507 125638 4559 125690
rect 7648 125638 7700 125690
rect 7712 125638 7764 125690
rect 7776 125638 7828 125690
rect 7840 125638 7892 125690
rect 2648 125094 2700 125146
rect 2712 125094 2764 125146
rect 2776 125094 2828 125146
rect 2840 125094 2892 125146
rect 5982 125094 6034 125146
rect 6046 125094 6098 125146
rect 6110 125094 6162 125146
rect 6174 125094 6226 125146
rect 4315 124550 4367 124602
rect 4379 124550 4431 124602
rect 4443 124550 4495 124602
rect 4507 124550 4559 124602
rect 7648 124550 7700 124602
rect 7712 124550 7764 124602
rect 7776 124550 7828 124602
rect 7840 124550 7892 124602
rect 2648 124006 2700 124058
rect 2712 124006 2764 124058
rect 2776 124006 2828 124058
rect 2840 124006 2892 124058
rect 5982 124006 6034 124058
rect 6046 124006 6098 124058
rect 6110 124006 6162 124058
rect 6174 124006 6226 124058
rect 4315 123462 4367 123514
rect 4379 123462 4431 123514
rect 4443 123462 4495 123514
rect 4507 123462 4559 123514
rect 7648 123462 7700 123514
rect 7712 123462 7764 123514
rect 7776 123462 7828 123514
rect 7840 123462 7892 123514
rect 2648 122918 2700 122970
rect 2712 122918 2764 122970
rect 2776 122918 2828 122970
rect 2840 122918 2892 122970
rect 5982 122918 6034 122970
rect 6046 122918 6098 122970
rect 6110 122918 6162 122970
rect 6174 122918 6226 122970
rect 4315 122374 4367 122426
rect 4379 122374 4431 122426
rect 4443 122374 4495 122426
rect 4507 122374 4559 122426
rect 7648 122374 7700 122426
rect 7712 122374 7764 122426
rect 7776 122374 7828 122426
rect 7840 122374 7892 122426
rect 2648 121830 2700 121882
rect 2712 121830 2764 121882
rect 2776 121830 2828 121882
rect 2840 121830 2892 121882
rect 5982 121830 6034 121882
rect 6046 121830 6098 121882
rect 6110 121830 6162 121882
rect 6174 121830 6226 121882
rect 4315 121286 4367 121338
rect 4379 121286 4431 121338
rect 4443 121286 4495 121338
rect 4507 121286 4559 121338
rect 7648 121286 7700 121338
rect 7712 121286 7764 121338
rect 7776 121286 7828 121338
rect 7840 121286 7892 121338
rect 2648 120742 2700 120794
rect 2712 120742 2764 120794
rect 2776 120742 2828 120794
rect 2840 120742 2892 120794
rect 5982 120742 6034 120794
rect 6046 120742 6098 120794
rect 6110 120742 6162 120794
rect 6174 120742 6226 120794
rect 4315 120198 4367 120250
rect 4379 120198 4431 120250
rect 4443 120198 4495 120250
rect 4507 120198 4559 120250
rect 7648 120198 7700 120250
rect 7712 120198 7764 120250
rect 7776 120198 7828 120250
rect 7840 120198 7892 120250
rect 2648 119654 2700 119706
rect 2712 119654 2764 119706
rect 2776 119654 2828 119706
rect 2840 119654 2892 119706
rect 5982 119654 6034 119706
rect 6046 119654 6098 119706
rect 6110 119654 6162 119706
rect 6174 119654 6226 119706
rect 4315 119110 4367 119162
rect 4379 119110 4431 119162
rect 4443 119110 4495 119162
rect 4507 119110 4559 119162
rect 7648 119110 7700 119162
rect 7712 119110 7764 119162
rect 7776 119110 7828 119162
rect 7840 119110 7892 119162
rect 2648 118566 2700 118618
rect 2712 118566 2764 118618
rect 2776 118566 2828 118618
rect 2840 118566 2892 118618
rect 5982 118566 6034 118618
rect 6046 118566 6098 118618
rect 6110 118566 6162 118618
rect 6174 118566 6226 118618
rect 4315 118022 4367 118074
rect 4379 118022 4431 118074
rect 4443 118022 4495 118074
rect 4507 118022 4559 118074
rect 7648 118022 7700 118074
rect 7712 118022 7764 118074
rect 7776 118022 7828 118074
rect 7840 118022 7892 118074
rect 2648 117478 2700 117530
rect 2712 117478 2764 117530
rect 2776 117478 2828 117530
rect 2840 117478 2892 117530
rect 5982 117478 6034 117530
rect 6046 117478 6098 117530
rect 6110 117478 6162 117530
rect 6174 117478 6226 117530
rect 4315 116934 4367 116986
rect 4379 116934 4431 116986
rect 4443 116934 4495 116986
rect 4507 116934 4559 116986
rect 7648 116934 7700 116986
rect 7712 116934 7764 116986
rect 7776 116934 7828 116986
rect 7840 116934 7892 116986
rect 2648 116390 2700 116442
rect 2712 116390 2764 116442
rect 2776 116390 2828 116442
rect 2840 116390 2892 116442
rect 5982 116390 6034 116442
rect 6046 116390 6098 116442
rect 6110 116390 6162 116442
rect 6174 116390 6226 116442
rect 4315 115846 4367 115898
rect 4379 115846 4431 115898
rect 4443 115846 4495 115898
rect 4507 115846 4559 115898
rect 7648 115846 7700 115898
rect 7712 115846 7764 115898
rect 7776 115846 7828 115898
rect 7840 115846 7892 115898
rect 2648 115302 2700 115354
rect 2712 115302 2764 115354
rect 2776 115302 2828 115354
rect 2840 115302 2892 115354
rect 5982 115302 6034 115354
rect 6046 115302 6098 115354
rect 6110 115302 6162 115354
rect 6174 115302 6226 115354
rect 4315 114758 4367 114810
rect 4379 114758 4431 114810
rect 4443 114758 4495 114810
rect 4507 114758 4559 114810
rect 7648 114758 7700 114810
rect 7712 114758 7764 114810
rect 7776 114758 7828 114810
rect 7840 114758 7892 114810
rect 2648 114214 2700 114266
rect 2712 114214 2764 114266
rect 2776 114214 2828 114266
rect 2840 114214 2892 114266
rect 5982 114214 6034 114266
rect 6046 114214 6098 114266
rect 6110 114214 6162 114266
rect 6174 114214 6226 114266
rect 4315 113670 4367 113722
rect 4379 113670 4431 113722
rect 4443 113670 4495 113722
rect 4507 113670 4559 113722
rect 7648 113670 7700 113722
rect 7712 113670 7764 113722
rect 7776 113670 7828 113722
rect 7840 113670 7892 113722
rect 2648 113126 2700 113178
rect 2712 113126 2764 113178
rect 2776 113126 2828 113178
rect 2840 113126 2892 113178
rect 5982 113126 6034 113178
rect 6046 113126 6098 113178
rect 6110 113126 6162 113178
rect 6174 113126 6226 113178
rect 4315 112582 4367 112634
rect 4379 112582 4431 112634
rect 4443 112582 4495 112634
rect 4507 112582 4559 112634
rect 7648 112582 7700 112634
rect 7712 112582 7764 112634
rect 7776 112582 7828 112634
rect 7840 112582 7892 112634
rect 2648 112038 2700 112090
rect 2712 112038 2764 112090
rect 2776 112038 2828 112090
rect 2840 112038 2892 112090
rect 5982 112038 6034 112090
rect 6046 112038 6098 112090
rect 6110 112038 6162 112090
rect 6174 112038 6226 112090
rect 4315 111494 4367 111546
rect 4379 111494 4431 111546
rect 4443 111494 4495 111546
rect 4507 111494 4559 111546
rect 7648 111494 7700 111546
rect 7712 111494 7764 111546
rect 7776 111494 7828 111546
rect 7840 111494 7892 111546
rect 2648 110950 2700 111002
rect 2712 110950 2764 111002
rect 2776 110950 2828 111002
rect 2840 110950 2892 111002
rect 5982 110950 6034 111002
rect 6046 110950 6098 111002
rect 6110 110950 6162 111002
rect 6174 110950 6226 111002
rect 4315 110406 4367 110458
rect 4379 110406 4431 110458
rect 4443 110406 4495 110458
rect 4507 110406 4559 110458
rect 7648 110406 7700 110458
rect 7712 110406 7764 110458
rect 7776 110406 7828 110458
rect 7840 110406 7892 110458
rect 2648 109862 2700 109914
rect 2712 109862 2764 109914
rect 2776 109862 2828 109914
rect 2840 109862 2892 109914
rect 5982 109862 6034 109914
rect 6046 109862 6098 109914
rect 6110 109862 6162 109914
rect 6174 109862 6226 109914
rect 4315 109318 4367 109370
rect 4379 109318 4431 109370
rect 4443 109318 4495 109370
rect 4507 109318 4559 109370
rect 7648 109318 7700 109370
rect 7712 109318 7764 109370
rect 7776 109318 7828 109370
rect 7840 109318 7892 109370
rect 2648 108774 2700 108826
rect 2712 108774 2764 108826
rect 2776 108774 2828 108826
rect 2840 108774 2892 108826
rect 5982 108774 6034 108826
rect 6046 108774 6098 108826
rect 6110 108774 6162 108826
rect 6174 108774 6226 108826
rect 4315 108230 4367 108282
rect 4379 108230 4431 108282
rect 4443 108230 4495 108282
rect 4507 108230 4559 108282
rect 7648 108230 7700 108282
rect 7712 108230 7764 108282
rect 7776 108230 7828 108282
rect 7840 108230 7892 108282
rect 2648 107686 2700 107738
rect 2712 107686 2764 107738
rect 2776 107686 2828 107738
rect 2840 107686 2892 107738
rect 5982 107686 6034 107738
rect 6046 107686 6098 107738
rect 6110 107686 6162 107738
rect 6174 107686 6226 107738
rect 4315 107142 4367 107194
rect 4379 107142 4431 107194
rect 4443 107142 4495 107194
rect 4507 107142 4559 107194
rect 7648 107142 7700 107194
rect 7712 107142 7764 107194
rect 7776 107142 7828 107194
rect 7840 107142 7892 107194
rect 2648 106598 2700 106650
rect 2712 106598 2764 106650
rect 2776 106598 2828 106650
rect 2840 106598 2892 106650
rect 5982 106598 6034 106650
rect 6046 106598 6098 106650
rect 6110 106598 6162 106650
rect 6174 106598 6226 106650
rect 4315 106054 4367 106106
rect 4379 106054 4431 106106
rect 4443 106054 4495 106106
rect 4507 106054 4559 106106
rect 7648 106054 7700 106106
rect 7712 106054 7764 106106
rect 7776 106054 7828 106106
rect 7840 106054 7892 106106
rect 2648 105510 2700 105562
rect 2712 105510 2764 105562
rect 2776 105510 2828 105562
rect 2840 105510 2892 105562
rect 5982 105510 6034 105562
rect 6046 105510 6098 105562
rect 6110 105510 6162 105562
rect 6174 105510 6226 105562
rect 4315 104966 4367 105018
rect 4379 104966 4431 105018
rect 4443 104966 4495 105018
rect 4507 104966 4559 105018
rect 7648 104966 7700 105018
rect 7712 104966 7764 105018
rect 7776 104966 7828 105018
rect 7840 104966 7892 105018
rect 2648 104422 2700 104474
rect 2712 104422 2764 104474
rect 2776 104422 2828 104474
rect 2840 104422 2892 104474
rect 5982 104422 6034 104474
rect 6046 104422 6098 104474
rect 6110 104422 6162 104474
rect 6174 104422 6226 104474
rect 4315 103878 4367 103930
rect 4379 103878 4431 103930
rect 4443 103878 4495 103930
rect 4507 103878 4559 103930
rect 7648 103878 7700 103930
rect 7712 103878 7764 103930
rect 7776 103878 7828 103930
rect 7840 103878 7892 103930
rect 2648 103334 2700 103386
rect 2712 103334 2764 103386
rect 2776 103334 2828 103386
rect 2840 103334 2892 103386
rect 5982 103334 6034 103386
rect 6046 103334 6098 103386
rect 6110 103334 6162 103386
rect 6174 103334 6226 103386
rect 4315 102790 4367 102842
rect 4379 102790 4431 102842
rect 4443 102790 4495 102842
rect 4507 102790 4559 102842
rect 7648 102790 7700 102842
rect 7712 102790 7764 102842
rect 7776 102790 7828 102842
rect 7840 102790 7892 102842
rect 2648 102246 2700 102298
rect 2712 102246 2764 102298
rect 2776 102246 2828 102298
rect 2840 102246 2892 102298
rect 5982 102246 6034 102298
rect 6046 102246 6098 102298
rect 6110 102246 6162 102298
rect 6174 102246 6226 102298
rect 4315 101702 4367 101754
rect 4379 101702 4431 101754
rect 4443 101702 4495 101754
rect 4507 101702 4559 101754
rect 7648 101702 7700 101754
rect 7712 101702 7764 101754
rect 7776 101702 7828 101754
rect 7840 101702 7892 101754
rect 2648 101158 2700 101210
rect 2712 101158 2764 101210
rect 2776 101158 2828 101210
rect 2840 101158 2892 101210
rect 5982 101158 6034 101210
rect 6046 101158 6098 101210
rect 6110 101158 6162 101210
rect 6174 101158 6226 101210
rect 4315 100614 4367 100666
rect 4379 100614 4431 100666
rect 4443 100614 4495 100666
rect 4507 100614 4559 100666
rect 7648 100614 7700 100666
rect 7712 100614 7764 100666
rect 7776 100614 7828 100666
rect 7840 100614 7892 100666
rect 2648 100070 2700 100122
rect 2712 100070 2764 100122
rect 2776 100070 2828 100122
rect 2840 100070 2892 100122
rect 5982 100070 6034 100122
rect 6046 100070 6098 100122
rect 6110 100070 6162 100122
rect 6174 100070 6226 100122
rect 4315 99526 4367 99578
rect 4379 99526 4431 99578
rect 4443 99526 4495 99578
rect 4507 99526 4559 99578
rect 7648 99526 7700 99578
rect 7712 99526 7764 99578
rect 7776 99526 7828 99578
rect 7840 99526 7892 99578
rect 2648 98982 2700 99034
rect 2712 98982 2764 99034
rect 2776 98982 2828 99034
rect 2840 98982 2892 99034
rect 5982 98982 6034 99034
rect 6046 98982 6098 99034
rect 6110 98982 6162 99034
rect 6174 98982 6226 99034
rect 4315 98438 4367 98490
rect 4379 98438 4431 98490
rect 4443 98438 4495 98490
rect 4507 98438 4559 98490
rect 7648 98438 7700 98490
rect 7712 98438 7764 98490
rect 7776 98438 7828 98490
rect 7840 98438 7892 98490
rect 2648 97894 2700 97946
rect 2712 97894 2764 97946
rect 2776 97894 2828 97946
rect 2840 97894 2892 97946
rect 5982 97894 6034 97946
rect 6046 97894 6098 97946
rect 6110 97894 6162 97946
rect 6174 97894 6226 97946
rect 4315 97350 4367 97402
rect 4379 97350 4431 97402
rect 4443 97350 4495 97402
rect 4507 97350 4559 97402
rect 7648 97350 7700 97402
rect 7712 97350 7764 97402
rect 7776 97350 7828 97402
rect 7840 97350 7892 97402
rect 2648 96806 2700 96858
rect 2712 96806 2764 96858
rect 2776 96806 2828 96858
rect 2840 96806 2892 96858
rect 5982 96806 6034 96858
rect 6046 96806 6098 96858
rect 6110 96806 6162 96858
rect 6174 96806 6226 96858
rect 4315 96262 4367 96314
rect 4379 96262 4431 96314
rect 4443 96262 4495 96314
rect 4507 96262 4559 96314
rect 7648 96262 7700 96314
rect 7712 96262 7764 96314
rect 7776 96262 7828 96314
rect 7840 96262 7892 96314
rect 2648 95718 2700 95770
rect 2712 95718 2764 95770
rect 2776 95718 2828 95770
rect 2840 95718 2892 95770
rect 5982 95718 6034 95770
rect 6046 95718 6098 95770
rect 6110 95718 6162 95770
rect 6174 95718 6226 95770
rect 4315 95174 4367 95226
rect 4379 95174 4431 95226
rect 4443 95174 4495 95226
rect 4507 95174 4559 95226
rect 7648 95174 7700 95226
rect 7712 95174 7764 95226
rect 7776 95174 7828 95226
rect 7840 95174 7892 95226
rect 2648 94630 2700 94682
rect 2712 94630 2764 94682
rect 2776 94630 2828 94682
rect 2840 94630 2892 94682
rect 5982 94630 6034 94682
rect 6046 94630 6098 94682
rect 6110 94630 6162 94682
rect 6174 94630 6226 94682
rect 4315 94086 4367 94138
rect 4379 94086 4431 94138
rect 4443 94086 4495 94138
rect 4507 94086 4559 94138
rect 7648 94086 7700 94138
rect 7712 94086 7764 94138
rect 7776 94086 7828 94138
rect 7840 94086 7892 94138
rect 2648 93542 2700 93594
rect 2712 93542 2764 93594
rect 2776 93542 2828 93594
rect 2840 93542 2892 93594
rect 5982 93542 6034 93594
rect 6046 93542 6098 93594
rect 6110 93542 6162 93594
rect 6174 93542 6226 93594
rect 4315 92998 4367 93050
rect 4379 92998 4431 93050
rect 4443 92998 4495 93050
rect 4507 92998 4559 93050
rect 7648 92998 7700 93050
rect 7712 92998 7764 93050
rect 7776 92998 7828 93050
rect 7840 92998 7892 93050
rect 2648 92454 2700 92506
rect 2712 92454 2764 92506
rect 2776 92454 2828 92506
rect 2840 92454 2892 92506
rect 5982 92454 6034 92506
rect 6046 92454 6098 92506
rect 6110 92454 6162 92506
rect 6174 92454 6226 92506
rect 4315 91910 4367 91962
rect 4379 91910 4431 91962
rect 4443 91910 4495 91962
rect 4507 91910 4559 91962
rect 7648 91910 7700 91962
rect 7712 91910 7764 91962
rect 7776 91910 7828 91962
rect 7840 91910 7892 91962
rect 2648 91366 2700 91418
rect 2712 91366 2764 91418
rect 2776 91366 2828 91418
rect 2840 91366 2892 91418
rect 5982 91366 6034 91418
rect 6046 91366 6098 91418
rect 6110 91366 6162 91418
rect 6174 91366 6226 91418
rect 4315 90822 4367 90874
rect 4379 90822 4431 90874
rect 4443 90822 4495 90874
rect 4507 90822 4559 90874
rect 7648 90822 7700 90874
rect 7712 90822 7764 90874
rect 7776 90822 7828 90874
rect 7840 90822 7892 90874
rect 2648 90278 2700 90330
rect 2712 90278 2764 90330
rect 2776 90278 2828 90330
rect 2840 90278 2892 90330
rect 5982 90278 6034 90330
rect 6046 90278 6098 90330
rect 6110 90278 6162 90330
rect 6174 90278 6226 90330
rect 4315 89734 4367 89786
rect 4379 89734 4431 89786
rect 4443 89734 4495 89786
rect 4507 89734 4559 89786
rect 7648 89734 7700 89786
rect 7712 89734 7764 89786
rect 7776 89734 7828 89786
rect 7840 89734 7892 89786
rect 2648 89190 2700 89242
rect 2712 89190 2764 89242
rect 2776 89190 2828 89242
rect 2840 89190 2892 89242
rect 5982 89190 6034 89242
rect 6046 89190 6098 89242
rect 6110 89190 6162 89242
rect 6174 89190 6226 89242
rect 4315 88646 4367 88698
rect 4379 88646 4431 88698
rect 4443 88646 4495 88698
rect 4507 88646 4559 88698
rect 7648 88646 7700 88698
rect 7712 88646 7764 88698
rect 7776 88646 7828 88698
rect 7840 88646 7892 88698
rect 2648 88102 2700 88154
rect 2712 88102 2764 88154
rect 2776 88102 2828 88154
rect 2840 88102 2892 88154
rect 5982 88102 6034 88154
rect 6046 88102 6098 88154
rect 6110 88102 6162 88154
rect 6174 88102 6226 88154
rect 4315 87558 4367 87610
rect 4379 87558 4431 87610
rect 4443 87558 4495 87610
rect 4507 87558 4559 87610
rect 7648 87558 7700 87610
rect 7712 87558 7764 87610
rect 7776 87558 7828 87610
rect 7840 87558 7892 87610
rect 2648 87014 2700 87066
rect 2712 87014 2764 87066
rect 2776 87014 2828 87066
rect 2840 87014 2892 87066
rect 5982 87014 6034 87066
rect 6046 87014 6098 87066
rect 6110 87014 6162 87066
rect 6174 87014 6226 87066
rect 4315 86470 4367 86522
rect 4379 86470 4431 86522
rect 4443 86470 4495 86522
rect 4507 86470 4559 86522
rect 7648 86470 7700 86522
rect 7712 86470 7764 86522
rect 7776 86470 7828 86522
rect 7840 86470 7892 86522
rect 2648 85926 2700 85978
rect 2712 85926 2764 85978
rect 2776 85926 2828 85978
rect 2840 85926 2892 85978
rect 5982 85926 6034 85978
rect 6046 85926 6098 85978
rect 6110 85926 6162 85978
rect 6174 85926 6226 85978
rect 4315 85382 4367 85434
rect 4379 85382 4431 85434
rect 4443 85382 4495 85434
rect 4507 85382 4559 85434
rect 7648 85382 7700 85434
rect 7712 85382 7764 85434
rect 7776 85382 7828 85434
rect 7840 85382 7892 85434
rect 2648 84838 2700 84890
rect 2712 84838 2764 84890
rect 2776 84838 2828 84890
rect 2840 84838 2892 84890
rect 5982 84838 6034 84890
rect 6046 84838 6098 84890
rect 6110 84838 6162 84890
rect 6174 84838 6226 84890
rect 4315 84294 4367 84346
rect 4379 84294 4431 84346
rect 4443 84294 4495 84346
rect 4507 84294 4559 84346
rect 7648 84294 7700 84346
rect 7712 84294 7764 84346
rect 7776 84294 7828 84346
rect 7840 84294 7892 84346
rect 2648 83750 2700 83802
rect 2712 83750 2764 83802
rect 2776 83750 2828 83802
rect 2840 83750 2892 83802
rect 5982 83750 6034 83802
rect 6046 83750 6098 83802
rect 6110 83750 6162 83802
rect 6174 83750 6226 83802
rect 4315 83206 4367 83258
rect 4379 83206 4431 83258
rect 4443 83206 4495 83258
rect 4507 83206 4559 83258
rect 7648 83206 7700 83258
rect 7712 83206 7764 83258
rect 7776 83206 7828 83258
rect 7840 83206 7892 83258
rect 2648 82662 2700 82714
rect 2712 82662 2764 82714
rect 2776 82662 2828 82714
rect 2840 82662 2892 82714
rect 5982 82662 6034 82714
rect 6046 82662 6098 82714
rect 6110 82662 6162 82714
rect 6174 82662 6226 82714
rect 4315 82118 4367 82170
rect 4379 82118 4431 82170
rect 4443 82118 4495 82170
rect 4507 82118 4559 82170
rect 7648 82118 7700 82170
rect 7712 82118 7764 82170
rect 7776 82118 7828 82170
rect 7840 82118 7892 82170
rect 2648 81574 2700 81626
rect 2712 81574 2764 81626
rect 2776 81574 2828 81626
rect 2840 81574 2892 81626
rect 5982 81574 6034 81626
rect 6046 81574 6098 81626
rect 6110 81574 6162 81626
rect 6174 81574 6226 81626
rect 4315 81030 4367 81082
rect 4379 81030 4431 81082
rect 4443 81030 4495 81082
rect 4507 81030 4559 81082
rect 7648 81030 7700 81082
rect 7712 81030 7764 81082
rect 7776 81030 7828 81082
rect 7840 81030 7892 81082
rect 2648 80486 2700 80538
rect 2712 80486 2764 80538
rect 2776 80486 2828 80538
rect 2840 80486 2892 80538
rect 5982 80486 6034 80538
rect 6046 80486 6098 80538
rect 6110 80486 6162 80538
rect 6174 80486 6226 80538
rect 4315 79942 4367 79994
rect 4379 79942 4431 79994
rect 4443 79942 4495 79994
rect 4507 79942 4559 79994
rect 7648 79942 7700 79994
rect 7712 79942 7764 79994
rect 7776 79942 7828 79994
rect 7840 79942 7892 79994
rect 2648 79398 2700 79450
rect 2712 79398 2764 79450
rect 2776 79398 2828 79450
rect 2840 79398 2892 79450
rect 5982 79398 6034 79450
rect 6046 79398 6098 79450
rect 6110 79398 6162 79450
rect 6174 79398 6226 79450
rect 4315 78854 4367 78906
rect 4379 78854 4431 78906
rect 4443 78854 4495 78906
rect 4507 78854 4559 78906
rect 7648 78854 7700 78906
rect 7712 78854 7764 78906
rect 7776 78854 7828 78906
rect 7840 78854 7892 78906
rect 2648 78310 2700 78362
rect 2712 78310 2764 78362
rect 2776 78310 2828 78362
rect 2840 78310 2892 78362
rect 5982 78310 6034 78362
rect 6046 78310 6098 78362
rect 6110 78310 6162 78362
rect 6174 78310 6226 78362
rect 4315 77766 4367 77818
rect 4379 77766 4431 77818
rect 4443 77766 4495 77818
rect 4507 77766 4559 77818
rect 7648 77766 7700 77818
rect 7712 77766 7764 77818
rect 7776 77766 7828 77818
rect 7840 77766 7892 77818
rect 2648 77222 2700 77274
rect 2712 77222 2764 77274
rect 2776 77222 2828 77274
rect 2840 77222 2892 77274
rect 5982 77222 6034 77274
rect 6046 77222 6098 77274
rect 6110 77222 6162 77274
rect 6174 77222 6226 77274
rect 4315 76678 4367 76730
rect 4379 76678 4431 76730
rect 4443 76678 4495 76730
rect 4507 76678 4559 76730
rect 7648 76678 7700 76730
rect 7712 76678 7764 76730
rect 7776 76678 7828 76730
rect 7840 76678 7892 76730
rect 2648 76134 2700 76186
rect 2712 76134 2764 76186
rect 2776 76134 2828 76186
rect 2840 76134 2892 76186
rect 5982 76134 6034 76186
rect 6046 76134 6098 76186
rect 6110 76134 6162 76186
rect 6174 76134 6226 76186
rect 4315 75590 4367 75642
rect 4379 75590 4431 75642
rect 4443 75590 4495 75642
rect 4507 75590 4559 75642
rect 7648 75590 7700 75642
rect 7712 75590 7764 75642
rect 7776 75590 7828 75642
rect 7840 75590 7892 75642
rect 2648 75046 2700 75098
rect 2712 75046 2764 75098
rect 2776 75046 2828 75098
rect 2840 75046 2892 75098
rect 5982 75046 6034 75098
rect 6046 75046 6098 75098
rect 6110 75046 6162 75098
rect 6174 75046 6226 75098
rect 4315 74502 4367 74554
rect 4379 74502 4431 74554
rect 4443 74502 4495 74554
rect 4507 74502 4559 74554
rect 7648 74502 7700 74554
rect 7712 74502 7764 74554
rect 7776 74502 7828 74554
rect 7840 74502 7892 74554
rect 2648 73958 2700 74010
rect 2712 73958 2764 74010
rect 2776 73958 2828 74010
rect 2840 73958 2892 74010
rect 5982 73958 6034 74010
rect 6046 73958 6098 74010
rect 6110 73958 6162 74010
rect 6174 73958 6226 74010
rect 4315 73414 4367 73466
rect 4379 73414 4431 73466
rect 4443 73414 4495 73466
rect 4507 73414 4559 73466
rect 7648 73414 7700 73466
rect 7712 73414 7764 73466
rect 7776 73414 7828 73466
rect 7840 73414 7892 73466
rect 2648 72870 2700 72922
rect 2712 72870 2764 72922
rect 2776 72870 2828 72922
rect 2840 72870 2892 72922
rect 5982 72870 6034 72922
rect 6046 72870 6098 72922
rect 6110 72870 6162 72922
rect 6174 72870 6226 72922
rect 4315 72326 4367 72378
rect 4379 72326 4431 72378
rect 4443 72326 4495 72378
rect 4507 72326 4559 72378
rect 7648 72326 7700 72378
rect 7712 72326 7764 72378
rect 7776 72326 7828 72378
rect 7840 72326 7892 72378
rect 112 72020 164 72072
rect 5632 72020 5684 72072
rect 5632 71884 5684 71936
rect 6736 71884 6788 71936
rect 2648 71782 2700 71834
rect 2712 71782 2764 71834
rect 2776 71782 2828 71834
rect 2840 71782 2892 71834
rect 5982 71782 6034 71834
rect 6046 71782 6098 71834
rect 6110 71782 6162 71834
rect 6174 71782 6226 71834
rect 4315 71238 4367 71290
rect 4379 71238 4431 71290
rect 4443 71238 4495 71290
rect 4507 71238 4559 71290
rect 7648 71238 7700 71290
rect 7712 71238 7764 71290
rect 7776 71238 7828 71290
rect 7840 71238 7892 71290
rect 2648 70694 2700 70746
rect 2712 70694 2764 70746
rect 2776 70694 2828 70746
rect 2840 70694 2892 70746
rect 5982 70694 6034 70746
rect 6046 70694 6098 70746
rect 6110 70694 6162 70746
rect 6174 70694 6226 70746
rect 4315 70150 4367 70202
rect 4379 70150 4431 70202
rect 4443 70150 4495 70202
rect 4507 70150 4559 70202
rect 7648 70150 7700 70202
rect 7712 70150 7764 70202
rect 7776 70150 7828 70202
rect 7840 70150 7892 70202
rect 2648 69606 2700 69658
rect 2712 69606 2764 69658
rect 2776 69606 2828 69658
rect 2840 69606 2892 69658
rect 5982 69606 6034 69658
rect 6046 69606 6098 69658
rect 6110 69606 6162 69658
rect 6174 69606 6226 69658
rect 4315 69062 4367 69114
rect 4379 69062 4431 69114
rect 4443 69062 4495 69114
rect 4507 69062 4559 69114
rect 7648 69062 7700 69114
rect 7712 69062 7764 69114
rect 7776 69062 7828 69114
rect 7840 69062 7892 69114
rect 2648 68518 2700 68570
rect 2712 68518 2764 68570
rect 2776 68518 2828 68570
rect 2840 68518 2892 68570
rect 5982 68518 6034 68570
rect 6046 68518 6098 68570
rect 6110 68518 6162 68570
rect 6174 68518 6226 68570
rect 4315 67974 4367 68026
rect 4379 67974 4431 68026
rect 4443 67974 4495 68026
rect 4507 67974 4559 68026
rect 7648 67974 7700 68026
rect 7712 67974 7764 68026
rect 7776 67974 7828 68026
rect 7840 67974 7892 68026
rect 2648 67430 2700 67482
rect 2712 67430 2764 67482
rect 2776 67430 2828 67482
rect 2840 67430 2892 67482
rect 5982 67430 6034 67482
rect 6046 67430 6098 67482
rect 6110 67430 6162 67482
rect 6174 67430 6226 67482
rect 4315 66886 4367 66938
rect 4379 66886 4431 66938
rect 4443 66886 4495 66938
rect 4507 66886 4559 66938
rect 7648 66886 7700 66938
rect 7712 66886 7764 66938
rect 7776 66886 7828 66938
rect 7840 66886 7892 66938
rect 2648 66342 2700 66394
rect 2712 66342 2764 66394
rect 2776 66342 2828 66394
rect 2840 66342 2892 66394
rect 5982 66342 6034 66394
rect 6046 66342 6098 66394
rect 6110 66342 6162 66394
rect 6174 66342 6226 66394
rect 4315 65798 4367 65850
rect 4379 65798 4431 65850
rect 4443 65798 4495 65850
rect 4507 65798 4559 65850
rect 7648 65798 7700 65850
rect 7712 65798 7764 65850
rect 7776 65798 7828 65850
rect 7840 65798 7892 65850
rect 2648 65254 2700 65306
rect 2712 65254 2764 65306
rect 2776 65254 2828 65306
rect 2840 65254 2892 65306
rect 5982 65254 6034 65306
rect 6046 65254 6098 65306
rect 6110 65254 6162 65306
rect 6174 65254 6226 65306
rect 4315 64710 4367 64762
rect 4379 64710 4431 64762
rect 4443 64710 4495 64762
rect 4507 64710 4559 64762
rect 7648 64710 7700 64762
rect 7712 64710 7764 64762
rect 7776 64710 7828 64762
rect 7840 64710 7892 64762
rect 2648 64166 2700 64218
rect 2712 64166 2764 64218
rect 2776 64166 2828 64218
rect 2840 64166 2892 64218
rect 5982 64166 6034 64218
rect 6046 64166 6098 64218
rect 6110 64166 6162 64218
rect 6174 64166 6226 64218
rect 4315 63622 4367 63674
rect 4379 63622 4431 63674
rect 4443 63622 4495 63674
rect 4507 63622 4559 63674
rect 7648 63622 7700 63674
rect 7712 63622 7764 63674
rect 7776 63622 7828 63674
rect 7840 63622 7892 63674
rect 2648 63078 2700 63130
rect 2712 63078 2764 63130
rect 2776 63078 2828 63130
rect 2840 63078 2892 63130
rect 5982 63078 6034 63130
rect 6046 63078 6098 63130
rect 6110 63078 6162 63130
rect 6174 63078 6226 63130
rect 4315 62534 4367 62586
rect 4379 62534 4431 62586
rect 4443 62534 4495 62586
rect 4507 62534 4559 62586
rect 7648 62534 7700 62586
rect 7712 62534 7764 62586
rect 7776 62534 7828 62586
rect 7840 62534 7892 62586
rect 2648 61990 2700 62042
rect 2712 61990 2764 62042
rect 2776 61990 2828 62042
rect 2840 61990 2892 62042
rect 5982 61990 6034 62042
rect 6046 61990 6098 62042
rect 6110 61990 6162 62042
rect 6174 61990 6226 62042
rect 4315 61446 4367 61498
rect 4379 61446 4431 61498
rect 4443 61446 4495 61498
rect 4507 61446 4559 61498
rect 7648 61446 7700 61498
rect 7712 61446 7764 61498
rect 7776 61446 7828 61498
rect 7840 61446 7892 61498
rect 2648 60902 2700 60954
rect 2712 60902 2764 60954
rect 2776 60902 2828 60954
rect 2840 60902 2892 60954
rect 5982 60902 6034 60954
rect 6046 60902 6098 60954
rect 6110 60902 6162 60954
rect 6174 60902 6226 60954
rect 4315 60358 4367 60410
rect 4379 60358 4431 60410
rect 4443 60358 4495 60410
rect 4507 60358 4559 60410
rect 7648 60358 7700 60410
rect 7712 60358 7764 60410
rect 7776 60358 7828 60410
rect 7840 60358 7892 60410
rect 2648 59814 2700 59866
rect 2712 59814 2764 59866
rect 2776 59814 2828 59866
rect 2840 59814 2892 59866
rect 5982 59814 6034 59866
rect 6046 59814 6098 59866
rect 6110 59814 6162 59866
rect 6174 59814 6226 59866
rect 4315 59270 4367 59322
rect 4379 59270 4431 59322
rect 4443 59270 4495 59322
rect 4507 59270 4559 59322
rect 7648 59270 7700 59322
rect 7712 59270 7764 59322
rect 7776 59270 7828 59322
rect 7840 59270 7892 59322
rect 2648 58726 2700 58778
rect 2712 58726 2764 58778
rect 2776 58726 2828 58778
rect 2840 58726 2892 58778
rect 5982 58726 6034 58778
rect 6046 58726 6098 58778
rect 6110 58726 6162 58778
rect 6174 58726 6226 58778
rect 4315 58182 4367 58234
rect 4379 58182 4431 58234
rect 4443 58182 4495 58234
rect 4507 58182 4559 58234
rect 7648 58182 7700 58234
rect 7712 58182 7764 58234
rect 7776 58182 7828 58234
rect 7840 58182 7892 58234
rect 2648 57638 2700 57690
rect 2712 57638 2764 57690
rect 2776 57638 2828 57690
rect 2840 57638 2892 57690
rect 5982 57638 6034 57690
rect 6046 57638 6098 57690
rect 6110 57638 6162 57690
rect 6174 57638 6226 57690
rect 4315 57094 4367 57146
rect 4379 57094 4431 57146
rect 4443 57094 4495 57146
rect 4507 57094 4559 57146
rect 7648 57094 7700 57146
rect 7712 57094 7764 57146
rect 7776 57094 7828 57146
rect 7840 57094 7892 57146
rect 2648 56550 2700 56602
rect 2712 56550 2764 56602
rect 2776 56550 2828 56602
rect 2840 56550 2892 56602
rect 5982 56550 6034 56602
rect 6046 56550 6098 56602
rect 6110 56550 6162 56602
rect 6174 56550 6226 56602
rect 4315 56006 4367 56058
rect 4379 56006 4431 56058
rect 4443 56006 4495 56058
rect 4507 56006 4559 56058
rect 7648 56006 7700 56058
rect 7712 56006 7764 56058
rect 7776 56006 7828 56058
rect 7840 56006 7892 56058
rect 2648 55462 2700 55514
rect 2712 55462 2764 55514
rect 2776 55462 2828 55514
rect 2840 55462 2892 55514
rect 5982 55462 6034 55514
rect 6046 55462 6098 55514
rect 6110 55462 6162 55514
rect 6174 55462 6226 55514
rect 4315 54918 4367 54970
rect 4379 54918 4431 54970
rect 4443 54918 4495 54970
rect 4507 54918 4559 54970
rect 7648 54918 7700 54970
rect 7712 54918 7764 54970
rect 7776 54918 7828 54970
rect 7840 54918 7892 54970
rect 2648 54374 2700 54426
rect 2712 54374 2764 54426
rect 2776 54374 2828 54426
rect 2840 54374 2892 54426
rect 5982 54374 6034 54426
rect 6046 54374 6098 54426
rect 6110 54374 6162 54426
rect 6174 54374 6226 54426
rect 4315 53830 4367 53882
rect 4379 53830 4431 53882
rect 4443 53830 4495 53882
rect 4507 53830 4559 53882
rect 7648 53830 7700 53882
rect 7712 53830 7764 53882
rect 7776 53830 7828 53882
rect 7840 53830 7892 53882
rect 2648 53286 2700 53338
rect 2712 53286 2764 53338
rect 2776 53286 2828 53338
rect 2840 53286 2892 53338
rect 5982 53286 6034 53338
rect 6046 53286 6098 53338
rect 6110 53286 6162 53338
rect 6174 53286 6226 53338
rect 4315 52742 4367 52794
rect 4379 52742 4431 52794
rect 4443 52742 4495 52794
rect 4507 52742 4559 52794
rect 7648 52742 7700 52794
rect 7712 52742 7764 52794
rect 7776 52742 7828 52794
rect 7840 52742 7892 52794
rect 2648 52198 2700 52250
rect 2712 52198 2764 52250
rect 2776 52198 2828 52250
rect 2840 52198 2892 52250
rect 5982 52198 6034 52250
rect 6046 52198 6098 52250
rect 6110 52198 6162 52250
rect 6174 52198 6226 52250
rect 4315 51654 4367 51706
rect 4379 51654 4431 51706
rect 4443 51654 4495 51706
rect 4507 51654 4559 51706
rect 7648 51654 7700 51706
rect 7712 51654 7764 51706
rect 7776 51654 7828 51706
rect 7840 51654 7892 51706
rect 2648 51110 2700 51162
rect 2712 51110 2764 51162
rect 2776 51110 2828 51162
rect 2840 51110 2892 51162
rect 5982 51110 6034 51162
rect 6046 51110 6098 51162
rect 6110 51110 6162 51162
rect 6174 51110 6226 51162
rect 8208 50940 8260 50992
rect 6736 50804 6788 50856
rect 4315 50566 4367 50618
rect 4379 50566 4431 50618
rect 4443 50566 4495 50618
rect 4507 50566 4559 50618
rect 7648 50566 7700 50618
rect 7712 50566 7764 50618
rect 7776 50566 7828 50618
rect 7840 50566 7892 50618
rect 2648 50022 2700 50074
rect 2712 50022 2764 50074
rect 2776 50022 2828 50074
rect 2840 50022 2892 50074
rect 5982 50022 6034 50074
rect 6046 50022 6098 50074
rect 6110 50022 6162 50074
rect 6174 50022 6226 50074
rect 4315 49478 4367 49530
rect 4379 49478 4431 49530
rect 4443 49478 4495 49530
rect 4507 49478 4559 49530
rect 7648 49478 7700 49530
rect 7712 49478 7764 49530
rect 7776 49478 7828 49530
rect 7840 49478 7892 49530
rect 2648 48934 2700 48986
rect 2712 48934 2764 48986
rect 2776 48934 2828 48986
rect 2840 48934 2892 48986
rect 5982 48934 6034 48986
rect 6046 48934 6098 48986
rect 6110 48934 6162 48986
rect 6174 48934 6226 48986
rect 4315 48390 4367 48442
rect 4379 48390 4431 48442
rect 4443 48390 4495 48442
rect 4507 48390 4559 48442
rect 7648 48390 7700 48442
rect 7712 48390 7764 48442
rect 7776 48390 7828 48442
rect 7840 48390 7892 48442
rect 2648 47846 2700 47898
rect 2712 47846 2764 47898
rect 2776 47846 2828 47898
rect 2840 47846 2892 47898
rect 5982 47846 6034 47898
rect 6046 47846 6098 47898
rect 6110 47846 6162 47898
rect 6174 47846 6226 47898
rect 4315 47302 4367 47354
rect 4379 47302 4431 47354
rect 4443 47302 4495 47354
rect 4507 47302 4559 47354
rect 7648 47302 7700 47354
rect 7712 47302 7764 47354
rect 7776 47302 7828 47354
rect 7840 47302 7892 47354
rect 2648 46758 2700 46810
rect 2712 46758 2764 46810
rect 2776 46758 2828 46810
rect 2840 46758 2892 46810
rect 5982 46758 6034 46810
rect 6046 46758 6098 46810
rect 6110 46758 6162 46810
rect 6174 46758 6226 46810
rect 4315 46214 4367 46266
rect 4379 46214 4431 46266
rect 4443 46214 4495 46266
rect 4507 46214 4559 46266
rect 7648 46214 7700 46266
rect 7712 46214 7764 46266
rect 7776 46214 7828 46266
rect 7840 46214 7892 46266
rect 2648 45670 2700 45722
rect 2712 45670 2764 45722
rect 2776 45670 2828 45722
rect 2840 45670 2892 45722
rect 5982 45670 6034 45722
rect 6046 45670 6098 45722
rect 6110 45670 6162 45722
rect 6174 45670 6226 45722
rect 4315 45126 4367 45178
rect 4379 45126 4431 45178
rect 4443 45126 4495 45178
rect 4507 45126 4559 45178
rect 7648 45126 7700 45178
rect 7712 45126 7764 45178
rect 7776 45126 7828 45178
rect 7840 45126 7892 45178
rect 2648 44582 2700 44634
rect 2712 44582 2764 44634
rect 2776 44582 2828 44634
rect 2840 44582 2892 44634
rect 5982 44582 6034 44634
rect 6046 44582 6098 44634
rect 6110 44582 6162 44634
rect 6174 44582 6226 44634
rect 4315 44038 4367 44090
rect 4379 44038 4431 44090
rect 4443 44038 4495 44090
rect 4507 44038 4559 44090
rect 7648 44038 7700 44090
rect 7712 44038 7764 44090
rect 7776 44038 7828 44090
rect 7840 44038 7892 44090
rect 2648 43494 2700 43546
rect 2712 43494 2764 43546
rect 2776 43494 2828 43546
rect 2840 43494 2892 43546
rect 5982 43494 6034 43546
rect 6046 43494 6098 43546
rect 6110 43494 6162 43546
rect 6174 43494 6226 43546
rect 4315 42950 4367 43002
rect 4379 42950 4431 43002
rect 4443 42950 4495 43002
rect 4507 42950 4559 43002
rect 7648 42950 7700 43002
rect 7712 42950 7764 43002
rect 7776 42950 7828 43002
rect 7840 42950 7892 43002
rect 2648 42406 2700 42458
rect 2712 42406 2764 42458
rect 2776 42406 2828 42458
rect 2840 42406 2892 42458
rect 5982 42406 6034 42458
rect 6046 42406 6098 42458
rect 6110 42406 6162 42458
rect 6174 42406 6226 42458
rect 4315 41862 4367 41914
rect 4379 41862 4431 41914
rect 4443 41862 4495 41914
rect 4507 41862 4559 41914
rect 7648 41862 7700 41914
rect 7712 41862 7764 41914
rect 7776 41862 7828 41914
rect 7840 41862 7892 41914
rect 2648 41318 2700 41370
rect 2712 41318 2764 41370
rect 2776 41318 2828 41370
rect 2840 41318 2892 41370
rect 5982 41318 6034 41370
rect 6046 41318 6098 41370
rect 6110 41318 6162 41370
rect 6174 41318 6226 41370
rect 4315 40774 4367 40826
rect 4379 40774 4431 40826
rect 4443 40774 4495 40826
rect 4507 40774 4559 40826
rect 7648 40774 7700 40826
rect 7712 40774 7764 40826
rect 7776 40774 7828 40826
rect 7840 40774 7892 40826
rect 2648 40230 2700 40282
rect 2712 40230 2764 40282
rect 2776 40230 2828 40282
rect 2840 40230 2892 40282
rect 5982 40230 6034 40282
rect 6046 40230 6098 40282
rect 6110 40230 6162 40282
rect 6174 40230 6226 40282
rect 4315 39686 4367 39738
rect 4379 39686 4431 39738
rect 4443 39686 4495 39738
rect 4507 39686 4559 39738
rect 7648 39686 7700 39738
rect 7712 39686 7764 39738
rect 7776 39686 7828 39738
rect 7840 39686 7892 39738
rect 2648 39142 2700 39194
rect 2712 39142 2764 39194
rect 2776 39142 2828 39194
rect 2840 39142 2892 39194
rect 5982 39142 6034 39194
rect 6046 39142 6098 39194
rect 6110 39142 6162 39194
rect 6174 39142 6226 39194
rect 4315 38598 4367 38650
rect 4379 38598 4431 38650
rect 4443 38598 4495 38650
rect 4507 38598 4559 38650
rect 7648 38598 7700 38650
rect 7712 38598 7764 38650
rect 7776 38598 7828 38650
rect 7840 38598 7892 38650
rect 2648 38054 2700 38106
rect 2712 38054 2764 38106
rect 2776 38054 2828 38106
rect 2840 38054 2892 38106
rect 5982 38054 6034 38106
rect 6046 38054 6098 38106
rect 6110 38054 6162 38106
rect 6174 38054 6226 38106
rect 4315 37510 4367 37562
rect 4379 37510 4431 37562
rect 4443 37510 4495 37562
rect 4507 37510 4559 37562
rect 7648 37510 7700 37562
rect 7712 37510 7764 37562
rect 7776 37510 7828 37562
rect 7840 37510 7892 37562
rect 2648 36966 2700 37018
rect 2712 36966 2764 37018
rect 2776 36966 2828 37018
rect 2840 36966 2892 37018
rect 5982 36966 6034 37018
rect 6046 36966 6098 37018
rect 6110 36966 6162 37018
rect 6174 36966 6226 37018
rect 4315 36422 4367 36474
rect 4379 36422 4431 36474
rect 4443 36422 4495 36474
rect 4507 36422 4559 36474
rect 7648 36422 7700 36474
rect 7712 36422 7764 36474
rect 7776 36422 7828 36474
rect 7840 36422 7892 36474
rect 2648 35878 2700 35930
rect 2712 35878 2764 35930
rect 2776 35878 2828 35930
rect 2840 35878 2892 35930
rect 5982 35878 6034 35930
rect 6046 35878 6098 35930
rect 6110 35878 6162 35930
rect 6174 35878 6226 35930
rect 4315 35334 4367 35386
rect 4379 35334 4431 35386
rect 4443 35334 4495 35386
rect 4507 35334 4559 35386
rect 7648 35334 7700 35386
rect 7712 35334 7764 35386
rect 7776 35334 7828 35386
rect 7840 35334 7892 35386
rect 2648 34790 2700 34842
rect 2712 34790 2764 34842
rect 2776 34790 2828 34842
rect 2840 34790 2892 34842
rect 5982 34790 6034 34842
rect 6046 34790 6098 34842
rect 6110 34790 6162 34842
rect 6174 34790 6226 34842
rect 4315 34246 4367 34298
rect 4379 34246 4431 34298
rect 4443 34246 4495 34298
rect 4507 34246 4559 34298
rect 7648 34246 7700 34298
rect 7712 34246 7764 34298
rect 7776 34246 7828 34298
rect 7840 34246 7892 34298
rect 2648 33702 2700 33754
rect 2712 33702 2764 33754
rect 2776 33702 2828 33754
rect 2840 33702 2892 33754
rect 5982 33702 6034 33754
rect 6046 33702 6098 33754
rect 6110 33702 6162 33754
rect 6174 33702 6226 33754
rect 4315 33158 4367 33210
rect 4379 33158 4431 33210
rect 4443 33158 4495 33210
rect 4507 33158 4559 33210
rect 7648 33158 7700 33210
rect 7712 33158 7764 33210
rect 7776 33158 7828 33210
rect 7840 33158 7892 33210
rect 2648 32614 2700 32666
rect 2712 32614 2764 32666
rect 2776 32614 2828 32666
rect 2840 32614 2892 32666
rect 5982 32614 6034 32666
rect 6046 32614 6098 32666
rect 6110 32614 6162 32666
rect 6174 32614 6226 32666
rect 4315 32070 4367 32122
rect 4379 32070 4431 32122
rect 4443 32070 4495 32122
rect 4507 32070 4559 32122
rect 7648 32070 7700 32122
rect 7712 32070 7764 32122
rect 7776 32070 7828 32122
rect 7840 32070 7892 32122
rect 2648 31526 2700 31578
rect 2712 31526 2764 31578
rect 2776 31526 2828 31578
rect 2840 31526 2892 31578
rect 5982 31526 6034 31578
rect 6046 31526 6098 31578
rect 6110 31526 6162 31578
rect 6174 31526 6226 31578
rect 4315 30982 4367 31034
rect 4379 30982 4431 31034
rect 4443 30982 4495 31034
rect 4507 30982 4559 31034
rect 7648 30982 7700 31034
rect 7712 30982 7764 31034
rect 7776 30982 7828 31034
rect 7840 30982 7892 31034
rect 2648 30438 2700 30490
rect 2712 30438 2764 30490
rect 2776 30438 2828 30490
rect 2840 30438 2892 30490
rect 5982 30438 6034 30490
rect 6046 30438 6098 30490
rect 6110 30438 6162 30490
rect 6174 30438 6226 30490
rect 4315 29894 4367 29946
rect 4379 29894 4431 29946
rect 4443 29894 4495 29946
rect 4507 29894 4559 29946
rect 7648 29894 7700 29946
rect 7712 29894 7764 29946
rect 7776 29894 7828 29946
rect 7840 29894 7892 29946
rect 2648 29350 2700 29402
rect 2712 29350 2764 29402
rect 2776 29350 2828 29402
rect 2840 29350 2892 29402
rect 5982 29350 6034 29402
rect 6046 29350 6098 29402
rect 6110 29350 6162 29402
rect 6174 29350 6226 29402
rect 4315 28806 4367 28858
rect 4379 28806 4431 28858
rect 4443 28806 4495 28858
rect 4507 28806 4559 28858
rect 7648 28806 7700 28858
rect 7712 28806 7764 28858
rect 7776 28806 7828 28858
rect 7840 28806 7892 28858
rect 2648 28262 2700 28314
rect 2712 28262 2764 28314
rect 2776 28262 2828 28314
rect 2840 28262 2892 28314
rect 5982 28262 6034 28314
rect 6046 28262 6098 28314
rect 6110 28262 6162 28314
rect 6174 28262 6226 28314
rect 4315 27718 4367 27770
rect 4379 27718 4431 27770
rect 4443 27718 4495 27770
rect 4507 27718 4559 27770
rect 7648 27718 7700 27770
rect 7712 27718 7764 27770
rect 7776 27718 7828 27770
rect 7840 27718 7892 27770
rect 2648 27174 2700 27226
rect 2712 27174 2764 27226
rect 2776 27174 2828 27226
rect 2840 27174 2892 27226
rect 5982 27174 6034 27226
rect 6046 27174 6098 27226
rect 6110 27174 6162 27226
rect 6174 27174 6226 27226
rect 4315 26630 4367 26682
rect 4379 26630 4431 26682
rect 4443 26630 4495 26682
rect 4507 26630 4559 26682
rect 7648 26630 7700 26682
rect 7712 26630 7764 26682
rect 7776 26630 7828 26682
rect 7840 26630 7892 26682
rect 2648 26086 2700 26138
rect 2712 26086 2764 26138
rect 2776 26086 2828 26138
rect 2840 26086 2892 26138
rect 5982 26086 6034 26138
rect 6046 26086 6098 26138
rect 6110 26086 6162 26138
rect 6174 26086 6226 26138
rect 4315 25542 4367 25594
rect 4379 25542 4431 25594
rect 4443 25542 4495 25594
rect 4507 25542 4559 25594
rect 7648 25542 7700 25594
rect 7712 25542 7764 25594
rect 7776 25542 7828 25594
rect 7840 25542 7892 25594
rect 2648 24998 2700 25050
rect 2712 24998 2764 25050
rect 2776 24998 2828 25050
rect 2840 24998 2892 25050
rect 5982 24998 6034 25050
rect 6046 24998 6098 25050
rect 6110 24998 6162 25050
rect 6174 24998 6226 25050
rect 4315 24454 4367 24506
rect 4379 24454 4431 24506
rect 4443 24454 4495 24506
rect 4507 24454 4559 24506
rect 7648 24454 7700 24506
rect 7712 24454 7764 24506
rect 7776 24454 7828 24506
rect 7840 24454 7892 24506
rect 2648 23910 2700 23962
rect 2712 23910 2764 23962
rect 2776 23910 2828 23962
rect 2840 23910 2892 23962
rect 5982 23910 6034 23962
rect 6046 23910 6098 23962
rect 6110 23910 6162 23962
rect 6174 23910 6226 23962
rect 4315 23366 4367 23418
rect 4379 23366 4431 23418
rect 4443 23366 4495 23418
rect 4507 23366 4559 23418
rect 7648 23366 7700 23418
rect 7712 23366 7764 23418
rect 7776 23366 7828 23418
rect 7840 23366 7892 23418
rect 2648 22822 2700 22874
rect 2712 22822 2764 22874
rect 2776 22822 2828 22874
rect 2840 22822 2892 22874
rect 5982 22822 6034 22874
rect 6046 22822 6098 22874
rect 6110 22822 6162 22874
rect 6174 22822 6226 22874
rect 4315 22278 4367 22330
rect 4379 22278 4431 22330
rect 4443 22278 4495 22330
rect 4507 22278 4559 22330
rect 7648 22278 7700 22330
rect 7712 22278 7764 22330
rect 7776 22278 7828 22330
rect 7840 22278 7892 22330
rect 2648 21734 2700 21786
rect 2712 21734 2764 21786
rect 2776 21734 2828 21786
rect 2840 21734 2892 21786
rect 5982 21734 6034 21786
rect 6046 21734 6098 21786
rect 6110 21734 6162 21786
rect 6174 21734 6226 21786
rect 4315 21190 4367 21242
rect 4379 21190 4431 21242
rect 4443 21190 4495 21242
rect 4507 21190 4559 21242
rect 7648 21190 7700 21242
rect 7712 21190 7764 21242
rect 7776 21190 7828 21242
rect 7840 21190 7892 21242
rect 2648 20646 2700 20698
rect 2712 20646 2764 20698
rect 2776 20646 2828 20698
rect 2840 20646 2892 20698
rect 5982 20646 6034 20698
rect 6046 20646 6098 20698
rect 6110 20646 6162 20698
rect 6174 20646 6226 20698
rect 4315 20102 4367 20154
rect 4379 20102 4431 20154
rect 4443 20102 4495 20154
rect 4507 20102 4559 20154
rect 7648 20102 7700 20154
rect 7712 20102 7764 20154
rect 7776 20102 7828 20154
rect 7840 20102 7892 20154
rect 2648 19558 2700 19610
rect 2712 19558 2764 19610
rect 2776 19558 2828 19610
rect 2840 19558 2892 19610
rect 5982 19558 6034 19610
rect 6046 19558 6098 19610
rect 6110 19558 6162 19610
rect 6174 19558 6226 19610
rect 4315 19014 4367 19066
rect 4379 19014 4431 19066
rect 4443 19014 4495 19066
rect 4507 19014 4559 19066
rect 7648 19014 7700 19066
rect 7712 19014 7764 19066
rect 7776 19014 7828 19066
rect 7840 19014 7892 19066
rect 2648 18470 2700 18522
rect 2712 18470 2764 18522
rect 2776 18470 2828 18522
rect 2840 18470 2892 18522
rect 5982 18470 6034 18522
rect 6046 18470 6098 18522
rect 6110 18470 6162 18522
rect 6174 18470 6226 18522
rect 4315 17926 4367 17978
rect 4379 17926 4431 17978
rect 4443 17926 4495 17978
rect 4507 17926 4559 17978
rect 7648 17926 7700 17978
rect 7712 17926 7764 17978
rect 7776 17926 7828 17978
rect 7840 17926 7892 17978
rect 2648 17382 2700 17434
rect 2712 17382 2764 17434
rect 2776 17382 2828 17434
rect 2840 17382 2892 17434
rect 5982 17382 6034 17434
rect 6046 17382 6098 17434
rect 6110 17382 6162 17434
rect 6174 17382 6226 17434
rect 4315 16838 4367 16890
rect 4379 16838 4431 16890
rect 4443 16838 4495 16890
rect 4507 16838 4559 16890
rect 7648 16838 7700 16890
rect 7712 16838 7764 16890
rect 7776 16838 7828 16890
rect 7840 16838 7892 16890
rect 2648 16294 2700 16346
rect 2712 16294 2764 16346
rect 2776 16294 2828 16346
rect 2840 16294 2892 16346
rect 5982 16294 6034 16346
rect 6046 16294 6098 16346
rect 6110 16294 6162 16346
rect 6174 16294 6226 16346
rect 4315 15750 4367 15802
rect 4379 15750 4431 15802
rect 4443 15750 4495 15802
rect 4507 15750 4559 15802
rect 7648 15750 7700 15802
rect 7712 15750 7764 15802
rect 7776 15750 7828 15802
rect 7840 15750 7892 15802
rect 2648 15206 2700 15258
rect 2712 15206 2764 15258
rect 2776 15206 2828 15258
rect 2840 15206 2892 15258
rect 5982 15206 6034 15258
rect 6046 15206 6098 15258
rect 6110 15206 6162 15258
rect 6174 15206 6226 15258
rect 4315 14662 4367 14714
rect 4379 14662 4431 14714
rect 4443 14662 4495 14714
rect 4507 14662 4559 14714
rect 7648 14662 7700 14714
rect 7712 14662 7764 14714
rect 7776 14662 7828 14714
rect 7840 14662 7892 14714
rect 2648 14118 2700 14170
rect 2712 14118 2764 14170
rect 2776 14118 2828 14170
rect 2840 14118 2892 14170
rect 5982 14118 6034 14170
rect 6046 14118 6098 14170
rect 6110 14118 6162 14170
rect 6174 14118 6226 14170
rect 4315 13574 4367 13626
rect 4379 13574 4431 13626
rect 4443 13574 4495 13626
rect 4507 13574 4559 13626
rect 7648 13574 7700 13626
rect 7712 13574 7764 13626
rect 7776 13574 7828 13626
rect 7840 13574 7892 13626
rect 2648 13030 2700 13082
rect 2712 13030 2764 13082
rect 2776 13030 2828 13082
rect 2840 13030 2892 13082
rect 5982 13030 6034 13082
rect 6046 13030 6098 13082
rect 6110 13030 6162 13082
rect 6174 13030 6226 13082
rect 4315 12486 4367 12538
rect 4379 12486 4431 12538
rect 4443 12486 4495 12538
rect 4507 12486 4559 12538
rect 7648 12486 7700 12538
rect 7712 12486 7764 12538
rect 7776 12486 7828 12538
rect 7840 12486 7892 12538
rect 2648 11942 2700 11994
rect 2712 11942 2764 11994
rect 2776 11942 2828 11994
rect 2840 11942 2892 11994
rect 5982 11942 6034 11994
rect 6046 11942 6098 11994
rect 6110 11942 6162 11994
rect 6174 11942 6226 11994
rect 4315 11398 4367 11450
rect 4379 11398 4431 11450
rect 4443 11398 4495 11450
rect 4507 11398 4559 11450
rect 7648 11398 7700 11450
rect 7712 11398 7764 11450
rect 7776 11398 7828 11450
rect 7840 11398 7892 11450
rect 2648 10854 2700 10906
rect 2712 10854 2764 10906
rect 2776 10854 2828 10906
rect 2840 10854 2892 10906
rect 5982 10854 6034 10906
rect 6046 10854 6098 10906
rect 6110 10854 6162 10906
rect 6174 10854 6226 10906
rect 4315 10310 4367 10362
rect 4379 10310 4431 10362
rect 4443 10310 4495 10362
rect 4507 10310 4559 10362
rect 7648 10310 7700 10362
rect 7712 10310 7764 10362
rect 7776 10310 7828 10362
rect 7840 10310 7892 10362
rect 2648 9766 2700 9818
rect 2712 9766 2764 9818
rect 2776 9766 2828 9818
rect 2840 9766 2892 9818
rect 5982 9766 6034 9818
rect 6046 9766 6098 9818
rect 6110 9766 6162 9818
rect 6174 9766 6226 9818
rect 4315 9222 4367 9274
rect 4379 9222 4431 9274
rect 4443 9222 4495 9274
rect 4507 9222 4559 9274
rect 7648 9222 7700 9274
rect 7712 9222 7764 9274
rect 7776 9222 7828 9274
rect 7840 9222 7892 9274
rect 2648 8678 2700 8730
rect 2712 8678 2764 8730
rect 2776 8678 2828 8730
rect 2840 8678 2892 8730
rect 5982 8678 6034 8730
rect 6046 8678 6098 8730
rect 6110 8678 6162 8730
rect 6174 8678 6226 8730
rect 4315 8134 4367 8186
rect 4379 8134 4431 8186
rect 4443 8134 4495 8186
rect 4507 8134 4559 8186
rect 7648 8134 7700 8186
rect 7712 8134 7764 8186
rect 7776 8134 7828 8186
rect 7840 8134 7892 8186
rect 2648 7590 2700 7642
rect 2712 7590 2764 7642
rect 2776 7590 2828 7642
rect 2840 7590 2892 7642
rect 5982 7590 6034 7642
rect 6046 7590 6098 7642
rect 6110 7590 6162 7642
rect 6174 7590 6226 7642
rect 4315 7046 4367 7098
rect 4379 7046 4431 7098
rect 4443 7046 4495 7098
rect 4507 7046 4559 7098
rect 7648 7046 7700 7098
rect 7712 7046 7764 7098
rect 7776 7046 7828 7098
rect 7840 7046 7892 7098
rect 2648 6502 2700 6554
rect 2712 6502 2764 6554
rect 2776 6502 2828 6554
rect 2840 6502 2892 6554
rect 5982 6502 6034 6554
rect 6046 6502 6098 6554
rect 6110 6502 6162 6554
rect 6174 6502 6226 6554
rect 4315 5958 4367 6010
rect 4379 5958 4431 6010
rect 4443 5958 4495 6010
rect 4507 5958 4559 6010
rect 7648 5958 7700 6010
rect 7712 5958 7764 6010
rect 7776 5958 7828 6010
rect 7840 5958 7892 6010
rect 2648 5414 2700 5466
rect 2712 5414 2764 5466
rect 2776 5414 2828 5466
rect 2840 5414 2892 5466
rect 5982 5414 6034 5466
rect 6046 5414 6098 5466
rect 6110 5414 6162 5466
rect 6174 5414 6226 5466
rect 4315 4870 4367 4922
rect 4379 4870 4431 4922
rect 4443 4870 4495 4922
rect 4507 4870 4559 4922
rect 7648 4870 7700 4922
rect 7712 4870 7764 4922
rect 7776 4870 7828 4922
rect 7840 4870 7892 4922
rect 2648 4326 2700 4378
rect 2712 4326 2764 4378
rect 2776 4326 2828 4378
rect 2840 4326 2892 4378
rect 5982 4326 6034 4378
rect 6046 4326 6098 4378
rect 6110 4326 6162 4378
rect 6174 4326 6226 4378
rect 4315 3782 4367 3834
rect 4379 3782 4431 3834
rect 4443 3782 4495 3834
rect 4507 3782 4559 3834
rect 7648 3782 7700 3834
rect 7712 3782 7764 3834
rect 7776 3782 7828 3834
rect 7840 3782 7892 3834
rect 2648 3238 2700 3290
rect 2712 3238 2764 3290
rect 2776 3238 2828 3290
rect 2840 3238 2892 3290
rect 5982 3238 6034 3290
rect 6046 3238 6098 3290
rect 6110 3238 6162 3290
rect 6174 3238 6226 3290
rect 4315 2694 4367 2746
rect 4379 2694 4431 2746
rect 4443 2694 4495 2746
rect 4507 2694 4559 2746
rect 7648 2694 7700 2746
rect 7712 2694 7764 2746
rect 7776 2694 7828 2746
rect 7840 2694 7892 2746
rect 2648 2150 2700 2202
rect 2712 2150 2764 2202
rect 2776 2150 2828 2202
rect 2840 2150 2892 2202
rect 5982 2150 6034 2202
rect 6046 2150 6098 2202
rect 6110 2150 6162 2202
rect 6174 2150 6226 2202
rect 8208 76 8260 128
rect 8944 76 8996 128
<< metal2 >>
rect 570 332580 626 333000
rect 1766 332602 1822 333000
rect 570 332528 572 332580
rect 624 332528 626 332580
rect 570 332520 626 332528
rect 1216 332580 1268 332586
rect 1216 332522 1268 332528
rect 1504 332574 1822 332602
rect 584 332491 612 332520
rect 1228 228342 1256 332522
rect 1504 229974 1532 332574
rect 1766 332520 1822 332574
rect 3054 332580 3110 333000
rect 3054 332528 3056 332580
rect 3108 332528 3110 332580
rect 3054 332520 3110 332528
rect 3884 332580 3936 332586
rect 3884 332522 3936 332528
rect 4250 332580 4306 333000
rect 5538 332602 5594 333000
rect 6826 332602 6882 333000
rect 8022 332602 8078 333000
rect 4250 332528 4252 332580
rect 4304 332528 4306 332580
rect 3068 332491 3096 332520
rect 2622 330780 2918 330800
rect 2678 330778 2702 330780
rect 2758 330778 2782 330780
rect 2838 330778 2862 330780
rect 2700 330726 2702 330778
rect 2764 330726 2776 330778
rect 2838 330726 2840 330778
rect 2678 330724 2702 330726
rect 2758 330724 2782 330726
rect 2838 330724 2862 330726
rect 2622 330704 2918 330724
rect 2622 329692 2918 329712
rect 2678 329690 2702 329692
rect 2758 329690 2782 329692
rect 2838 329690 2862 329692
rect 2700 329638 2702 329690
rect 2764 329638 2776 329690
rect 2838 329638 2840 329690
rect 2678 329636 2702 329638
rect 2758 329636 2782 329638
rect 2838 329636 2862 329638
rect 2622 329616 2918 329636
rect 2622 328604 2918 328624
rect 2678 328602 2702 328604
rect 2758 328602 2782 328604
rect 2838 328602 2862 328604
rect 2700 328550 2702 328602
rect 2764 328550 2776 328602
rect 2838 328550 2840 328602
rect 2678 328548 2702 328550
rect 2758 328548 2782 328550
rect 2838 328548 2862 328550
rect 2622 328528 2918 328548
rect 2622 327516 2918 327536
rect 2678 327514 2702 327516
rect 2758 327514 2782 327516
rect 2838 327514 2862 327516
rect 2700 327462 2702 327514
rect 2764 327462 2776 327514
rect 2838 327462 2840 327514
rect 2678 327460 2702 327462
rect 2758 327460 2782 327462
rect 2838 327460 2862 327462
rect 2622 327440 2918 327460
rect 2622 326428 2918 326448
rect 2678 326426 2702 326428
rect 2758 326426 2782 326428
rect 2838 326426 2862 326428
rect 2700 326374 2702 326426
rect 2764 326374 2776 326426
rect 2838 326374 2840 326426
rect 2678 326372 2702 326374
rect 2758 326372 2782 326374
rect 2838 326372 2862 326374
rect 2622 326352 2918 326372
rect 2622 325340 2918 325360
rect 2678 325338 2702 325340
rect 2758 325338 2782 325340
rect 2838 325338 2862 325340
rect 2700 325286 2702 325338
rect 2764 325286 2776 325338
rect 2838 325286 2840 325338
rect 2678 325284 2702 325286
rect 2758 325284 2782 325286
rect 2838 325284 2862 325286
rect 2622 325264 2918 325284
rect 2622 324252 2918 324272
rect 2678 324250 2702 324252
rect 2758 324250 2782 324252
rect 2838 324250 2862 324252
rect 2700 324198 2702 324250
rect 2764 324198 2776 324250
rect 2838 324198 2840 324250
rect 2678 324196 2702 324198
rect 2758 324196 2782 324198
rect 2838 324196 2862 324198
rect 2622 324176 2918 324196
rect 2622 323164 2918 323184
rect 2678 323162 2702 323164
rect 2758 323162 2782 323164
rect 2838 323162 2862 323164
rect 2700 323110 2702 323162
rect 2764 323110 2776 323162
rect 2838 323110 2840 323162
rect 2678 323108 2702 323110
rect 2758 323108 2782 323110
rect 2838 323108 2862 323110
rect 2622 323088 2918 323108
rect 2622 322076 2918 322096
rect 2678 322074 2702 322076
rect 2758 322074 2782 322076
rect 2838 322074 2862 322076
rect 2700 322022 2702 322074
rect 2764 322022 2776 322074
rect 2838 322022 2840 322074
rect 2678 322020 2702 322022
rect 2758 322020 2782 322022
rect 2838 322020 2862 322022
rect 2622 322000 2918 322020
rect 2622 320988 2918 321008
rect 2678 320986 2702 320988
rect 2758 320986 2782 320988
rect 2838 320986 2862 320988
rect 2700 320934 2702 320986
rect 2764 320934 2776 320986
rect 2838 320934 2840 320986
rect 2678 320932 2702 320934
rect 2758 320932 2782 320934
rect 2838 320932 2862 320934
rect 2622 320912 2918 320932
rect 2622 319900 2918 319920
rect 2678 319898 2702 319900
rect 2758 319898 2782 319900
rect 2838 319898 2862 319900
rect 2700 319846 2702 319898
rect 2764 319846 2776 319898
rect 2838 319846 2840 319898
rect 2678 319844 2702 319846
rect 2758 319844 2782 319846
rect 2838 319844 2862 319846
rect 2622 319824 2918 319844
rect 2622 318812 2918 318832
rect 2678 318810 2702 318812
rect 2758 318810 2782 318812
rect 2838 318810 2862 318812
rect 2700 318758 2702 318810
rect 2764 318758 2776 318810
rect 2838 318758 2840 318810
rect 2678 318756 2702 318758
rect 2758 318756 2782 318758
rect 2838 318756 2862 318758
rect 2622 318736 2918 318756
rect 2622 317724 2918 317744
rect 2678 317722 2702 317724
rect 2758 317722 2782 317724
rect 2838 317722 2862 317724
rect 2700 317670 2702 317722
rect 2764 317670 2776 317722
rect 2838 317670 2840 317722
rect 2678 317668 2702 317670
rect 2758 317668 2782 317670
rect 2838 317668 2862 317670
rect 2622 317648 2918 317668
rect 2622 316636 2918 316656
rect 2678 316634 2702 316636
rect 2758 316634 2782 316636
rect 2838 316634 2862 316636
rect 2700 316582 2702 316634
rect 2764 316582 2776 316634
rect 2838 316582 2840 316634
rect 2678 316580 2702 316582
rect 2758 316580 2782 316582
rect 2838 316580 2862 316582
rect 2622 316560 2918 316580
rect 2622 315548 2918 315568
rect 2678 315546 2702 315548
rect 2758 315546 2782 315548
rect 2838 315546 2862 315548
rect 2700 315494 2702 315546
rect 2764 315494 2776 315546
rect 2838 315494 2840 315546
rect 2678 315492 2702 315494
rect 2758 315492 2782 315494
rect 2838 315492 2862 315494
rect 2622 315472 2918 315492
rect 2622 314460 2918 314480
rect 2678 314458 2702 314460
rect 2758 314458 2782 314460
rect 2838 314458 2862 314460
rect 2700 314406 2702 314458
rect 2764 314406 2776 314458
rect 2838 314406 2840 314458
rect 2678 314404 2702 314406
rect 2758 314404 2782 314406
rect 2838 314404 2862 314406
rect 2622 314384 2918 314404
rect 2622 313372 2918 313392
rect 2678 313370 2702 313372
rect 2758 313370 2782 313372
rect 2838 313370 2862 313372
rect 2700 313318 2702 313370
rect 2764 313318 2776 313370
rect 2838 313318 2840 313370
rect 2678 313316 2702 313318
rect 2758 313316 2782 313318
rect 2838 313316 2862 313318
rect 2622 313296 2918 313316
rect 2622 312284 2918 312304
rect 2678 312282 2702 312284
rect 2758 312282 2782 312284
rect 2838 312282 2862 312284
rect 2700 312230 2702 312282
rect 2764 312230 2776 312282
rect 2838 312230 2840 312282
rect 2678 312228 2702 312230
rect 2758 312228 2782 312230
rect 2838 312228 2862 312230
rect 2622 312208 2918 312228
rect 2622 311196 2918 311216
rect 2678 311194 2702 311196
rect 2758 311194 2782 311196
rect 2838 311194 2862 311196
rect 2700 311142 2702 311194
rect 2764 311142 2776 311194
rect 2838 311142 2840 311194
rect 2678 311140 2702 311142
rect 2758 311140 2782 311142
rect 2838 311140 2862 311142
rect 2622 311120 2918 311140
rect 2622 310108 2918 310128
rect 2678 310106 2702 310108
rect 2758 310106 2782 310108
rect 2838 310106 2862 310108
rect 2700 310054 2702 310106
rect 2764 310054 2776 310106
rect 2838 310054 2840 310106
rect 2678 310052 2702 310054
rect 2758 310052 2782 310054
rect 2838 310052 2862 310054
rect 2622 310032 2918 310052
rect 2622 309020 2918 309040
rect 2678 309018 2702 309020
rect 2758 309018 2782 309020
rect 2838 309018 2862 309020
rect 2700 308966 2702 309018
rect 2764 308966 2776 309018
rect 2838 308966 2840 309018
rect 2678 308964 2702 308966
rect 2758 308964 2782 308966
rect 2838 308964 2862 308966
rect 2622 308944 2918 308964
rect 2226 308680 2282 308689
rect 2226 308615 2282 308624
rect 2240 244730 2268 308615
rect 2622 307932 2918 307952
rect 2678 307930 2702 307932
rect 2758 307930 2782 307932
rect 2838 307930 2862 307932
rect 2700 307878 2702 307930
rect 2764 307878 2776 307930
rect 2838 307878 2840 307930
rect 2678 307876 2702 307878
rect 2758 307876 2782 307878
rect 2838 307876 2862 307878
rect 2622 307856 2918 307876
rect 2622 306844 2918 306864
rect 2678 306842 2702 306844
rect 2758 306842 2782 306844
rect 2838 306842 2862 306844
rect 2700 306790 2702 306842
rect 2764 306790 2776 306842
rect 2838 306790 2840 306842
rect 2678 306788 2702 306790
rect 2758 306788 2782 306790
rect 2838 306788 2862 306790
rect 2622 306768 2918 306788
rect 2622 305756 2918 305776
rect 2678 305754 2702 305756
rect 2758 305754 2782 305756
rect 2838 305754 2862 305756
rect 2700 305702 2702 305754
rect 2764 305702 2776 305754
rect 2838 305702 2840 305754
rect 2678 305700 2702 305702
rect 2758 305700 2782 305702
rect 2838 305700 2862 305702
rect 2622 305680 2918 305700
rect 2622 304668 2918 304688
rect 2678 304666 2702 304668
rect 2758 304666 2782 304668
rect 2838 304666 2862 304668
rect 2700 304614 2702 304666
rect 2764 304614 2776 304666
rect 2838 304614 2840 304666
rect 2678 304612 2702 304614
rect 2758 304612 2782 304614
rect 2838 304612 2862 304614
rect 2622 304592 2918 304612
rect 2622 303580 2918 303600
rect 2678 303578 2702 303580
rect 2758 303578 2782 303580
rect 2838 303578 2862 303580
rect 2700 303526 2702 303578
rect 2764 303526 2776 303578
rect 2838 303526 2840 303578
rect 2678 303524 2702 303526
rect 2758 303524 2782 303526
rect 2838 303524 2862 303526
rect 2622 303504 2918 303524
rect 2622 302492 2918 302512
rect 2678 302490 2702 302492
rect 2758 302490 2782 302492
rect 2838 302490 2862 302492
rect 2700 302438 2702 302490
rect 2764 302438 2776 302490
rect 2838 302438 2840 302490
rect 2678 302436 2702 302438
rect 2758 302436 2782 302438
rect 2838 302436 2862 302438
rect 2622 302416 2918 302436
rect 2622 301404 2918 301424
rect 2678 301402 2702 301404
rect 2758 301402 2782 301404
rect 2838 301402 2862 301404
rect 2700 301350 2702 301402
rect 2764 301350 2776 301402
rect 2838 301350 2840 301402
rect 2678 301348 2702 301350
rect 2758 301348 2782 301350
rect 2838 301348 2862 301350
rect 2622 301328 2918 301348
rect 2622 300316 2918 300336
rect 2678 300314 2702 300316
rect 2758 300314 2782 300316
rect 2838 300314 2862 300316
rect 2700 300262 2702 300314
rect 2764 300262 2776 300314
rect 2838 300262 2840 300314
rect 2678 300260 2702 300262
rect 2758 300260 2782 300262
rect 2838 300260 2862 300262
rect 2622 300240 2918 300260
rect 2622 299228 2918 299248
rect 2678 299226 2702 299228
rect 2758 299226 2782 299228
rect 2838 299226 2862 299228
rect 2700 299174 2702 299226
rect 2764 299174 2776 299226
rect 2838 299174 2840 299226
rect 2678 299172 2702 299174
rect 2758 299172 2782 299174
rect 2838 299172 2862 299174
rect 2622 299152 2918 299172
rect 2622 298140 2918 298160
rect 2678 298138 2702 298140
rect 2758 298138 2782 298140
rect 2838 298138 2862 298140
rect 2700 298086 2702 298138
rect 2764 298086 2776 298138
rect 2838 298086 2840 298138
rect 2678 298084 2702 298086
rect 2758 298084 2782 298086
rect 2838 298084 2862 298086
rect 2622 298064 2918 298084
rect 2622 297052 2918 297072
rect 2678 297050 2702 297052
rect 2758 297050 2782 297052
rect 2838 297050 2862 297052
rect 2700 296998 2702 297050
rect 2764 296998 2776 297050
rect 2838 296998 2840 297050
rect 2678 296996 2702 296998
rect 2758 296996 2782 296998
rect 2838 296996 2862 296998
rect 2622 296976 2918 296996
rect 2622 295964 2918 295984
rect 2678 295962 2702 295964
rect 2758 295962 2782 295964
rect 2838 295962 2862 295964
rect 2700 295910 2702 295962
rect 2764 295910 2776 295962
rect 2838 295910 2840 295962
rect 2678 295908 2702 295910
rect 2758 295908 2782 295910
rect 2838 295908 2862 295910
rect 2622 295888 2918 295908
rect 2622 294876 2918 294896
rect 2678 294874 2702 294876
rect 2758 294874 2782 294876
rect 2838 294874 2862 294876
rect 2700 294822 2702 294874
rect 2764 294822 2776 294874
rect 2838 294822 2840 294874
rect 2678 294820 2702 294822
rect 2758 294820 2782 294822
rect 2838 294820 2862 294822
rect 2622 294800 2918 294820
rect 2622 293788 2918 293808
rect 2678 293786 2702 293788
rect 2758 293786 2782 293788
rect 2838 293786 2862 293788
rect 2700 293734 2702 293786
rect 2764 293734 2776 293786
rect 2838 293734 2840 293786
rect 2678 293732 2702 293734
rect 2758 293732 2782 293734
rect 2838 293732 2862 293734
rect 2622 293712 2918 293732
rect 2622 292700 2918 292720
rect 2678 292698 2702 292700
rect 2758 292698 2782 292700
rect 2838 292698 2862 292700
rect 2700 292646 2702 292698
rect 2764 292646 2776 292698
rect 2838 292646 2840 292698
rect 2678 292644 2702 292646
rect 2758 292644 2782 292646
rect 2838 292644 2862 292646
rect 2622 292624 2918 292644
rect 2622 291612 2918 291632
rect 2678 291610 2702 291612
rect 2758 291610 2782 291612
rect 2838 291610 2862 291612
rect 2700 291558 2702 291610
rect 2764 291558 2776 291610
rect 2838 291558 2840 291610
rect 2678 291556 2702 291558
rect 2758 291556 2782 291558
rect 2838 291556 2862 291558
rect 2622 291536 2918 291556
rect 2622 290524 2918 290544
rect 2678 290522 2702 290524
rect 2758 290522 2782 290524
rect 2838 290522 2862 290524
rect 2700 290470 2702 290522
rect 2764 290470 2776 290522
rect 2838 290470 2840 290522
rect 2678 290468 2702 290470
rect 2758 290468 2782 290470
rect 2838 290468 2862 290470
rect 2622 290448 2918 290468
rect 2622 289436 2918 289456
rect 2678 289434 2702 289436
rect 2758 289434 2782 289436
rect 2838 289434 2862 289436
rect 2700 289382 2702 289434
rect 2764 289382 2776 289434
rect 2838 289382 2840 289434
rect 2678 289380 2702 289382
rect 2758 289380 2782 289382
rect 2838 289380 2862 289382
rect 2622 289360 2918 289380
rect 2622 288348 2918 288368
rect 2678 288346 2702 288348
rect 2758 288346 2782 288348
rect 2838 288346 2862 288348
rect 2700 288294 2702 288346
rect 2764 288294 2776 288346
rect 2838 288294 2840 288346
rect 2678 288292 2702 288294
rect 2758 288292 2782 288294
rect 2838 288292 2862 288294
rect 2622 288272 2918 288292
rect 2622 287260 2918 287280
rect 2678 287258 2702 287260
rect 2758 287258 2782 287260
rect 2838 287258 2862 287260
rect 2700 287206 2702 287258
rect 2764 287206 2776 287258
rect 2838 287206 2840 287258
rect 2678 287204 2702 287206
rect 2758 287204 2782 287206
rect 2838 287204 2862 287206
rect 2622 287184 2918 287204
rect 2622 286172 2918 286192
rect 2678 286170 2702 286172
rect 2758 286170 2782 286172
rect 2838 286170 2862 286172
rect 2700 286118 2702 286170
rect 2764 286118 2776 286170
rect 2838 286118 2840 286170
rect 2678 286116 2702 286118
rect 2758 286116 2782 286118
rect 2838 286116 2862 286118
rect 2622 286096 2918 286116
rect 2622 285084 2918 285104
rect 2678 285082 2702 285084
rect 2758 285082 2782 285084
rect 2838 285082 2862 285084
rect 2700 285030 2702 285082
rect 2764 285030 2776 285082
rect 2838 285030 2840 285082
rect 2678 285028 2702 285030
rect 2758 285028 2782 285030
rect 2838 285028 2862 285030
rect 2622 285008 2918 285028
rect 2622 283996 2918 284016
rect 2678 283994 2702 283996
rect 2758 283994 2782 283996
rect 2838 283994 2862 283996
rect 2700 283942 2702 283994
rect 2764 283942 2776 283994
rect 2838 283942 2840 283994
rect 2678 283940 2702 283942
rect 2758 283940 2782 283942
rect 2838 283940 2862 283942
rect 2622 283920 2918 283940
rect 2622 282908 2918 282928
rect 2678 282906 2702 282908
rect 2758 282906 2782 282908
rect 2838 282906 2862 282908
rect 2700 282854 2702 282906
rect 2764 282854 2776 282906
rect 2838 282854 2840 282906
rect 2678 282852 2702 282854
rect 2758 282852 2782 282854
rect 2838 282852 2862 282854
rect 2622 282832 2918 282852
rect 2622 281820 2918 281840
rect 2678 281818 2702 281820
rect 2758 281818 2782 281820
rect 2838 281818 2862 281820
rect 2700 281766 2702 281818
rect 2764 281766 2776 281818
rect 2838 281766 2840 281818
rect 2678 281764 2702 281766
rect 2758 281764 2782 281766
rect 2838 281764 2862 281766
rect 2622 281744 2918 281764
rect 2622 280732 2918 280752
rect 2678 280730 2702 280732
rect 2758 280730 2782 280732
rect 2838 280730 2862 280732
rect 2700 280678 2702 280730
rect 2764 280678 2776 280730
rect 2838 280678 2840 280730
rect 2678 280676 2702 280678
rect 2758 280676 2782 280678
rect 2838 280676 2862 280678
rect 2622 280656 2918 280676
rect 2622 279644 2918 279664
rect 2678 279642 2702 279644
rect 2758 279642 2782 279644
rect 2838 279642 2862 279644
rect 2700 279590 2702 279642
rect 2764 279590 2776 279642
rect 2838 279590 2840 279642
rect 2678 279588 2702 279590
rect 2758 279588 2782 279590
rect 2838 279588 2862 279590
rect 2622 279568 2918 279588
rect 2622 278556 2918 278576
rect 2678 278554 2702 278556
rect 2758 278554 2782 278556
rect 2838 278554 2862 278556
rect 2700 278502 2702 278554
rect 2764 278502 2776 278554
rect 2838 278502 2840 278554
rect 2678 278500 2702 278502
rect 2758 278500 2782 278502
rect 2838 278500 2862 278502
rect 2622 278480 2918 278500
rect 2622 277468 2918 277488
rect 2678 277466 2702 277468
rect 2758 277466 2782 277468
rect 2838 277466 2862 277468
rect 2700 277414 2702 277466
rect 2764 277414 2776 277466
rect 2838 277414 2840 277466
rect 2678 277412 2702 277414
rect 2758 277412 2782 277414
rect 2838 277412 2862 277414
rect 2622 277392 2918 277412
rect 2622 276380 2918 276400
rect 2678 276378 2702 276380
rect 2758 276378 2782 276380
rect 2838 276378 2862 276380
rect 2700 276326 2702 276378
rect 2764 276326 2776 276378
rect 2838 276326 2840 276378
rect 2678 276324 2702 276326
rect 2758 276324 2782 276326
rect 2838 276324 2862 276326
rect 2622 276304 2918 276324
rect 2622 275292 2918 275312
rect 2678 275290 2702 275292
rect 2758 275290 2782 275292
rect 2838 275290 2862 275292
rect 2700 275238 2702 275290
rect 2764 275238 2776 275290
rect 2838 275238 2840 275290
rect 2678 275236 2702 275238
rect 2758 275236 2782 275238
rect 2838 275236 2862 275238
rect 2622 275216 2918 275236
rect 2622 274204 2918 274224
rect 2678 274202 2702 274204
rect 2758 274202 2782 274204
rect 2838 274202 2862 274204
rect 2700 274150 2702 274202
rect 2764 274150 2776 274202
rect 2838 274150 2840 274202
rect 2678 274148 2702 274150
rect 2758 274148 2782 274150
rect 2838 274148 2862 274150
rect 2622 274128 2918 274148
rect 2622 273116 2918 273136
rect 2678 273114 2702 273116
rect 2758 273114 2782 273116
rect 2838 273114 2862 273116
rect 2700 273062 2702 273114
rect 2764 273062 2776 273114
rect 2838 273062 2840 273114
rect 2678 273060 2702 273062
rect 2758 273060 2782 273062
rect 2838 273060 2862 273062
rect 2622 273040 2918 273060
rect 2622 272028 2918 272048
rect 2678 272026 2702 272028
rect 2758 272026 2782 272028
rect 2838 272026 2862 272028
rect 2700 271974 2702 272026
rect 2764 271974 2776 272026
rect 2838 271974 2840 272026
rect 2678 271972 2702 271974
rect 2758 271972 2782 271974
rect 2838 271972 2862 271974
rect 2622 271952 2918 271972
rect 2622 270940 2918 270960
rect 2678 270938 2702 270940
rect 2758 270938 2782 270940
rect 2838 270938 2862 270940
rect 2700 270886 2702 270938
rect 2764 270886 2776 270938
rect 2838 270886 2840 270938
rect 2678 270884 2702 270886
rect 2758 270884 2782 270886
rect 2838 270884 2862 270886
rect 2622 270864 2918 270884
rect 2622 269852 2918 269872
rect 2678 269850 2702 269852
rect 2758 269850 2782 269852
rect 2838 269850 2862 269852
rect 2700 269798 2702 269850
rect 2764 269798 2776 269850
rect 2838 269798 2840 269850
rect 2678 269796 2702 269798
rect 2758 269796 2782 269798
rect 2838 269796 2862 269798
rect 2622 269776 2918 269796
rect 2622 268764 2918 268784
rect 2678 268762 2702 268764
rect 2758 268762 2782 268764
rect 2838 268762 2862 268764
rect 2700 268710 2702 268762
rect 2764 268710 2776 268762
rect 2838 268710 2840 268762
rect 2678 268708 2702 268710
rect 2758 268708 2782 268710
rect 2838 268708 2862 268710
rect 2622 268688 2918 268708
rect 2622 267676 2918 267696
rect 2678 267674 2702 267676
rect 2758 267674 2782 267676
rect 2838 267674 2862 267676
rect 2700 267622 2702 267674
rect 2764 267622 2776 267674
rect 2838 267622 2840 267674
rect 2678 267620 2702 267622
rect 2758 267620 2782 267622
rect 2838 267620 2862 267622
rect 2622 267600 2918 267620
rect 2622 266588 2918 266608
rect 2678 266586 2702 266588
rect 2758 266586 2782 266588
rect 2838 266586 2862 266588
rect 2700 266534 2702 266586
rect 2764 266534 2776 266586
rect 2838 266534 2840 266586
rect 2678 266532 2702 266534
rect 2758 266532 2782 266534
rect 2838 266532 2862 266534
rect 2622 266512 2918 266532
rect 2622 265500 2918 265520
rect 2678 265498 2702 265500
rect 2758 265498 2782 265500
rect 2838 265498 2862 265500
rect 2700 265446 2702 265498
rect 2764 265446 2776 265498
rect 2838 265446 2840 265498
rect 2678 265444 2702 265446
rect 2758 265444 2782 265446
rect 2838 265444 2862 265446
rect 2622 265424 2918 265444
rect 2622 264412 2918 264432
rect 2678 264410 2702 264412
rect 2758 264410 2782 264412
rect 2838 264410 2862 264412
rect 2700 264358 2702 264410
rect 2764 264358 2776 264410
rect 2838 264358 2840 264410
rect 2678 264356 2702 264358
rect 2758 264356 2782 264358
rect 2838 264356 2862 264358
rect 2622 264336 2918 264356
rect 2622 263324 2918 263344
rect 2678 263322 2702 263324
rect 2758 263322 2782 263324
rect 2838 263322 2862 263324
rect 2700 263270 2702 263322
rect 2764 263270 2776 263322
rect 2838 263270 2840 263322
rect 2678 263268 2702 263270
rect 2758 263268 2782 263270
rect 2838 263268 2862 263270
rect 2622 263248 2918 263268
rect 2622 262236 2918 262256
rect 2678 262234 2702 262236
rect 2758 262234 2782 262236
rect 2838 262234 2862 262236
rect 2700 262182 2702 262234
rect 2764 262182 2776 262234
rect 2838 262182 2840 262234
rect 2678 262180 2702 262182
rect 2758 262180 2782 262182
rect 2838 262180 2862 262182
rect 2622 262160 2918 262180
rect 2502 261352 2558 261361
rect 2502 261287 2558 261296
rect 2228 244724 2280 244730
rect 2228 244666 2280 244672
rect 2516 237522 2544 261287
rect 2622 261148 2918 261168
rect 2678 261146 2702 261148
rect 2758 261146 2782 261148
rect 2838 261146 2862 261148
rect 2700 261094 2702 261146
rect 2764 261094 2776 261146
rect 2838 261094 2840 261146
rect 2678 261092 2702 261094
rect 2758 261092 2782 261094
rect 2838 261092 2862 261094
rect 2622 261072 2918 261092
rect 2622 260060 2918 260080
rect 2678 260058 2702 260060
rect 2758 260058 2782 260060
rect 2838 260058 2862 260060
rect 2700 260006 2702 260058
rect 2764 260006 2776 260058
rect 2838 260006 2840 260058
rect 2678 260004 2702 260006
rect 2758 260004 2782 260006
rect 2838 260004 2862 260006
rect 2622 259984 2918 260004
rect 2622 258972 2918 258992
rect 2678 258970 2702 258972
rect 2758 258970 2782 258972
rect 2838 258970 2862 258972
rect 2700 258918 2702 258970
rect 2764 258918 2776 258970
rect 2838 258918 2840 258970
rect 2678 258916 2702 258918
rect 2758 258916 2782 258918
rect 2838 258916 2862 258918
rect 2622 258896 2918 258916
rect 2622 257884 2918 257904
rect 2678 257882 2702 257884
rect 2758 257882 2782 257884
rect 2838 257882 2862 257884
rect 2700 257830 2702 257882
rect 2764 257830 2776 257882
rect 2838 257830 2840 257882
rect 2678 257828 2702 257830
rect 2758 257828 2782 257830
rect 2838 257828 2862 257830
rect 2622 257808 2918 257828
rect 2622 256796 2918 256816
rect 2678 256794 2702 256796
rect 2758 256794 2782 256796
rect 2838 256794 2862 256796
rect 2700 256742 2702 256794
rect 2764 256742 2776 256794
rect 2838 256742 2840 256794
rect 2678 256740 2702 256742
rect 2758 256740 2782 256742
rect 2838 256740 2862 256742
rect 2622 256720 2918 256740
rect 2622 255708 2918 255728
rect 2678 255706 2702 255708
rect 2758 255706 2782 255708
rect 2838 255706 2862 255708
rect 2700 255654 2702 255706
rect 2764 255654 2776 255706
rect 2838 255654 2840 255706
rect 2678 255652 2702 255654
rect 2758 255652 2782 255654
rect 2838 255652 2862 255654
rect 2622 255632 2918 255652
rect 2622 254620 2918 254640
rect 2678 254618 2702 254620
rect 2758 254618 2782 254620
rect 2838 254618 2862 254620
rect 2700 254566 2702 254618
rect 2764 254566 2776 254618
rect 2838 254566 2840 254618
rect 2678 254564 2702 254566
rect 2758 254564 2782 254566
rect 2838 254564 2862 254566
rect 2622 254544 2918 254564
rect 2622 253532 2918 253552
rect 2678 253530 2702 253532
rect 2758 253530 2782 253532
rect 2838 253530 2862 253532
rect 2700 253478 2702 253530
rect 2764 253478 2776 253530
rect 2838 253478 2840 253530
rect 2678 253476 2702 253478
rect 2758 253476 2782 253478
rect 2838 253476 2862 253478
rect 2622 253456 2918 253476
rect 2622 252444 2918 252464
rect 2678 252442 2702 252444
rect 2758 252442 2782 252444
rect 2838 252442 2862 252444
rect 2700 252390 2702 252442
rect 2764 252390 2776 252442
rect 2838 252390 2840 252442
rect 2678 252388 2702 252390
rect 2758 252388 2782 252390
rect 2838 252388 2862 252390
rect 2622 252368 2918 252388
rect 2622 251356 2918 251376
rect 2678 251354 2702 251356
rect 2758 251354 2782 251356
rect 2838 251354 2862 251356
rect 2700 251302 2702 251354
rect 2764 251302 2776 251354
rect 2838 251302 2840 251354
rect 2678 251300 2702 251302
rect 2758 251300 2782 251302
rect 2838 251300 2862 251302
rect 2622 251280 2918 251300
rect 2622 250268 2918 250288
rect 2678 250266 2702 250268
rect 2758 250266 2782 250268
rect 2838 250266 2862 250268
rect 2700 250214 2702 250266
rect 2764 250214 2776 250266
rect 2838 250214 2840 250266
rect 2678 250212 2702 250214
rect 2758 250212 2782 250214
rect 2838 250212 2862 250214
rect 2622 250192 2918 250212
rect 2622 249180 2918 249200
rect 2678 249178 2702 249180
rect 2758 249178 2782 249180
rect 2838 249178 2862 249180
rect 2700 249126 2702 249178
rect 2764 249126 2776 249178
rect 2838 249126 2840 249178
rect 2678 249124 2702 249126
rect 2758 249124 2782 249126
rect 2838 249124 2862 249126
rect 2622 249104 2918 249124
rect 2622 248092 2918 248112
rect 2678 248090 2702 248092
rect 2758 248090 2782 248092
rect 2838 248090 2862 248092
rect 2700 248038 2702 248090
rect 2764 248038 2776 248090
rect 2838 248038 2840 248090
rect 2678 248036 2702 248038
rect 2758 248036 2782 248038
rect 2838 248036 2862 248038
rect 2622 248016 2918 248036
rect 2622 247004 2918 247024
rect 2678 247002 2702 247004
rect 2758 247002 2782 247004
rect 2838 247002 2862 247004
rect 2700 246950 2702 247002
rect 2764 246950 2776 247002
rect 2838 246950 2840 247002
rect 2678 246948 2702 246950
rect 2758 246948 2782 246950
rect 2838 246948 2862 246950
rect 2622 246928 2918 246948
rect 2622 245916 2918 245936
rect 2678 245914 2702 245916
rect 2758 245914 2782 245916
rect 2838 245914 2862 245916
rect 2700 245862 2702 245914
rect 2764 245862 2776 245914
rect 2838 245862 2840 245914
rect 2678 245860 2702 245862
rect 2758 245860 2782 245862
rect 2838 245860 2862 245862
rect 2622 245840 2918 245860
rect 2622 244828 2918 244848
rect 2678 244826 2702 244828
rect 2758 244826 2782 244828
rect 2838 244826 2862 244828
rect 2700 244774 2702 244826
rect 2764 244774 2776 244826
rect 2838 244774 2840 244826
rect 2678 244772 2702 244774
rect 2758 244772 2782 244774
rect 2838 244772 2862 244774
rect 2622 244752 2918 244772
rect 3516 244384 3568 244390
rect 3516 244326 3568 244332
rect 2622 243740 2918 243760
rect 2678 243738 2702 243740
rect 2758 243738 2782 243740
rect 2838 243738 2862 243740
rect 2700 243686 2702 243738
rect 2764 243686 2776 243738
rect 2838 243686 2840 243738
rect 2678 243684 2702 243686
rect 2758 243684 2782 243686
rect 2838 243684 2862 243686
rect 2622 243664 2918 243684
rect 2622 242652 2918 242672
rect 2678 242650 2702 242652
rect 2758 242650 2782 242652
rect 2838 242650 2862 242652
rect 2700 242598 2702 242650
rect 2764 242598 2776 242650
rect 2838 242598 2840 242650
rect 2678 242596 2702 242598
rect 2758 242596 2782 242598
rect 2838 242596 2862 242598
rect 2622 242576 2918 242596
rect 2622 241564 2918 241584
rect 2678 241562 2702 241564
rect 2758 241562 2782 241564
rect 2838 241562 2862 241564
rect 2700 241510 2702 241562
rect 2764 241510 2776 241562
rect 2838 241510 2840 241562
rect 2678 241508 2702 241510
rect 2758 241508 2782 241510
rect 2838 241508 2862 241510
rect 2622 241488 2918 241508
rect 2622 240476 2918 240496
rect 2678 240474 2702 240476
rect 2758 240474 2782 240476
rect 2838 240474 2862 240476
rect 2700 240422 2702 240474
rect 2764 240422 2776 240474
rect 2838 240422 2840 240474
rect 2678 240420 2702 240422
rect 2758 240420 2782 240422
rect 2838 240420 2862 240422
rect 2622 240400 2918 240420
rect 2622 239388 2918 239408
rect 2678 239386 2702 239388
rect 2758 239386 2782 239388
rect 2838 239386 2862 239388
rect 2700 239334 2702 239386
rect 2764 239334 2776 239386
rect 2838 239334 2840 239386
rect 2678 239332 2702 239334
rect 2758 239332 2782 239334
rect 2838 239332 2862 239334
rect 2622 239312 2918 239332
rect 2622 238300 2918 238320
rect 2678 238298 2702 238300
rect 2758 238298 2782 238300
rect 2838 238298 2862 238300
rect 2700 238246 2702 238298
rect 2764 238246 2776 238298
rect 2838 238246 2840 238298
rect 2678 238244 2702 238246
rect 2758 238244 2782 238246
rect 2838 238244 2862 238246
rect 2622 238224 2918 238244
rect 2504 237516 2556 237522
rect 2504 237458 2556 237464
rect 2516 237114 2544 237458
rect 2964 237448 3016 237454
rect 2964 237390 3016 237396
rect 2622 237212 2918 237232
rect 2678 237210 2702 237212
rect 2758 237210 2782 237212
rect 2838 237210 2862 237212
rect 2700 237158 2702 237210
rect 2764 237158 2776 237210
rect 2838 237158 2840 237210
rect 2678 237156 2702 237158
rect 2758 237156 2782 237158
rect 2838 237156 2862 237158
rect 2622 237136 2918 237156
rect 2504 237108 2556 237114
rect 2504 237050 2556 237056
rect 2976 236774 3004 237390
rect 3528 237318 3556 244326
rect 3516 237312 3568 237318
rect 3516 237254 3568 237260
rect 2964 236768 3016 236774
rect 2964 236710 3016 236716
rect 2622 236124 2918 236144
rect 2678 236122 2702 236124
rect 2758 236122 2782 236124
rect 2838 236122 2862 236124
rect 2700 236070 2702 236122
rect 2764 236070 2776 236122
rect 2838 236070 2840 236122
rect 2678 236068 2702 236070
rect 2758 236068 2782 236070
rect 2838 236068 2862 236070
rect 2622 236048 2918 236068
rect 2622 235036 2918 235056
rect 2678 235034 2702 235036
rect 2758 235034 2782 235036
rect 2838 235034 2862 235036
rect 2700 234982 2702 235034
rect 2764 234982 2776 235034
rect 2838 234982 2840 235034
rect 2678 234980 2702 234982
rect 2758 234980 2782 234982
rect 2838 234980 2862 234982
rect 2622 234960 2918 234980
rect 2622 233948 2918 233968
rect 2678 233946 2702 233948
rect 2758 233946 2782 233948
rect 2838 233946 2862 233948
rect 2700 233894 2702 233946
rect 2764 233894 2776 233946
rect 2838 233894 2840 233946
rect 2678 233892 2702 233894
rect 2758 233892 2782 233894
rect 2838 233892 2862 233894
rect 2622 233872 2918 233892
rect 2622 232860 2918 232880
rect 2678 232858 2702 232860
rect 2758 232858 2782 232860
rect 2838 232858 2862 232860
rect 2700 232806 2702 232858
rect 2764 232806 2776 232858
rect 2838 232806 2840 232858
rect 2678 232804 2702 232806
rect 2758 232804 2782 232806
rect 2838 232804 2862 232806
rect 2622 232784 2918 232804
rect 2964 232552 3016 232558
rect 2964 232494 3016 232500
rect 2976 231878 3004 232494
rect 2964 231872 3016 231878
rect 2964 231814 3016 231820
rect 2622 231772 2918 231792
rect 2678 231770 2702 231772
rect 2758 231770 2782 231772
rect 2838 231770 2862 231772
rect 2700 231718 2702 231770
rect 2764 231718 2776 231770
rect 2838 231718 2840 231770
rect 2678 231716 2702 231718
rect 2758 231716 2782 231718
rect 2838 231716 2862 231718
rect 2622 231696 2918 231716
rect 2622 230684 2918 230704
rect 2678 230682 2702 230684
rect 2758 230682 2782 230684
rect 2838 230682 2862 230684
rect 2700 230630 2702 230682
rect 2764 230630 2776 230682
rect 2838 230630 2840 230682
rect 2678 230628 2702 230630
rect 2758 230628 2782 230630
rect 2838 230628 2862 230630
rect 2622 230608 2918 230628
rect 2412 230240 2464 230246
rect 2412 230182 2464 230188
rect 1492 229968 1544 229974
rect 1492 229910 1544 229916
rect 1504 228818 1532 229910
rect 2424 229362 2452 230182
rect 2504 229696 2556 229702
rect 2504 229638 2556 229644
rect 2412 229356 2464 229362
rect 2412 229298 2464 229304
rect 2412 229152 2464 229158
rect 2412 229094 2464 229100
rect 1492 228812 1544 228818
rect 1492 228754 1544 228760
rect 1504 228410 1532 228754
rect 2424 228750 2452 229094
rect 2516 228886 2544 229638
rect 2622 229596 2918 229616
rect 2678 229594 2702 229596
rect 2758 229594 2782 229596
rect 2838 229594 2862 229596
rect 2700 229542 2702 229594
rect 2764 229542 2776 229594
rect 2838 229542 2840 229594
rect 2678 229540 2702 229542
rect 2758 229540 2782 229542
rect 2838 229540 2862 229542
rect 2622 229520 2918 229540
rect 2504 228880 2556 228886
rect 2504 228822 2556 228828
rect 1768 228744 1820 228750
rect 1768 228686 1820 228692
rect 2412 228744 2464 228750
rect 2412 228686 2464 228692
rect 1492 228404 1544 228410
rect 1492 228346 1544 228352
rect 1216 228336 1268 228342
rect 1216 228278 1268 228284
rect 1780 228070 1808 228686
rect 2412 228608 2464 228614
rect 2516 228596 2544 228822
rect 2464 228568 2544 228596
rect 2412 228550 2464 228556
rect 2044 228404 2096 228410
rect 2044 228346 2096 228352
rect 1768 228064 1820 228070
rect 1768 228006 1820 228012
rect 1780 224602 1808 228006
rect 2056 227730 2084 228346
rect 2320 228064 2372 228070
rect 2320 228006 2372 228012
rect 2044 227724 2096 227730
rect 2044 227666 2096 227672
rect 2056 227322 2084 227666
rect 2332 227322 2360 228006
rect 2044 227316 2096 227322
rect 2044 227258 2096 227264
rect 2320 227316 2372 227322
rect 2320 227258 2372 227264
rect 2332 227186 2360 227258
rect 2320 227180 2372 227186
rect 2320 227122 2372 227128
rect 2332 226642 2360 227122
rect 2424 226710 2452 228550
rect 2622 228508 2918 228528
rect 2678 228506 2702 228508
rect 2758 228506 2782 228508
rect 2838 228506 2862 228508
rect 2700 228454 2702 228506
rect 2764 228454 2776 228506
rect 2838 228454 2840 228506
rect 2678 228452 2702 228454
rect 2758 228452 2782 228454
rect 2838 228452 2862 228454
rect 2622 228432 2918 228452
rect 2976 228274 3004 231814
rect 3424 230376 3476 230382
rect 3424 230318 3476 230324
rect 3436 230042 3464 230318
rect 3424 230036 3476 230042
rect 3424 229978 3476 229984
rect 3056 229764 3108 229770
rect 3056 229706 3108 229712
rect 3068 228954 3096 229706
rect 3436 229498 3464 229978
rect 3424 229492 3476 229498
rect 3424 229434 3476 229440
rect 3436 229294 3464 229434
rect 3424 229288 3476 229294
rect 3424 229230 3476 229236
rect 3436 228954 3464 229230
rect 3056 228948 3108 228954
rect 3056 228890 3108 228896
rect 3424 228948 3476 228954
rect 3424 228890 3476 228896
rect 2964 228268 3016 228274
rect 2964 228210 3016 228216
rect 3068 228206 3096 228890
rect 3148 228744 3200 228750
rect 3148 228686 3200 228692
rect 3056 228200 3108 228206
rect 3056 228142 3108 228148
rect 2964 228132 3016 228138
rect 2964 228074 3016 228080
rect 2976 227866 3004 228074
rect 2964 227860 3016 227866
rect 2964 227802 3016 227808
rect 3068 227526 3096 228142
rect 3056 227520 3108 227526
rect 3056 227462 3108 227468
rect 2622 227420 2918 227440
rect 2678 227418 2702 227420
rect 2758 227418 2782 227420
rect 2838 227418 2862 227420
rect 2700 227366 2702 227418
rect 2764 227366 2776 227418
rect 2838 227366 2840 227418
rect 2678 227364 2702 227366
rect 2758 227364 2782 227366
rect 2838 227364 2862 227366
rect 2622 227344 2918 227364
rect 3056 226976 3108 226982
rect 3056 226918 3108 226924
rect 2412 226704 2464 226710
rect 2412 226646 2464 226652
rect 2320 226636 2372 226642
rect 2320 226578 2372 226584
rect 2332 226234 2360 226578
rect 2622 226332 2918 226352
rect 2678 226330 2702 226332
rect 2758 226330 2782 226332
rect 2838 226330 2862 226332
rect 2700 226278 2702 226330
rect 2764 226278 2776 226330
rect 2838 226278 2840 226330
rect 2678 226276 2702 226278
rect 2758 226276 2782 226278
rect 2838 226276 2862 226278
rect 2622 226256 2918 226276
rect 2320 226228 2372 226234
rect 2320 226170 2372 226176
rect 1768 224596 1820 224602
rect 1768 224538 1820 224544
rect 2332 224058 2360 226170
rect 2622 225244 2918 225264
rect 2678 225242 2702 225244
rect 2758 225242 2782 225244
rect 2838 225242 2862 225244
rect 2700 225190 2702 225242
rect 2764 225190 2776 225242
rect 2838 225190 2840 225242
rect 2678 225188 2702 225190
rect 2758 225188 2782 225190
rect 2838 225188 2862 225190
rect 2622 225168 2918 225188
rect 2504 224596 2556 224602
rect 2504 224538 2556 224544
rect 2320 224052 2372 224058
rect 2320 223994 2372 224000
rect 2516 223854 2544 224538
rect 2622 224156 2918 224176
rect 2678 224154 2702 224156
rect 2758 224154 2782 224156
rect 2838 224154 2862 224156
rect 2700 224102 2702 224154
rect 2764 224102 2776 224154
rect 2838 224102 2840 224154
rect 2678 224100 2702 224102
rect 2758 224100 2782 224102
rect 2838 224100 2862 224102
rect 2622 224080 2918 224100
rect 2964 223916 3016 223922
rect 2964 223858 3016 223864
rect 2504 223848 2556 223854
rect 2504 223790 2556 223796
rect 2516 221882 2544 223790
rect 2622 223068 2918 223088
rect 2678 223066 2702 223068
rect 2758 223066 2782 223068
rect 2838 223066 2862 223068
rect 2700 223014 2702 223066
rect 2764 223014 2776 223066
rect 2838 223014 2840 223066
rect 2678 223012 2702 223014
rect 2758 223012 2782 223014
rect 2838 223012 2862 223014
rect 2622 222992 2918 223012
rect 2622 221980 2918 222000
rect 2678 221978 2702 221980
rect 2758 221978 2782 221980
rect 2838 221978 2862 221980
rect 2700 221926 2702 221978
rect 2764 221926 2776 221978
rect 2838 221926 2840 221978
rect 2678 221924 2702 221926
rect 2758 221924 2782 221926
rect 2838 221924 2862 221926
rect 2622 221904 2918 221924
rect 2976 221882 3004 223858
rect 3068 223786 3096 226918
rect 3160 226234 3188 228686
rect 3240 228336 3292 228342
rect 3240 228278 3292 228284
rect 3252 228070 3280 228278
rect 3240 228064 3292 228070
rect 3240 228006 3292 228012
rect 3252 227118 3280 228006
rect 3436 227866 3464 228890
rect 3424 227860 3476 227866
rect 3424 227802 3476 227808
rect 3332 227520 3384 227526
rect 3332 227462 3384 227468
rect 3240 227112 3292 227118
rect 3240 227054 3292 227060
rect 3148 226228 3200 226234
rect 3148 226170 3200 226176
rect 3240 223848 3292 223854
rect 3240 223790 3292 223796
rect 3056 223780 3108 223786
rect 3056 223722 3108 223728
rect 3148 223712 3200 223718
rect 3148 223654 3200 223660
rect 3056 223508 3108 223514
rect 3056 223450 3108 223456
rect 3068 222426 3096 223450
rect 3056 222420 3108 222426
rect 3056 222362 3108 222368
rect 2504 221876 2556 221882
rect 2504 221818 2556 221824
rect 2964 221876 3016 221882
rect 2964 221818 3016 221824
rect 2516 221678 2544 221818
rect 2504 221672 2556 221678
rect 2504 221614 2556 221620
rect 2976 221610 3004 221818
rect 3068 221746 3096 222362
rect 3056 221740 3108 221746
rect 3056 221682 3108 221688
rect 2964 221604 3016 221610
rect 2964 221546 3016 221552
rect 1400 220992 1452 220998
rect 1400 220934 1452 220940
rect 110 214024 166 214033
rect 110 213959 166 213968
rect 124 212090 152 213959
rect 112 212084 164 212090
rect 112 212026 164 212032
rect 20 209568 72 209574
rect 20 209510 72 209516
rect 32 118833 60 209510
rect 18 118824 74 118833
rect 18 118759 74 118768
rect 112 72072 164 72078
rect 112 72014 164 72020
rect 124 71233 152 72014
rect 110 71224 166 71233
rect 110 71159 166 71168
rect 1412 4154 1440 220934
rect 2622 220892 2918 220912
rect 2678 220890 2702 220892
rect 2758 220890 2782 220892
rect 2838 220890 2862 220892
rect 2700 220838 2702 220890
rect 2764 220838 2776 220890
rect 2838 220838 2840 220890
rect 2678 220836 2702 220838
rect 2758 220836 2782 220838
rect 2838 220836 2862 220838
rect 2622 220816 2918 220836
rect 2622 219804 2918 219824
rect 2678 219802 2702 219804
rect 2758 219802 2782 219804
rect 2838 219802 2862 219804
rect 2700 219750 2702 219802
rect 2764 219750 2776 219802
rect 2838 219750 2840 219802
rect 2678 219748 2702 219750
rect 2758 219748 2782 219750
rect 2838 219748 2862 219750
rect 2622 219728 2918 219748
rect 2622 218716 2918 218736
rect 2678 218714 2702 218716
rect 2758 218714 2782 218716
rect 2838 218714 2862 218716
rect 2700 218662 2702 218714
rect 2764 218662 2776 218714
rect 2838 218662 2840 218714
rect 2678 218660 2702 218662
rect 2758 218660 2782 218662
rect 2838 218660 2862 218662
rect 2622 218640 2918 218660
rect 2622 217628 2918 217648
rect 2678 217626 2702 217628
rect 2758 217626 2782 217628
rect 2838 217626 2862 217628
rect 2700 217574 2702 217626
rect 2764 217574 2776 217626
rect 2838 217574 2840 217626
rect 2678 217572 2702 217574
rect 2758 217572 2782 217574
rect 2838 217572 2862 217574
rect 2622 217552 2918 217572
rect 2622 216540 2918 216560
rect 2678 216538 2702 216540
rect 2758 216538 2782 216540
rect 2838 216538 2862 216540
rect 2700 216486 2702 216538
rect 2764 216486 2776 216538
rect 2838 216486 2840 216538
rect 2678 216484 2702 216486
rect 2758 216484 2782 216486
rect 2838 216484 2862 216486
rect 2622 216464 2918 216484
rect 2622 215452 2918 215472
rect 2678 215450 2702 215452
rect 2758 215450 2782 215452
rect 2838 215450 2862 215452
rect 2700 215398 2702 215450
rect 2764 215398 2776 215450
rect 2838 215398 2840 215450
rect 2678 215396 2702 215398
rect 2758 215396 2782 215398
rect 2838 215396 2862 215398
rect 2622 215376 2918 215396
rect 2622 214364 2918 214384
rect 2678 214362 2702 214364
rect 2758 214362 2782 214364
rect 2838 214362 2862 214364
rect 2700 214310 2702 214362
rect 2764 214310 2776 214362
rect 2838 214310 2840 214362
rect 2678 214308 2702 214310
rect 2758 214308 2782 214310
rect 2838 214308 2862 214310
rect 2622 214288 2918 214308
rect 2622 213276 2918 213296
rect 2678 213274 2702 213276
rect 2758 213274 2782 213276
rect 2838 213274 2862 213276
rect 2700 213222 2702 213274
rect 2764 213222 2776 213274
rect 2838 213222 2840 213274
rect 2678 213220 2702 213222
rect 2758 213220 2782 213222
rect 2838 213220 2862 213222
rect 2622 213200 2918 213220
rect 2622 212188 2918 212208
rect 2678 212186 2702 212188
rect 2758 212186 2782 212188
rect 2838 212186 2862 212188
rect 2700 212134 2702 212186
rect 2764 212134 2776 212186
rect 2838 212134 2840 212186
rect 2678 212132 2702 212134
rect 2758 212132 2782 212134
rect 2838 212132 2862 212134
rect 2622 212112 2918 212132
rect 2622 211100 2918 211120
rect 2678 211098 2702 211100
rect 2758 211098 2782 211100
rect 2838 211098 2862 211100
rect 2700 211046 2702 211098
rect 2764 211046 2776 211098
rect 2838 211046 2840 211098
rect 2678 211044 2702 211046
rect 2758 211044 2782 211046
rect 2838 211044 2862 211046
rect 2622 211024 2918 211044
rect 2622 210012 2918 210032
rect 2678 210010 2702 210012
rect 2758 210010 2782 210012
rect 2838 210010 2862 210012
rect 2700 209958 2702 210010
rect 2764 209958 2776 210010
rect 2838 209958 2840 210010
rect 2678 209956 2702 209958
rect 2758 209956 2782 209958
rect 2838 209956 2862 209958
rect 2622 209936 2918 209956
rect 2964 209704 3016 209710
rect 2964 209646 3016 209652
rect 2976 209030 3004 209646
rect 2964 209024 3016 209030
rect 2964 208966 3016 208972
rect 2622 208924 2918 208944
rect 2678 208922 2702 208924
rect 2758 208922 2782 208924
rect 2838 208922 2862 208924
rect 2700 208870 2702 208922
rect 2764 208870 2776 208922
rect 2838 208870 2840 208922
rect 2678 208868 2702 208870
rect 2758 208868 2782 208870
rect 2838 208868 2862 208870
rect 2622 208848 2918 208868
rect 3160 208690 3188 223654
rect 3252 221814 3280 223790
rect 3240 221808 3292 221814
rect 3240 221750 3292 221756
rect 3344 221610 3372 227462
rect 3436 227118 3464 227802
rect 3424 227112 3476 227118
rect 3424 227054 3476 227060
rect 3436 226778 3464 227054
rect 3424 226772 3476 226778
rect 3424 226714 3476 226720
rect 3436 223854 3464 226714
rect 3424 223848 3476 223854
rect 3424 223790 3476 223796
rect 3436 223514 3464 223790
rect 3424 223508 3476 223514
rect 3424 223450 3476 223456
rect 3332 221604 3384 221610
rect 3332 221546 3384 221552
rect 3344 220998 3372 221546
rect 3332 220992 3384 220998
rect 3332 220934 3384 220940
rect 3332 215008 3384 215014
rect 3332 214950 3384 214956
rect 3148 208684 3200 208690
rect 3148 208626 3200 208632
rect 2964 208548 3016 208554
rect 2964 208490 3016 208496
rect 2622 207836 2918 207856
rect 2678 207834 2702 207836
rect 2758 207834 2782 207836
rect 2838 207834 2862 207836
rect 2700 207782 2702 207834
rect 2764 207782 2776 207834
rect 2838 207782 2840 207834
rect 2678 207780 2702 207782
rect 2758 207780 2782 207782
rect 2838 207780 2862 207782
rect 2622 207760 2918 207780
rect 2622 206748 2918 206768
rect 2678 206746 2702 206748
rect 2758 206746 2782 206748
rect 2838 206746 2862 206748
rect 2700 206694 2702 206746
rect 2764 206694 2776 206746
rect 2838 206694 2840 206746
rect 2678 206692 2702 206694
rect 2758 206692 2782 206694
rect 2838 206692 2862 206694
rect 2622 206672 2918 206692
rect 2622 205660 2918 205680
rect 2678 205658 2702 205660
rect 2758 205658 2782 205660
rect 2838 205658 2862 205660
rect 2700 205606 2702 205658
rect 2764 205606 2776 205658
rect 2838 205606 2840 205658
rect 2678 205604 2702 205606
rect 2758 205604 2782 205606
rect 2838 205604 2862 205606
rect 2622 205584 2918 205604
rect 2622 204572 2918 204592
rect 2678 204570 2702 204572
rect 2758 204570 2782 204572
rect 2838 204570 2862 204572
rect 2700 204518 2702 204570
rect 2764 204518 2776 204570
rect 2838 204518 2840 204570
rect 2678 204516 2702 204518
rect 2758 204516 2782 204518
rect 2838 204516 2862 204518
rect 2622 204496 2918 204516
rect 2622 203484 2918 203504
rect 2678 203482 2702 203484
rect 2758 203482 2782 203484
rect 2838 203482 2862 203484
rect 2700 203430 2702 203482
rect 2764 203430 2776 203482
rect 2838 203430 2840 203482
rect 2678 203428 2702 203430
rect 2758 203428 2782 203430
rect 2838 203428 2862 203430
rect 2622 203408 2918 203428
rect 2622 202396 2918 202416
rect 2678 202394 2702 202396
rect 2758 202394 2782 202396
rect 2838 202394 2862 202396
rect 2700 202342 2702 202394
rect 2764 202342 2776 202394
rect 2838 202342 2840 202394
rect 2678 202340 2702 202342
rect 2758 202340 2782 202342
rect 2838 202340 2862 202342
rect 2622 202320 2918 202340
rect 2622 201308 2918 201328
rect 2678 201306 2702 201308
rect 2758 201306 2782 201308
rect 2838 201306 2862 201308
rect 2700 201254 2702 201306
rect 2764 201254 2776 201306
rect 2838 201254 2840 201306
rect 2678 201252 2702 201254
rect 2758 201252 2782 201254
rect 2838 201252 2862 201254
rect 2622 201232 2918 201252
rect 2622 200220 2918 200240
rect 2678 200218 2702 200220
rect 2758 200218 2782 200220
rect 2838 200218 2862 200220
rect 2700 200166 2702 200218
rect 2764 200166 2776 200218
rect 2838 200166 2840 200218
rect 2678 200164 2702 200166
rect 2758 200164 2782 200166
rect 2838 200164 2862 200166
rect 2622 200144 2918 200164
rect 2622 199132 2918 199152
rect 2678 199130 2702 199132
rect 2758 199130 2782 199132
rect 2838 199130 2862 199132
rect 2700 199078 2702 199130
rect 2764 199078 2776 199130
rect 2838 199078 2840 199130
rect 2678 199076 2702 199078
rect 2758 199076 2782 199078
rect 2838 199076 2862 199078
rect 2622 199056 2918 199076
rect 2622 198044 2918 198064
rect 2678 198042 2702 198044
rect 2758 198042 2782 198044
rect 2838 198042 2862 198044
rect 2700 197990 2702 198042
rect 2764 197990 2776 198042
rect 2838 197990 2840 198042
rect 2678 197988 2702 197990
rect 2758 197988 2782 197990
rect 2838 197988 2862 197990
rect 2622 197968 2918 197988
rect 2622 196956 2918 196976
rect 2678 196954 2702 196956
rect 2758 196954 2782 196956
rect 2838 196954 2862 196956
rect 2700 196902 2702 196954
rect 2764 196902 2776 196954
rect 2838 196902 2840 196954
rect 2678 196900 2702 196902
rect 2758 196900 2782 196902
rect 2838 196900 2862 196902
rect 2622 196880 2918 196900
rect 2622 195868 2918 195888
rect 2678 195866 2702 195868
rect 2758 195866 2782 195868
rect 2838 195866 2862 195868
rect 2700 195814 2702 195866
rect 2764 195814 2776 195866
rect 2838 195814 2840 195866
rect 2678 195812 2702 195814
rect 2758 195812 2782 195814
rect 2838 195812 2862 195814
rect 2622 195792 2918 195812
rect 2622 194780 2918 194800
rect 2678 194778 2702 194780
rect 2758 194778 2782 194780
rect 2838 194778 2862 194780
rect 2700 194726 2702 194778
rect 2764 194726 2776 194778
rect 2838 194726 2840 194778
rect 2678 194724 2702 194726
rect 2758 194724 2782 194726
rect 2838 194724 2862 194726
rect 2622 194704 2918 194724
rect 2622 193692 2918 193712
rect 2678 193690 2702 193692
rect 2758 193690 2782 193692
rect 2838 193690 2862 193692
rect 2700 193638 2702 193690
rect 2764 193638 2776 193690
rect 2838 193638 2840 193690
rect 2678 193636 2702 193638
rect 2758 193636 2782 193638
rect 2838 193636 2862 193638
rect 2622 193616 2918 193636
rect 2622 192604 2918 192624
rect 2678 192602 2702 192604
rect 2758 192602 2782 192604
rect 2838 192602 2862 192604
rect 2700 192550 2702 192602
rect 2764 192550 2776 192602
rect 2838 192550 2840 192602
rect 2678 192548 2702 192550
rect 2758 192548 2782 192550
rect 2838 192548 2862 192550
rect 2622 192528 2918 192548
rect 2622 191516 2918 191536
rect 2678 191514 2702 191516
rect 2758 191514 2782 191516
rect 2838 191514 2862 191516
rect 2700 191462 2702 191514
rect 2764 191462 2776 191514
rect 2838 191462 2840 191514
rect 2678 191460 2702 191462
rect 2758 191460 2782 191462
rect 2838 191460 2862 191462
rect 2622 191440 2918 191460
rect 2622 190428 2918 190448
rect 2678 190426 2702 190428
rect 2758 190426 2782 190428
rect 2838 190426 2862 190428
rect 2700 190374 2702 190426
rect 2764 190374 2776 190426
rect 2838 190374 2840 190426
rect 2678 190372 2702 190374
rect 2758 190372 2782 190374
rect 2838 190372 2862 190374
rect 2622 190352 2918 190372
rect 2622 189340 2918 189360
rect 2678 189338 2702 189340
rect 2758 189338 2782 189340
rect 2838 189338 2862 189340
rect 2700 189286 2702 189338
rect 2764 189286 2776 189338
rect 2838 189286 2840 189338
rect 2678 189284 2702 189286
rect 2758 189284 2782 189286
rect 2838 189284 2862 189286
rect 2622 189264 2918 189284
rect 2622 188252 2918 188272
rect 2678 188250 2702 188252
rect 2758 188250 2782 188252
rect 2838 188250 2862 188252
rect 2700 188198 2702 188250
rect 2764 188198 2776 188250
rect 2838 188198 2840 188250
rect 2678 188196 2702 188198
rect 2758 188196 2782 188198
rect 2838 188196 2862 188198
rect 2622 188176 2918 188196
rect 2622 187164 2918 187184
rect 2678 187162 2702 187164
rect 2758 187162 2782 187164
rect 2838 187162 2862 187164
rect 2700 187110 2702 187162
rect 2764 187110 2776 187162
rect 2838 187110 2840 187162
rect 2678 187108 2702 187110
rect 2758 187108 2782 187110
rect 2838 187108 2862 187110
rect 2622 187088 2918 187108
rect 2622 186076 2918 186096
rect 2678 186074 2702 186076
rect 2758 186074 2782 186076
rect 2838 186074 2862 186076
rect 2700 186022 2702 186074
rect 2764 186022 2776 186074
rect 2838 186022 2840 186074
rect 2678 186020 2702 186022
rect 2758 186020 2782 186022
rect 2838 186020 2862 186022
rect 2622 186000 2918 186020
rect 2622 184988 2918 185008
rect 2678 184986 2702 184988
rect 2758 184986 2782 184988
rect 2838 184986 2862 184988
rect 2700 184934 2702 184986
rect 2764 184934 2776 184986
rect 2838 184934 2840 184986
rect 2678 184932 2702 184934
rect 2758 184932 2782 184934
rect 2838 184932 2862 184934
rect 2622 184912 2918 184932
rect 2622 183900 2918 183920
rect 2678 183898 2702 183900
rect 2758 183898 2782 183900
rect 2838 183898 2862 183900
rect 2700 183846 2702 183898
rect 2764 183846 2776 183898
rect 2838 183846 2840 183898
rect 2678 183844 2702 183846
rect 2758 183844 2782 183846
rect 2838 183844 2862 183846
rect 2622 183824 2918 183844
rect 2622 182812 2918 182832
rect 2678 182810 2702 182812
rect 2758 182810 2782 182812
rect 2838 182810 2862 182812
rect 2700 182758 2702 182810
rect 2764 182758 2776 182810
rect 2838 182758 2840 182810
rect 2678 182756 2702 182758
rect 2758 182756 2782 182758
rect 2838 182756 2862 182758
rect 2622 182736 2918 182756
rect 2622 181724 2918 181744
rect 2678 181722 2702 181724
rect 2758 181722 2782 181724
rect 2838 181722 2862 181724
rect 2700 181670 2702 181722
rect 2764 181670 2776 181722
rect 2838 181670 2840 181722
rect 2678 181668 2702 181670
rect 2758 181668 2782 181670
rect 2838 181668 2862 181670
rect 2622 181648 2918 181668
rect 2622 180636 2918 180656
rect 2678 180634 2702 180636
rect 2758 180634 2782 180636
rect 2838 180634 2862 180636
rect 2700 180582 2702 180634
rect 2764 180582 2776 180634
rect 2838 180582 2840 180634
rect 2678 180580 2702 180582
rect 2758 180580 2782 180582
rect 2838 180580 2862 180582
rect 2622 180560 2918 180580
rect 2622 179548 2918 179568
rect 2678 179546 2702 179548
rect 2758 179546 2782 179548
rect 2838 179546 2862 179548
rect 2700 179494 2702 179546
rect 2764 179494 2776 179546
rect 2838 179494 2840 179546
rect 2678 179492 2702 179494
rect 2758 179492 2782 179494
rect 2838 179492 2862 179494
rect 2622 179472 2918 179492
rect 2622 178460 2918 178480
rect 2678 178458 2702 178460
rect 2758 178458 2782 178460
rect 2838 178458 2862 178460
rect 2700 178406 2702 178458
rect 2764 178406 2776 178458
rect 2838 178406 2840 178458
rect 2678 178404 2702 178406
rect 2758 178404 2782 178406
rect 2838 178404 2862 178406
rect 2622 178384 2918 178404
rect 2622 177372 2918 177392
rect 2678 177370 2702 177372
rect 2758 177370 2782 177372
rect 2838 177370 2862 177372
rect 2700 177318 2702 177370
rect 2764 177318 2776 177370
rect 2838 177318 2840 177370
rect 2678 177316 2702 177318
rect 2758 177316 2782 177318
rect 2838 177316 2862 177318
rect 2622 177296 2918 177316
rect 2622 176284 2918 176304
rect 2678 176282 2702 176284
rect 2758 176282 2782 176284
rect 2838 176282 2862 176284
rect 2700 176230 2702 176282
rect 2764 176230 2776 176282
rect 2838 176230 2840 176282
rect 2678 176228 2702 176230
rect 2758 176228 2782 176230
rect 2838 176228 2862 176230
rect 2622 176208 2918 176228
rect 2622 175196 2918 175216
rect 2678 175194 2702 175196
rect 2758 175194 2782 175196
rect 2838 175194 2862 175196
rect 2700 175142 2702 175194
rect 2764 175142 2776 175194
rect 2838 175142 2840 175194
rect 2678 175140 2702 175142
rect 2758 175140 2782 175142
rect 2838 175140 2862 175142
rect 2622 175120 2918 175140
rect 2622 174108 2918 174128
rect 2678 174106 2702 174108
rect 2758 174106 2782 174108
rect 2838 174106 2862 174108
rect 2700 174054 2702 174106
rect 2764 174054 2776 174106
rect 2838 174054 2840 174106
rect 2678 174052 2702 174054
rect 2758 174052 2782 174054
rect 2838 174052 2862 174054
rect 2622 174032 2918 174052
rect 2622 173020 2918 173040
rect 2678 173018 2702 173020
rect 2758 173018 2782 173020
rect 2838 173018 2862 173020
rect 2700 172966 2702 173018
rect 2764 172966 2776 173018
rect 2838 172966 2840 173018
rect 2678 172964 2702 172966
rect 2758 172964 2782 172966
rect 2838 172964 2862 172966
rect 2622 172944 2918 172964
rect 2622 171932 2918 171952
rect 2678 171930 2702 171932
rect 2758 171930 2782 171932
rect 2838 171930 2862 171932
rect 2700 171878 2702 171930
rect 2764 171878 2776 171930
rect 2838 171878 2840 171930
rect 2678 171876 2702 171878
rect 2758 171876 2782 171878
rect 2838 171876 2862 171878
rect 2622 171856 2918 171876
rect 2622 170844 2918 170864
rect 2678 170842 2702 170844
rect 2758 170842 2782 170844
rect 2838 170842 2862 170844
rect 2700 170790 2702 170842
rect 2764 170790 2776 170842
rect 2838 170790 2840 170842
rect 2678 170788 2702 170790
rect 2758 170788 2782 170790
rect 2838 170788 2862 170790
rect 2622 170768 2918 170788
rect 2622 169756 2918 169776
rect 2678 169754 2702 169756
rect 2758 169754 2782 169756
rect 2838 169754 2862 169756
rect 2700 169702 2702 169754
rect 2764 169702 2776 169754
rect 2838 169702 2840 169754
rect 2678 169700 2702 169702
rect 2758 169700 2782 169702
rect 2838 169700 2862 169702
rect 2622 169680 2918 169700
rect 2622 168668 2918 168688
rect 2678 168666 2702 168668
rect 2758 168666 2782 168668
rect 2838 168666 2862 168668
rect 2700 168614 2702 168666
rect 2764 168614 2776 168666
rect 2838 168614 2840 168666
rect 2678 168612 2702 168614
rect 2758 168612 2782 168614
rect 2838 168612 2862 168614
rect 2622 168592 2918 168612
rect 2622 167580 2918 167600
rect 2678 167578 2702 167580
rect 2758 167578 2782 167580
rect 2838 167578 2862 167580
rect 2700 167526 2702 167578
rect 2764 167526 2776 167578
rect 2838 167526 2840 167578
rect 2678 167524 2702 167526
rect 2758 167524 2782 167526
rect 2838 167524 2862 167526
rect 2622 167504 2918 167524
rect 2622 166492 2918 166512
rect 2678 166490 2702 166492
rect 2758 166490 2782 166492
rect 2838 166490 2862 166492
rect 2700 166438 2702 166490
rect 2764 166438 2776 166490
rect 2838 166438 2840 166490
rect 2678 166436 2702 166438
rect 2758 166436 2782 166438
rect 2838 166436 2862 166438
rect 2622 166416 2918 166436
rect 2622 165404 2918 165424
rect 2678 165402 2702 165404
rect 2758 165402 2782 165404
rect 2838 165402 2862 165404
rect 2700 165350 2702 165402
rect 2764 165350 2776 165402
rect 2838 165350 2840 165402
rect 2678 165348 2702 165350
rect 2758 165348 2782 165350
rect 2838 165348 2862 165350
rect 2622 165328 2918 165348
rect 2622 164316 2918 164336
rect 2678 164314 2702 164316
rect 2758 164314 2782 164316
rect 2838 164314 2862 164316
rect 2700 164262 2702 164314
rect 2764 164262 2776 164314
rect 2838 164262 2840 164314
rect 2678 164260 2702 164262
rect 2758 164260 2782 164262
rect 2838 164260 2862 164262
rect 2622 164240 2918 164260
rect 2622 163228 2918 163248
rect 2678 163226 2702 163228
rect 2758 163226 2782 163228
rect 2838 163226 2862 163228
rect 2700 163174 2702 163226
rect 2764 163174 2776 163226
rect 2838 163174 2840 163226
rect 2678 163172 2702 163174
rect 2758 163172 2782 163174
rect 2838 163172 2862 163174
rect 2622 163152 2918 163172
rect 2622 162140 2918 162160
rect 2678 162138 2702 162140
rect 2758 162138 2782 162140
rect 2838 162138 2862 162140
rect 2700 162086 2702 162138
rect 2764 162086 2776 162138
rect 2838 162086 2840 162138
rect 2678 162084 2702 162086
rect 2758 162084 2782 162086
rect 2838 162084 2862 162086
rect 2622 162064 2918 162084
rect 2622 161052 2918 161072
rect 2678 161050 2702 161052
rect 2758 161050 2782 161052
rect 2838 161050 2862 161052
rect 2700 160998 2702 161050
rect 2764 160998 2776 161050
rect 2838 160998 2840 161050
rect 2678 160996 2702 160998
rect 2758 160996 2782 160998
rect 2838 160996 2862 160998
rect 2622 160976 2918 160996
rect 2622 159964 2918 159984
rect 2678 159962 2702 159964
rect 2758 159962 2782 159964
rect 2838 159962 2862 159964
rect 2700 159910 2702 159962
rect 2764 159910 2776 159962
rect 2838 159910 2840 159962
rect 2678 159908 2702 159910
rect 2758 159908 2782 159910
rect 2838 159908 2862 159910
rect 2622 159888 2918 159908
rect 2622 158876 2918 158896
rect 2678 158874 2702 158876
rect 2758 158874 2782 158876
rect 2838 158874 2862 158876
rect 2700 158822 2702 158874
rect 2764 158822 2776 158874
rect 2838 158822 2840 158874
rect 2678 158820 2702 158822
rect 2758 158820 2782 158822
rect 2838 158820 2862 158822
rect 2622 158800 2918 158820
rect 2622 157788 2918 157808
rect 2678 157786 2702 157788
rect 2758 157786 2782 157788
rect 2838 157786 2862 157788
rect 2700 157734 2702 157786
rect 2764 157734 2776 157786
rect 2838 157734 2840 157786
rect 2678 157732 2702 157734
rect 2758 157732 2782 157734
rect 2838 157732 2862 157734
rect 2622 157712 2918 157732
rect 2622 156700 2918 156720
rect 2678 156698 2702 156700
rect 2758 156698 2782 156700
rect 2838 156698 2862 156700
rect 2700 156646 2702 156698
rect 2764 156646 2776 156698
rect 2838 156646 2840 156698
rect 2678 156644 2702 156646
rect 2758 156644 2782 156646
rect 2838 156644 2862 156646
rect 2622 156624 2918 156644
rect 2622 155612 2918 155632
rect 2678 155610 2702 155612
rect 2758 155610 2782 155612
rect 2838 155610 2862 155612
rect 2700 155558 2702 155610
rect 2764 155558 2776 155610
rect 2838 155558 2840 155610
rect 2678 155556 2702 155558
rect 2758 155556 2782 155558
rect 2838 155556 2862 155558
rect 2622 155536 2918 155556
rect 2622 154524 2918 154544
rect 2678 154522 2702 154524
rect 2758 154522 2782 154524
rect 2838 154522 2862 154524
rect 2700 154470 2702 154522
rect 2764 154470 2776 154522
rect 2838 154470 2840 154522
rect 2678 154468 2702 154470
rect 2758 154468 2782 154470
rect 2838 154468 2862 154470
rect 2622 154448 2918 154468
rect 2622 153436 2918 153456
rect 2678 153434 2702 153436
rect 2758 153434 2782 153436
rect 2838 153434 2862 153436
rect 2700 153382 2702 153434
rect 2764 153382 2776 153434
rect 2838 153382 2840 153434
rect 2678 153380 2702 153382
rect 2758 153380 2782 153382
rect 2838 153380 2862 153382
rect 2622 153360 2918 153380
rect 2622 152348 2918 152368
rect 2678 152346 2702 152348
rect 2758 152346 2782 152348
rect 2838 152346 2862 152348
rect 2700 152294 2702 152346
rect 2764 152294 2776 152346
rect 2838 152294 2840 152346
rect 2678 152292 2702 152294
rect 2758 152292 2782 152294
rect 2838 152292 2862 152294
rect 2622 152272 2918 152292
rect 2622 151260 2918 151280
rect 2678 151258 2702 151260
rect 2758 151258 2782 151260
rect 2838 151258 2862 151260
rect 2700 151206 2702 151258
rect 2764 151206 2776 151258
rect 2838 151206 2840 151258
rect 2678 151204 2702 151206
rect 2758 151204 2782 151206
rect 2838 151204 2862 151206
rect 2622 151184 2918 151204
rect 2622 150172 2918 150192
rect 2678 150170 2702 150172
rect 2758 150170 2782 150172
rect 2838 150170 2862 150172
rect 2700 150118 2702 150170
rect 2764 150118 2776 150170
rect 2838 150118 2840 150170
rect 2678 150116 2702 150118
rect 2758 150116 2782 150118
rect 2838 150116 2862 150118
rect 2622 150096 2918 150116
rect 2622 149084 2918 149104
rect 2678 149082 2702 149084
rect 2758 149082 2782 149084
rect 2838 149082 2862 149084
rect 2700 149030 2702 149082
rect 2764 149030 2776 149082
rect 2838 149030 2840 149082
rect 2678 149028 2702 149030
rect 2758 149028 2782 149030
rect 2838 149028 2862 149030
rect 2622 149008 2918 149028
rect 2622 147996 2918 148016
rect 2678 147994 2702 147996
rect 2758 147994 2782 147996
rect 2838 147994 2862 147996
rect 2700 147942 2702 147994
rect 2764 147942 2776 147994
rect 2838 147942 2840 147994
rect 2678 147940 2702 147942
rect 2758 147940 2782 147942
rect 2838 147940 2862 147942
rect 2622 147920 2918 147940
rect 2622 146908 2918 146928
rect 2678 146906 2702 146908
rect 2758 146906 2782 146908
rect 2838 146906 2862 146908
rect 2700 146854 2702 146906
rect 2764 146854 2776 146906
rect 2838 146854 2840 146906
rect 2678 146852 2702 146854
rect 2758 146852 2782 146854
rect 2838 146852 2862 146854
rect 2622 146832 2918 146852
rect 2622 145820 2918 145840
rect 2678 145818 2702 145820
rect 2758 145818 2782 145820
rect 2838 145818 2862 145820
rect 2700 145766 2702 145818
rect 2764 145766 2776 145818
rect 2838 145766 2840 145818
rect 2678 145764 2702 145766
rect 2758 145764 2782 145766
rect 2838 145764 2862 145766
rect 2622 145744 2918 145764
rect 2622 144732 2918 144752
rect 2678 144730 2702 144732
rect 2758 144730 2782 144732
rect 2838 144730 2862 144732
rect 2700 144678 2702 144730
rect 2764 144678 2776 144730
rect 2838 144678 2840 144730
rect 2678 144676 2702 144678
rect 2758 144676 2782 144678
rect 2838 144676 2862 144678
rect 2622 144656 2918 144676
rect 2622 143644 2918 143664
rect 2678 143642 2702 143644
rect 2758 143642 2782 143644
rect 2838 143642 2862 143644
rect 2700 143590 2702 143642
rect 2764 143590 2776 143642
rect 2838 143590 2840 143642
rect 2678 143588 2702 143590
rect 2758 143588 2782 143590
rect 2838 143588 2862 143590
rect 2622 143568 2918 143588
rect 2622 142556 2918 142576
rect 2678 142554 2702 142556
rect 2758 142554 2782 142556
rect 2838 142554 2862 142556
rect 2700 142502 2702 142554
rect 2764 142502 2776 142554
rect 2838 142502 2840 142554
rect 2678 142500 2702 142502
rect 2758 142500 2782 142502
rect 2838 142500 2862 142502
rect 2622 142480 2918 142500
rect 2622 141468 2918 141488
rect 2678 141466 2702 141468
rect 2758 141466 2782 141468
rect 2838 141466 2862 141468
rect 2700 141414 2702 141466
rect 2764 141414 2776 141466
rect 2838 141414 2840 141466
rect 2678 141412 2702 141414
rect 2758 141412 2782 141414
rect 2838 141412 2862 141414
rect 2622 141392 2918 141412
rect 2622 140380 2918 140400
rect 2678 140378 2702 140380
rect 2758 140378 2782 140380
rect 2838 140378 2862 140380
rect 2700 140326 2702 140378
rect 2764 140326 2776 140378
rect 2838 140326 2840 140378
rect 2678 140324 2702 140326
rect 2758 140324 2782 140326
rect 2838 140324 2862 140326
rect 2622 140304 2918 140324
rect 2622 139292 2918 139312
rect 2678 139290 2702 139292
rect 2758 139290 2782 139292
rect 2838 139290 2862 139292
rect 2700 139238 2702 139290
rect 2764 139238 2776 139290
rect 2838 139238 2840 139290
rect 2678 139236 2702 139238
rect 2758 139236 2782 139238
rect 2838 139236 2862 139238
rect 2622 139216 2918 139236
rect 2622 138204 2918 138224
rect 2678 138202 2702 138204
rect 2758 138202 2782 138204
rect 2838 138202 2862 138204
rect 2700 138150 2702 138202
rect 2764 138150 2776 138202
rect 2838 138150 2840 138202
rect 2678 138148 2702 138150
rect 2758 138148 2782 138150
rect 2838 138148 2862 138150
rect 2622 138128 2918 138148
rect 2622 137116 2918 137136
rect 2678 137114 2702 137116
rect 2758 137114 2782 137116
rect 2838 137114 2862 137116
rect 2700 137062 2702 137114
rect 2764 137062 2776 137114
rect 2838 137062 2840 137114
rect 2678 137060 2702 137062
rect 2758 137060 2782 137062
rect 2838 137060 2862 137062
rect 2622 137040 2918 137060
rect 2622 136028 2918 136048
rect 2678 136026 2702 136028
rect 2758 136026 2782 136028
rect 2838 136026 2862 136028
rect 2700 135974 2702 136026
rect 2764 135974 2776 136026
rect 2838 135974 2840 136026
rect 2678 135972 2702 135974
rect 2758 135972 2782 135974
rect 2838 135972 2862 135974
rect 2622 135952 2918 135972
rect 2622 134940 2918 134960
rect 2678 134938 2702 134940
rect 2758 134938 2782 134940
rect 2838 134938 2862 134940
rect 2700 134886 2702 134938
rect 2764 134886 2776 134938
rect 2838 134886 2840 134938
rect 2678 134884 2702 134886
rect 2758 134884 2782 134886
rect 2838 134884 2862 134886
rect 2622 134864 2918 134884
rect 2622 133852 2918 133872
rect 2678 133850 2702 133852
rect 2758 133850 2782 133852
rect 2838 133850 2862 133852
rect 2700 133798 2702 133850
rect 2764 133798 2776 133850
rect 2838 133798 2840 133850
rect 2678 133796 2702 133798
rect 2758 133796 2782 133798
rect 2838 133796 2862 133798
rect 2622 133776 2918 133796
rect 2622 132764 2918 132784
rect 2678 132762 2702 132764
rect 2758 132762 2782 132764
rect 2838 132762 2862 132764
rect 2700 132710 2702 132762
rect 2764 132710 2776 132762
rect 2838 132710 2840 132762
rect 2678 132708 2702 132710
rect 2758 132708 2782 132710
rect 2838 132708 2862 132710
rect 2622 132688 2918 132708
rect 2622 131676 2918 131696
rect 2678 131674 2702 131676
rect 2758 131674 2782 131676
rect 2838 131674 2862 131676
rect 2700 131622 2702 131674
rect 2764 131622 2776 131674
rect 2838 131622 2840 131674
rect 2678 131620 2702 131622
rect 2758 131620 2782 131622
rect 2838 131620 2862 131622
rect 2622 131600 2918 131620
rect 2622 130588 2918 130608
rect 2678 130586 2702 130588
rect 2758 130586 2782 130588
rect 2838 130586 2862 130588
rect 2700 130534 2702 130586
rect 2764 130534 2776 130586
rect 2838 130534 2840 130586
rect 2678 130532 2702 130534
rect 2758 130532 2782 130534
rect 2838 130532 2862 130534
rect 2622 130512 2918 130532
rect 2622 129500 2918 129520
rect 2678 129498 2702 129500
rect 2758 129498 2782 129500
rect 2838 129498 2862 129500
rect 2700 129446 2702 129498
rect 2764 129446 2776 129498
rect 2838 129446 2840 129498
rect 2678 129444 2702 129446
rect 2758 129444 2782 129446
rect 2838 129444 2862 129446
rect 2622 129424 2918 129444
rect 2622 128412 2918 128432
rect 2678 128410 2702 128412
rect 2758 128410 2782 128412
rect 2838 128410 2862 128412
rect 2700 128358 2702 128410
rect 2764 128358 2776 128410
rect 2838 128358 2840 128410
rect 2678 128356 2702 128358
rect 2758 128356 2782 128358
rect 2838 128356 2862 128358
rect 2622 128336 2918 128356
rect 2622 127324 2918 127344
rect 2678 127322 2702 127324
rect 2758 127322 2782 127324
rect 2838 127322 2862 127324
rect 2700 127270 2702 127322
rect 2764 127270 2776 127322
rect 2838 127270 2840 127322
rect 2678 127268 2702 127270
rect 2758 127268 2782 127270
rect 2838 127268 2862 127270
rect 2622 127248 2918 127268
rect 2622 126236 2918 126256
rect 2678 126234 2702 126236
rect 2758 126234 2782 126236
rect 2838 126234 2862 126236
rect 2700 126182 2702 126234
rect 2764 126182 2776 126234
rect 2838 126182 2840 126234
rect 2678 126180 2702 126182
rect 2758 126180 2782 126182
rect 2838 126180 2862 126182
rect 2622 126160 2918 126180
rect 2622 125148 2918 125168
rect 2678 125146 2702 125148
rect 2758 125146 2782 125148
rect 2838 125146 2862 125148
rect 2700 125094 2702 125146
rect 2764 125094 2776 125146
rect 2838 125094 2840 125146
rect 2678 125092 2702 125094
rect 2758 125092 2782 125094
rect 2838 125092 2862 125094
rect 2622 125072 2918 125092
rect 2622 124060 2918 124080
rect 2678 124058 2702 124060
rect 2758 124058 2782 124060
rect 2838 124058 2862 124060
rect 2700 124006 2702 124058
rect 2764 124006 2776 124058
rect 2838 124006 2840 124058
rect 2678 124004 2702 124006
rect 2758 124004 2782 124006
rect 2838 124004 2862 124006
rect 2622 123984 2918 124004
rect 2622 122972 2918 122992
rect 2678 122970 2702 122972
rect 2758 122970 2782 122972
rect 2838 122970 2862 122972
rect 2700 122918 2702 122970
rect 2764 122918 2776 122970
rect 2838 122918 2840 122970
rect 2678 122916 2702 122918
rect 2758 122916 2782 122918
rect 2838 122916 2862 122918
rect 2622 122896 2918 122916
rect 2622 121884 2918 121904
rect 2678 121882 2702 121884
rect 2758 121882 2782 121884
rect 2838 121882 2862 121884
rect 2700 121830 2702 121882
rect 2764 121830 2776 121882
rect 2838 121830 2840 121882
rect 2678 121828 2702 121830
rect 2758 121828 2782 121830
rect 2838 121828 2862 121830
rect 2622 121808 2918 121828
rect 2622 120796 2918 120816
rect 2678 120794 2702 120796
rect 2758 120794 2782 120796
rect 2838 120794 2862 120796
rect 2700 120742 2702 120794
rect 2764 120742 2776 120794
rect 2838 120742 2840 120794
rect 2678 120740 2702 120742
rect 2758 120740 2782 120742
rect 2838 120740 2862 120742
rect 2622 120720 2918 120740
rect 2622 119708 2918 119728
rect 2678 119706 2702 119708
rect 2758 119706 2782 119708
rect 2838 119706 2862 119708
rect 2700 119654 2702 119706
rect 2764 119654 2776 119706
rect 2838 119654 2840 119706
rect 2678 119652 2702 119654
rect 2758 119652 2782 119654
rect 2838 119652 2862 119654
rect 2622 119632 2918 119652
rect 2622 118620 2918 118640
rect 2678 118618 2702 118620
rect 2758 118618 2782 118620
rect 2838 118618 2862 118620
rect 2700 118566 2702 118618
rect 2764 118566 2776 118618
rect 2838 118566 2840 118618
rect 2678 118564 2702 118566
rect 2758 118564 2782 118566
rect 2838 118564 2862 118566
rect 2622 118544 2918 118564
rect 2622 117532 2918 117552
rect 2678 117530 2702 117532
rect 2758 117530 2782 117532
rect 2838 117530 2862 117532
rect 2700 117478 2702 117530
rect 2764 117478 2776 117530
rect 2838 117478 2840 117530
rect 2678 117476 2702 117478
rect 2758 117476 2782 117478
rect 2838 117476 2862 117478
rect 2622 117456 2918 117476
rect 2622 116444 2918 116464
rect 2678 116442 2702 116444
rect 2758 116442 2782 116444
rect 2838 116442 2862 116444
rect 2700 116390 2702 116442
rect 2764 116390 2776 116442
rect 2838 116390 2840 116442
rect 2678 116388 2702 116390
rect 2758 116388 2782 116390
rect 2838 116388 2862 116390
rect 2622 116368 2918 116388
rect 2622 115356 2918 115376
rect 2678 115354 2702 115356
rect 2758 115354 2782 115356
rect 2838 115354 2862 115356
rect 2700 115302 2702 115354
rect 2764 115302 2776 115354
rect 2838 115302 2840 115354
rect 2678 115300 2702 115302
rect 2758 115300 2782 115302
rect 2838 115300 2862 115302
rect 2622 115280 2918 115300
rect 2622 114268 2918 114288
rect 2678 114266 2702 114268
rect 2758 114266 2782 114268
rect 2838 114266 2862 114268
rect 2700 114214 2702 114266
rect 2764 114214 2776 114266
rect 2838 114214 2840 114266
rect 2678 114212 2702 114214
rect 2758 114212 2782 114214
rect 2838 114212 2862 114214
rect 2622 114192 2918 114212
rect 2622 113180 2918 113200
rect 2678 113178 2702 113180
rect 2758 113178 2782 113180
rect 2838 113178 2862 113180
rect 2700 113126 2702 113178
rect 2764 113126 2776 113178
rect 2838 113126 2840 113178
rect 2678 113124 2702 113126
rect 2758 113124 2782 113126
rect 2838 113124 2862 113126
rect 2622 113104 2918 113124
rect 2622 112092 2918 112112
rect 2678 112090 2702 112092
rect 2758 112090 2782 112092
rect 2838 112090 2862 112092
rect 2700 112038 2702 112090
rect 2764 112038 2776 112090
rect 2838 112038 2840 112090
rect 2678 112036 2702 112038
rect 2758 112036 2782 112038
rect 2838 112036 2862 112038
rect 2622 112016 2918 112036
rect 2622 111004 2918 111024
rect 2678 111002 2702 111004
rect 2758 111002 2782 111004
rect 2838 111002 2862 111004
rect 2700 110950 2702 111002
rect 2764 110950 2776 111002
rect 2838 110950 2840 111002
rect 2678 110948 2702 110950
rect 2758 110948 2782 110950
rect 2838 110948 2862 110950
rect 2622 110928 2918 110948
rect 2622 109916 2918 109936
rect 2678 109914 2702 109916
rect 2758 109914 2782 109916
rect 2838 109914 2862 109916
rect 2700 109862 2702 109914
rect 2764 109862 2776 109914
rect 2838 109862 2840 109914
rect 2678 109860 2702 109862
rect 2758 109860 2782 109862
rect 2838 109860 2862 109862
rect 2622 109840 2918 109860
rect 2622 108828 2918 108848
rect 2678 108826 2702 108828
rect 2758 108826 2782 108828
rect 2838 108826 2862 108828
rect 2700 108774 2702 108826
rect 2764 108774 2776 108826
rect 2838 108774 2840 108826
rect 2678 108772 2702 108774
rect 2758 108772 2782 108774
rect 2838 108772 2862 108774
rect 2622 108752 2918 108772
rect 2622 107740 2918 107760
rect 2678 107738 2702 107740
rect 2758 107738 2782 107740
rect 2838 107738 2862 107740
rect 2700 107686 2702 107738
rect 2764 107686 2776 107738
rect 2838 107686 2840 107738
rect 2678 107684 2702 107686
rect 2758 107684 2782 107686
rect 2838 107684 2862 107686
rect 2622 107664 2918 107684
rect 2622 106652 2918 106672
rect 2678 106650 2702 106652
rect 2758 106650 2782 106652
rect 2838 106650 2862 106652
rect 2700 106598 2702 106650
rect 2764 106598 2776 106650
rect 2838 106598 2840 106650
rect 2678 106596 2702 106598
rect 2758 106596 2782 106598
rect 2838 106596 2862 106598
rect 2622 106576 2918 106596
rect 2622 105564 2918 105584
rect 2678 105562 2702 105564
rect 2758 105562 2782 105564
rect 2838 105562 2862 105564
rect 2700 105510 2702 105562
rect 2764 105510 2776 105562
rect 2838 105510 2840 105562
rect 2678 105508 2702 105510
rect 2758 105508 2782 105510
rect 2838 105508 2862 105510
rect 2622 105488 2918 105508
rect 2622 104476 2918 104496
rect 2678 104474 2702 104476
rect 2758 104474 2782 104476
rect 2838 104474 2862 104476
rect 2700 104422 2702 104474
rect 2764 104422 2776 104474
rect 2838 104422 2840 104474
rect 2678 104420 2702 104422
rect 2758 104420 2782 104422
rect 2838 104420 2862 104422
rect 2622 104400 2918 104420
rect 2622 103388 2918 103408
rect 2678 103386 2702 103388
rect 2758 103386 2782 103388
rect 2838 103386 2862 103388
rect 2700 103334 2702 103386
rect 2764 103334 2776 103386
rect 2838 103334 2840 103386
rect 2678 103332 2702 103334
rect 2758 103332 2782 103334
rect 2838 103332 2862 103334
rect 2622 103312 2918 103332
rect 2622 102300 2918 102320
rect 2678 102298 2702 102300
rect 2758 102298 2782 102300
rect 2838 102298 2862 102300
rect 2700 102246 2702 102298
rect 2764 102246 2776 102298
rect 2838 102246 2840 102298
rect 2678 102244 2702 102246
rect 2758 102244 2782 102246
rect 2838 102244 2862 102246
rect 2622 102224 2918 102244
rect 2622 101212 2918 101232
rect 2678 101210 2702 101212
rect 2758 101210 2782 101212
rect 2838 101210 2862 101212
rect 2700 101158 2702 101210
rect 2764 101158 2776 101210
rect 2838 101158 2840 101210
rect 2678 101156 2702 101158
rect 2758 101156 2782 101158
rect 2838 101156 2862 101158
rect 2622 101136 2918 101156
rect 2622 100124 2918 100144
rect 2678 100122 2702 100124
rect 2758 100122 2782 100124
rect 2838 100122 2862 100124
rect 2700 100070 2702 100122
rect 2764 100070 2776 100122
rect 2838 100070 2840 100122
rect 2678 100068 2702 100070
rect 2758 100068 2782 100070
rect 2838 100068 2862 100070
rect 2622 100048 2918 100068
rect 2622 99036 2918 99056
rect 2678 99034 2702 99036
rect 2758 99034 2782 99036
rect 2838 99034 2862 99036
rect 2700 98982 2702 99034
rect 2764 98982 2776 99034
rect 2838 98982 2840 99034
rect 2678 98980 2702 98982
rect 2758 98980 2782 98982
rect 2838 98980 2862 98982
rect 2622 98960 2918 98980
rect 2622 97948 2918 97968
rect 2678 97946 2702 97948
rect 2758 97946 2782 97948
rect 2838 97946 2862 97948
rect 2700 97894 2702 97946
rect 2764 97894 2776 97946
rect 2838 97894 2840 97946
rect 2678 97892 2702 97894
rect 2758 97892 2782 97894
rect 2838 97892 2862 97894
rect 2622 97872 2918 97892
rect 2622 96860 2918 96880
rect 2678 96858 2702 96860
rect 2758 96858 2782 96860
rect 2838 96858 2862 96860
rect 2700 96806 2702 96858
rect 2764 96806 2776 96858
rect 2838 96806 2840 96858
rect 2678 96804 2702 96806
rect 2758 96804 2782 96806
rect 2838 96804 2862 96806
rect 2622 96784 2918 96804
rect 2622 95772 2918 95792
rect 2678 95770 2702 95772
rect 2758 95770 2782 95772
rect 2838 95770 2862 95772
rect 2700 95718 2702 95770
rect 2764 95718 2776 95770
rect 2838 95718 2840 95770
rect 2678 95716 2702 95718
rect 2758 95716 2782 95718
rect 2838 95716 2862 95718
rect 2622 95696 2918 95716
rect 2622 94684 2918 94704
rect 2678 94682 2702 94684
rect 2758 94682 2782 94684
rect 2838 94682 2862 94684
rect 2700 94630 2702 94682
rect 2764 94630 2776 94682
rect 2838 94630 2840 94682
rect 2678 94628 2702 94630
rect 2758 94628 2782 94630
rect 2838 94628 2862 94630
rect 2622 94608 2918 94628
rect 2622 93596 2918 93616
rect 2678 93594 2702 93596
rect 2758 93594 2782 93596
rect 2838 93594 2862 93596
rect 2700 93542 2702 93594
rect 2764 93542 2776 93594
rect 2838 93542 2840 93594
rect 2678 93540 2702 93542
rect 2758 93540 2782 93542
rect 2838 93540 2862 93542
rect 2622 93520 2918 93540
rect 2622 92508 2918 92528
rect 2678 92506 2702 92508
rect 2758 92506 2782 92508
rect 2838 92506 2862 92508
rect 2700 92454 2702 92506
rect 2764 92454 2776 92506
rect 2838 92454 2840 92506
rect 2678 92452 2702 92454
rect 2758 92452 2782 92454
rect 2838 92452 2862 92454
rect 2622 92432 2918 92452
rect 2622 91420 2918 91440
rect 2678 91418 2702 91420
rect 2758 91418 2782 91420
rect 2838 91418 2862 91420
rect 2700 91366 2702 91418
rect 2764 91366 2776 91418
rect 2838 91366 2840 91418
rect 2678 91364 2702 91366
rect 2758 91364 2782 91366
rect 2838 91364 2862 91366
rect 2622 91344 2918 91364
rect 2622 90332 2918 90352
rect 2678 90330 2702 90332
rect 2758 90330 2782 90332
rect 2838 90330 2862 90332
rect 2700 90278 2702 90330
rect 2764 90278 2776 90330
rect 2838 90278 2840 90330
rect 2678 90276 2702 90278
rect 2758 90276 2782 90278
rect 2838 90276 2862 90278
rect 2622 90256 2918 90276
rect 2622 89244 2918 89264
rect 2678 89242 2702 89244
rect 2758 89242 2782 89244
rect 2838 89242 2862 89244
rect 2700 89190 2702 89242
rect 2764 89190 2776 89242
rect 2838 89190 2840 89242
rect 2678 89188 2702 89190
rect 2758 89188 2782 89190
rect 2838 89188 2862 89190
rect 2622 89168 2918 89188
rect 2622 88156 2918 88176
rect 2678 88154 2702 88156
rect 2758 88154 2782 88156
rect 2838 88154 2862 88156
rect 2700 88102 2702 88154
rect 2764 88102 2776 88154
rect 2838 88102 2840 88154
rect 2678 88100 2702 88102
rect 2758 88100 2782 88102
rect 2838 88100 2862 88102
rect 2622 88080 2918 88100
rect 2622 87068 2918 87088
rect 2678 87066 2702 87068
rect 2758 87066 2782 87068
rect 2838 87066 2862 87068
rect 2700 87014 2702 87066
rect 2764 87014 2776 87066
rect 2838 87014 2840 87066
rect 2678 87012 2702 87014
rect 2758 87012 2782 87014
rect 2838 87012 2862 87014
rect 2622 86992 2918 87012
rect 2622 85980 2918 86000
rect 2678 85978 2702 85980
rect 2758 85978 2782 85980
rect 2838 85978 2862 85980
rect 2700 85926 2702 85978
rect 2764 85926 2776 85978
rect 2838 85926 2840 85978
rect 2678 85924 2702 85926
rect 2758 85924 2782 85926
rect 2838 85924 2862 85926
rect 2622 85904 2918 85924
rect 2622 84892 2918 84912
rect 2678 84890 2702 84892
rect 2758 84890 2782 84892
rect 2838 84890 2862 84892
rect 2700 84838 2702 84890
rect 2764 84838 2776 84890
rect 2838 84838 2840 84890
rect 2678 84836 2702 84838
rect 2758 84836 2782 84838
rect 2838 84836 2862 84838
rect 2622 84816 2918 84836
rect 2622 83804 2918 83824
rect 2678 83802 2702 83804
rect 2758 83802 2782 83804
rect 2838 83802 2862 83804
rect 2700 83750 2702 83802
rect 2764 83750 2776 83802
rect 2838 83750 2840 83802
rect 2678 83748 2702 83750
rect 2758 83748 2782 83750
rect 2838 83748 2862 83750
rect 2622 83728 2918 83748
rect 2622 82716 2918 82736
rect 2678 82714 2702 82716
rect 2758 82714 2782 82716
rect 2838 82714 2862 82716
rect 2700 82662 2702 82714
rect 2764 82662 2776 82714
rect 2838 82662 2840 82714
rect 2678 82660 2702 82662
rect 2758 82660 2782 82662
rect 2838 82660 2862 82662
rect 2622 82640 2918 82660
rect 2622 81628 2918 81648
rect 2678 81626 2702 81628
rect 2758 81626 2782 81628
rect 2838 81626 2862 81628
rect 2700 81574 2702 81626
rect 2764 81574 2776 81626
rect 2838 81574 2840 81626
rect 2678 81572 2702 81574
rect 2758 81572 2782 81574
rect 2838 81572 2862 81574
rect 2622 81552 2918 81572
rect 2622 80540 2918 80560
rect 2678 80538 2702 80540
rect 2758 80538 2782 80540
rect 2838 80538 2862 80540
rect 2700 80486 2702 80538
rect 2764 80486 2776 80538
rect 2838 80486 2840 80538
rect 2678 80484 2702 80486
rect 2758 80484 2782 80486
rect 2838 80484 2862 80486
rect 2622 80464 2918 80484
rect 2622 79452 2918 79472
rect 2678 79450 2702 79452
rect 2758 79450 2782 79452
rect 2838 79450 2862 79452
rect 2700 79398 2702 79450
rect 2764 79398 2776 79450
rect 2838 79398 2840 79450
rect 2678 79396 2702 79398
rect 2758 79396 2782 79398
rect 2838 79396 2862 79398
rect 2622 79376 2918 79396
rect 2622 78364 2918 78384
rect 2678 78362 2702 78364
rect 2758 78362 2782 78364
rect 2838 78362 2862 78364
rect 2700 78310 2702 78362
rect 2764 78310 2776 78362
rect 2838 78310 2840 78362
rect 2678 78308 2702 78310
rect 2758 78308 2782 78310
rect 2838 78308 2862 78310
rect 2622 78288 2918 78308
rect 2622 77276 2918 77296
rect 2678 77274 2702 77276
rect 2758 77274 2782 77276
rect 2838 77274 2862 77276
rect 2700 77222 2702 77274
rect 2764 77222 2776 77274
rect 2838 77222 2840 77274
rect 2678 77220 2702 77222
rect 2758 77220 2782 77222
rect 2838 77220 2862 77222
rect 2622 77200 2918 77220
rect 2622 76188 2918 76208
rect 2678 76186 2702 76188
rect 2758 76186 2782 76188
rect 2838 76186 2862 76188
rect 2700 76134 2702 76186
rect 2764 76134 2776 76186
rect 2838 76134 2840 76186
rect 2678 76132 2702 76134
rect 2758 76132 2782 76134
rect 2838 76132 2862 76134
rect 2622 76112 2918 76132
rect 2622 75100 2918 75120
rect 2678 75098 2702 75100
rect 2758 75098 2782 75100
rect 2838 75098 2862 75100
rect 2700 75046 2702 75098
rect 2764 75046 2776 75098
rect 2838 75046 2840 75098
rect 2678 75044 2702 75046
rect 2758 75044 2782 75046
rect 2838 75044 2862 75046
rect 2622 75024 2918 75044
rect 2622 74012 2918 74032
rect 2678 74010 2702 74012
rect 2758 74010 2782 74012
rect 2838 74010 2862 74012
rect 2700 73958 2702 74010
rect 2764 73958 2776 74010
rect 2838 73958 2840 74010
rect 2678 73956 2702 73958
rect 2758 73956 2782 73958
rect 2838 73956 2862 73958
rect 2622 73936 2918 73956
rect 2622 72924 2918 72944
rect 2678 72922 2702 72924
rect 2758 72922 2782 72924
rect 2838 72922 2862 72924
rect 2700 72870 2702 72922
rect 2764 72870 2776 72922
rect 2838 72870 2840 72922
rect 2678 72868 2702 72870
rect 2758 72868 2782 72870
rect 2838 72868 2862 72870
rect 2622 72848 2918 72868
rect 2622 71836 2918 71856
rect 2678 71834 2702 71836
rect 2758 71834 2782 71836
rect 2838 71834 2862 71836
rect 2700 71782 2702 71834
rect 2764 71782 2776 71834
rect 2838 71782 2840 71834
rect 2678 71780 2702 71782
rect 2758 71780 2782 71782
rect 2838 71780 2862 71782
rect 2622 71760 2918 71780
rect 2622 70748 2918 70768
rect 2678 70746 2702 70748
rect 2758 70746 2782 70748
rect 2838 70746 2862 70748
rect 2700 70694 2702 70746
rect 2764 70694 2776 70746
rect 2838 70694 2840 70746
rect 2678 70692 2702 70694
rect 2758 70692 2782 70694
rect 2838 70692 2862 70694
rect 2622 70672 2918 70692
rect 2622 69660 2918 69680
rect 2678 69658 2702 69660
rect 2758 69658 2782 69660
rect 2838 69658 2862 69660
rect 2700 69606 2702 69658
rect 2764 69606 2776 69658
rect 2838 69606 2840 69658
rect 2678 69604 2702 69606
rect 2758 69604 2782 69606
rect 2838 69604 2862 69606
rect 2622 69584 2918 69604
rect 2622 68572 2918 68592
rect 2678 68570 2702 68572
rect 2758 68570 2782 68572
rect 2838 68570 2862 68572
rect 2700 68518 2702 68570
rect 2764 68518 2776 68570
rect 2838 68518 2840 68570
rect 2678 68516 2702 68518
rect 2758 68516 2782 68518
rect 2838 68516 2862 68518
rect 2622 68496 2918 68516
rect 2622 67484 2918 67504
rect 2678 67482 2702 67484
rect 2758 67482 2782 67484
rect 2838 67482 2862 67484
rect 2700 67430 2702 67482
rect 2764 67430 2776 67482
rect 2838 67430 2840 67482
rect 2678 67428 2702 67430
rect 2758 67428 2782 67430
rect 2838 67428 2862 67430
rect 2622 67408 2918 67428
rect 2622 66396 2918 66416
rect 2678 66394 2702 66396
rect 2758 66394 2782 66396
rect 2838 66394 2862 66396
rect 2700 66342 2702 66394
rect 2764 66342 2776 66394
rect 2838 66342 2840 66394
rect 2678 66340 2702 66342
rect 2758 66340 2782 66342
rect 2838 66340 2862 66342
rect 2622 66320 2918 66340
rect 2622 65308 2918 65328
rect 2678 65306 2702 65308
rect 2758 65306 2782 65308
rect 2838 65306 2862 65308
rect 2700 65254 2702 65306
rect 2764 65254 2776 65306
rect 2838 65254 2840 65306
rect 2678 65252 2702 65254
rect 2758 65252 2782 65254
rect 2838 65252 2862 65254
rect 2622 65232 2918 65252
rect 2622 64220 2918 64240
rect 2678 64218 2702 64220
rect 2758 64218 2782 64220
rect 2838 64218 2862 64220
rect 2700 64166 2702 64218
rect 2764 64166 2776 64218
rect 2838 64166 2840 64218
rect 2678 64164 2702 64166
rect 2758 64164 2782 64166
rect 2838 64164 2862 64166
rect 2622 64144 2918 64164
rect 2622 63132 2918 63152
rect 2678 63130 2702 63132
rect 2758 63130 2782 63132
rect 2838 63130 2862 63132
rect 2700 63078 2702 63130
rect 2764 63078 2776 63130
rect 2838 63078 2840 63130
rect 2678 63076 2702 63078
rect 2758 63076 2782 63078
rect 2838 63076 2862 63078
rect 2622 63056 2918 63076
rect 2622 62044 2918 62064
rect 2678 62042 2702 62044
rect 2758 62042 2782 62044
rect 2838 62042 2862 62044
rect 2700 61990 2702 62042
rect 2764 61990 2776 62042
rect 2838 61990 2840 62042
rect 2678 61988 2702 61990
rect 2758 61988 2782 61990
rect 2838 61988 2862 61990
rect 2622 61968 2918 61988
rect 2622 60956 2918 60976
rect 2678 60954 2702 60956
rect 2758 60954 2782 60956
rect 2838 60954 2862 60956
rect 2700 60902 2702 60954
rect 2764 60902 2776 60954
rect 2838 60902 2840 60954
rect 2678 60900 2702 60902
rect 2758 60900 2782 60902
rect 2838 60900 2862 60902
rect 2622 60880 2918 60900
rect 2622 59868 2918 59888
rect 2678 59866 2702 59868
rect 2758 59866 2782 59868
rect 2838 59866 2862 59868
rect 2700 59814 2702 59866
rect 2764 59814 2776 59866
rect 2838 59814 2840 59866
rect 2678 59812 2702 59814
rect 2758 59812 2782 59814
rect 2838 59812 2862 59814
rect 2622 59792 2918 59812
rect 2622 58780 2918 58800
rect 2678 58778 2702 58780
rect 2758 58778 2782 58780
rect 2838 58778 2862 58780
rect 2700 58726 2702 58778
rect 2764 58726 2776 58778
rect 2838 58726 2840 58778
rect 2678 58724 2702 58726
rect 2758 58724 2782 58726
rect 2838 58724 2862 58726
rect 2622 58704 2918 58724
rect 2622 57692 2918 57712
rect 2678 57690 2702 57692
rect 2758 57690 2782 57692
rect 2838 57690 2862 57692
rect 2700 57638 2702 57690
rect 2764 57638 2776 57690
rect 2838 57638 2840 57690
rect 2678 57636 2702 57638
rect 2758 57636 2782 57638
rect 2838 57636 2862 57638
rect 2622 57616 2918 57636
rect 2622 56604 2918 56624
rect 2678 56602 2702 56604
rect 2758 56602 2782 56604
rect 2838 56602 2862 56604
rect 2700 56550 2702 56602
rect 2764 56550 2776 56602
rect 2838 56550 2840 56602
rect 2678 56548 2702 56550
rect 2758 56548 2782 56550
rect 2838 56548 2862 56550
rect 2622 56528 2918 56548
rect 2622 55516 2918 55536
rect 2678 55514 2702 55516
rect 2758 55514 2782 55516
rect 2838 55514 2862 55516
rect 2700 55462 2702 55514
rect 2764 55462 2776 55514
rect 2838 55462 2840 55514
rect 2678 55460 2702 55462
rect 2758 55460 2782 55462
rect 2838 55460 2862 55462
rect 2622 55440 2918 55460
rect 2622 54428 2918 54448
rect 2678 54426 2702 54428
rect 2758 54426 2782 54428
rect 2838 54426 2862 54428
rect 2700 54374 2702 54426
rect 2764 54374 2776 54426
rect 2838 54374 2840 54426
rect 2678 54372 2702 54374
rect 2758 54372 2782 54374
rect 2838 54372 2862 54374
rect 2622 54352 2918 54372
rect 2622 53340 2918 53360
rect 2678 53338 2702 53340
rect 2758 53338 2782 53340
rect 2838 53338 2862 53340
rect 2700 53286 2702 53338
rect 2764 53286 2776 53338
rect 2838 53286 2840 53338
rect 2678 53284 2702 53286
rect 2758 53284 2782 53286
rect 2838 53284 2862 53286
rect 2622 53264 2918 53284
rect 2622 52252 2918 52272
rect 2678 52250 2702 52252
rect 2758 52250 2782 52252
rect 2838 52250 2862 52252
rect 2700 52198 2702 52250
rect 2764 52198 2776 52250
rect 2838 52198 2840 52250
rect 2678 52196 2702 52198
rect 2758 52196 2782 52198
rect 2838 52196 2862 52198
rect 2622 52176 2918 52196
rect 2622 51164 2918 51184
rect 2678 51162 2702 51164
rect 2758 51162 2782 51164
rect 2838 51162 2862 51164
rect 2700 51110 2702 51162
rect 2764 51110 2776 51162
rect 2838 51110 2840 51162
rect 2678 51108 2702 51110
rect 2758 51108 2782 51110
rect 2838 51108 2862 51110
rect 2622 51088 2918 51108
rect 2622 50076 2918 50096
rect 2678 50074 2702 50076
rect 2758 50074 2782 50076
rect 2838 50074 2862 50076
rect 2700 50022 2702 50074
rect 2764 50022 2776 50074
rect 2838 50022 2840 50074
rect 2678 50020 2702 50022
rect 2758 50020 2782 50022
rect 2838 50020 2862 50022
rect 2622 50000 2918 50020
rect 2622 48988 2918 49008
rect 2678 48986 2702 48988
rect 2758 48986 2782 48988
rect 2838 48986 2862 48988
rect 2700 48934 2702 48986
rect 2764 48934 2776 48986
rect 2838 48934 2840 48986
rect 2678 48932 2702 48934
rect 2758 48932 2782 48934
rect 2838 48932 2862 48934
rect 2622 48912 2918 48932
rect 2622 47900 2918 47920
rect 2678 47898 2702 47900
rect 2758 47898 2782 47900
rect 2838 47898 2862 47900
rect 2700 47846 2702 47898
rect 2764 47846 2776 47898
rect 2838 47846 2840 47898
rect 2678 47844 2702 47846
rect 2758 47844 2782 47846
rect 2838 47844 2862 47846
rect 2622 47824 2918 47844
rect 2622 46812 2918 46832
rect 2678 46810 2702 46812
rect 2758 46810 2782 46812
rect 2838 46810 2862 46812
rect 2700 46758 2702 46810
rect 2764 46758 2776 46810
rect 2838 46758 2840 46810
rect 2678 46756 2702 46758
rect 2758 46756 2782 46758
rect 2838 46756 2862 46758
rect 2622 46736 2918 46756
rect 2622 45724 2918 45744
rect 2678 45722 2702 45724
rect 2758 45722 2782 45724
rect 2838 45722 2862 45724
rect 2700 45670 2702 45722
rect 2764 45670 2776 45722
rect 2838 45670 2840 45722
rect 2678 45668 2702 45670
rect 2758 45668 2782 45670
rect 2838 45668 2862 45670
rect 2622 45648 2918 45668
rect 2622 44636 2918 44656
rect 2678 44634 2702 44636
rect 2758 44634 2782 44636
rect 2838 44634 2862 44636
rect 2700 44582 2702 44634
rect 2764 44582 2776 44634
rect 2838 44582 2840 44634
rect 2678 44580 2702 44582
rect 2758 44580 2782 44582
rect 2838 44580 2862 44582
rect 2622 44560 2918 44580
rect 2622 43548 2918 43568
rect 2678 43546 2702 43548
rect 2758 43546 2782 43548
rect 2838 43546 2862 43548
rect 2700 43494 2702 43546
rect 2764 43494 2776 43546
rect 2838 43494 2840 43546
rect 2678 43492 2702 43494
rect 2758 43492 2782 43494
rect 2838 43492 2862 43494
rect 2622 43472 2918 43492
rect 2622 42460 2918 42480
rect 2678 42458 2702 42460
rect 2758 42458 2782 42460
rect 2838 42458 2862 42460
rect 2700 42406 2702 42458
rect 2764 42406 2776 42458
rect 2838 42406 2840 42458
rect 2678 42404 2702 42406
rect 2758 42404 2782 42406
rect 2838 42404 2862 42406
rect 2622 42384 2918 42404
rect 2622 41372 2918 41392
rect 2678 41370 2702 41372
rect 2758 41370 2782 41372
rect 2838 41370 2862 41372
rect 2700 41318 2702 41370
rect 2764 41318 2776 41370
rect 2838 41318 2840 41370
rect 2678 41316 2702 41318
rect 2758 41316 2782 41318
rect 2838 41316 2862 41318
rect 2622 41296 2918 41316
rect 2622 40284 2918 40304
rect 2678 40282 2702 40284
rect 2758 40282 2782 40284
rect 2838 40282 2862 40284
rect 2700 40230 2702 40282
rect 2764 40230 2776 40282
rect 2838 40230 2840 40282
rect 2678 40228 2702 40230
rect 2758 40228 2782 40230
rect 2838 40228 2862 40230
rect 2622 40208 2918 40228
rect 2622 39196 2918 39216
rect 2678 39194 2702 39196
rect 2758 39194 2782 39196
rect 2838 39194 2862 39196
rect 2700 39142 2702 39194
rect 2764 39142 2776 39194
rect 2838 39142 2840 39194
rect 2678 39140 2702 39142
rect 2758 39140 2782 39142
rect 2838 39140 2862 39142
rect 2622 39120 2918 39140
rect 2622 38108 2918 38128
rect 2678 38106 2702 38108
rect 2758 38106 2782 38108
rect 2838 38106 2862 38108
rect 2700 38054 2702 38106
rect 2764 38054 2776 38106
rect 2838 38054 2840 38106
rect 2678 38052 2702 38054
rect 2758 38052 2782 38054
rect 2838 38052 2862 38054
rect 2622 38032 2918 38052
rect 2622 37020 2918 37040
rect 2678 37018 2702 37020
rect 2758 37018 2782 37020
rect 2838 37018 2862 37020
rect 2700 36966 2702 37018
rect 2764 36966 2776 37018
rect 2838 36966 2840 37018
rect 2678 36964 2702 36966
rect 2758 36964 2782 36966
rect 2838 36964 2862 36966
rect 2622 36944 2918 36964
rect 2622 35932 2918 35952
rect 2678 35930 2702 35932
rect 2758 35930 2782 35932
rect 2838 35930 2862 35932
rect 2700 35878 2702 35930
rect 2764 35878 2776 35930
rect 2838 35878 2840 35930
rect 2678 35876 2702 35878
rect 2758 35876 2782 35878
rect 2838 35876 2862 35878
rect 2622 35856 2918 35876
rect 2622 34844 2918 34864
rect 2678 34842 2702 34844
rect 2758 34842 2782 34844
rect 2838 34842 2862 34844
rect 2700 34790 2702 34842
rect 2764 34790 2776 34842
rect 2838 34790 2840 34842
rect 2678 34788 2702 34790
rect 2758 34788 2782 34790
rect 2838 34788 2862 34790
rect 2622 34768 2918 34788
rect 2622 33756 2918 33776
rect 2678 33754 2702 33756
rect 2758 33754 2782 33756
rect 2838 33754 2862 33756
rect 2700 33702 2702 33754
rect 2764 33702 2776 33754
rect 2838 33702 2840 33754
rect 2678 33700 2702 33702
rect 2758 33700 2782 33702
rect 2838 33700 2862 33702
rect 2622 33680 2918 33700
rect 2622 32668 2918 32688
rect 2678 32666 2702 32668
rect 2758 32666 2782 32668
rect 2838 32666 2862 32668
rect 2700 32614 2702 32666
rect 2764 32614 2776 32666
rect 2838 32614 2840 32666
rect 2678 32612 2702 32614
rect 2758 32612 2782 32614
rect 2838 32612 2862 32614
rect 2622 32592 2918 32612
rect 2622 31580 2918 31600
rect 2678 31578 2702 31580
rect 2758 31578 2782 31580
rect 2838 31578 2862 31580
rect 2700 31526 2702 31578
rect 2764 31526 2776 31578
rect 2838 31526 2840 31578
rect 2678 31524 2702 31526
rect 2758 31524 2782 31526
rect 2838 31524 2862 31526
rect 2622 31504 2918 31524
rect 2622 30492 2918 30512
rect 2678 30490 2702 30492
rect 2758 30490 2782 30492
rect 2838 30490 2862 30492
rect 2700 30438 2702 30490
rect 2764 30438 2776 30490
rect 2838 30438 2840 30490
rect 2678 30436 2702 30438
rect 2758 30436 2782 30438
rect 2838 30436 2862 30438
rect 2622 30416 2918 30436
rect 2622 29404 2918 29424
rect 2678 29402 2702 29404
rect 2758 29402 2782 29404
rect 2838 29402 2862 29404
rect 2700 29350 2702 29402
rect 2764 29350 2776 29402
rect 2838 29350 2840 29402
rect 2678 29348 2702 29350
rect 2758 29348 2782 29350
rect 2838 29348 2862 29350
rect 2622 29328 2918 29348
rect 2622 28316 2918 28336
rect 2678 28314 2702 28316
rect 2758 28314 2782 28316
rect 2838 28314 2862 28316
rect 2700 28262 2702 28314
rect 2764 28262 2776 28314
rect 2838 28262 2840 28314
rect 2678 28260 2702 28262
rect 2758 28260 2782 28262
rect 2838 28260 2862 28262
rect 2622 28240 2918 28260
rect 2622 27228 2918 27248
rect 2678 27226 2702 27228
rect 2758 27226 2782 27228
rect 2838 27226 2862 27228
rect 2700 27174 2702 27226
rect 2764 27174 2776 27226
rect 2838 27174 2840 27226
rect 2678 27172 2702 27174
rect 2758 27172 2782 27174
rect 2838 27172 2862 27174
rect 2622 27152 2918 27172
rect 2622 26140 2918 26160
rect 2678 26138 2702 26140
rect 2758 26138 2782 26140
rect 2838 26138 2862 26140
rect 2700 26086 2702 26138
rect 2764 26086 2776 26138
rect 2838 26086 2840 26138
rect 2678 26084 2702 26086
rect 2758 26084 2782 26086
rect 2838 26084 2862 26086
rect 2622 26064 2918 26084
rect 2622 25052 2918 25072
rect 2678 25050 2702 25052
rect 2758 25050 2782 25052
rect 2838 25050 2862 25052
rect 2700 24998 2702 25050
rect 2764 24998 2776 25050
rect 2838 24998 2840 25050
rect 2678 24996 2702 24998
rect 2758 24996 2782 24998
rect 2838 24996 2862 24998
rect 2622 24976 2918 24996
rect 2622 23964 2918 23984
rect 2678 23962 2702 23964
rect 2758 23962 2782 23964
rect 2838 23962 2862 23964
rect 2700 23910 2702 23962
rect 2764 23910 2776 23962
rect 2838 23910 2840 23962
rect 2678 23908 2702 23910
rect 2758 23908 2782 23910
rect 2838 23908 2862 23910
rect 2622 23888 2918 23908
rect 2622 22876 2918 22896
rect 2678 22874 2702 22876
rect 2758 22874 2782 22876
rect 2838 22874 2862 22876
rect 2700 22822 2702 22874
rect 2764 22822 2776 22874
rect 2838 22822 2840 22874
rect 2678 22820 2702 22822
rect 2758 22820 2782 22822
rect 2838 22820 2862 22822
rect 2622 22800 2918 22820
rect 2622 21788 2918 21808
rect 2678 21786 2702 21788
rect 2758 21786 2782 21788
rect 2838 21786 2862 21788
rect 2700 21734 2702 21786
rect 2764 21734 2776 21786
rect 2838 21734 2840 21786
rect 2678 21732 2702 21734
rect 2758 21732 2782 21734
rect 2838 21732 2862 21734
rect 2622 21712 2918 21732
rect 2622 20700 2918 20720
rect 2678 20698 2702 20700
rect 2758 20698 2782 20700
rect 2838 20698 2862 20700
rect 2700 20646 2702 20698
rect 2764 20646 2776 20698
rect 2838 20646 2840 20698
rect 2678 20644 2702 20646
rect 2758 20644 2782 20646
rect 2838 20644 2862 20646
rect 2622 20624 2918 20644
rect 2622 19612 2918 19632
rect 2678 19610 2702 19612
rect 2758 19610 2782 19612
rect 2838 19610 2862 19612
rect 2700 19558 2702 19610
rect 2764 19558 2776 19610
rect 2838 19558 2840 19610
rect 2678 19556 2702 19558
rect 2758 19556 2782 19558
rect 2838 19556 2862 19558
rect 2622 19536 2918 19556
rect 2622 18524 2918 18544
rect 2678 18522 2702 18524
rect 2758 18522 2782 18524
rect 2838 18522 2862 18524
rect 2700 18470 2702 18522
rect 2764 18470 2776 18522
rect 2838 18470 2840 18522
rect 2678 18468 2702 18470
rect 2758 18468 2782 18470
rect 2838 18468 2862 18470
rect 2622 18448 2918 18468
rect 2622 17436 2918 17456
rect 2678 17434 2702 17436
rect 2758 17434 2782 17436
rect 2838 17434 2862 17436
rect 2700 17382 2702 17434
rect 2764 17382 2776 17434
rect 2838 17382 2840 17434
rect 2678 17380 2702 17382
rect 2758 17380 2782 17382
rect 2838 17380 2862 17382
rect 2622 17360 2918 17380
rect 2622 16348 2918 16368
rect 2678 16346 2702 16348
rect 2758 16346 2782 16348
rect 2838 16346 2862 16348
rect 2700 16294 2702 16346
rect 2764 16294 2776 16346
rect 2838 16294 2840 16346
rect 2678 16292 2702 16294
rect 2758 16292 2782 16294
rect 2838 16292 2862 16294
rect 2622 16272 2918 16292
rect 2622 15260 2918 15280
rect 2678 15258 2702 15260
rect 2758 15258 2782 15260
rect 2838 15258 2862 15260
rect 2700 15206 2702 15258
rect 2764 15206 2776 15258
rect 2838 15206 2840 15258
rect 2678 15204 2702 15206
rect 2758 15204 2782 15206
rect 2838 15204 2862 15206
rect 2622 15184 2918 15204
rect 2622 14172 2918 14192
rect 2678 14170 2702 14172
rect 2758 14170 2782 14172
rect 2838 14170 2862 14172
rect 2700 14118 2702 14170
rect 2764 14118 2776 14170
rect 2838 14118 2840 14170
rect 2678 14116 2702 14118
rect 2758 14116 2782 14118
rect 2838 14116 2862 14118
rect 2622 14096 2918 14116
rect 2622 13084 2918 13104
rect 2678 13082 2702 13084
rect 2758 13082 2782 13084
rect 2838 13082 2862 13084
rect 2700 13030 2702 13082
rect 2764 13030 2776 13082
rect 2838 13030 2840 13082
rect 2678 13028 2702 13030
rect 2758 13028 2782 13030
rect 2838 13028 2862 13030
rect 2622 13008 2918 13028
rect 2622 11996 2918 12016
rect 2678 11994 2702 11996
rect 2758 11994 2782 11996
rect 2838 11994 2862 11996
rect 2700 11942 2702 11994
rect 2764 11942 2776 11994
rect 2838 11942 2840 11994
rect 2678 11940 2702 11942
rect 2758 11940 2782 11942
rect 2838 11940 2862 11942
rect 2622 11920 2918 11940
rect 2622 10908 2918 10928
rect 2678 10906 2702 10908
rect 2758 10906 2782 10908
rect 2838 10906 2862 10908
rect 2700 10854 2702 10906
rect 2764 10854 2776 10906
rect 2838 10854 2840 10906
rect 2678 10852 2702 10854
rect 2758 10852 2782 10854
rect 2838 10852 2862 10854
rect 2622 10832 2918 10852
rect 2622 9820 2918 9840
rect 2678 9818 2702 9820
rect 2758 9818 2782 9820
rect 2838 9818 2862 9820
rect 2700 9766 2702 9818
rect 2764 9766 2776 9818
rect 2838 9766 2840 9818
rect 2678 9764 2702 9766
rect 2758 9764 2782 9766
rect 2838 9764 2862 9766
rect 2622 9744 2918 9764
rect 2622 8732 2918 8752
rect 2678 8730 2702 8732
rect 2758 8730 2782 8732
rect 2838 8730 2862 8732
rect 2700 8678 2702 8730
rect 2764 8678 2776 8730
rect 2838 8678 2840 8730
rect 2678 8676 2702 8678
rect 2758 8676 2782 8678
rect 2838 8676 2862 8678
rect 2622 8656 2918 8676
rect 2622 7644 2918 7664
rect 2678 7642 2702 7644
rect 2758 7642 2782 7644
rect 2838 7642 2862 7644
rect 2700 7590 2702 7642
rect 2764 7590 2776 7642
rect 2838 7590 2840 7642
rect 2678 7588 2702 7590
rect 2758 7588 2782 7590
rect 2838 7588 2862 7590
rect 2622 7568 2918 7588
rect 2622 6556 2918 6576
rect 2678 6554 2702 6556
rect 2758 6554 2782 6556
rect 2838 6554 2862 6556
rect 2700 6502 2702 6554
rect 2764 6502 2776 6554
rect 2838 6502 2840 6554
rect 2678 6500 2702 6502
rect 2758 6500 2782 6502
rect 2838 6500 2862 6502
rect 2622 6480 2918 6500
rect 2622 5468 2918 5488
rect 2678 5466 2702 5468
rect 2758 5466 2782 5468
rect 2838 5466 2862 5468
rect 2700 5414 2702 5466
rect 2764 5414 2776 5466
rect 2838 5414 2840 5466
rect 2678 5412 2702 5414
rect 2758 5412 2782 5414
rect 2838 5412 2862 5414
rect 2622 5392 2918 5412
rect 2622 4380 2918 4400
rect 2678 4378 2702 4380
rect 2758 4378 2782 4380
rect 2838 4378 2862 4380
rect 2700 4326 2702 4378
rect 2764 4326 2776 4378
rect 2838 4326 2840 4378
rect 2678 4324 2702 4326
rect 2758 4324 2782 4326
rect 2838 4324 2862 4326
rect 2622 4304 2918 4324
rect 1320 4126 1440 4154
rect 938 82 994 480
rect 1320 82 1348 4126
rect 2622 3292 2918 3312
rect 2678 3290 2702 3292
rect 2758 3290 2782 3292
rect 2838 3290 2862 3292
rect 2700 3238 2702 3290
rect 2764 3238 2776 3290
rect 2838 3238 2840 3290
rect 2678 3236 2702 3238
rect 2758 3236 2782 3238
rect 2838 3236 2862 3238
rect 2622 3216 2918 3236
rect 2622 2204 2918 2224
rect 2678 2202 2702 2204
rect 2758 2202 2782 2204
rect 2838 2202 2862 2204
rect 2700 2150 2702 2202
rect 2764 2150 2776 2202
rect 2838 2150 2840 2202
rect 2678 2148 2702 2150
rect 2758 2148 2782 2150
rect 2838 2148 2862 2150
rect 2622 2128 2918 2148
rect 938 54 1348 82
rect 2870 82 2926 480
rect 2976 82 3004 208490
rect 3160 208282 3188 208626
rect 3344 208554 3372 214950
rect 3332 208548 3384 208554
rect 3332 208490 3384 208496
rect 3148 208276 3200 208282
rect 3148 208218 3200 208224
rect 3422 165880 3478 165889
rect 3422 165815 3478 165824
rect 3436 158234 3464 165815
rect 3424 158228 3476 158234
rect 3424 158170 3476 158176
rect 3528 150385 3556 237254
rect 3792 236768 3844 236774
rect 3792 236710 3844 236716
rect 3700 233776 3752 233782
rect 3700 233718 3752 233724
rect 3608 229220 3660 229226
rect 3608 229162 3660 229168
rect 3620 227526 3648 229162
rect 3608 227520 3660 227526
rect 3608 227462 3660 227468
rect 3620 227050 3648 227462
rect 3608 227044 3660 227050
rect 3608 226986 3660 226992
rect 3712 226334 3740 233718
rect 3804 232762 3832 236710
rect 3792 232756 3844 232762
rect 3792 232698 3844 232704
rect 3792 230784 3844 230790
rect 3792 230726 3844 230732
rect 3804 230382 3832 230726
rect 3792 230376 3844 230382
rect 3792 230318 3844 230324
rect 3804 229974 3832 230318
rect 3792 229968 3844 229974
rect 3792 229910 3844 229916
rect 3804 229702 3832 229910
rect 3792 229696 3844 229702
rect 3792 229638 3844 229644
rect 3804 229294 3832 229638
rect 3792 229288 3844 229294
rect 3792 229230 3844 229236
rect 3712 226306 3832 226334
rect 3700 221604 3752 221610
rect 3700 221546 3752 221552
rect 3712 215218 3740 221546
rect 3700 215212 3752 215218
rect 3700 215154 3752 215160
rect 3712 214810 3740 215154
rect 3700 214804 3752 214810
rect 3700 214746 3752 214752
rect 3700 209024 3752 209030
rect 3700 208966 3752 208972
rect 3712 208826 3740 208966
rect 3700 208820 3752 208826
rect 3700 208762 3752 208768
rect 3514 150376 3570 150385
rect 3514 150311 3570 150320
rect 3804 24313 3832 226306
rect 3896 210798 3924 332522
rect 4250 332520 4306 332528
rect 5448 332580 5500 332586
rect 5448 332522 5500 332528
rect 5538 332574 5672 332602
rect 4264 332491 4292 332520
rect 4289 330236 4585 330256
rect 4345 330234 4369 330236
rect 4425 330234 4449 330236
rect 4505 330234 4529 330236
rect 4367 330182 4369 330234
rect 4431 330182 4443 330234
rect 4505 330182 4507 330234
rect 4345 330180 4369 330182
rect 4425 330180 4449 330182
rect 4505 330180 4529 330182
rect 4289 330160 4585 330180
rect 4289 329148 4585 329168
rect 4345 329146 4369 329148
rect 4425 329146 4449 329148
rect 4505 329146 4529 329148
rect 4367 329094 4369 329146
rect 4431 329094 4443 329146
rect 4505 329094 4507 329146
rect 4345 329092 4369 329094
rect 4425 329092 4449 329094
rect 4505 329092 4529 329094
rect 4289 329072 4585 329092
rect 4289 328060 4585 328080
rect 4345 328058 4369 328060
rect 4425 328058 4449 328060
rect 4505 328058 4529 328060
rect 4367 328006 4369 328058
rect 4431 328006 4443 328058
rect 4505 328006 4507 328058
rect 4345 328004 4369 328006
rect 4425 328004 4449 328006
rect 4505 328004 4529 328006
rect 4289 327984 4585 328004
rect 4289 326972 4585 326992
rect 4345 326970 4369 326972
rect 4425 326970 4449 326972
rect 4505 326970 4529 326972
rect 4367 326918 4369 326970
rect 4431 326918 4443 326970
rect 4505 326918 4507 326970
rect 4345 326916 4369 326918
rect 4425 326916 4449 326918
rect 4505 326916 4529 326918
rect 4289 326896 4585 326916
rect 4289 325884 4585 325904
rect 4345 325882 4369 325884
rect 4425 325882 4449 325884
rect 4505 325882 4529 325884
rect 4367 325830 4369 325882
rect 4431 325830 4443 325882
rect 4505 325830 4507 325882
rect 4345 325828 4369 325830
rect 4425 325828 4449 325830
rect 4505 325828 4529 325830
rect 4289 325808 4585 325828
rect 4289 324796 4585 324816
rect 4345 324794 4369 324796
rect 4425 324794 4449 324796
rect 4505 324794 4529 324796
rect 4367 324742 4369 324794
rect 4431 324742 4443 324794
rect 4505 324742 4507 324794
rect 4345 324740 4369 324742
rect 4425 324740 4449 324742
rect 4505 324740 4529 324742
rect 4289 324720 4585 324740
rect 4289 323708 4585 323728
rect 4345 323706 4369 323708
rect 4425 323706 4449 323708
rect 4505 323706 4529 323708
rect 4367 323654 4369 323706
rect 4431 323654 4443 323706
rect 4505 323654 4507 323706
rect 4345 323652 4369 323654
rect 4425 323652 4449 323654
rect 4505 323652 4529 323654
rect 4289 323632 4585 323652
rect 4289 322620 4585 322640
rect 4345 322618 4369 322620
rect 4425 322618 4449 322620
rect 4505 322618 4529 322620
rect 4367 322566 4369 322618
rect 4431 322566 4443 322618
rect 4505 322566 4507 322618
rect 4345 322564 4369 322566
rect 4425 322564 4449 322566
rect 4505 322564 4529 322566
rect 4289 322544 4585 322564
rect 4289 321532 4585 321552
rect 4345 321530 4369 321532
rect 4425 321530 4449 321532
rect 4505 321530 4529 321532
rect 4367 321478 4369 321530
rect 4431 321478 4443 321530
rect 4505 321478 4507 321530
rect 4345 321476 4369 321478
rect 4425 321476 4449 321478
rect 4505 321476 4529 321478
rect 4289 321456 4585 321476
rect 4289 320444 4585 320464
rect 4345 320442 4369 320444
rect 4425 320442 4449 320444
rect 4505 320442 4529 320444
rect 4367 320390 4369 320442
rect 4431 320390 4443 320442
rect 4505 320390 4507 320442
rect 4345 320388 4369 320390
rect 4425 320388 4449 320390
rect 4505 320388 4529 320390
rect 4289 320368 4585 320388
rect 4289 319356 4585 319376
rect 4345 319354 4369 319356
rect 4425 319354 4449 319356
rect 4505 319354 4529 319356
rect 4367 319302 4369 319354
rect 4431 319302 4443 319354
rect 4505 319302 4507 319354
rect 4345 319300 4369 319302
rect 4425 319300 4449 319302
rect 4505 319300 4529 319302
rect 4289 319280 4585 319300
rect 4289 318268 4585 318288
rect 4345 318266 4369 318268
rect 4425 318266 4449 318268
rect 4505 318266 4529 318268
rect 4367 318214 4369 318266
rect 4431 318214 4443 318266
rect 4505 318214 4507 318266
rect 4345 318212 4369 318214
rect 4425 318212 4449 318214
rect 4505 318212 4529 318214
rect 4289 318192 4585 318212
rect 4289 317180 4585 317200
rect 4345 317178 4369 317180
rect 4425 317178 4449 317180
rect 4505 317178 4529 317180
rect 4367 317126 4369 317178
rect 4431 317126 4443 317178
rect 4505 317126 4507 317178
rect 4345 317124 4369 317126
rect 4425 317124 4449 317126
rect 4505 317124 4529 317126
rect 4289 317104 4585 317124
rect 4289 316092 4585 316112
rect 4345 316090 4369 316092
rect 4425 316090 4449 316092
rect 4505 316090 4529 316092
rect 4367 316038 4369 316090
rect 4431 316038 4443 316090
rect 4505 316038 4507 316090
rect 4345 316036 4369 316038
rect 4425 316036 4449 316038
rect 4505 316036 4529 316038
rect 4289 316016 4585 316036
rect 4289 315004 4585 315024
rect 4345 315002 4369 315004
rect 4425 315002 4449 315004
rect 4505 315002 4529 315004
rect 4367 314950 4369 315002
rect 4431 314950 4443 315002
rect 4505 314950 4507 315002
rect 4345 314948 4369 314950
rect 4425 314948 4449 314950
rect 4505 314948 4529 314950
rect 4289 314928 4585 314948
rect 4289 313916 4585 313936
rect 4345 313914 4369 313916
rect 4425 313914 4449 313916
rect 4505 313914 4529 313916
rect 4367 313862 4369 313914
rect 4431 313862 4443 313914
rect 4505 313862 4507 313914
rect 4345 313860 4369 313862
rect 4425 313860 4449 313862
rect 4505 313860 4529 313862
rect 4289 313840 4585 313860
rect 4289 312828 4585 312848
rect 4345 312826 4369 312828
rect 4425 312826 4449 312828
rect 4505 312826 4529 312828
rect 4367 312774 4369 312826
rect 4431 312774 4443 312826
rect 4505 312774 4507 312826
rect 4345 312772 4369 312774
rect 4425 312772 4449 312774
rect 4505 312772 4529 312774
rect 4289 312752 4585 312772
rect 4289 311740 4585 311760
rect 4345 311738 4369 311740
rect 4425 311738 4449 311740
rect 4505 311738 4529 311740
rect 4367 311686 4369 311738
rect 4431 311686 4443 311738
rect 4505 311686 4507 311738
rect 4345 311684 4369 311686
rect 4425 311684 4449 311686
rect 4505 311684 4529 311686
rect 4289 311664 4585 311684
rect 4289 310652 4585 310672
rect 4345 310650 4369 310652
rect 4425 310650 4449 310652
rect 4505 310650 4529 310652
rect 4367 310598 4369 310650
rect 4431 310598 4443 310650
rect 4505 310598 4507 310650
rect 4345 310596 4369 310598
rect 4425 310596 4449 310598
rect 4505 310596 4529 310598
rect 4289 310576 4585 310596
rect 4289 309564 4585 309584
rect 4345 309562 4369 309564
rect 4425 309562 4449 309564
rect 4505 309562 4529 309564
rect 4367 309510 4369 309562
rect 4431 309510 4443 309562
rect 4505 309510 4507 309562
rect 4345 309508 4369 309510
rect 4425 309508 4449 309510
rect 4505 309508 4529 309510
rect 4289 309488 4585 309508
rect 4289 308476 4585 308496
rect 4345 308474 4369 308476
rect 4425 308474 4449 308476
rect 4505 308474 4529 308476
rect 4367 308422 4369 308474
rect 4431 308422 4443 308474
rect 4505 308422 4507 308474
rect 4345 308420 4369 308422
rect 4425 308420 4449 308422
rect 4505 308420 4529 308422
rect 4289 308400 4585 308420
rect 4289 307388 4585 307408
rect 4345 307386 4369 307388
rect 4425 307386 4449 307388
rect 4505 307386 4529 307388
rect 4367 307334 4369 307386
rect 4431 307334 4443 307386
rect 4505 307334 4507 307386
rect 4345 307332 4369 307334
rect 4425 307332 4449 307334
rect 4505 307332 4529 307334
rect 4289 307312 4585 307332
rect 4289 306300 4585 306320
rect 4345 306298 4369 306300
rect 4425 306298 4449 306300
rect 4505 306298 4529 306300
rect 4367 306246 4369 306298
rect 4431 306246 4443 306298
rect 4505 306246 4507 306298
rect 4345 306244 4369 306246
rect 4425 306244 4449 306246
rect 4505 306244 4529 306246
rect 4289 306224 4585 306244
rect 4289 305212 4585 305232
rect 4345 305210 4369 305212
rect 4425 305210 4449 305212
rect 4505 305210 4529 305212
rect 4367 305158 4369 305210
rect 4431 305158 4443 305210
rect 4505 305158 4507 305210
rect 4345 305156 4369 305158
rect 4425 305156 4449 305158
rect 4505 305156 4529 305158
rect 4289 305136 4585 305156
rect 4289 304124 4585 304144
rect 4345 304122 4369 304124
rect 4425 304122 4449 304124
rect 4505 304122 4529 304124
rect 4367 304070 4369 304122
rect 4431 304070 4443 304122
rect 4505 304070 4507 304122
rect 4345 304068 4369 304070
rect 4425 304068 4449 304070
rect 4505 304068 4529 304070
rect 4289 304048 4585 304068
rect 4289 303036 4585 303056
rect 4345 303034 4369 303036
rect 4425 303034 4449 303036
rect 4505 303034 4529 303036
rect 4367 302982 4369 303034
rect 4431 302982 4443 303034
rect 4505 302982 4507 303034
rect 4345 302980 4369 302982
rect 4425 302980 4449 302982
rect 4505 302980 4529 302982
rect 4289 302960 4585 302980
rect 4289 301948 4585 301968
rect 4345 301946 4369 301948
rect 4425 301946 4449 301948
rect 4505 301946 4529 301948
rect 4367 301894 4369 301946
rect 4431 301894 4443 301946
rect 4505 301894 4507 301946
rect 4345 301892 4369 301894
rect 4425 301892 4449 301894
rect 4505 301892 4529 301894
rect 4289 301872 4585 301892
rect 4289 300860 4585 300880
rect 4345 300858 4369 300860
rect 4425 300858 4449 300860
rect 4505 300858 4529 300860
rect 4367 300806 4369 300858
rect 4431 300806 4443 300858
rect 4505 300806 4507 300858
rect 4345 300804 4369 300806
rect 4425 300804 4449 300806
rect 4505 300804 4529 300806
rect 4289 300784 4585 300804
rect 4289 299772 4585 299792
rect 4345 299770 4369 299772
rect 4425 299770 4449 299772
rect 4505 299770 4529 299772
rect 4367 299718 4369 299770
rect 4431 299718 4443 299770
rect 4505 299718 4507 299770
rect 4345 299716 4369 299718
rect 4425 299716 4449 299718
rect 4505 299716 4529 299718
rect 4289 299696 4585 299716
rect 4289 298684 4585 298704
rect 4345 298682 4369 298684
rect 4425 298682 4449 298684
rect 4505 298682 4529 298684
rect 4367 298630 4369 298682
rect 4431 298630 4443 298682
rect 4505 298630 4507 298682
rect 4345 298628 4369 298630
rect 4425 298628 4449 298630
rect 4505 298628 4529 298630
rect 4289 298608 4585 298628
rect 4289 297596 4585 297616
rect 4345 297594 4369 297596
rect 4425 297594 4449 297596
rect 4505 297594 4529 297596
rect 4367 297542 4369 297594
rect 4431 297542 4443 297594
rect 4505 297542 4507 297594
rect 4345 297540 4369 297542
rect 4425 297540 4449 297542
rect 4505 297540 4529 297542
rect 4289 297520 4585 297540
rect 4289 296508 4585 296528
rect 4345 296506 4369 296508
rect 4425 296506 4449 296508
rect 4505 296506 4529 296508
rect 4367 296454 4369 296506
rect 4431 296454 4443 296506
rect 4505 296454 4507 296506
rect 4345 296452 4369 296454
rect 4425 296452 4449 296454
rect 4505 296452 4529 296454
rect 4289 296432 4585 296452
rect 4289 295420 4585 295440
rect 4345 295418 4369 295420
rect 4425 295418 4449 295420
rect 4505 295418 4529 295420
rect 4367 295366 4369 295418
rect 4431 295366 4443 295418
rect 4505 295366 4507 295418
rect 4345 295364 4369 295366
rect 4425 295364 4449 295366
rect 4505 295364 4529 295366
rect 4289 295344 4585 295364
rect 4289 294332 4585 294352
rect 4345 294330 4369 294332
rect 4425 294330 4449 294332
rect 4505 294330 4529 294332
rect 4367 294278 4369 294330
rect 4431 294278 4443 294330
rect 4505 294278 4507 294330
rect 4345 294276 4369 294278
rect 4425 294276 4449 294278
rect 4505 294276 4529 294278
rect 4289 294256 4585 294276
rect 4289 293244 4585 293264
rect 4345 293242 4369 293244
rect 4425 293242 4449 293244
rect 4505 293242 4529 293244
rect 4367 293190 4369 293242
rect 4431 293190 4443 293242
rect 4505 293190 4507 293242
rect 4345 293188 4369 293190
rect 4425 293188 4449 293190
rect 4505 293188 4529 293190
rect 4289 293168 4585 293188
rect 4289 292156 4585 292176
rect 4345 292154 4369 292156
rect 4425 292154 4449 292156
rect 4505 292154 4529 292156
rect 4367 292102 4369 292154
rect 4431 292102 4443 292154
rect 4505 292102 4507 292154
rect 4345 292100 4369 292102
rect 4425 292100 4449 292102
rect 4505 292100 4529 292102
rect 4289 292080 4585 292100
rect 4289 291068 4585 291088
rect 4345 291066 4369 291068
rect 4425 291066 4449 291068
rect 4505 291066 4529 291068
rect 4367 291014 4369 291066
rect 4431 291014 4443 291066
rect 4505 291014 4507 291066
rect 4345 291012 4369 291014
rect 4425 291012 4449 291014
rect 4505 291012 4529 291014
rect 4289 290992 4585 291012
rect 4289 289980 4585 290000
rect 4345 289978 4369 289980
rect 4425 289978 4449 289980
rect 4505 289978 4529 289980
rect 4367 289926 4369 289978
rect 4431 289926 4443 289978
rect 4505 289926 4507 289978
rect 4345 289924 4369 289926
rect 4425 289924 4449 289926
rect 4505 289924 4529 289926
rect 4289 289904 4585 289924
rect 4289 288892 4585 288912
rect 4345 288890 4369 288892
rect 4425 288890 4449 288892
rect 4505 288890 4529 288892
rect 4367 288838 4369 288890
rect 4431 288838 4443 288890
rect 4505 288838 4507 288890
rect 4345 288836 4369 288838
rect 4425 288836 4449 288838
rect 4505 288836 4529 288838
rect 4289 288816 4585 288836
rect 4289 287804 4585 287824
rect 4345 287802 4369 287804
rect 4425 287802 4449 287804
rect 4505 287802 4529 287804
rect 4367 287750 4369 287802
rect 4431 287750 4443 287802
rect 4505 287750 4507 287802
rect 4345 287748 4369 287750
rect 4425 287748 4449 287750
rect 4505 287748 4529 287750
rect 4289 287728 4585 287748
rect 4289 286716 4585 286736
rect 4345 286714 4369 286716
rect 4425 286714 4449 286716
rect 4505 286714 4529 286716
rect 4367 286662 4369 286714
rect 4431 286662 4443 286714
rect 4505 286662 4507 286714
rect 4345 286660 4369 286662
rect 4425 286660 4449 286662
rect 4505 286660 4529 286662
rect 4289 286640 4585 286660
rect 4289 285628 4585 285648
rect 4345 285626 4369 285628
rect 4425 285626 4449 285628
rect 4505 285626 4529 285628
rect 4367 285574 4369 285626
rect 4431 285574 4443 285626
rect 4505 285574 4507 285626
rect 4345 285572 4369 285574
rect 4425 285572 4449 285574
rect 4505 285572 4529 285574
rect 4289 285552 4585 285572
rect 4289 284540 4585 284560
rect 4345 284538 4369 284540
rect 4425 284538 4449 284540
rect 4505 284538 4529 284540
rect 4367 284486 4369 284538
rect 4431 284486 4443 284538
rect 4505 284486 4507 284538
rect 4345 284484 4369 284486
rect 4425 284484 4449 284486
rect 4505 284484 4529 284486
rect 4289 284464 4585 284484
rect 4289 283452 4585 283472
rect 4345 283450 4369 283452
rect 4425 283450 4449 283452
rect 4505 283450 4529 283452
rect 4367 283398 4369 283450
rect 4431 283398 4443 283450
rect 4505 283398 4507 283450
rect 4345 283396 4369 283398
rect 4425 283396 4449 283398
rect 4505 283396 4529 283398
rect 4289 283376 4585 283396
rect 4289 282364 4585 282384
rect 4345 282362 4369 282364
rect 4425 282362 4449 282364
rect 4505 282362 4529 282364
rect 4367 282310 4369 282362
rect 4431 282310 4443 282362
rect 4505 282310 4507 282362
rect 4345 282308 4369 282310
rect 4425 282308 4449 282310
rect 4505 282308 4529 282310
rect 4289 282288 4585 282308
rect 4289 281276 4585 281296
rect 4345 281274 4369 281276
rect 4425 281274 4449 281276
rect 4505 281274 4529 281276
rect 4367 281222 4369 281274
rect 4431 281222 4443 281274
rect 4505 281222 4507 281274
rect 4345 281220 4369 281222
rect 4425 281220 4449 281222
rect 4505 281220 4529 281222
rect 4289 281200 4585 281220
rect 4289 280188 4585 280208
rect 4345 280186 4369 280188
rect 4425 280186 4449 280188
rect 4505 280186 4529 280188
rect 4367 280134 4369 280186
rect 4431 280134 4443 280186
rect 4505 280134 4507 280186
rect 4345 280132 4369 280134
rect 4425 280132 4449 280134
rect 4505 280132 4529 280134
rect 4289 280112 4585 280132
rect 4289 279100 4585 279120
rect 4345 279098 4369 279100
rect 4425 279098 4449 279100
rect 4505 279098 4529 279100
rect 4367 279046 4369 279098
rect 4431 279046 4443 279098
rect 4505 279046 4507 279098
rect 4345 279044 4369 279046
rect 4425 279044 4449 279046
rect 4505 279044 4529 279046
rect 4289 279024 4585 279044
rect 4289 278012 4585 278032
rect 4345 278010 4369 278012
rect 4425 278010 4449 278012
rect 4505 278010 4529 278012
rect 4367 277958 4369 278010
rect 4431 277958 4443 278010
rect 4505 277958 4507 278010
rect 4345 277956 4369 277958
rect 4425 277956 4449 277958
rect 4505 277956 4529 277958
rect 4289 277936 4585 277956
rect 4289 276924 4585 276944
rect 4345 276922 4369 276924
rect 4425 276922 4449 276924
rect 4505 276922 4529 276924
rect 4367 276870 4369 276922
rect 4431 276870 4443 276922
rect 4505 276870 4507 276922
rect 4345 276868 4369 276870
rect 4425 276868 4449 276870
rect 4505 276868 4529 276870
rect 4289 276848 4585 276868
rect 4289 275836 4585 275856
rect 4345 275834 4369 275836
rect 4425 275834 4449 275836
rect 4505 275834 4529 275836
rect 4367 275782 4369 275834
rect 4431 275782 4443 275834
rect 4505 275782 4507 275834
rect 4345 275780 4369 275782
rect 4425 275780 4449 275782
rect 4505 275780 4529 275782
rect 4289 275760 4585 275780
rect 4289 274748 4585 274768
rect 4345 274746 4369 274748
rect 4425 274746 4449 274748
rect 4505 274746 4529 274748
rect 4367 274694 4369 274746
rect 4431 274694 4443 274746
rect 4505 274694 4507 274746
rect 4345 274692 4369 274694
rect 4425 274692 4449 274694
rect 4505 274692 4529 274694
rect 4289 274672 4585 274692
rect 4289 273660 4585 273680
rect 4345 273658 4369 273660
rect 4425 273658 4449 273660
rect 4505 273658 4529 273660
rect 4367 273606 4369 273658
rect 4431 273606 4443 273658
rect 4505 273606 4507 273658
rect 4345 273604 4369 273606
rect 4425 273604 4449 273606
rect 4505 273604 4529 273606
rect 4289 273584 4585 273604
rect 4289 272572 4585 272592
rect 4345 272570 4369 272572
rect 4425 272570 4449 272572
rect 4505 272570 4529 272572
rect 4367 272518 4369 272570
rect 4431 272518 4443 272570
rect 4505 272518 4507 272570
rect 4345 272516 4369 272518
rect 4425 272516 4449 272518
rect 4505 272516 4529 272518
rect 4289 272496 4585 272516
rect 4289 271484 4585 271504
rect 4345 271482 4369 271484
rect 4425 271482 4449 271484
rect 4505 271482 4529 271484
rect 4367 271430 4369 271482
rect 4431 271430 4443 271482
rect 4505 271430 4507 271482
rect 4345 271428 4369 271430
rect 4425 271428 4449 271430
rect 4505 271428 4529 271430
rect 4289 271408 4585 271428
rect 4289 270396 4585 270416
rect 4345 270394 4369 270396
rect 4425 270394 4449 270396
rect 4505 270394 4529 270396
rect 4367 270342 4369 270394
rect 4431 270342 4443 270394
rect 4505 270342 4507 270394
rect 4345 270340 4369 270342
rect 4425 270340 4449 270342
rect 4505 270340 4529 270342
rect 4289 270320 4585 270340
rect 4289 269308 4585 269328
rect 4345 269306 4369 269308
rect 4425 269306 4449 269308
rect 4505 269306 4529 269308
rect 4367 269254 4369 269306
rect 4431 269254 4443 269306
rect 4505 269254 4507 269306
rect 4345 269252 4369 269254
rect 4425 269252 4449 269254
rect 4505 269252 4529 269254
rect 4289 269232 4585 269252
rect 4289 268220 4585 268240
rect 4345 268218 4369 268220
rect 4425 268218 4449 268220
rect 4505 268218 4529 268220
rect 4367 268166 4369 268218
rect 4431 268166 4443 268218
rect 4505 268166 4507 268218
rect 4345 268164 4369 268166
rect 4425 268164 4449 268166
rect 4505 268164 4529 268166
rect 4289 268144 4585 268164
rect 4289 267132 4585 267152
rect 4345 267130 4369 267132
rect 4425 267130 4449 267132
rect 4505 267130 4529 267132
rect 4367 267078 4369 267130
rect 4431 267078 4443 267130
rect 4505 267078 4507 267130
rect 4345 267076 4369 267078
rect 4425 267076 4449 267078
rect 4505 267076 4529 267078
rect 4289 267056 4585 267076
rect 4289 266044 4585 266064
rect 4345 266042 4369 266044
rect 4425 266042 4449 266044
rect 4505 266042 4529 266044
rect 4367 265990 4369 266042
rect 4431 265990 4443 266042
rect 4505 265990 4507 266042
rect 4345 265988 4369 265990
rect 4425 265988 4449 265990
rect 4505 265988 4529 265990
rect 4289 265968 4585 265988
rect 4289 264956 4585 264976
rect 4345 264954 4369 264956
rect 4425 264954 4449 264956
rect 4505 264954 4529 264956
rect 4367 264902 4369 264954
rect 4431 264902 4443 264954
rect 4505 264902 4507 264954
rect 4345 264900 4369 264902
rect 4425 264900 4449 264902
rect 4505 264900 4529 264902
rect 4289 264880 4585 264900
rect 4289 263868 4585 263888
rect 4345 263866 4369 263868
rect 4425 263866 4449 263868
rect 4505 263866 4529 263868
rect 4367 263814 4369 263866
rect 4431 263814 4443 263866
rect 4505 263814 4507 263866
rect 4345 263812 4369 263814
rect 4425 263812 4449 263814
rect 4505 263812 4529 263814
rect 4289 263792 4585 263812
rect 4289 262780 4585 262800
rect 4345 262778 4369 262780
rect 4425 262778 4449 262780
rect 4505 262778 4529 262780
rect 4367 262726 4369 262778
rect 4431 262726 4443 262778
rect 4505 262726 4507 262778
rect 4345 262724 4369 262726
rect 4425 262724 4449 262726
rect 4505 262724 4529 262726
rect 4289 262704 4585 262724
rect 4289 261692 4585 261712
rect 4345 261690 4369 261692
rect 4425 261690 4449 261692
rect 4505 261690 4529 261692
rect 4367 261638 4369 261690
rect 4431 261638 4443 261690
rect 4505 261638 4507 261690
rect 4345 261636 4369 261638
rect 4425 261636 4449 261638
rect 4505 261636 4529 261638
rect 4289 261616 4585 261636
rect 4289 260604 4585 260624
rect 4345 260602 4369 260604
rect 4425 260602 4449 260604
rect 4505 260602 4529 260604
rect 4367 260550 4369 260602
rect 4431 260550 4443 260602
rect 4505 260550 4507 260602
rect 4345 260548 4369 260550
rect 4425 260548 4449 260550
rect 4505 260548 4529 260550
rect 4289 260528 4585 260548
rect 4289 259516 4585 259536
rect 4345 259514 4369 259516
rect 4425 259514 4449 259516
rect 4505 259514 4529 259516
rect 4367 259462 4369 259514
rect 4431 259462 4443 259514
rect 4505 259462 4507 259514
rect 4345 259460 4369 259462
rect 4425 259460 4449 259462
rect 4505 259460 4529 259462
rect 4289 259440 4585 259460
rect 4289 258428 4585 258448
rect 4345 258426 4369 258428
rect 4425 258426 4449 258428
rect 4505 258426 4529 258428
rect 4367 258374 4369 258426
rect 4431 258374 4443 258426
rect 4505 258374 4507 258426
rect 4345 258372 4369 258374
rect 4425 258372 4449 258374
rect 4505 258372 4529 258374
rect 4289 258352 4585 258372
rect 4289 257340 4585 257360
rect 4345 257338 4369 257340
rect 4425 257338 4449 257340
rect 4505 257338 4529 257340
rect 4367 257286 4369 257338
rect 4431 257286 4443 257338
rect 4505 257286 4507 257338
rect 4345 257284 4369 257286
rect 4425 257284 4449 257286
rect 4505 257284 4529 257286
rect 4289 257264 4585 257284
rect 4289 256252 4585 256272
rect 4345 256250 4369 256252
rect 4425 256250 4449 256252
rect 4505 256250 4529 256252
rect 4367 256198 4369 256250
rect 4431 256198 4443 256250
rect 4505 256198 4507 256250
rect 4345 256196 4369 256198
rect 4425 256196 4449 256198
rect 4505 256196 4529 256198
rect 4289 256176 4585 256196
rect 4289 255164 4585 255184
rect 4345 255162 4369 255164
rect 4425 255162 4449 255164
rect 4505 255162 4529 255164
rect 4367 255110 4369 255162
rect 4431 255110 4443 255162
rect 4505 255110 4507 255162
rect 4345 255108 4369 255110
rect 4425 255108 4449 255110
rect 4505 255108 4529 255110
rect 4289 255088 4585 255108
rect 4289 254076 4585 254096
rect 4345 254074 4369 254076
rect 4425 254074 4449 254076
rect 4505 254074 4529 254076
rect 4367 254022 4369 254074
rect 4431 254022 4443 254074
rect 4505 254022 4507 254074
rect 4345 254020 4369 254022
rect 4425 254020 4449 254022
rect 4505 254020 4529 254022
rect 4289 254000 4585 254020
rect 4289 252988 4585 253008
rect 4345 252986 4369 252988
rect 4425 252986 4449 252988
rect 4505 252986 4529 252988
rect 4367 252934 4369 252986
rect 4431 252934 4443 252986
rect 4505 252934 4507 252986
rect 4345 252932 4369 252934
rect 4425 252932 4449 252934
rect 4505 252932 4529 252934
rect 4289 252912 4585 252932
rect 4289 251900 4585 251920
rect 4345 251898 4369 251900
rect 4425 251898 4449 251900
rect 4505 251898 4529 251900
rect 4367 251846 4369 251898
rect 4431 251846 4443 251898
rect 4505 251846 4507 251898
rect 4345 251844 4369 251846
rect 4425 251844 4449 251846
rect 4505 251844 4529 251846
rect 4289 251824 4585 251844
rect 4289 250812 4585 250832
rect 4345 250810 4369 250812
rect 4425 250810 4449 250812
rect 4505 250810 4529 250812
rect 4367 250758 4369 250810
rect 4431 250758 4443 250810
rect 4505 250758 4507 250810
rect 4345 250756 4369 250758
rect 4425 250756 4449 250758
rect 4505 250756 4529 250758
rect 4289 250736 4585 250756
rect 4289 249724 4585 249744
rect 4345 249722 4369 249724
rect 4425 249722 4449 249724
rect 4505 249722 4529 249724
rect 4367 249670 4369 249722
rect 4431 249670 4443 249722
rect 4505 249670 4507 249722
rect 4345 249668 4369 249670
rect 4425 249668 4449 249670
rect 4505 249668 4529 249670
rect 4289 249648 4585 249668
rect 4289 248636 4585 248656
rect 4345 248634 4369 248636
rect 4425 248634 4449 248636
rect 4505 248634 4529 248636
rect 4367 248582 4369 248634
rect 4431 248582 4443 248634
rect 4505 248582 4507 248634
rect 4345 248580 4369 248582
rect 4425 248580 4449 248582
rect 4505 248580 4529 248582
rect 4289 248560 4585 248580
rect 4289 247548 4585 247568
rect 4345 247546 4369 247548
rect 4425 247546 4449 247548
rect 4505 247546 4529 247548
rect 4367 247494 4369 247546
rect 4431 247494 4443 247546
rect 4505 247494 4507 247546
rect 4345 247492 4369 247494
rect 4425 247492 4449 247494
rect 4505 247492 4529 247494
rect 4289 247472 4585 247492
rect 4289 246460 4585 246480
rect 4345 246458 4369 246460
rect 4425 246458 4449 246460
rect 4505 246458 4529 246460
rect 4367 246406 4369 246458
rect 4431 246406 4443 246458
rect 4505 246406 4507 246458
rect 4345 246404 4369 246406
rect 4425 246404 4449 246406
rect 4505 246404 4529 246406
rect 4289 246384 4585 246404
rect 4289 245372 4585 245392
rect 4345 245370 4369 245372
rect 4425 245370 4449 245372
rect 4505 245370 4529 245372
rect 4367 245318 4369 245370
rect 4431 245318 4443 245370
rect 4505 245318 4507 245370
rect 4345 245316 4369 245318
rect 4425 245316 4449 245318
rect 4505 245316 4529 245318
rect 4289 245296 4585 245316
rect 4289 244284 4585 244304
rect 4345 244282 4369 244284
rect 4425 244282 4449 244284
rect 4505 244282 4529 244284
rect 4367 244230 4369 244282
rect 4431 244230 4443 244282
rect 4505 244230 4507 244282
rect 4345 244228 4369 244230
rect 4425 244228 4449 244230
rect 4505 244228 4529 244230
rect 4289 244208 4585 244228
rect 4289 243196 4585 243216
rect 4345 243194 4369 243196
rect 4425 243194 4449 243196
rect 4505 243194 4529 243196
rect 4367 243142 4369 243194
rect 4431 243142 4443 243194
rect 4505 243142 4507 243194
rect 4345 243140 4369 243142
rect 4425 243140 4449 243142
rect 4505 243140 4529 243142
rect 4289 243120 4585 243140
rect 4289 242108 4585 242128
rect 4345 242106 4369 242108
rect 4425 242106 4449 242108
rect 4505 242106 4529 242108
rect 4367 242054 4369 242106
rect 4431 242054 4443 242106
rect 4505 242054 4507 242106
rect 4345 242052 4369 242054
rect 4425 242052 4449 242054
rect 4505 242052 4529 242054
rect 4289 242032 4585 242052
rect 4289 241020 4585 241040
rect 4345 241018 4369 241020
rect 4425 241018 4449 241020
rect 4505 241018 4529 241020
rect 4367 240966 4369 241018
rect 4431 240966 4443 241018
rect 4505 240966 4507 241018
rect 4345 240964 4369 240966
rect 4425 240964 4449 240966
rect 4505 240964 4529 240966
rect 4289 240944 4585 240964
rect 4289 239932 4585 239952
rect 4345 239930 4369 239932
rect 4425 239930 4449 239932
rect 4505 239930 4529 239932
rect 4367 239878 4369 239930
rect 4431 239878 4443 239930
rect 4505 239878 4507 239930
rect 4345 239876 4369 239878
rect 4425 239876 4449 239878
rect 4505 239876 4529 239878
rect 4289 239856 4585 239876
rect 4289 238844 4585 238864
rect 4345 238842 4369 238844
rect 4425 238842 4449 238844
rect 4505 238842 4529 238844
rect 4367 238790 4369 238842
rect 4431 238790 4443 238842
rect 4505 238790 4507 238842
rect 4345 238788 4369 238790
rect 4425 238788 4449 238790
rect 4505 238788 4529 238790
rect 4289 238768 4585 238788
rect 4289 237756 4585 237776
rect 4345 237754 4369 237756
rect 4425 237754 4449 237756
rect 4505 237754 4529 237756
rect 4367 237702 4369 237754
rect 4431 237702 4443 237754
rect 4505 237702 4507 237754
rect 4345 237700 4369 237702
rect 4425 237700 4449 237702
rect 4505 237700 4529 237702
rect 4289 237680 4585 237700
rect 4289 236668 4585 236688
rect 4345 236666 4369 236668
rect 4425 236666 4449 236668
rect 4505 236666 4529 236668
rect 4367 236614 4369 236666
rect 4431 236614 4443 236666
rect 4505 236614 4507 236666
rect 4345 236612 4369 236614
rect 4425 236612 4449 236614
rect 4505 236612 4529 236614
rect 4289 236592 4585 236612
rect 4289 235580 4585 235600
rect 4345 235578 4369 235580
rect 4425 235578 4449 235580
rect 4505 235578 4529 235580
rect 4367 235526 4369 235578
rect 4431 235526 4443 235578
rect 4505 235526 4507 235578
rect 4345 235524 4369 235526
rect 4425 235524 4449 235526
rect 4505 235524 4529 235526
rect 4289 235504 4585 235524
rect 4289 234492 4585 234512
rect 4345 234490 4369 234492
rect 4425 234490 4449 234492
rect 4505 234490 4529 234492
rect 4367 234438 4369 234490
rect 4431 234438 4443 234490
rect 4505 234438 4507 234490
rect 4345 234436 4369 234438
rect 4425 234436 4449 234438
rect 4505 234436 4529 234438
rect 4289 234416 4585 234436
rect 4160 234320 4212 234326
rect 4160 234262 4212 234268
rect 3976 234184 4028 234190
rect 3976 234126 4028 234132
rect 3988 233510 4016 234126
rect 4172 233510 4200 234262
rect 4988 234048 5040 234054
rect 4988 233990 5040 233996
rect 5000 233714 5028 233990
rect 4988 233708 5040 233714
rect 4988 233650 5040 233656
rect 4712 233640 4764 233646
rect 4712 233582 4764 233588
rect 3976 233504 4028 233510
rect 3976 233446 4028 233452
rect 4160 233504 4212 233510
rect 4160 233446 4212 233452
rect 3988 230246 4016 233446
rect 4172 232490 4200 233446
rect 4289 233404 4585 233424
rect 4345 233402 4369 233404
rect 4425 233402 4449 233404
rect 4505 233402 4529 233404
rect 4367 233350 4369 233402
rect 4431 233350 4443 233402
rect 4505 233350 4507 233402
rect 4345 233348 4369 233350
rect 4425 233348 4449 233350
rect 4505 233348 4529 233350
rect 4289 233328 4585 233348
rect 4724 233306 4752 233582
rect 5000 233306 5028 233650
rect 5356 233504 5408 233510
rect 5356 233446 5408 233452
rect 4712 233300 4764 233306
rect 4712 233242 4764 233248
rect 4988 233300 5040 233306
rect 4988 233242 5040 233248
rect 4068 232484 4120 232490
rect 4068 232426 4120 232432
rect 4160 232484 4212 232490
rect 4160 232426 4212 232432
rect 4080 231062 4108 232426
rect 4289 232316 4585 232336
rect 4345 232314 4369 232316
rect 4425 232314 4449 232316
rect 4505 232314 4529 232316
rect 4367 232262 4369 232314
rect 4431 232262 4443 232314
rect 4505 232262 4507 232314
rect 4345 232260 4369 232262
rect 4425 232260 4449 232262
rect 4505 232260 4529 232262
rect 4289 232240 4585 232260
rect 4289 231228 4585 231248
rect 4345 231226 4369 231228
rect 4425 231226 4449 231228
rect 4505 231226 4529 231228
rect 4367 231174 4369 231226
rect 4431 231174 4443 231226
rect 4505 231174 4507 231226
rect 4345 231172 4369 231174
rect 4425 231172 4449 231174
rect 4505 231172 4529 231174
rect 4289 231152 4585 231172
rect 5368 231130 5396 233446
rect 4712 231124 4764 231130
rect 4712 231066 4764 231072
rect 5356 231124 5408 231130
rect 5356 231066 5408 231072
rect 4068 231056 4120 231062
rect 4068 230998 4120 231004
rect 4068 230512 4120 230518
rect 4068 230454 4120 230460
rect 3976 230240 4028 230246
rect 3976 230182 4028 230188
rect 4080 229906 4108 230454
rect 4724 230246 4752 231066
rect 4988 230920 5040 230926
rect 4988 230862 5040 230868
rect 5000 230246 5028 230862
rect 4712 230240 4764 230246
rect 4712 230182 4764 230188
rect 4988 230240 5040 230246
rect 4988 230182 5040 230188
rect 4289 230140 4585 230160
rect 4345 230138 4369 230140
rect 4425 230138 4449 230140
rect 4505 230138 4529 230140
rect 4367 230086 4369 230138
rect 4431 230086 4443 230138
rect 4505 230086 4507 230138
rect 4345 230084 4369 230086
rect 4425 230084 4449 230086
rect 4505 230084 4529 230086
rect 4289 230064 4585 230084
rect 4068 229900 4120 229906
rect 4068 229842 4120 229848
rect 4080 229158 4108 229842
rect 4620 229832 4672 229838
rect 4620 229774 4672 229780
rect 4068 229152 4120 229158
rect 4068 229094 4120 229100
rect 4289 229052 4585 229072
rect 4345 229050 4369 229052
rect 4425 229050 4449 229052
rect 4505 229050 4529 229052
rect 4367 228998 4369 229050
rect 4431 228998 4443 229050
rect 4505 228998 4507 229050
rect 4345 228996 4369 228998
rect 4425 228996 4449 228998
rect 4505 228996 4529 228998
rect 4289 228976 4585 228996
rect 4289 227964 4585 227984
rect 4345 227962 4369 227964
rect 4425 227962 4449 227964
rect 4505 227962 4529 227964
rect 4367 227910 4369 227962
rect 4431 227910 4443 227962
rect 4505 227910 4507 227962
rect 4345 227908 4369 227910
rect 4425 227908 4449 227910
rect 4505 227908 4529 227910
rect 4289 227888 4585 227908
rect 4068 226976 4120 226982
rect 4068 226918 4120 226924
rect 4080 225554 4108 226918
rect 4289 226876 4585 226896
rect 4345 226874 4369 226876
rect 4425 226874 4449 226876
rect 4505 226874 4529 226876
rect 4367 226822 4369 226874
rect 4431 226822 4443 226874
rect 4505 226822 4507 226874
rect 4345 226820 4369 226822
rect 4425 226820 4449 226822
rect 4505 226820 4529 226822
rect 4289 226800 4585 226820
rect 4632 226642 4660 229774
rect 4724 226778 4752 230182
rect 5000 229362 5028 230182
rect 5080 229900 5132 229906
rect 5080 229842 5132 229848
rect 5092 229430 5120 229842
rect 5356 229764 5408 229770
rect 5356 229706 5408 229712
rect 5368 229498 5396 229706
rect 5356 229492 5408 229498
rect 5356 229434 5408 229440
rect 5080 229424 5132 229430
rect 5080 229366 5132 229372
rect 4988 229356 5040 229362
rect 4988 229298 5040 229304
rect 4804 229152 4856 229158
rect 4804 229094 4856 229100
rect 4816 228818 4844 229094
rect 4804 228812 4856 228818
rect 4804 228754 4856 228760
rect 4816 228070 4844 228754
rect 4804 228064 4856 228070
rect 4804 228006 4856 228012
rect 4712 226772 4764 226778
rect 4712 226714 4764 226720
rect 4620 226636 4672 226642
rect 4620 226578 4672 226584
rect 4632 226234 4660 226578
rect 4620 226228 4672 226234
rect 4620 226170 4672 226176
rect 4724 225962 4752 226714
rect 4712 225956 4764 225962
rect 4712 225898 4764 225904
rect 4289 225788 4585 225808
rect 4345 225786 4369 225788
rect 4425 225786 4449 225788
rect 4505 225786 4529 225788
rect 4367 225734 4369 225786
rect 4431 225734 4443 225786
rect 4505 225734 4507 225786
rect 4345 225732 4369 225734
rect 4425 225732 4449 225734
rect 4505 225732 4529 225734
rect 4289 225712 4585 225732
rect 4724 225690 4752 225898
rect 4712 225684 4764 225690
rect 4712 225626 4764 225632
rect 4068 225548 4120 225554
rect 4068 225490 4120 225496
rect 4080 225146 4108 225490
rect 4068 225140 4120 225146
rect 4068 225082 4120 225088
rect 4724 225078 4752 225626
rect 3976 225072 4028 225078
rect 3976 225014 4028 225020
rect 4712 225072 4764 225078
rect 4712 225014 4764 225020
rect 3988 215014 4016 225014
rect 4289 224700 4585 224720
rect 4345 224698 4369 224700
rect 4425 224698 4449 224700
rect 4505 224698 4529 224700
rect 4367 224646 4369 224698
rect 4431 224646 4443 224698
rect 4505 224646 4507 224698
rect 4345 224644 4369 224646
rect 4425 224644 4449 224646
rect 4505 224644 4529 224646
rect 4289 224624 4585 224644
rect 4289 223612 4585 223632
rect 4345 223610 4369 223612
rect 4425 223610 4449 223612
rect 4505 223610 4529 223612
rect 4367 223558 4369 223610
rect 4431 223558 4443 223610
rect 4505 223558 4507 223610
rect 4345 223556 4369 223558
rect 4425 223556 4449 223558
rect 4505 223556 4529 223558
rect 4289 223536 4585 223556
rect 4289 222524 4585 222544
rect 4345 222522 4369 222524
rect 4425 222522 4449 222524
rect 4505 222522 4529 222524
rect 4367 222470 4369 222522
rect 4431 222470 4443 222522
rect 4505 222470 4507 222522
rect 4345 222468 4369 222470
rect 4425 222468 4449 222470
rect 4505 222468 4529 222470
rect 4289 222448 4585 222468
rect 4289 221436 4585 221456
rect 4345 221434 4369 221436
rect 4425 221434 4449 221436
rect 4505 221434 4529 221436
rect 4367 221382 4369 221434
rect 4431 221382 4443 221434
rect 4505 221382 4507 221434
rect 4345 221380 4369 221382
rect 4425 221380 4449 221382
rect 4505 221380 4529 221382
rect 4289 221360 4585 221380
rect 4289 220348 4585 220368
rect 4345 220346 4369 220348
rect 4425 220346 4449 220348
rect 4505 220346 4529 220348
rect 4367 220294 4369 220346
rect 4431 220294 4443 220346
rect 4505 220294 4507 220346
rect 4345 220292 4369 220294
rect 4425 220292 4449 220294
rect 4505 220292 4529 220294
rect 4289 220272 4585 220292
rect 4289 219260 4585 219280
rect 4345 219258 4369 219260
rect 4425 219258 4449 219260
rect 4505 219258 4529 219260
rect 4367 219206 4369 219258
rect 4431 219206 4443 219258
rect 4505 219206 4507 219258
rect 4345 219204 4369 219206
rect 4425 219204 4449 219206
rect 4505 219204 4529 219206
rect 4289 219184 4585 219204
rect 4289 218172 4585 218192
rect 4345 218170 4369 218172
rect 4425 218170 4449 218172
rect 4505 218170 4529 218172
rect 4367 218118 4369 218170
rect 4431 218118 4443 218170
rect 4505 218118 4507 218170
rect 4345 218116 4369 218118
rect 4425 218116 4449 218118
rect 4505 218116 4529 218118
rect 4289 218096 4585 218116
rect 4289 217084 4585 217104
rect 4345 217082 4369 217084
rect 4425 217082 4449 217084
rect 4505 217082 4529 217084
rect 4367 217030 4369 217082
rect 4431 217030 4443 217082
rect 4505 217030 4507 217082
rect 4345 217028 4369 217030
rect 4425 217028 4449 217030
rect 4505 217028 4529 217030
rect 4289 217008 4585 217028
rect 4289 215996 4585 216016
rect 4345 215994 4369 215996
rect 4425 215994 4449 215996
rect 4505 215994 4529 215996
rect 4367 215942 4369 215994
rect 4431 215942 4443 215994
rect 4505 215942 4507 215994
rect 4345 215940 4369 215942
rect 4425 215940 4449 215942
rect 4505 215940 4529 215942
rect 4289 215920 4585 215940
rect 3976 215008 4028 215014
rect 3976 214950 4028 214956
rect 4620 215008 4672 215014
rect 4620 214950 4672 214956
rect 4289 214908 4585 214928
rect 4345 214906 4369 214908
rect 4425 214906 4449 214908
rect 4505 214906 4529 214908
rect 4367 214854 4369 214906
rect 4431 214854 4443 214906
rect 4505 214854 4507 214906
rect 4345 214852 4369 214854
rect 4425 214852 4449 214854
rect 4505 214852 4529 214854
rect 4289 214832 4585 214852
rect 4289 213820 4585 213840
rect 4345 213818 4369 213820
rect 4425 213818 4449 213820
rect 4505 213818 4529 213820
rect 4367 213766 4369 213818
rect 4431 213766 4443 213818
rect 4505 213766 4507 213818
rect 4345 213764 4369 213766
rect 4425 213764 4449 213766
rect 4505 213764 4529 213766
rect 4289 213744 4585 213764
rect 4289 212732 4585 212752
rect 4345 212730 4369 212732
rect 4425 212730 4449 212732
rect 4505 212730 4529 212732
rect 4367 212678 4369 212730
rect 4431 212678 4443 212730
rect 4505 212678 4507 212730
rect 4345 212676 4369 212678
rect 4425 212676 4449 212678
rect 4505 212676 4529 212678
rect 4289 212656 4585 212676
rect 4632 211954 4660 214950
rect 4620 211948 4672 211954
rect 4620 211890 4672 211896
rect 4289 211644 4585 211664
rect 4345 211642 4369 211644
rect 4425 211642 4449 211644
rect 4505 211642 4529 211644
rect 4367 211590 4369 211642
rect 4431 211590 4443 211642
rect 4505 211590 4507 211642
rect 4345 211588 4369 211590
rect 4425 211588 4449 211590
rect 4505 211588 4529 211590
rect 4289 211568 4585 211588
rect 4632 211546 4660 211890
rect 4620 211540 4672 211546
rect 4620 211482 4672 211488
rect 3884 210792 3936 210798
rect 3884 210734 3936 210740
rect 3896 209914 3924 210734
rect 4289 210556 4585 210576
rect 4345 210554 4369 210556
rect 4425 210554 4449 210556
rect 4505 210554 4529 210556
rect 4367 210502 4369 210554
rect 4431 210502 4443 210554
rect 4505 210502 4507 210554
rect 4345 210500 4369 210502
rect 4425 210500 4449 210502
rect 4505 210500 4529 210502
rect 4289 210480 4585 210500
rect 3884 209908 3936 209914
rect 3884 209850 3936 209856
rect 4289 209468 4585 209488
rect 4345 209466 4369 209468
rect 4425 209466 4449 209468
rect 4505 209466 4529 209468
rect 4367 209414 4369 209466
rect 4431 209414 4443 209466
rect 4505 209414 4507 209466
rect 4345 209412 4369 209414
rect 4425 209412 4449 209414
rect 4505 209412 4529 209414
rect 4289 209392 4585 209412
rect 4289 208380 4585 208400
rect 4345 208378 4369 208380
rect 4425 208378 4449 208380
rect 4505 208378 4529 208380
rect 4367 208326 4369 208378
rect 4431 208326 4443 208378
rect 4505 208326 4507 208378
rect 4345 208324 4369 208326
rect 4425 208324 4449 208326
rect 4505 208324 4529 208326
rect 4289 208304 4585 208324
rect 4289 207292 4585 207312
rect 4345 207290 4369 207292
rect 4425 207290 4449 207292
rect 4505 207290 4529 207292
rect 4367 207238 4369 207290
rect 4431 207238 4443 207290
rect 4505 207238 4507 207290
rect 4345 207236 4369 207238
rect 4425 207236 4449 207238
rect 4505 207236 4529 207238
rect 4289 207216 4585 207236
rect 4289 206204 4585 206224
rect 4345 206202 4369 206204
rect 4425 206202 4449 206204
rect 4505 206202 4529 206204
rect 4367 206150 4369 206202
rect 4431 206150 4443 206202
rect 4505 206150 4507 206202
rect 4345 206148 4369 206150
rect 4425 206148 4449 206150
rect 4505 206148 4529 206150
rect 4289 206128 4585 206148
rect 4289 205116 4585 205136
rect 4345 205114 4369 205116
rect 4425 205114 4449 205116
rect 4505 205114 4529 205116
rect 4367 205062 4369 205114
rect 4431 205062 4443 205114
rect 4505 205062 4507 205114
rect 4345 205060 4369 205062
rect 4425 205060 4449 205062
rect 4505 205060 4529 205062
rect 4289 205040 4585 205060
rect 4289 204028 4585 204048
rect 4345 204026 4369 204028
rect 4425 204026 4449 204028
rect 4505 204026 4529 204028
rect 4367 203974 4369 204026
rect 4431 203974 4443 204026
rect 4505 203974 4507 204026
rect 4345 203972 4369 203974
rect 4425 203972 4449 203974
rect 4505 203972 4529 203974
rect 4289 203952 4585 203972
rect 4289 202940 4585 202960
rect 4345 202938 4369 202940
rect 4425 202938 4449 202940
rect 4505 202938 4529 202940
rect 4367 202886 4369 202938
rect 4431 202886 4443 202938
rect 4505 202886 4507 202938
rect 4345 202884 4369 202886
rect 4425 202884 4449 202886
rect 4505 202884 4529 202886
rect 4289 202864 4585 202884
rect 4289 201852 4585 201872
rect 4345 201850 4369 201852
rect 4425 201850 4449 201852
rect 4505 201850 4529 201852
rect 4367 201798 4369 201850
rect 4431 201798 4443 201850
rect 4505 201798 4507 201850
rect 4345 201796 4369 201798
rect 4425 201796 4449 201798
rect 4505 201796 4529 201798
rect 4289 201776 4585 201796
rect 4289 200764 4585 200784
rect 4345 200762 4369 200764
rect 4425 200762 4449 200764
rect 4505 200762 4529 200764
rect 4367 200710 4369 200762
rect 4431 200710 4443 200762
rect 4505 200710 4507 200762
rect 4345 200708 4369 200710
rect 4425 200708 4449 200710
rect 4505 200708 4529 200710
rect 4289 200688 4585 200708
rect 4289 199676 4585 199696
rect 4345 199674 4369 199676
rect 4425 199674 4449 199676
rect 4505 199674 4529 199676
rect 4367 199622 4369 199674
rect 4431 199622 4443 199674
rect 4505 199622 4507 199674
rect 4345 199620 4369 199622
rect 4425 199620 4449 199622
rect 4505 199620 4529 199622
rect 4289 199600 4585 199620
rect 4289 198588 4585 198608
rect 4345 198586 4369 198588
rect 4425 198586 4449 198588
rect 4505 198586 4529 198588
rect 4367 198534 4369 198586
rect 4431 198534 4443 198586
rect 4505 198534 4507 198586
rect 4345 198532 4369 198534
rect 4425 198532 4449 198534
rect 4505 198532 4529 198534
rect 4289 198512 4585 198532
rect 4289 197500 4585 197520
rect 4345 197498 4369 197500
rect 4425 197498 4449 197500
rect 4505 197498 4529 197500
rect 4367 197446 4369 197498
rect 4431 197446 4443 197498
rect 4505 197446 4507 197498
rect 4345 197444 4369 197446
rect 4425 197444 4449 197446
rect 4505 197444 4529 197446
rect 4289 197424 4585 197444
rect 4289 196412 4585 196432
rect 4345 196410 4369 196412
rect 4425 196410 4449 196412
rect 4505 196410 4529 196412
rect 4367 196358 4369 196410
rect 4431 196358 4443 196410
rect 4505 196358 4507 196410
rect 4345 196356 4369 196358
rect 4425 196356 4449 196358
rect 4505 196356 4529 196358
rect 4289 196336 4585 196356
rect 4289 195324 4585 195344
rect 4345 195322 4369 195324
rect 4425 195322 4449 195324
rect 4505 195322 4529 195324
rect 4367 195270 4369 195322
rect 4431 195270 4443 195322
rect 4505 195270 4507 195322
rect 4345 195268 4369 195270
rect 4425 195268 4449 195270
rect 4505 195268 4529 195270
rect 4289 195248 4585 195268
rect 4289 194236 4585 194256
rect 4345 194234 4369 194236
rect 4425 194234 4449 194236
rect 4505 194234 4529 194236
rect 4367 194182 4369 194234
rect 4431 194182 4443 194234
rect 4505 194182 4507 194234
rect 4345 194180 4369 194182
rect 4425 194180 4449 194182
rect 4505 194180 4529 194182
rect 4289 194160 4585 194180
rect 4289 193148 4585 193168
rect 4345 193146 4369 193148
rect 4425 193146 4449 193148
rect 4505 193146 4529 193148
rect 4367 193094 4369 193146
rect 4431 193094 4443 193146
rect 4505 193094 4507 193146
rect 4345 193092 4369 193094
rect 4425 193092 4449 193094
rect 4505 193092 4529 193094
rect 4289 193072 4585 193092
rect 4289 192060 4585 192080
rect 4345 192058 4369 192060
rect 4425 192058 4449 192060
rect 4505 192058 4529 192060
rect 4367 192006 4369 192058
rect 4431 192006 4443 192058
rect 4505 192006 4507 192058
rect 4345 192004 4369 192006
rect 4425 192004 4449 192006
rect 4505 192004 4529 192006
rect 4289 191984 4585 192004
rect 4289 190972 4585 190992
rect 4345 190970 4369 190972
rect 4425 190970 4449 190972
rect 4505 190970 4529 190972
rect 4367 190918 4369 190970
rect 4431 190918 4443 190970
rect 4505 190918 4507 190970
rect 4345 190916 4369 190918
rect 4425 190916 4449 190918
rect 4505 190916 4529 190918
rect 4289 190896 4585 190916
rect 4289 189884 4585 189904
rect 4345 189882 4369 189884
rect 4425 189882 4449 189884
rect 4505 189882 4529 189884
rect 4367 189830 4369 189882
rect 4431 189830 4443 189882
rect 4505 189830 4507 189882
rect 4345 189828 4369 189830
rect 4425 189828 4449 189830
rect 4505 189828 4529 189830
rect 4289 189808 4585 189828
rect 4289 188796 4585 188816
rect 4345 188794 4369 188796
rect 4425 188794 4449 188796
rect 4505 188794 4529 188796
rect 4367 188742 4369 188794
rect 4431 188742 4443 188794
rect 4505 188742 4507 188794
rect 4345 188740 4369 188742
rect 4425 188740 4449 188742
rect 4505 188740 4529 188742
rect 4289 188720 4585 188740
rect 4289 187708 4585 187728
rect 4345 187706 4369 187708
rect 4425 187706 4449 187708
rect 4505 187706 4529 187708
rect 4367 187654 4369 187706
rect 4431 187654 4443 187706
rect 4505 187654 4507 187706
rect 4345 187652 4369 187654
rect 4425 187652 4449 187654
rect 4505 187652 4529 187654
rect 4289 187632 4585 187652
rect 4289 186620 4585 186640
rect 4345 186618 4369 186620
rect 4425 186618 4449 186620
rect 4505 186618 4529 186620
rect 4367 186566 4369 186618
rect 4431 186566 4443 186618
rect 4505 186566 4507 186618
rect 4345 186564 4369 186566
rect 4425 186564 4449 186566
rect 4505 186564 4529 186566
rect 4289 186544 4585 186564
rect 4289 185532 4585 185552
rect 4345 185530 4369 185532
rect 4425 185530 4449 185532
rect 4505 185530 4529 185532
rect 4367 185478 4369 185530
rect 4431 185478 4443 185530
rect 4505 185478 4507 185530
rect 4345 185476 4369 185478
rect 4425 185476 4449 185478
rect 4505 185476 4529 185478
rect 4289 185456 4585 185476
rect 4289 184444 4585 184464
rect 4345 184442 4369 184444
rect 4425 184442 4449 184444
rect 4505 184442 4529 184444
rect 4367 184390 4369 184442
rect 4431 184390 4443 184442
rect 4505 184390 4507 184442
rect 4345 184388 4369 184390
rect 4425 184388 4449 184390
rect 4505 184388 4529 184390
rect 4289 184368 4585 184388
rect 4289 183356 4585 183376
rect 4345 183354 4369 183356
rect 4425 183354 4449 183356
rect 4505 183354 4529 183356
rect 4367 183302 4369 183354
rect 4431 183302 4443 183354
rect 4505 183302 4507 183354
rect 4345 183300 4369 183302
rect 4425 183300 4449 183302
rect 4505 183300 4529 183302
rect 4289 183280 4585 183300
rect 4289 182268 4585 182288
rect 4345 182266 4369 182268
rect 4425 182266 4449 182268
rect 4505 182266 4529 182268
rect 4367 182214 4369 182266
rect 4431 182214 4443 182266
rect 4505 182214 4507 182266
rect 4345 182212 4369 182214
rect 4425 182212 4449 182214
rect 4505 182212 4529 182214
rect 4289 182192 4585 182212
rect 4289 181180 4585 181200
rect 4345 181178 4369 181180
rect 4425 181178 4449 181180
rect 4505 181178 4529 181180
rect 4367 181126 4369 181178
rect 4431 181126 4443 181178
rect 4505 181126 4507 181178
rect 4345 181124 4369 181126
rect 4425 181124 4449 181126
rect 4505 181124 4529 181126
rect 4289 181104 4585 181124
rect 4289 180092 4585 180112
rect 4345 180090 4369 180092
rect 4425 180090 4449 180092
rect 4505 180090 4529 180092
rect 4367 180038 4369 180090
rect 4431 180038 4443 180090
rect 4505 180038 4507 180090
rect 4345 180036 4369 180038
rect 4425 180036 4449 180038
rect 4505 180036 4529 180038
rect 4289 180016 4585 180036
rect 4289 179004 4585 179024
rect 4345 179002 4369 179004
rect 4425 179002 4449 179004
rect 4505 179002 4529 179004
rect 4367 178950 4369 179002
rect 4431 178950 4443 179002
rect 4505 178950 4507 179002
rect 4345 178948 4369 178950
rect 4425 178948 4449 178950
rect 4505 178948 4529 178950
rect 4289 178928 4585 178948
rect 4289 177916 4585 177936
rect 4345 177914 4369 177916
rect 4425 177914 4449 177916
rect 4505 177914 4529 177916
rect 4367 177862 4369 177914
rect 4431 177862 4443 177914
rect 4505 177862 4507 177914
rect 4345 177860 4369 177862
rect 4425 177860 4449 177862
rect 4505 177860 4529 177862
rect 4289 177840 4585 177860
rect 4289 176828 4585 176848
rect 4345 176826 4369 176828
rect 4425 176826 4449 176828
rect 4505 176826 4529 176828
rect 4367 176774 4369 176826
rect 4431 176774 4443 176826
rect 4505 176774 4507 176826
rect 4345 176772 4369 176774
rect 4425 176772 4449 176774
rect 4505 176772 4529 176774
rect 4289 176752 4585 176772
rect 4289 175740 4585 175760
rect 4345 175738 4369 175740
rect 4425 175738 4449 175740
rect 4505 175738 4529 175740
rect 4367 175686 4369 175738
rect 4431 175686 4443 175738
rect 4505 175686 4507 175738
rect 4345 175684 4369 175686
rect 4425 175684 4449 175686
rect 4505 175684 4529 175686
rect 4289 175664 4585 175684
rect 4289 174652 4585 174672
rect 4345 174650 4369 174652
rect 4425 174650 4449 174652
rect 4505 174650 4529 174652
rect 4367 174598 4369 174650
rect 4431 174598 4443 174650
rect 4505 174598 4507 174650
rect 4345 174596 4369 174598
rect 4425 174596 4449 174598
rect 4505 174596 4529 174598
rect 4289 174576 4585 174596
rect 4289 173564 4585 173584
rect 4345 173562 4369 173564
rect 4425 173562 4449 173564
rect 4505 173562 4529 173564
rect 4367 173510 4369 173562
rect 4431 173510 4443 173562
rect 4505 173510 4507 173562
rect 4345 173508 4369 173510
rect 4425 173508 4449 173510
rect 4505 173508 4529 173510
rect 4289 173488 4585 173508
rect 4289 172476 4585 172496
rect 4345 172474 4369 172476
rect 4425 172474 4449 172476
rect 4505 172474 4529 172476
rect 4367 172422 4369 172474
rect 4431 172422 4443 172474
rect 4505 172422 4507 172474
rect 4345 172420 4369 172422
rect 4425 172420 4449 172422
rect 4505 172420 4529 172422
rect 4289 172400 4585 172420
rect 4289 171388 4585 171408
rect 4345 171386 4369 171388
rect 4425 171386 4449 171388
rect 4505 171386 4529 171388
rect 4367 171334 4369 171386
rect 4431 171334 4443 171386
rect 4505 171334 4507 171386
rect 4345 171332 4369 171334
rect 4425 171332 4449 171334
rect 4505 171332 4529 171334
rect 4289 171312 4585 171332
rect 4289 170300 4585 170320
rect 4345 170298 4369 170300
rect 4425 170298 4449 170300
rect 4505 170298 4529 170300
rect 4367 170246 4369 170298
rect 4431 170246 4443 170298
rect 4505 170246 4507 170298
rect 4345 170244 4369 170246
rect 4425 170244 4449 170246
rect 4505 170244 4529 170246
rect 4289 170224 4585 170244
rect 4289 169212 4585 169232
rect 4345 169210 4369 169212
rect 4425 169210 4449 169212
rect 4505 169210 4529 169212
rect 4367 169158 4369 169210
rect 4431 169158 4443 169210
rect 4505 169158 4507 169210
rect 4345 169156 4369 169158
rect 4425 169156 4449 169158
rect 4505 169156 4529 169158
rect 4289 169136 4585 169156
rect 4289 168124 4585 168144
rect 4345 168122 4369 168124
rect 4425 168122 4449 168124
rect 4505 168122 4529 168124
rect 4367 168070 4369 168122
rect 4431 168070 4443 168122
rect 4505 168070 4507 168122
rect 4345 168068 4369 168070
rect 4425 168068 4449 168070
rect 4505 168068 4529 168070
rect 4289 168048 4585 168068
rect 4289 167036 4585 167056
rect 4345 167034 4369 167036
rect 4425 167034 4449 167036
rect 4505 167034 4529 167036
rect 4367 166982 4369 167034
rect 4431 166982 4443 167034
rect 4505 166982 4507 167034
rect 4345 166980 4369 166982
rect 4425 166980 4449 166982
rect 4505 166980 4529 166982
rect 4289 166960 4585 166980
rect 4289 165948 4585 165968
rect 4345 165946 4369 165948
rect 4425 165946 4449 165948
rect 4505 165946 4529 165948
rect 4367 165894 4369 165946
rect 4431 165894 4443 165946
rect 4505 165894 4507 165946
rect 4345 165892 4369 165894
rect 4425 165892 4449 165894
rect 4505 165892 4529 165894
rect 4289 165872 4585 165892
rect 4289 164860 4585 164880
rect 4345 164858 4369 164860
rect 4425 164858 4449 164860
rect 4505 164858 4529 164860
rect 4367 164806 4369 164858
rect 4431 164806 4443 164858
rect 4505 164806 4507 164858
rect 4345 164804 4369 164806
rect 4425 164804 4449 164806
rect 4505 164804 4529 164806
rect 4289 164784 4585 164804
rect 4289 163772 4585 163792
rect 4345 163770 4369 163772
rect 4425 163770 4449 163772
rect 4505 163770 4529 163772
rect 4367 163718 4369 163770
rect 4431 163718 4443 163770
rect 4505 163718 4507 163770
rect 4345 163716 4369 163718
rect 4425 163716 4449 163718
rect 4505 163716 4529 163718
rect 4289 163696 4585 163716
rect 4289 162684 4585 162704
rect 4345 162682 4369 162684
rect 4425 162682 4449 162684
rect 4505 162682 4529 162684
rect 4367 162630 4369 162682
rect 4431 162630 4443 162682
rect 4505 162630 4507 162682
rect 4345 162628 4369 162630
rect 4425 162628 4449 162630
rect 4505 162628 4529 162630
rect 4289 162608 4585 162628
rect 4289 161596 4585 161616
rect 4345 161594 4369 161596
rect 4425 161594 4449 161596
rect 4505 161594 4529 161596
rect 4367 161542 4369 161594
rect 4431 161542 4443 161594
rect 4505 161542 4507 161594
rect 4345 161540 4369 161542
rect 4425 161540 4449 161542
rect 4505 161540 4529 161542
rect 4289 161520 4585 161540
rect 4289 160508 4585 160528
rect 4345 160506 4369 160508
rect 4425 160506 4449 160508
rect 4505 160506 4529 160508
rect 4367 160454 4369 160506
rect 4431 160454 4443 160506
rect 4505 160454 4507 160506
rect 4345 160452 4369 160454
rect 4425 160452 4449 160454
rect 4505 160452 4529 160454
rect 4289 160432 4585 160452
rect 4289 159420 4585 159440
rect 4345 159418 4369 159420
rect 4425 159418 4449 159420
rect 4505 159418 4529 159420
rect 4367 159366 4369 159418
rect 4431 159366 4443 159418
rect 4505 159366 4507 159418
rect 4345 159364 4369 159366
rect 4425 159364 4449 159366
rect 4505 159364 4529 159366
rect 4289 159344 4585 159364
rect 4289 158332 4585 158352
rect 4345 158330 4369 158332
rect 4425 158330 4449 158332
rect 4505 158330 4529 158332
rect 4367 158278 4369 158330
rect 4431 158278 4443 158330
rect 4505 158278 4507 158330
rect 4345 158276 4369 158278
rect 4425 158276 4449 158278
rect 4505 158276 4529 158278
rect 4289 158256 4585 158276
rect 4068 158092 4120 158098
rect 4068 158034 4120 158040
rect 4080 157690 4108 158034
rect 4068 157684 4120 157690
rect 4068 157626 4120 157632
rect 4289 157244 4585 157264
rect 4345 157242 4369 157244
rect 4425 157242 4449 157244
rect 4505 157242 4529 157244
rect 4367 157190 4369 157242
rect 4431 157190 4443 157242
rect 4505 157190 4507 157242
rect 4345 157188 4369 157190
rect 4425 157188 4449 157190
rect 4505 157188 4529 157190
rect 4289 157168 4585 157188
rect 4289 156156 4585 156176
rect 4345 156154 4369 156156
rect 4425 156154 4449 156156
rect 4505 156154 4529 156156
rect 4367 156102 4369 156154
rect 4431 156102 4443 156154
rect 4505 156102 4507 156154
rect 4345 156100 4369 156102
rect 4425 156100 4449 156102
rect 4505 156100 4529 156102
rect 4289 156080 4585 156100
rect 4289 155068 4585 155088
rect 4345 155066 4369 155068
rect 4425 155066 4449 155068
rect 4505 155066 4529 155068
rect 4367 155014 4369 155066
rect 4431 155014 4443 155066
rect 4505 155014 4507 155066
rect 4345 155012 4369 155014
rect 4425 155012 4449 155014
rect 4505 155012 4529 155014
rect 4289 154992 4585 155012
rect 4289 153980 4585 154000
rect 4345 153978 4369 153980
rect 4425 153978 4449 153980
rect 4505 153978 4529 153980
rect 4367 153926 4369 153978
rect 4431 153926 4443 153978
rect 4505 153926 4507 153978
rect 4345 153924 4369 153926
rect 4425 153924 4449 153926
rect 4505 153924 4529 153926
rect 4289 153904 4585 153924
rect 4289 152892 4585 152912
rect 4345 152890 4369 152892
rect 4425 152890 4449 152892
rect 4505 152890 4529 152892
rect 4367 152838 4369 152890
rect 4431 152838 4443 152890
rect 4505 152838 4507 152890
rect 4345 152836 4369 152838
rect 4425 152836 4449 152838
rect 4505 152836 4529 152838
rect 4289 152816 4585 152836
rect 4289 151804 4585 151824
rect 4345 151802 4369 151804
rect 4425 151802 4449 151804
rect 4505 151802 4529 151804
rect 4367 151750 4369 151802
rect 4431 151750 4443 151802
rect 4505 151750 4507 151802
rect 4345 151748 4369 151750
rect 4425 151748 4449 151750
rect 4505 151748 4529 151750
rect 4289 151728 4585 151748
rect 4289 150716 4585 150736
rect 4345 150714 4369 150716
rect 4425 150714 4449 150716
rect 4505 150714 4529 150716
rect 4367 150662 4369 150714
rect 4431 150662 4443 150714
rect 4505 150662 4507 150714
rect 4345 150660 4369 150662
rect 4425 150660 4449 150662
rect 4505 150660 4529 150662
rect 4289 150640 4585 150660
rect 4289 149628 4585 149648
rect 4345 149626 4369 149628
rect 4425 149626 4449 149628
rect 4505 149626 4529 149628
rect 4367 149574 4369 149626
rect 4431 149574 4443 149626
rect 4505 149574 4507 149626
rect 4345 149572 4369 149574
rect 4425 149572 4449 149574
rect 4505 149572 4529 149574
rect 4289 149552 4585 149572
rect 4289 148540 4585 148560
rect 4345 148538 4369 148540
rect 4425 148538 4449 148540
rect 4505 148538 4529 148540
rect 4367 148486 4369 148538
rect 4431 148486 4443 148538
rect 4505 148486 4507 148538
rect 4345 148484 4369 148486
rect 4425 148484 4449 148486
rect 4505 148484 4529 148486
rect 4289 148464 4585 148484
rect 4289 147452 4585 147472
rect 4345 147450 4369 147452
rect 4425 147450 4449 147452
rect 4505 147450 4529 147452
rect 4367 147398 4369 147450
rect 4431 147398 4443 147450
rect 4505 147398 4507 147450
rect 4345 147396 4369 147398
rect 4425 147396 4449 147398
rect 4505 147396 4529 147398
rect 4289 147376 4585 147396
rect 4289 146364 4585 146384
rect 4345 146362 4369 146364
rect 4425 146362 4449 146364
rect 4505 146362 4529 146364
rect 4367 146310 4369 146362
rect 4431 146310 4443 146362
rect 4505 146310 4507 146362
rect 4345 146308 4369 146310
rect 4425 146308 4449 146310
rect 4505 146308 4529 146310
rect 4289 146288 4585 146308
rect 4289 145276 4585 145296
rect 4345 145274 4369 145276
rect 4425 145274 4449 145276
rect 4505 145274 4529 145276
rect 4367 145222 4369 145274
rect 4431 145222 4443 145274
rect 4505 145222 4507 145274
rect 4345 145220 4369 145222
rect 4425 145220 4449 145222
rect 4505 145220 4529 145222
rect 4289 145200 4585 145220
rect 4289 144188 4585 144208
rect 4345 144186 4369 144188
rect 4425 144186 4449 144188
rect 4505 144186 4529 144188
rect 4367 144134 4369 144186
rect 4431 144134 4443 144186
rect 4505 144134 4507 144186
rect 4345 144132 4369 144134
rect 4425 144132 4449 144134
rect 4505 144132 4529 144134
rect 4289 144112 4585 144132
rect 4289 143100 4585 143120
rect 4345 143098 4369 143100
rect 4425 143098 4449 143100
rect 4505 143098 4529 143100
rect 4367 143046 4369 143098
rect 4431 143046 4443 143098
rect 4505 143046 4507 143098
rect 4345 143044 4369 143046
rect 4425 143044 4449 143046
rect 4505 143044 4529 143046
rect 4289 143024 4585 143044
rect 4289 142012 4585 142032
rect 4345 142010 4369 142012
rect 4425 142010 4449 142012
rect 4505 142010 4529 142012
rect 4367 141958 4369 142010
rect 4431 141958 4443 142010
rect 4505 141958 4507 142010
rect 4345 141956 4369 141958
rect 4425 141956 4449 141958
rect 4505 141956 4529 141958
rect 4289 141936 4585 141956
rect 4289 140924 4585 140944
rect 4345 140922 4369 140924
rect 4425 140922 4449 140924
rect 4505 140922 4529 140924
rect 4367 140870 4369 140922
rect 4431 140870 4443 140922
rect 4505 140870 4507 140922
rect 4345 140868 4369 140870
rect 4425 140868 4449 140870
rect 4505 140868 4529 140870
rect 4289 140848 4585 140868
rect 4289 139836 4585 139856
rect 4345 139834 4369 139836
rect 4425 139834 4449 139836
rect 4505 139834 4529 139836
rect 4367 139782 4369 139834
rect 4431 139782 4443 139834
rect 4505 139782 4507 139834
rect 4345 139780 4369 139782
rect 4425 139780 4449 139782
rect 4505 139780 4529 139782
rect 4289 139760 4585 139780
rect 4289 138748 4585 138768
rect 4345 138746 4369 138748
rect 4425 138746 4449 138748
rect 4505 138746 4529 138748
rect 4367 138694 4369 138746
rect 4431 138694 4443 138746
rect 4505 138694 4507 138746
rect 4345 138692 4369 138694
rect 4425 138692 4449 138694
rect 4505 138692 4529 138694
rect 4289 138672 4585 138692
rect 4289 137660 4585 137680
rect 4345 137658 4369 137660
rect 4425 137658 4449 137660
rect 4505 137658 4529 137660
rect 4367 137606 4369 137658
rect 4431 137606 4443 137658
rect 4505 137606 4507 137658
rect 4345 137604 4369 137606
rect 4425 137604 4449 137606
rect 4505 137604 4529 137606
rect 4289 137584 4585 137604
rect 4289 136572 4585 136592
rect 4345 136570 4369 136572
rect 4425 136570 4449 136572
rect 4505 136570 4529 136572
rect 4367 136518 4369 136570
rect 4431 136518 4443 136570
rect 4505 136518 4507 136570
rect 4345 136516 4369 136518
rect 4425 136516 4449 136518
rect 4505 136516 4529 136518
rect 4289 136496 4585 136516
rect 4289 135484 4585 135504
rect 4345 135482 4369 135484
rect 4425 135482 4449 135484
rect 4505 135482 4529 135484
rect 4367 135430 4369 135482
rect 4431 135430 4443 135482
rect 4505 135430 4507 135482
rect 4345 135428 4369 135430
rect 4425 135428 4449 135430
rect 4505 135428 4529 135430
rect 4289 135408 4585 135428
rect 4289 134396 4585 134416
rect 4345 134394 4369 134396
rect 4425 134394 4449 134396
rect 4505 134394 4529 134396
rect 4367 134342 4369 134394
rect 4431 134342 4443 134394
rect 4505 134342 4507 134394
rect 4345 134340 4369 134342
rect 4425 134340 4449 134342
rect 4505 134340 4529 134342
rect 4289 134320 4585 134340
rect 4289 133308 4585 133328
rect 4345 133306 4369 133308
rect 4425 133306 4449 133308
rect 4505 133306 4529 133308
rect 4367 133254 4369 133306
rect 4431 133254 4443 133306
rect 4505 133254 4507 133306
rect 4345 133252 4369 133254
rect 4425 133252 4449 133254
rect 4505 133252 4529 133254
rect 4289 133232 4585 133252
rect 4289 132220 4585 132240
rect 4345 132218 4369 132220
rect 4425 132218 4449 132220
rect 4505 132218 4529 132220
rect 4367 132166 4369 132218
rect 4431 132166 4443 132218
rect 4505 132166 4507 132218
rect 4345 132164 4369 132166
rect 4425 132164 4449 132166
rect 4505 132164 4529 132166
rect 4289 132144 4585 132164
rect 4289 131132 4585 131152
rect 4345 131130 4369 131132
rect 4425 131130 4449 131132
rect 4505 131130 4529 131132
rect 4367 131078 4369 131130
rect 4431 131078 4443 131130
rect 4505 131078 4507 131130
rect 4345 131076 4369 131078
rect 4425 131076 4449 131078
rect 4505 131076 4529 131078
rect 4289 131056 4585 131076
rect 4289 130044 4585 130064
rect 4345 130042 4369 130044
rect 4425 130042 4449 130044
rect 4505 130042 4529 130044
rect 4367 129990 4369 130042
rect 4431 129990 4443 130042
rect 4505 129990 4507 130042
rect 4345 129988 4369 129990
rect 4425 129988 4449 129990
rect 4505 129988 4529 129990
rect 4289 129968 4585 129988
rect 4289 128956 4585 128976
rect 4345 128954 4369 128956
rect 4425 128954 4449 128956
rect 4505 128954 4529 128956
rect 4367 128902 4369 128954
rect 4431 128902 4443 128954
rect 4505 128902 4507 128954
rect 4345 128900 4369 128902
rect 4425 128900 4449 128902
rect 4505 128900 4529 128902
rect 4289 128880 4585 128900
rect 4289 127868 4585 127888
rect 4345 127866 4369 127868
rect 4425 127866 4449 127868
rect 4505 127866 4529 127868
rect 4367 127814 4369 127866
rect 4431 127814 4443 127866
rect 4505 127814 4507 127866
rect 4345 127812 4369 127814
rect 4425 127812 4449 127814
rect 4505 127812 4529 127814
rect 4289 127792 4585 127812
rect 4289 126780 4585 126800
rect 4345 126778 4369 126780
rect 4425 126778 4449 126780
rect 4505 126778 4529 126780
rect 4367 126726 4369 126778
rect 4431 126726 4443 126778
rect 4505 126726 4507 126778
rect 4345 126724 4369 126726
rect 4425 126724 4449 126726
rect 4505 126724 4529 126726
rect 4289 126704 4585 126724
rect 4289 125692 4585 125712
rect 4345 125690 4369 125692
rect 4425 125690 4449 125692
rect 4505 125690 4529 125692
rect 4367 125638 4369 125690
rect 4431 125638 4443 125690
rect 4505 125638 4507 125690
rect 4345 125636 4369 125638
rect 4425 125636 4449 125638
rect 4505 125636 4529 125638
rect 4289 125616 4585 125636
rect 4289 124604 4585 124624
rect 4345 124602 4369 124604
rect 4425 124602 4449 124604
rect 4505 124602 4529 124604
rect 4367 124550 4369 124602
rect 4431 124550 4443 124602
rect 4505 124550 4507 124602
rect 4345 124548 4369 124550
rect 4425 124548 4449 124550
rect 4505 124548 4529 124550
rect 4289 124528 4585 124548
rect 4289 123516 4585 123536
rect 4345 123514 4369 123516
rect 4425 123514 4449 123516
rect 4505 123514 4529 123516
rect 4367 123462 4369 123514
rect 4431 123462 4443 123514
rect 4505 123462 4507 123514
rect 4345 123460 4369 123462
rect 4425 123460 4449 123462
rect 4505 123460 4529 123462
rect 4289 123440 4585 123460
rect 4289 122428 4585 122448
rect 4345 122426 4369 122428
rect 4425 122426 4449 122428
rect 4505 122426 4529 122428
rect 4367 122374 4369 122426
rect 4431 122374 4443 122426
rect 4505 122374 4507 122426
rect 4345 122372 4369 122374
rect 4425 122372 4449 122374
rect 4505 122372 4529 122374
rect 4289 122352 4585 122372
rect 4289 121340 4585 121360
rect 4345 121338 4369 121340
rect 4425 121338 4449 121340
rect 4505 121338 4529 121340
rect 4367 121286 4369 121338
rect 4431 121286 4443 121338
rect 4505 121286 4507 121338
rect 4345 121284 4369 121286
rect 4425 121284 4449 121286
rect 4505 121284 4529 121286
rect 4289 121264 4585 121284
rect 4289 120252 4585 120272
rect 4345 120250 4369 120252
rect 4425 120250 4449 120252
rect 4505 120250 4529 120252
rect 4367 120198 4369 120250
rect 4431 120198 4443 120250
rect 4505 120198 4507 120250
rect 4345 120196 4369 120198
rect 4425 120196 4449 120198
rect 4505 120196 4529 120198
rect 4289 120176 4585 120196
rect 4289 119164 4585 119184
rect 4345 119162 4369 119164
rect 4425 119162 4449 119164
rect 4505 119162 4529 119164
rect 4367 119110 4369 119162
rect 4431 119110 4443 119162
rect 4505 119110 4507 119162
rect 4345 119108 4369 119110
rect 4425 119108 4449 119110
rect 4505 119108 4529 119110
rect 4289 119088 4585 119108
rect 4289 118076 4585 118096
rect 4345 118074 4369 118076
rect 4425 118074 4449 118076
rect 4505 118074 4529 118076
rect 4367 118022 4369 118074
rect 4431 118022 4443 118074
rect 4505 118022 4507 118074
rect 4345 118020 4369 118022
rect 4425 118020 4449 118022
rect 4505 118020 4529 118022
rect 4289 118000 4585 118020
rect 4289 116988 4585 117008
rect 4345 116986 4369 116988
rect 4425 116986 4449 116988
rect 4505 116986 4529 116988
rect 4367 116934 4369 116986
rect 4431 116934 4443 116986
rect 4505 116934 4507 116986
rect 4345 116932 4369 116934
rect 4425 116932 4449 116934
rect 4505 116932 4529 116934
rect 4289 116912 4585 116932
rect 4289 115900 4585 115920
rect 4345 115898 4369 115900
rect 4425 115898 4449 115900
rect 4505 115898 4529 115900
rect 4367 115846 4369 115898
rect 4431 115846 4443 115898
rect 4505 115846 4507 115898
rect 4345 115844 4369 115846
rect 4425 115844 4449 115846
rect 4505 115844 4529 115846
rect 4289 115824 4585 115844
rect 4289 114812 4585 114832
rect 4345 114810 4369 114812
rect 4425 114810 4449 114812
rect 4505 114810 4529 114812
rect 4367 114758 4369 114810
rect 4431 114758 4443 114810
rect 4505 114758 4507 114810
rect 4345 114756 4369 114758
rect 4425 114756 4449 114758
rect 4505 114756 4529 114758
rect 4289 114736 4585 114756
rect 4289 113724 4585 113744
rect 4345 113722 4369 113724
rect 4425 113722 4449 113724
rect 4505 113722 4529 113724
rect 4367 113670 4369 113722
rect 4431 113670 4443 113722
rect 4505 113670 4507 113722
rect 4345 113668 4369 113670
rect 4425 113668 4449 113670
rect 4505 113668 4529 113670
rect 4289 113648 4585 113668
rect 4289 112636 4585 112656
rect 4345 112634 4369 112636
rect 4425 112634 4449 112636
rect 4505 112634 4529 112636
rect 4367 112582 4369 112634
rect 4431 112582 4443 112634
rect 4505 112582 4507 112634
rect 4345 112580 4369 112582
rect 4425 112580 4449 112582
rect 4505 112580 4529 112582
rect 4289 112560 4585 112580
rect 4289 111548 4585 111568
rect 4345 111546 4369 111548
rect 4425 111546 4449 111548
rect 4505 111546 4529 111548
rect 4367 111494 4369 111546
rect 4431 111494 4443 111546
rect 4505 111494 4507 111546
rect 4345 111492 4369 111494
rect 4425 111492 4449 111494
rect 4505 111492 4529 111494
rect 4289 111472 4585 111492
rect 4289 110460 4585 110480
rect 4345 110458 4369 110460
rect 4425 110458 4449 110460
rect 4505 110458 4529 110460
rect 4367 110406 4369 110458
rect 4431 110406 4443 110458
rect 4505 110406 4507 110458
rect 4345 110404 4369 110406
rect 4425 110404 4449 110406
rect 4505 110404 4529 110406
rect 4289 110384 4585 110404
rect 4289 109372 4585 109392
rect 4345 109370 4369 109372
rect 4425 109370 4449 109372
rect 4505 109370 4529 109372
rect 4367 109318 4369 109370
rect 4431 109318 4443 109370
rect 4505 109318 4507 109370
rect 4345 109316 4369 109318
rect 4425 109316 4449 109318
rect 4505 109316 4529 109318
rect 4289 109296 4585 109316
rect 4289 108284 4585 108304
rect 4345 108282 4369 108284
rect 4425 108282 4449 108284
rect 4505 108282 4529 108284
rect 4367 108230 4369 108282
rect 4431 108230 4443 108282
rect 4505 108230 4507 108282
rect 4345 108228 4369 108230
rect 4425 108228 4449 108230
rect 4505 108228 4529 108230
rect 4289 108208 4585 108228
rect 4289 107196 4585 107216
rect 4345 107194 4369 107196
rect 4425 107194 4449 107196
rect 4505 107194 4529 107196
rect 4367 107142 4369 107194
rect 4431 107142 4443 107194
rect 4505 107142 4507 107194
rect 4345 107140 4369 107142
rect 4425 107140 4449 107142
rect 4505 107140 4529 107142
rect 4289 107120 4585 107140
rect 4289 106108 4585 106128
rect 4345 106106 4369 106108
rect 4425 106106 4449 106108
rect 4505 106106 4529 106108
rect 4367 106054 4369 106106
rect 4431 106054 4443 106106
rect 4505 106054 4507 106106
rect 4345 106052 4369 106054
rect 4425 106052 4449 106054
rect 4505 106052 4529 106054
rect 4289 106032 4585 106052
rect 4289 105020 4585 105040
rect 4345 105018 4369 105020
rect 4425 105018 4449 105020
rect 4505 105018 4529 105020
rect 4367 104966 4369 105018
rect 4431 104966 4443 105018
rect 4505 104966 4507 105018
rect 4345 104964 4369 104966
rect 4425 104964 4449 104966
rect 4505 104964 4529 104966
rect 4289 104944 4585 104964
rect 4289 103932 4585 103952
rect 4345 103930 4369 103932
rect 4425 103930 4449 103932
rect 4505 103930 4529 103932
rect 4367 103878 4369 103930
rect 4431 103878 4443 103930
rect 4505 103878 4507 103930
rect 4345 103876 4369 103878
rect 4425 103876 4449 103878
rect 4505 103876 4529 103878
rect 4289 103856 4585 103876
rect 4289 102844 4585 102864
rect 4345 102842 4369 102844
rect 4425 102842 4449 102844
rect 4505 102842 4529 102844
rect 4367 102790 4369 102842
rect 4431 102790 4443 102842
rect 4505 102790 4507 102842
rect 4345 102788 4369 102790
rect 4425 102788 4449 102790
rect 4505 102788 4529 102790
rect 4289 102768 4585 102788
rect 4289 101756 4585 101776
rect 4345 101754 4369 101756
rect 4425 101754 4449 101756
rect 4505 101754 4529 101756
rect 4367 101702 4369 101754
rect 4431 101702 4443 101754
rect 4505 101702 4507 101754
rect 4345 101700 4369 101702
rect 4425 101700 4449 101702
rect 4505 101700 4529 101702
rect 4289 101680 4585 101700
rect 4289 100668 4585 100688
rect 4345 100666 4369 100668
rect 4425 100666 4449 100668
rect 4505 100666 4529 100668
rect 4367 100614 4369 100666
rect 4431 100614 4443 100666
rect 4505 100614 4507 100666
rect 4345 100612 4369 100614
rect 4425 100612 4449 100614
rect 4505 100612 4529 100614
rect 4289 100592 4585 100612
rect 4289 99580 4585 99600
rect 4345 99578 4369 99580
rect 4425 99578 4449 99580
rect 4505 99578 4529 99580
rect 4367 99526 4369 99578
rect 4431 99526 4443 99578
rect 4505 99526 4507 99578
rect 4345 99524 4369 99526
rect 4425 99524 4449 99526
rect 4505 99524 4529 99526
rect 4289 99504 4585 99524
rect 4289 98492 4585 98512
rect 4345 98490 4369 98492
rect 4425 98490 4449 98492
rect 4505 98490 4529 98492
rect 4367 98438 4369 98490
rect 4431 98438 4443 98490
rect 4505 98438 4507 98490
rect 4345 98436 4369 98438
rect 4425 98436 4449 98438
rect 4505 98436 4529 98438
rect 4289 98416 4585 98436
rect 4289 97404 4585 97424
rect 4345 97402 4369 97404
rect 4425 97402 4449 97404
rect 4505 97402 4529 97404
rect 4367 97350 4369 97402
rect 4431 97350 4443 97402
rect 4505 97350 4507 97402
rect 4345 97348 4369 97350
rect 4425 97348 4449 97350
rect 4505 97348 4529 97350
rect 4289 97328 4585 97348
rect 4289 96316 4585 96336
rect 4345 96314 4369 96316
rect 4425 96314 4449 96316
rect 4505 96314 4529 96316
rect 4367 96262 4369 96314
rect 4431 96262 4443 96314
rect 4505 96262 4507 96314
rect 4345 96260 4369 96262
rect 4425 96260 4449 96262
rect 4505 96260 4529 96262
rect 4289 96240 4585 96260
rect 4289 95228 4585 95248
rect 4345 95226 4369 95228
rect 4425 95226 4449 95228
rect 4505 95226 4529 95228
rect 4367 95174 4369 95226
rect 4431 95174 4443 95226
rect 4505 95174 4507 95226
rect 4345 95172 4369 95174
rect 4425 95172 4449 95174
rect 4505 95172 4529 95174
rect 4289 95152 4585 95172
rect 4289 94140 4585 94160
rect 4345 94138 4369 94140
rect 4425 94138 4449 94140
rect 4505 94138 4529 94140
rect 4367 94086 4369 94138
rect 4431 94086 4443 94138
rect 4505 94086 4507 94138
rect 4345 94084 4369 94086
rect 4425 94084 4449 94086
rect 4505 94084 4529 94086
rect 4289 94064 4585 94084
rect 4289 93052 4585 93072
rect 4345 93050 4369 93052
rect 4425 93050 4449 93052
rect 4505 93050 4529 93052
rect 4367 92998 4369 93050
rect 4431 92998 4443 93050
rect 4505 92998 4507 93050
rect 4345 92996 4369 92998
rect 4425 92996 4449 92998
rect 4505 92996 4529 92998
rect 4289 92976 4585 92996
rect 4289 91964 4585 91984
rect 4345 91962 4369 91964
rect 4425 91962 4449 91964
rect 4505 91962 4529 91964
rect 4367 91910 4369 91962
rect 4431 91910 4443 91962
rect 4505 91910 4507 91962
rect 4345 91908 4369 91910
rect 4425 91908 4449 91910
rect 4505 91908 4529 91910
rect 4289 91888 4585 91908
rect 4289 90876 4585 90896
rect 4345 90874 4369 90876
rect 4425 90874 4449 90876
rect 4505 90874 4529 90876
rect 4367 90822 4369 90874
rect 4431 90822 4443 90874
rect 4505 90822 4507 90874
rect 4345 90820 4369 90822
rect 4425 90820 4449 90822
rect 4505 90820 4529 90822
rect 4289 90800 4585 90820
rect 4289 89788 4585 89808
rect 4345 89786 4369 89788
rect 4425 89786 4449 89788
rect 4505 89786 4529 89788
rect 4367 89734 4369 89786
rect 4431 89734 4443 89786
rect 4505 89734 4507 89786
rect 4345 89732 4369 89734
rect 4425 89732 4449 89734
rect 4505 89732 4529 89734
rect 4289 89712 4585 89732
rect 4289 88700 4585 88720
rect 4345 88698 4369 88700
rect 4425 88698 4449 88700
rect 4505 88698 4529 88700
rect 4367 88646 4369 88698
rect 4431 88646 4443 88698
rect 4505 88646 4507 88698
rect 4345 88644 4369 88646
rect 4425 88644 4449 88646
rect 4505 88644 4529 88646
rect 4289 88624 4585 88644
rect 4289 87612 4585 87632
rect 4345 87610 4369 87612
rect 4425 87610 4449 87612
rect 4505 87610 4529 87612
rect 4367 87558 4369 87610
rect 4431 87558 4443 87610
rect 4505 87558 4507 87610
rect 4345 87556 4369 87558
rect 4425 87556 4449 87558
rect 4505 87556 4529 87558
rect 4289 87536 4585 87556
rect 4289 86524 4585 86544
rect 4345 86522 4369 86524
rect 4425 86522 4449 86524
rect 4505 86522 4529 86524
rect 4367 86470 4369 86522
rect 4431 86470 4443 86522
rect 4505 86470 4507 86522
rect 4345 86468 4369 86470
rect 4425 86468 4449 86470
rect 4505 86468 4529 86470
rect 4289 86448 4585 86468
rect 4289 85436 4585 85456
rect 4345 85434 4369 85436
rect 4425 85434 4449 85436
rect 4505 85434 4529 85436
rect 4367 85382 4369 85434
rect 4431 85382 4443 85434
rect 4505 85382 4507 85434
rect 4345 85380 4369 85382
rect 4425 85380 4449 85382
rect 4505 85380 4529 85382
rect 4289 85360 4585 85380
rect 4289 84348 4585 84368
rect 4345 84346 4369 84348
rect 4425 84346 4449 84348
rect 4505 84346 4529 84348
rect 4367 84294 4369 84346
rect 4431 84294 4443 84346
rect 4505 84294 4507 84346
rect 4345 84292 4369 84294
rect 4425 84292 4449 84294
rect 4505 84292 4529 84294
rect 4289 84272 4585 84292
rect 4289 83260 4585 83280
rect 4345 83258 4369 83260
rect 4425 83258 4449 83260
rect 4505 83258 4529 83260
rect 4367 83206 4369 83258
rect 4431 83206 4443 83258
rect 4505 83206 4507 83258
rect 4345 83204 4369 83206
rect 4425 83204 4449 83206
rect 4505 83204 4529 83206
rect 4289 83184 4585 83204
rect 4289 82172 4585 82192
rect 4345 82170 4369 82172
rect 4425 82170 4449 82172
rect 4505 82170 4529 82172
rect 4367 82118 4369 82170
rect 4431 82118 4443 82170
rect 4505 82118 4507 82170
rect 4345 82116 4369 82118
rect 4425 82116 4449 82118
rect 4505 82116 4529 82118
rect 4289 82096 4585 82116
rect 4289 81084 4585 81104
rect 4345 81082 4369 81084
rect 4425 81082 4449 81084
rect 4505 81082 4529 81084
rect 4367 81030 4369 81082
rect 4431 81030 4443 81082
rect 4505 81030 4507 81082
rect 4345 81028 4369 81030
rect 4425 81028 4449 81030
rect 4505 81028 4529 81030
rect 4289 81008 4585 81028
rect 4289 79996 4585 80016
rect 4345 79994 4369 79996
rect 4425 79994 4449 79996
rect 4505 79994 4529 79996
rect 4367 79942 4369 79994
rect 4431 79942 4443 79994
rect 4505 79942 4507 79994
rect 4345 79940 4369 79942
rect 4425 79940 4449 79942
rect 4505 79940 4529 79942
rect 4289 79920 4585 79940
rect 4289 78908 4585 78928
rect 4345 78906 4369 78908
rect 4425 78906 4449 78908
rect 4505 78906 4529 78908
rect 4367 78854 4369 78906
rect 4431 78854 4443 78906
rect 4505 78854 4507 78906
rect 4345 78852 4369 78854
rect 4425 78852 4449 78854
rect 4505 78852 4529 78854
rect 4289 78832 4585 78852
rect 4289 77820 4585 77840
rect 4345 77818 4369 77820
rect 4425 77818 4449 77820
rect 4505 77818 4529 77820
rect 4367 77766 4369 77818
rect 4431 77766 4443 77818
rect 4505 77766 4507 77818
rect 4345 77764 4369 77766
rect 4425 77764 4449 77766
rect 4505 77764 4529 77766
rect 4289 77744 4585 77764
rect 4289 76732 4585 76752
rect 4345 76730 4369 76732
rect 4425 76730 4449 76732
rect 4505 76730 4529 76732
rect 4367 76678 4369 76730
rect 4431 76678 4443 76730
rect 4505 76678 4507 76730
rect 4345 76676 4369 76678
rect 4425 76676 4449 76678
rect 4505 76676 4529 76678
rect 4289 76656 4585 76676
rect 4289 75644 4585 75664
rect 4345 75642 4369 75644
rect 4425 75642 4449 75644
rect 4505 75642 4529 75644
rect 4367 75590 4369 75642
rect 4431 75590 4443 75642
rect 4505 75590 4507 75642
rect 4345 75588 4369 75590
rect 4425 75588 4449 75590
rect 4505 75588 4529 75590
rect 4289 75568 4585 75588
rect 4289 74556 4585 74576
rect 4345 74554 4369 74556
rect 4425 74554 4449 74556
rect 4505 74554 4529 74556
rect 4367 74502 4369 74554
rect 4431 74502 4443 74554
rect 4505 74502 4507 74554
rect 4345 74500 4369 74502
rect 4425 74500 4449 74502
rect 4505 74500 4529 74502
rect 4289 74480 4585 74500
rect 4289 73468 4585 73488
rect 4345 73466 4369 73468
rect 4425 73466 4449 73468
rect 4505 73466 4529 73468
rect 4367 73414 4369 73466
rect 4431 73414 4443 73466
rect 4505 73414 4507 73466
rect 4345 73412 4369 73414
rect 4425 73412 4449 73414
rect 4505 73412 4529 73414
rect 4289 73392 4585 73412
rect 4289 72380 4585 72400
rect 4345 72378 4369 72380
rect 4425 72378 4449 72380
rect 4505 72378 4529 72380
rect 4367 72326 4369 72378
rect 4431 72326 4443 72378
rect 4505 72326 4507 72378
rect 4345 72324 4369 72326
rect 4425 72324 4449 72326
rect 4505 72324 4529 72326
rect 4289 72304 4585 72324
rect 4289 71292 4585 71312
rect 4345 71290 4369 71292
rect 4425 71290 4449 71292
rect 4505 71290 4529 71292
rect 4367 71238 4369 71290
rect 4431 71238 4443 71290
rect 4505 71238 4507 71290
rect 4345 71236 4369 71238
rect 4425 71236 4449 71238
rect 4505 71236 4529 71238
rect 4289 71216 4585 71236
rect 4289 70204 4585 70224
rect 4345 70202 4369 70204
rect 4425 70202 4449 70204
rect 4505 70202 4529 70204
rect 4367 70150 4369 70202
rect 4431 70150 4443 70202
rect 4505 70150 4507 70202
rect 4345 70148 4369 70150
rect 4425 70148 4449 70150
rect 4505 70148 4529 70150
rect 4289 70128 4585 70148
rect 4289 69116 4585 69136
rect 4345 69114 4369 69116
rect 4425 69114 4449 69116
rect 4505 69114 4529 69116
rect 4367 69062 4369 69114
rect 4431 69062 4443 69114
rect 4505 69062 4507 69114
rect 4345 69060 4369 69062
rect 4425 69060 4449 69062
rect 4505 69060 4529 69062
rect 4289 69040 4585 69060
rect 4289 68028 4585 68048
rect 4345 68026 4369 68028
rect 4425 68026 4449 68028
rect 4505 68026 4529 68028
rect 4367 67974 4369 68026
rect 4431 67974 4443 68026
rect 4505 67974 4507 68026
rect 4345 67972 4369 67974
rect 4425 67972 4449 67974
rect 4505 67972 4529 67974
rect 4289 67952 4585 67972
rect 4289 66940 4585 66960
rect 4345 66938 4369 66940
rect 4425 66938 4449 66940
rect 4505 66938 4529 66940
rect 4367 66886 4369 66938
rect 4431 66886 4443 66938
rect 4505 66886 4507 66938
rect 4345 66884 4369 66886
rect 4425 66884 4449 66886
rect 4505 66884 4529 66886
rect 4289 66864 4585 66884
rect 4289 65852 4585 65872
rect 4345 65850 4369 65852
rect 4425 65850 4449 65852
rect 4505 65850 4529 65852
rect 4367 65798 4369 65850
rect 4431 65798 4443 65850
rect 4505 65798 4507 65850
rect 4345 65796 4369 65798
rect 4425 65796 4449 65798
rect 4505 65796 4529 65798
rect 4289 65776 4585 65796
rect 4289 64764 4585 64784
rect 4345 64762 4369 64764
rect 4425 64762 4449 64764
rect 4505 64762 4529 64764
rect 4367 64710 4369 64762
rect 4431 64710 4443 64762
rect 4505 64710 4507 64762
rect 4345 64708 4369 64710
rect 4425 64708 4449 64710
rect 4505 64708 4529 64710
rect 4289 64688 4585 64708
rect 4289 63676 4585 63696
rect 4345 63674 4369 63676
rect 4425 63674 4449 63676
rect 4505 63674 4529 63676
rect 4367 63622 4369 63674
rect 4431 63622 4443 63674
rect 4505 63622 4507 63674
rect 4345 63620 4369 63622
rect 4425 63620 4449 63622
rect 4505 63620 4529 63622
rect 4289 63600 4585 63620
rect 4289 62588 4585 62608
rect 4345 62586 4369 62588
rect 4425 62586 4449 62588
rect 4505 62586 4529 62588
rect 4367 62534 4369 62586
rect 4431 62534 4443 62586
rect 4505 62534 4507 62586
rect 4345 62532 4369 62534
rect 4425 62532 4449 62534
rect 4505 62532 4529 62534
rect 4289 62512 4585 62532
rect 4289 61500 4585 61520
rect 4345 61498 4369 61500
rect 4425 61498 4449 61500
rect 4505 61498 4529 61500
rect 4367 61446 4369 61498
rect 4431 61446 4443 61498
rect 4505 61446 4507 61498
rect 4345 61444 4369 61446
rect 4425 61444 4449 61446
rect 4505 61444 4529 61446
rect 4289 61424 4585 61444
rect 4289 60412 4585 60432
rect 4345 60410 4369 60412
rect 4425 60410 4449 60412
rect 4505 60410 4529 60412
rect 4367 60358 4369 60410
rect 4431 60358 4443 60410
rect 4505 60358 4507 60410
rect 4345 60356 4369 60358
rect 4425 60356 4449 60358
rect 4505 60356 4529 60358
rect 4289 60336 4585 60356
rect 4289 59324 4585 59344
rect 4345 59322 4369 59324
rect 4425 59322 4449 59324
rect 4505 59322 4529 59324
rect 4367 59270 4369 59322
rect 4431 59270 4443 59322
rect 4505 59270 4507 59322
rect 4345 59268 4369 59270
rect 4425 59268 4449 59270
rect 4505 59268 4529 59270
rect 4289 59248 4585 59268
rect 4289 58236 4585 58256
rect 4345 58234 4369 58236
rect 4425 58234 4449 58236
rect 4505 58234 4529 58236
rect 4367 58182 4369 58234
rect 4431 58182 4443 58234
rect 4505 58182 4507 58234
rect 4345 58180 4369 58182
rect 4425 58180 4449 58182
rect 4505 58180 4529 58182
rect 4289 58160 4585 58180
rect 4289 57148 4585 57168
rect 4345 57146 4369 57148
rect 4425 57146 4449 57148
rect 4505 57146 4529 57148
rect 4367 57094 4369 57146
rect 4431 57094 4443 57146
rect 4505 57094 4507 57146
rect 4345 57092 4369 57094
rect 4425 57092 4449 57094
rect 4505 57092 4529 57094
rect 4289 57072 4585 57092
rect 4289 56060 4585 56080
rect 4345 56058 4369 56060
rect 4425 56058 4449 56060
rect 4505 56058 4529 56060
rect 4367 56006 4369 56058
rect 4431 56006 4443 56058
rect 4505 56006 4507 56058
rect 4345 56004 4369 56006
rect 4425 56004 4449 56006
rect 4505 56004 4529 56006
rect 4289 55984 4585 56004
rect 4289 54972 4585 54992
rect 4345 54970 4369 54972
rect 4425 54970 4449 54972
rect 4505 54970 4529 54972
rect 4367 54918 4369 54970
rect 4431 54918 4443 54970
rect 4505 54918 4507 54970
rect 4345 54916 4369 54918
rect 4425 54916 4449 54918
rect 4505 54916 4529 54918
rect 4289 54896 4585 54916
rect 4289 53884 4585 53904
rect 4345 53882 4369 53884
rect 4425 53882 4449 53884
rect 4505 53882 4529 53884
rect 4367 53830 4369 53882
rect 4431 53830 4443 53882
rect 4505 53830 4507 53882
rect 4345 53828 4369 53830
rect 4425 53828 4449 53830
rect 4505 53828 4529 53830
rect 4289 53808 4585 53828
rect 4289 52796 4585 52816
rect 4345 52794 4369 52796
rect 4425 52794 4449 52796
rect 4505 52794 4529 52796
rect 4367 52742 4369 52794
rect 4431 52742 4443 52794
rect 4505 52742 4507 52794
rect 4345 52740 4369 52742
rect 4425 52740 4449 52742
rect 4505 52740 4529 52742
rect 4289 52720 4585 52740
rect 4289 51708 4585 51728
rect 4345 51706 4369 51708
rect 4425 51706 4449 51708
rect 4505 51706 4529 51708
rect 4367 51654 4369 51706
rect 4431 51654 4443 51706
rect 4505 51654 4507 51706
rect 4345 51652 4369 51654
rect 4425 51652 4449 51654
rect 4505 51652 4529 51654
rect 4289 51632 4585 51652
rect 4289 50620 4585 50640
rect 4345 50618 4369 50620
rect 4425 50618 4449 50620
rect 4505 50618 4529 50620
rect 4367 50566 4369 50618
rect 4431 50566 4443 50618
rect 4505 50566 4507 50618
rect 4345 50564 4369 50566
rect 4425 50564 4449 50566
rect 4505 50564 4529 50566
rect 4289 50544 4585 50564
rect 4289 49532 4585 49552
rect 4345 49530 4369 49532
rect 4425 49530 4449 49532
rect 4505 49530 4529 49532
rect 4367 49478 4369 49530
rect 4431 49478 4443 49530
rect 4505 49478 4507 49530
rect 4345 49476 4369 49478
rect 4425 49476 4449 49478
rect 4505 49476 4529 49478
rect 4289 49456 4585 49476
rect 4289 48444 4585 48464
rect 4345 48442 4369 48444
rect 4425 48442 4449 48444
rect 4505 48442 4529 48444
rect 4367 48390 4369 48442
rect 4431 48390 4443 48442
rect 4505 48390 4507 48442
rect 4345 48388 4369 48390
rect 4425 48388 4449 48390
rect 4505 48388 4529 48390
rect 4289 48368 4585 48388
rect 4289 47356 4585 47376
rect 4345 47354 4369 47356
rect 4425 47354 4449 47356
rect 4505 47354 4529 47356
rect 4367 47302 4369 47354
rect 4431 47302 4443 47354
rect 4505 47302 4507 47354
rect 4345 47300 4369 47302
rect 4425 47300 4449 47302
rect 4505 47300 4529 47302
rect 4289 47280 4585 47300
rect 4289 46268 4585 46288
rect 4345 46266 4369 46268
rect 4425 46266 4449 46268
rect 4505 46266 4529 46268
rect 4367 46214 4369 46266
rect 4431 46214 4443 46266
rect 4505 46214 4507 46266
rect 4345 46212 4369 46214
rect 4425 46212 4449 46214
rect 4505 46212 4529 46214
rect 4289 46192 4585 46212
rect 4289 45180 4585 45200
rect 4345 45178 4369 45180
rect 4425 45178 4449 45180
rect 4505 45178 4529 45180
rect 4367 45126 4369 45178
rect 4431 45126 4443 45178
rect 4505 45126 4507 45178
rect 4345 45124 4369 45126
rect 4425 45124 4449 45126
rect 4505 45124 4529 45126
rect 4289 45104 4585 45124
rect 4289 44092 4585 44112
rect 4345 44090 4369 44092
rect 4425 44090 4449 44092
rect 4505 44090 4529 44092
rect 4367 44038 4369 44090
rect 4431 44038 4443 44090
rect 4505 44038 4507 44090
rect 4345 44036 4369 44038
rect 4425 44036 4449 44038
rect 4505 44036 4529 44038
rect 4289 44016 4585 44036
rect 4289 43004 4585 43024
rect 4345 43002 4369 43004
rect 4425 43002 4449 43004
rect 4505 43002 4529 43004
rect 4367 42950 4369 43002
rect 4431 42950 4443 43002
rect 4505 42950 4507 43002
rect 4345 42948 4369 42950
rect 4425 42948 4449 42950
rect 4505 42948 4529 42950
rect 4289 42928 4585 42948
rect 4289 41916 4585 41936
rect 4345 41914 4369 41916
rect 4425 41914 4449 41916
rect 4505 41914 4529 41916
rect 4367 41862 4369 41914
rect 4431 41862 4443 41914
rect 4505 41862 4507 41914
rect 4345 41860 4369 41862
rect 4425 41860 4449 41862
rect 4505 41860 4529 41862
rect 4289 41840 4585 41860
rect 4289 40828 4585 40848
rect 4345 40826 4369 40828
rect 4425 40826 4449 40828
rect 4505 40826 4529 40828
rect 4367 40774 4369 40826
rect 4431 40774 4443 40826
rect 4505 40774 4507 40826
rect 4345 40772 4369 40774
rect 4425 40772 4449 40774
rect 4505 40772 4529 40774
rect 4289 40752 4585 40772
rect 4289 39740 4585 39760
rect 4345 39738 4369 39740
rect 4425 39738 4449 39740
rect 4505 39738 4529 39740
rect 4367 39686 4369 39738
rect 4431 39686 4443 39738
rect 4505 39686 4507 39738
rect 4345 39684 4369 39686
rect 4425 39684 4449 39686
rect 4505 39684 4529 39686
rect 4289 39664 4585 39684
rect 4289 38652 4585 38672
rect 4345 38650 4369 38652
rect 4425 38650 4449 38652
rect 4505 38650 4529 38652
rect 4367 38598 4369 38650
rect 4431 38598 4443 38650
rect 4505 38598 4507 38650
rect 4345 38596 4369 38598
rect 4425 38596 4449 38598
rect 4505 38596 4529 38598
rect 4289 38576 4585 38596
rect 4289 37564 4585 37584
rect 4345 37562 4369 37564
rect 4425 37562 4449 37564
rect 4505 37562 4529 37564
rect 4367 37510 4369 37562
rect 4431 37510 4443 37562
rect 4505 37510 4507 37562
rect 4345 37508 4369 37510
rect 4425 37508 4449 37510
rect 4505 37508 4529 37510
rect 4289 37488 4585 37508
rect 4289 36476 4585 36496
rect 4345 36474 4369 36476
rect 4425 36474 4449 36476
rect 4505 36474 4529 36476
rect 4367 36422 4369 36474
rect 4431 36422 4443 36474
rect 4505 36422 4507 36474
rect 4345 36420 4369 36422
rect 4425 36420 4449 36422
rect 4505 36420 4529 36422
rect 4289 36400 4585 36420
rect 4289 35388 4585 35408
rect 4345 35386 4369 35388
rect 4425 35386 4449 35388
rect 4505 35386 4529 35388
rect 4367 35334 4369 35386
rect 4431 35334 4443 35386
rect 4505 35334 4507 35386
rect 4345 35332 4369 35334
rect 4425 35332 4449 35334
rect 4505 35332 4529 35334
rect 4289 35312 4585 35332
rect 4289 34300 4585 34320
rect 4345 34298 4369 34300
rect 4425 34298 4449 34300
rect 4505 34298 4529 34300
rect 4367 34246 4369 34298
rect 4431 34246 4443 34298
rect 4505 34246 4507 34298
rect 4345 34244 4369 34246
rect 4425 34244 4449 34246
rect 4505 34244 4529 34246
rect 4289 34224 4585 34244
rect 4289 33212 4585 33232
rect 4345 33210 4369 33212
rect 4425 33210 4449 33212
rect 4505 33210 4529 33212
rect 4367 33158 4369 33210
rect 4431 33158 4443 33210
rect 4505 33158 4507 33210
rect 4345 33156 4369 33158
rect 4425 33156 4449 33158
rect 4505 33156 4529 33158
rect 4289 33136 4585 33156
rect 4289 32124 4585 32144
rect 4345 32122 4369 32124
rect 4425 32122 4449 32124
rect 4505 32122 4529 32124
rect 4367 32070 4369 32122
rect 4431 32070 4443 32122
rect 4505 32070 4507 32122
rect 4345 32068 4369 32070
rect 4425 32068 4449 32070
rect 4505 32068 4529 32070
rect 4289 32048 4585 32068
rect 4289 31036 4585 31056
rect 4345 31034 4369 31036
rect 4425 31034 4449 31036
rect 4505 31034 4529 31036
rect 4367 30982 4369 31034
rect 4431 30982 4443 31034
rect 4505 30982 4507 31034
rect 4345 30980 4369 30982
rect 4425 30980 4449 30982
rect 4505 30980 4529 30982
rect 4289 30960 4585 30980
rect 4289 29948 4585 29968
rect 4345 29946 4369 29948
rect 4425 29946 4449 29948
rect 4505 29946 4529 29948
rect 4367 29894 4369 29946
rect 4431 29894 4443 29946
rect 4505 29894 4507 29946
rect 4345 29892 4369 29894
rect 4425 29892 4449 29894
rect 4505 29892 4529 29894
rect 4289 29872 4585 29892
rect 4289 28860 4585 28880
rect 4345 28858 4369 28860
rect 4425 28858 4449 28860
rect 4505 28858 4529 28860
rect 4367 28806 4369 28858
rect 4431 28806 4443 28858
rect 4505 28806 4507 28858
rect 4345 28804 4369 28806
rect 4425 28804 4449 28806
rect 4505 28804 4529 28806
rect 4289 28784 4585 28804
rect 4289 27772 4585 27792
rect 4345 27770 4369 27772
rect 4425 27770 4449 27772
rect 4505 27770 4529 27772
rect 4367 27718 4369 27770
rect 4431 27718 4443 27770
rect 4505 27718 4507 27770
rect 4345 27716 4369 27718
rect 4425 27716 4449 27718
rect 4505 27716 4529 27718
rect 4289 27696 4585 27716
rect 4289 26684 4585 26704
rect 4345 26682 4369 26684
rect 4425 26682 4449 26684
rect 4505 26682 4529 26684
rect 4367 26630 4369 26682
rect 4431 26630 4443 26682
rect 4505 26630 4507 26682
rect 4345 26628 4369 26630
rect 4425 26628 4449 26630
rect 4505 26628 4529 26630
rect 4289 26608 4585 26628
rect 4289 25596 4585 25616
rect 4345 25594 4369 25596
rect 4425 25594 4449 25596
rect 4505 25594 4529 25596
rect 4367 25542 4369 25594
rect 4431 25542 4443 25594
rect 4505 25542 4507 25594
rect 4345 25540 4369 25542
rect 4425 25540 4449 25542
rect 4505 25540 4529 25542
rect 4289 25520 4585 25540
rect 4289 24508 4585 24528
rect 4345 24506 4369 24508
rect 4425 24506 4449 24508
rect 4505 24506 4529 24508
rect 4367 24454 4369 24506
rect 4431 24454 4443 24506
rect 4505 24454 4507 24506
rect 4345 24452 4369 24454
rect 4425 24452 4449 24454
rect 4505 24452 4529 24454
rect 4289 24432 4585 24452
rect 3790 24304 3846 24313
rect 3790 24239 3846 24248
rect 4289 23420 4585 23440
rect 4345 23418 4369 23420
rect 4425 23418 4449 23420
rect 4505 23418 4529 23420
rect 4367 23366 4369 23418
rect 4431 23366 4443 23418
rect 4505 23366 4507 23418
rect 4345 23364 4369 23366
rect 4425 23364 4449 23366
rect 4505 23364 4529 23366
rect 4289 23344 4585 23364
rect 4289 22332 4585 22352
rect 4345 22330 4369 22332
rect 4425 22330 4449 22332
rect 4505 22330 4529 22332
rect 4367 22278 4369 22330
rect 4431 22278 4443 22330
rect 4505 22278 4507 22330
rect 4345 22276 4369 22278
rect 4425 22276 4449 22278
rect 4505 22276 4529 22278
rect 4289 22256 4585 22276
rect 4289 21244 4585 21264
rect 4345 21242 4369 21244
rect 4425 21242 4449 21244
rect 4505 21242 4529 21244
rect 4367 21190 4369 21242
rect 4431 21190 4443 21242
rect 4505 21190 4507 21242
rect 4345 21188 4369 21190
rect 4425 21188 4449 21190
rect 4505 21188 4529 21190
rect 4289 21168 4585 21188
rect 4289 20156 4585 20176
rect 4345 20154 4369 20156
rect 4425 20154 4449 20156
rect 4505 20154 4529 20156
rect 4367 20102 4369 20154
rect 4431 20102 4443 20154
rect 4505 20102 4507 20154
rect 4345 20100 4369 20102
rect 4425 20100 4449 20102
rect 4505 20100 4529 20102
rect 4289 20080 4585 20100
rect 4289 19068 4585 19088
rect 4345 19066 4369 19068
rect 4425 19066 4449 19068
rect 4505 19066 4529 19068
rect 4367 19014 4369 19066
rect 4431 19014 4443 19066
rect 4505 19014 4507 19066
rect 4345 19012 4369 19014
rect 4425 19012 4449 19014
rect 4505 19012 4529 19014
rect 4289 18992 4585 19012
rect 4289 17980 4585 18000
rect 4345 17978 4369 17980
rect 4425 17978 4449 17980
rect 4505 17978 4529 17980
rect 4367 17926 4369 17978
rect 4431 17926 4443 17978
rect 4505 17926 4507 17978
rect 4345 17924 4369 17926
rect 4425 17924 4449 17926
rect 4505 17924 4529 17926
rect 4289 17904 4585 17924
rect 4816 17241 4844 228006
rect 5356 225344 5408 225350
rect 5356 225286 5408 225292
rect 5368 224398 5396 225286
rect 5460 224466 5488 332522
rect 5538 332520 5594 332574
rect 5644 322934 5672 332574
rect 6748 332574 6882 332602
rect 5956 330780 6252 330800
rect 6012 330778 6036 330780
rect 6092 330778 6116 330780
rect 6172 330778 6196 330780
rect 6034 330726 6036 330778
rect 6098 330726 6110 330778
rect 6172 330726 6174 330778
rect 6012 330724 6036 330726
rect 6092 330724 6116 330726
rect 6172 330724 6196 330726
rect 5956 330704 6252 330724
rect 5956 329692 6252 329712
rect 6012 329690 6036 329692
rect 6092 329690 6116 329692
rect 6172 329690 6196 329692
rect 6034 329638 6036 329690
rect 6098 329638 6110 329690
rect 6172 329638 6174 329690
rect 6012 329636 6036 329638
rect 6092 329636 6116 329638
rect 6172 329636 6196 329638
rect 5956 329616 6252 329636
rect 5956 328604 6252 328624
rect 6012 328602 6036 328604
rect 6092 328602 6116 328604
rect 6172 328602 6196 328604
rect 6034 328550 6036 328602
rect 6098 328550 6110 328602
rect 6172 328550 6174 328602
rect 6012 328548 6036 328550
rect 6092 328548 6116 328550
rect 6172 328548 6196 328550
rect 5956 328528 6252 328548
rect 5956 327516 6252 327536
rect 6012 327514 6036 327516
rect 6092 327514 6116 327516
rect 6172 327514 6196 327516
rect 6034 327462 6036 327514
rect 6098 327462 6110 327514
rect 6172 327462 6174 327514
rect 6012 327460 6036 327462
rect 6092 327460 6116 327462
rect 6172 327460 6196 327462
rect 5956 327440 6252 327460
rect 5956 326428 6252 326448
rect 6012 326426 6036 326428
rect 6092 326426 6116 326428
rect 6172 326426 6196 326428
rect 6034 326374 6036 326426
rect 6098 326374 6110 326426
rect 6172 326374 6174 326426
rect 6012 326372 6036 326374
rect 6092 326372 6116 326374
rect 6172 326372 6196 326374
rect 5956 326352 6252 326372
rect 5956 325340 6252 325360
rect 6012 325338 6036 325340
rect 6092 325338 6116 325340
rect 6172 325338 6196 325340
rect 6034 325286 6036 325338
rect 6098 325286 6110 325338
rect 6172 325286 6174 325338
rect 6012 325284 6036 325286
rect 6092 325284 6116 325286
rect 6172 325284 6196 325286
rect 5956 325264 6252 325284
rect 5956 324252 6252 324272
rect 6012 324250 6036 324252
rect 6092 324250 6116 324252
rect 6172 324250 6196 324252
rect 6034 324198 6036 324250
rect 6098 324198 6110 324250
rect 6172 324198 6174 324250
rect 6012 324196 6036 324198
rect 6092 324196 6116 324198
rect 6172 324196 6196 324198
rect 5956 324176 6252 324196
rect 5956 323164 6252 323184
rect 6012 323162 6036 323164
rect 6092 323162 6116 323164
rect 6172 323162 6196 323164
rect 6034 323110 6036 323162
rect 6098 323110 6110 323162
rect 6172 323110 6174 323162
rect 6012 323108 6036 323110
rect 6092 323108 6116 323110
rect 6172 323108 6196 323110
rect 5956 323088 6252 323108
rect 5552 322906 5672 322934
rect 5552 233646 5580 322906
rect 5956 322076 6252 322096
rect 6012 322074 6036 322076
rect 6092 322074 6116 322076
rect 6172 322074 6196 322076
rect 6034 322022 6036 322074
rect 6098 322022 6110 322074
rect 6172 322022 6174 322074
rect 6012 322020 6036 322022
rect 6092 322020 6116 322022
rect 6172 322020 6196 322022
rect 5956 322000 6252 322020
rect 5956 320988 6252 321008
rect 6012 320986 6036 320988
rect 6092 320986 6116 320988
rect 6172 320986 6196 320988
rect 6034 320934 6036 320986
rect 6098 320934 6110 320986
rect 6172 320934 6174 320986
rect 6012 320932 6036 320934
rect 6092 320932 6116 320934
rect 6172 320932 6196 320934
rect 5956 320912 6252 320932
rect 5956 319900 6252 319920
rect 6012 319898 6036 319900
rect 6092 319898 6116 319900
rect 6172 319898 6196 319900
rect 6034 319846 6036 319898
rect 6098 319846 6110 319898
rect 6172 319846 6174 319898
rect 6012 319844 6036 319846
rect 6092 319844 6116 319846
rect 6172 319844 6196 319846
rect 5956 319824 6252 319844
rect 5956 318812 6252 318832
rect 6012 318810 6036 318812
rect 6092 318810 6116 318812
rect 6172 318810 6196 318812
rect 6034 318758 6036 318810
rect 6098 318758 6110 318810
rect 6172 318758 6174 318810
rect 6012 318756 6036 318758
rect 6092 318756 6116 318758
rect 6172 318756 6196 318758
rect 5956 318736 6252 318756
rect 5956 317724 6252 317744
rect 6012 317722 6036 317724
rect 6092 317722 6116 317724
rect 6172 317722 6196 317724
rect 6034 317670 6036 317722
rect 6098 317670 6110 317722
rect 6172 317670 6174 317722
rect 6012 317668 6036 317670
rect 6092 317668 6116 317670
rect 6172 317668 6196 317670
rect 5956 317648 6252 317668
rect 5956 316636 6252 316656
rect 6012 316634 6036 316636
rect 6092 316634 6116 316636
rect 6172 316634 6196 316636
rect 6034 316582 6036 316634
rect 6098 316582 6110 316634
rect 6172 316582 6174 316634
rect 6012 316580 6036 316582
rect 6092 316580 6116 316582
rect 6172 316580 6196 316582
rect 5956 316560 6252 316580
rect 5956 315548 6252 315568
rect 6012 315546 6036 315548
rect 6092 315546 6116 315548
rect 6172 315546 6196 315548
rect 6034 315494 6036 315546
rect 6098 315494 6110 315546
rect 6172 315494 6174 315546
rect 6012 315492 6036 315494
rect 6092 315492 6116 315494
rect 6172 315492 6196 315494
rect 5956 315472 6252 315492
rect 5956 314460 6252 314480
rect 6012 314458 6036 314460
rect 6092 314458 6116 314460
rect 6172 314458 6196 314460
rect 6034 314406 6036 314458
rect 6098 314406 6110 314458
rect 6172 314406 6174 314458
rect 6012 314404 6036 314406
rect 6092 314404 6116 314406
rect 6172 314404 6196 314406
rect 5956 314384 6252 314404
rect 5956 313372 6252 313392
rect 6012 313370 6036 313372
rect 6092 313370 6116 313372
rect 6172 313370 6196 313372
rect 6034 313318 6036 313370
rect 6098 313318 6110 313370
rect 6172 313318 6174 313370
rect 6012 313316 6036 313318
rect 6092 313316 6116 313318
rect 6172 313316 6196 313318
rect 5956 313296 6252 313316
rect 5956 312284 6252 312304
rect 6012 312282 6036 312284
rect 6092 312282 6116 312284
rect 6172 312282 6196 312284
rect 6034 312230 6036 312282
rect 6098 312230 6110 312282
rect 6172 312230 6174 312282
rect 6012 312228 6036 312230
rect 6092 312228 6116 312230
rect 6172 312228 6196 312230
rect 5956 312208 6252 312228
rect 5956 311196 6252 311216
rect 6012 311194 6036 311196
rect 6092 311194 6116 311196
rect 6172 311194 6196 311196
rect 6034 311142 6036 311194
rect 6098 311142 6110 311194
rect 6172 311142 6174 311194
rect 6012 311140 6036 311142
rect 6092 311140 6116 311142
rect 6172 311140 6196 311142
rect 5956 311120 6252 311140
rect 5956 310108 6252 310128
rect 6012 310106 6036 310108
rect 6092 310106 6116 310108
rect 6172 310106 6196 310108
rect 6034 310054 6036 310106
rect 6098 310054 6110 310106
rect 6172 310054 6174 310106
rect 6012 310052 6036 310054
rect 6092 310052 6116 310054
rect 6172 310052 6196 310054
rect 5956 310032 6252 310052
rect 5956 309020 6252 309040
rect 6012 309018 6036 309020
rect 6092 309018 6116 309020
rect 6172 309018 6196 309020
rect 6034 308966 6036 309018
rect 6098 308966 6110 309018
rect 6172 308966 6174 309018
rect 6012 308964 6036 308966
rect 6092 308964 6116 308966
rect 6172 308964 6196 308966
rect 5956 308944 6252 308964
rect 5956 307932 6252 307952
rect 6012 307930 6036 307932
rect 6092 307930 6116 307932
rect 6172 307930 6196 307932
rect 6034 307878 6036 307930
rect 6098 307878 6110 307930
rect 6172 307878 6174 307930
rect 6012 307876 6036 307878
rect 6092 307876 6116 307878
rect 6172 307876 6196 307878
rect 5956 307856 6252 307876
rect 5956 306844 6252 306864
rect 6012 306842 6036 306844
rect 6092 306842 6116 306844
rect 6172 306842 6196 306844
rect 6034 306790 6036 306842
rect 6098 306790 6110 306842
rect 6172 306790 6174 306842
rect 6012 306788 6036 306790
rect 6092 306788 6116 306790
rect 6172 306788 6196 306790
rect 5956 306768 6252 306788
rect 5956 305756 6252 305776
rect 6012 305754 6036 305756
rect 6092 305754 6116 305756
rect 6172 305754 6196 305756
rect 6034 305702 6036 305754
rect 6098 305702 6110 305754
rect 6172 305702 6174 305754
rect 6012 305700 6036 305702
rect 6092 305700 6116 305702
rect 6172 305700 6196 305702
rect 5956 305680 6252 305700
rect 5956 304668 6252 304688
rect 6012 304666 6036 304668
rect 6092 304666 6116 304668
rect 6172 304666 6196 304668
rect 6034 304614 6036 304666
rect 6098 304614 6110 304666
rect 6172 304614 6174 304666
rect 6012 304612 6036 304614
rect 6092 304612 6116 304614
rect 6172 304612 6196 304614
rect 5956 304592 6252 304612
rect 5956 303580 6252 303600
rect 6012 303578 6036 303580
rect 6092 303578 6116 303580
rect 6172 303578 6196 303580
rect 6034 303526 6036 303578
rect 6098 303526 6110 303578
rect 6172 303526 6174 303578
rect 6012 303524 6036 303526
rect 6092 303524 6116 303526
rect 6172 303524 6196 303526
rect 5956 303504 6252 303524
rect 5956 302492 6252 302512
rect 6012 302490 6036 302492
rect 6092 302490 6116 302492
rect 6172 302490 6196 302492
rect 6034 302438 6036 302490
rect 6098 302438 6110 302490
rect 6172 302438 6174 302490
rect 6012 302436 6036 302438
rect 6092 302436 6116 302438
rect 6172 302436 6196 302438
rect 5956 302416 6252 302436
rect 5956 301404 6252 301424
rect 6012 301402 6036 301404
rect 6092 301402 6116 301404
rect 6172 301402 6196 301404
rect 6034 301350 6036 301402
rect 6098 301350 6110 301402
rect 6172 301350 6174 301402
rect 6012 301348 6036 301350
rect 6092 301348 6116 301350
rect 6172 301348 6196 301350
rect 5956 301328 6252 301348
rect 5956 300316 6252 300336
rect 6012 300314 6036 300316
rect 6092 300314 6116 300316
rect 6172 300314 6196 300316
rect 6034 300262 6036 300314
rect 6098 300262 6110 300314
rect 6172 300262 6174 300314
rect 6012 300260 6036 300262
rect 6092 300260 6116 300262
rect 6172 300260 6196 300262
rect 5956 300240 6252 300260
rect 5956 299228 6252 299248
rect 6012 299226 6036 299228
rect 6092 299226 6116 299228
rect 6172 299226 6196 299228
rect 6034 299174 6036 299226
rect 6098 299174 6110 299226
rect 6172 299174 6174 299226
rect 6012 299172 6036 299174
rect 6092 299172 6116 299174
rect 6172 299172 6196 299174
rect 5956 299152 6252 299172
rect 5956 298140 6252 298160
rect 6012 298138 6036 298140
rect 6092 298138 6116 298140
rect 6172 298138 6196 298140
rect 6034 298086 6036 298138
rect 6098 298086 6110 298138
rect 6172 298086 6174 298138
rect 6012 298084 6036 298086
rect 6092 298084 6116 298086
rect 6172 298084 6196 298086
rect 5956 298064 6252 298084
rect 5956 297052 6252 297072
rect 6012 297050 6036 297052
rect 6092 297050 6116 297052
rect 6172 297050 6196 297052
rect 6034 296998 6036 297050
rect 6098 296998 6110 297050
rect 6172 296998 6174 297050
rect 6012 296996 6036 296998
rect 6092 296996 6116 296998
rect 6172 296996 6196 296998
rect 5956 296976 6252 296996
rect 5956 295964 6252 295984
rect 6012 295962 6036 295964
rect 6092 295962 6116 295964
rect 6172 295962 6196 295964
rect 6034 295910 6036 295962
rect 6098 295910 6110 295962
rect 6172 295910 6174 295962
rect 6012 295908 6036 295910
rect 6092 295908 6116 295910
rect 6172 295908 6196 295910
rect 5956 295888 6252 295908
rect 5956 294876 6252 294896
rect 6012 294874 6036 294876
rect 6092 294874 6116 294876
rect 6172 294874 6196 294876
rect 6034 294822 6036 294874
rect 6098 294822 6110 294874
rect 6172 294822 6174 294874
rect 6012 294820 6036 294822
rect 6092 294820 6116 294822
rect 6172 294820 6196 294822
rect 5956 294800 6252 294820
rect 5956 293788 6252 293808
rect 6012 293786 6036 293788
rect 6092 293786 6116 293788
rect 6172 293786 6196 293788
rect 6034 293734 6036 293786
rect 6098 293734 6110 293786
rect 6172 293734 6174 293786
rect 6012 293732 6036 293734
rect 6092 293732 6116 293734
rect 6172 293732 6196 293734
rect 5956 293712 6252 293732
rect 5956 292700 6252 292720
rect 6012 292698 6036 292700
rect 6092 292698 6116 292700
rect 6172 292698 6196 292700
rect 6034 292646 6036 292698
rect 6098 292646 6110 292698
rect 6172 292646 6174 292698
rect 6012 292644 6036 292646
rect 6092 292644 6116 292646
rect 6172 292644 6196 292646
rect 5956 292624 6252 292644
rect 5956 291612 6252 291632
rect 6012 291610 6036 291612
rect 6092 291610 6116 291612
rect 6172 291610 6196 291612
rect 6034 291558 6036 291610
rect 6098 291558 6110 291610
rect 6172 291558 6174 291610
rect 6012 291556 6036 291558
rect 6092 291556 6116 291558
rect 6172 291556 6196 291558
rect 5956 291536 6252 291556
rect 5956 290524 6252 290544
rect 6012 290522 6036 290524
rect 6092 290522 6116 290524
rect 6172 290522 6196 290524
rect 6034 290470 6036 290522
rect 6098 290470 6110 290522
rect 6172 290470 6174 290522
rect 6012 290468 6036 290470
rect 6092 290468 6116 290470
rect 6172 290468 6196 290470
rect 5956 290448 6252 290468
rect 5956 289436 6252 289456
rect 6012 289434 6036 289436
rect 6092 289434 6116 289436
rect 6172 289434 6196 289436
rect 6034 289382 6036 289434
rect 6098 289382 6110 289434
rect 6172 289382 6174 289434
rect 6012 289380 6036 289382
rect 6092 289380 6116 289382
rect 6172 289380 6196 289382
rect 5956 289360 6252 289380
rect 5956 288348 6252 288368
rect 6012 288346 6036 288348
rect 6092 288346 6116 288348
rect 6172 288346 6196 288348
rect 6034 288294 6036 288346
rect 6098 288294 6110 288346
rect 6172 288294 6174 288346
rect 6012 288292 6036 288294
rect 6092 288292 6116 288294
rect 6172 288292 6196 288294
rect 5956 288272 6252 288292
rect 5956 287260 6252 287280
rect 6012 287258 6036 287260
rect 6092 287258 6116 287260
rect 6172 287258 6196 287260
rect 6034 287206 6036 287258
rect 6098 287206 6110 287258
rect 6172 287206 6174 287258
rect 6012 287204 6036 287206
rect 6092 287204 6116 287206
rect 6172 287204 6196 287206
rect 5956 287184 6252 287204
rect 5956 286172 6252 286192
rect 6012 286170 6036 286172
rect 6092 286170 6116 286172
rect 6172 286170 6196 286172
rect 6034 286118 6036 286170
rect 6098 286118 6110 286170
rect 6172 286118 6174 286170
rect 6012 286116 6036 286118
rect 6092 286116 6116 286118
rect 6172 286116 6196 286118
rect 5956 286096 6252 286116
rect 5956 285084 6252 285104
rect 6012 285082 6036 285084
rect 6092 285082 6116 285084
rect 6172 285082 6196 285084
rect 6034 285030 6036 285082
rect 6098 285030 6110 285082
rect 6172 285030 6174 285082
rect 6012 285028 6036 285030
rect 6092 285028 6116 285030
rect 6172 285028 6196 285030
rect 5956 285008 6252 285028
rect 5956 283996 6252 284016
rect 6012 283994 6036 283996
rect 6092 283994 6116 283996
rect 6172 283994 6196 283996
rect 6034 283942 6036 283994
rect 6098 283942 6110 283994
rect 6172 283942 6174 283994
rect 6012 283940 6036 283942
rect 6092 283940 6116 283942
rect 6172 283940 6196 283942
rect 5956 283920 6252 283940
rect 5956 282908 6252 282928
rect 6012 282906 6036 282908
rect 6092 282906 6116 282908
rect 6172 282906 6196 282908
rect 6034 282854 6036 282906
rect 6098 282854 6110 282906
rect 6172 282854 6174 282906
rect 6012 282852 6036 282854
rect 6092 282852 6116 282854
rect 6172 282852 6196 282854
rect 5956 282832 6252 282852
rect 6274 282568 6330 282577
rect 6274 282503 6330 282512
rect 5956 281820 6252 281840
rect 6012 281818 6036 281820
rect 6092 281818 6116 281820
rect 6172 281818 6196 281820
rect 6034 281766 6036 281818
rect 6098 281766 6110 281818
rect 6172 281766 6174 281818
rect 6012 281764 6036 281766
rect 6092 281764 6116 281766
rect 6172 281764 6196 281766
rect 5956 281744 6252 281764
rect 5956 280732 6252 280752
rect 6012 280730 6036 280732
rect 6092 280730 6116 280732
rect 6172 280730 6196 280732
rect 6034 280678 6036 280730
rect 6098 280678 6110 280730
rect 6172 280678 6174 280730
rect 6012 280676 6036 280678
rect 6092 280676 6116 280678
rect 6172 280676 6196 280678
rect 5956 280656 6252 280676
rect 5956 279644 6252 279664
rect 6012 279642 6036 279644
rect 6092 279642 6116 279644
rect 6172 279642 6196 279644
rect 6034 279590 6036 279642
rect 6098 279590 6110 279642
rect 6172 279590 6174 279642
rect 6012 279588 6036 279590
rect 6092 279588 6116 279590
rect 6172 279588 6196 279590
rect 5956 279568 6252 279588
rect 5956 278556 6252 278576
rect 6012 278554 6036 278556
rect 6092 278554 6116 278556
rect 6172 278554 6196 278556
rect 6034 278502 6036 278554
rect 6098 278502 6110 278554
rect 6172 278502 6174 278554
rect 6012 278500 6036 278502
rect 6092 278500 6116 278502
rect 6172 278500 6196 278502
rect 5956 278480 6252 278500
rect 5956 277468 6252 277488
rect 6012 277466 6036 277468
rect 6092 277466 6116 277468
rect 6172 277466 6196 277468
rect 6034 277414 6036 277466
rect 6098 277414 6110 277466
rect 6172 277414 6174 277466
rect 6012 277412 6036 277414
rect 6092 277412 6116 277414
rect 6172 277412 6196 277414
rect 5956 277392 6252 277412
rect 5956 276380 6252 276400
rect 6012 276378 6036 276380
rect 6092 276378 6116 276380
rect 6172 276378 6196 276380
rect 6034 276326 6036 276378
rect 6098 276326 6110 276378
rect 6172 276326 6174 276378
rect 6012 276324 6036 276326
rect 6092 276324 6116 276326
rect 6172 276324 6196 276326
rect 5956 276304 6252 276324
rect 5956 275292 6252 275312
rect 6012 275290 6036 275292
rect 6092 275290 6116 275292
rect 6172 275290 6196 275292
rect 6034 275238 6036 275290
rect 6098 275238 6110 275290
rect 6172 275238 6174 275290
rect 6012 275236 6036 275238
rect 6092 275236 6116 275238
rect 6172 275236 6196 275238
rect 5956 275216 6252 275236
rect 5956 274204 6252 274224
rect 6012 274202 6036 274204
rect 6092 274202 6116 274204
rect 6172 274202 6196 274204
rect 6034 274150 6036 274202
rect 6098 274150 6110 274202
rect 6172 274150 6174 274202
rect 6012 274148 6036 274150
rect 6092 274148 6116 274150
rect 6172 274148 6196 274150
rect 5956 274128 6252 274148
rect 5956 273116 6252 273136
rect 6012 273114 6036 273116
rect 6092 273114 6116 273116
rect 6172 273114 6196 273116
rect 6034 273062 6036 273114
rect 6098 273062 6110 273114
rect 6172 273062 6174 273114
rect 6012 273060 6036 273062
rect 6092 273060 6116 273062
rect 6172 273060 6196 273062
rect 5956 273040 6252 273060
rect 5956 272028 6252 272048
rect 6012 272026 6036 272028
rect 6092 272026 6116 272028
rect 6172 272026 6196 272028
rect 6034 271974 6036 272026
rect 6098 271974 6110 272026
rect 6172 271974 6174 272026
rect 6012 271972 6036 271974
rect 6092 271972 6116 271974
rect 6172 271972 6196 271974
rect 5956 271952 6252 271972
rect 5956 270940 6252 270960
rect 6012 270938 6036 270940
rect 6092 270938 6116 270940
rect 6172 270938 6196 270940
rect 6034 270886 6036 270938
rect 6098 270886 6110 270938
rect 6172 270886 6174 270938
rect 6012 270884 6036 270886
rect 6092 270884 6116 270886
rect 6172 270884 6196 270886
rect 5956 270864 6252 270884
rect 5956 269852 6252 269872
rect 6012 269850 6036 269852
rect 6092 269850 6116 269852
rect 6172 269850 6196 269852
rect 6034 269798 6036 269850
rect 6098 269798 6110 269850
rect 6172 269798 6174 269850
rect 6012 269796 6036 269798
rect 6092 269796 6116 269798
rect 6172 269796 6196 269798
rect 5956 269776 6252 269796
rect 5956 268764 6252 268784
rect 6012 268762 6036 268764
rect 6092 268762 6116 268764
rect 6172 268762 6196 268764
rect 6034 268710 6036 268762
rect 6098 268710 6110 268762
rect 6172 268710 6174 268762
rect 6012 268708 6036 268710
rect 6092 268708 6116 268710
rect 6172 268708 6196 268710
rect 5956 268688 6252 268708
rect 5956 267676 6252 267696
rect 6012 267674 6036 267676
rect 6092 267674 6116 267676
rect 6172 267674 6196 267676
rect 6034 267622 6036 267674
rect 6098 267622 6110 267674
rect 6172 267622 6174 267674
rect 6012 267620 6036 267622
rect 6092 267620 6116 267622
rect 6172 267620 6196 267622
rect 5956 267600 6252 267620
rect 5956 266588 6252 266608
rect 6012 266586 6036 266588
rect 6092 266586 6116 266588
rect 6172 266586 6196 266588
rect 6034 266534 6036 266586
rect 6098 266534 6110 266586
rect 6172 266534 6174 266586
rect 6012 266532 6036 266534
rect 6092 266532 6116 266534
rect 6172 266532 6196 266534
rect 5956 266512 6252 266532
rect 5956 265500 6252 265520
rect 6012 265498 6036 265500
rect 6092 265498 6116 265500
rect 6172 265498 6196 265500
rect 6034 265446 6036 265498
rect 6098 265446 6110 265498
rect 6172 265446 6174 265498
rect 6012 265444 6036 265446
rect 6092 265444 6116 265446
rect 6172 265444 6196 265446
rect 5956 265424 6252 265444
rect 5956 264412 6252 264432
rect 6012 264410 6036 264412
rect 6092 264410 6116 264412
rect 6172 264410 6196 264412
rect 6034 264358 6036 264410
rect 6098 264358 6110 264410
rect 6172 264358 6174 264410
rect 6012 264356 6036 264358
rect 6092 264356 6116 264358
rect 6172 264356 6196 264358
rect 5956 264336 6252 264356
rect 5956 263324 6252 263344
rect 6012 263322 6036 263324
rect 6092 263322 6116 263324
rect 6172 263322 6196 263324
rect 6034 263270 6036 263322
rect 6098 263270 6110 263322
rect 6172 263270 6174 263322
rect 6012 263268 6036 263270
rect 6092 263268 6116 263270
rect 6172 263268 6196 263270
rect 5956 263248 6252 263268
rect 5956 262236 6252 262256
rect 6012 262234 6036 262236
rect 6092 262234 6116 262236
rect 6172 262234 6196 262236
rect 6034 262182 6036 262234
rect 6098 262182 6110 262234
rect 6172 262182 6174 262234
rect 6012 262180 6036 262182
rect 6092 262180 6116 262182
rect 6172 262180 6196 262182
rect 5956 262160 6252 262180
rect 5956 261148 6252 261168
rect 6012 261146 6036 261148
rect 6092 261146 6116 261148
rect 6172 261146 6196 261148
rect 6034 261094 6036 261146
rect 6098 261094 6110 261146
rect 6172 261094 6174 261146
rect 6012 261092 6036 261094
rect 6092 261092 6116 261094
rect 6172 261092 6196 261094
rect 5956 261072 6252 261092
rect 5956 260060 6252 260080
rect 6012 260058 6036 260060
rect 6092 260058 6116 260060
rect 6172 260058 6196 260060
rect 6034 260006 6036 260058
rect 6098 260006 6110 260058
rect 6172 260006 6174 260058
rect 6012 260004 6036 260006
rect 6092 260004 6116 260006
rect 6172 260004 6196 260006
rect 5956 259984 6252 260004
rect 5956 258972 6252 258992
rect 6012 258970 6036 258972
rect 6092 258970 6116 258972
rect 6172 258970 6196 258972
rect 6034 258918 6036 258970
rect 6098 258918 6110 258970
rect 6172 258918 6174 258970
rect 6012 258916 6036 258918
rect 6092 258916 6116 258918
rect 6172 258916 6196 258918
rect 5956 258896 6252 258916
rect 5956 257884 6252 257904
rect 6012 257882 6036 257884
rect 6092 257882 6116 257884
rect 6172 257882 6196 257884
rect 6034 257830 6036 257882
rect 6098 257830 6110 257882
rect 6172 257830 6174 257882
rect 6012 257828 6036 257830
rect 6092 257828 6116 257830
rect 6172 257828 6196 257830
rect 5956 257808 6252 257828
rect 5956 256796 6252 256816
rect 6012 256794 6036 256796
rect 6092 256794 6116 256796
rect 6172 256794 6196 256796
rect 6034 256742 6036 256794
rect 6098 256742 6110 256794
rect 6172 256742 6174 256794
rect 6012 256740 6036 256742
rect 6092 256740 6116 256742
rect 6172 256740 6196 256742
rect 5956 256720 6252 256740
rect 5956 255708 6252 255728
rect 6012 255706 6036 255708
rect 6092 255706 6116 255708
rect 6172 255706 6196 255708
rect 6034 255654 6036 255706
rect 6098 255654 6110 255706
rect 6172 255654 6174 255706
rect 6012 255652 6036 255654
rect 6092 255652 6116 255654
rect 6172 255652 6196 255654
rect 5956 255632 6252 255652
rect 5956 254620 6252 254640
rect 6012 254618 6036 254620
rect 6092 254618 6116 254620
rect 6172 254618 6196 254620
rect 6034 254566 6036 254618
rect 6098 254566 6110 254618
rect 6172 254566 6174 254618
rect 6012 254564 6036 254566
rect 6092 254564 6116 254566
rect 6172 254564 6196 254566
rect 5956 254544 6252 254564
rect 5956 253532 6252 253552
rect 6012 253530 6036 253532
rect 6092 253530 6116 253532
rect 6172 253530 6196 253532
rect 6034 253478 6036 253530
rect 6098 253478 6110 253530
rect 6172 253478 6174 253530
rect 6012 253476 6036 253478
rect 6092 253476 6116 253478
rect 6172 253476 6196 253478
rect 5956 253456 6252 253476
rect 5956 252444 6252 252464
rect 6012 252442 6036 252444
rect 6092 252442 6116 252444
rect 6172 252442 6196 252444
rect 6034 252390 6036 252442
rect 6098 252390 6110 252442
rect 6172 252390 6174 252442
rect 6012 252388 6036 252390
rect 6092 252388 6116 252390
rect 6172 252388 6196 252390
rect 5956 252368 6252 252388
rect 5956 251356 6252 251376
rect 6012 251354 6036 251356
rect 6092 251354 6116 251356
rect 6172 251354 6196 251356
rect 6034 251302 6036 251354
rect 6098 251302 6110 251354
rect 6172 251302 6174 251354
rect 6012 251300 6036 251302
rect 6092 251300 6116 251302
rect 6172 251300 6196 251302
rect 5956 251280 6252 251300
rect 5956 250268 6252 250288
rect 6012 250266 6036 250268
rect 6092 250266 6116 250268
rect 6172 250266 6196 250268
rect 6034 250214 6036 250266
rect 6098 250214 6110 250266
rect 6172 250214 6174 250266
rect 6012 250212 6036 250214
rect 6092 250212 6116 250214
rect 6172 250212 6196 250214
rect 5956 250192 6252 250212
rect 5956 249180 6252 249200
rect 6012 249178 6036 249180
rect 6092 249178 6116 249180
rect 6172 249178 6196 249180
rect 6034 249126 6036 249178
rect 6098 249126 6110 249178
rect 6172 249126 6174 249178
rect 6012 249124 6036 249126
rect 6092 249124 6116 249126
rect 6172 249124 6196 249126
rect 5956 249104 6252 249124
rect 5956 248092 6252 248112
rect 6012 248090 6036 248092
rect 6092 248090 6116 248092
rect 6172 248090 6196 248092
rect 6034 248038 6036 248090
rect 6098 248038 6110 248090
rect 6172 248038 6174 248090
rect 6012 248036 6036 248038
rect 6092 248036 6116 248038
rect 6172 248036 6196 248038
rect 5956 248016 6252 248036
rect 5956 247004 6252 247024
rect 6012 247002 6036 247004
rect 6092 247002 6116 247004
rect 6172 247002 6196 247004
rect 6034 246950 6036 247002
rect 6098 246950 6110 247002
rect 6172 246950 6174 247002
rect 6012 246948 6036 246950
rect 6092 246948 6116 246950
rect 6172 246948 6196 246950
rect 5956 246928 6252 246948
rect 5956 245916 6252 245936
rect 6012 245914 6036 245916
rect 6092 245914 6116 245916
rect 6172 245914 6196 245916
rect 6034 245862 6036 245914
rect 6098 245862 6110 245914
rect 6172 245862 6174 245914
rect 6012 245860 6036 245862
rect 6092 245860 6116 245862
rect 6172 245860 6196 245862
rect 5956 245840 6252 245860
rect 5956 244828 6252 244848
rect 6012 244826 6036 244828
rect 6092 244826 6116 244828
rect 6172 244826 6196 244828
rect 6034 244774 6036 244826
rect 6098 244774 6110 244826
rect 6172 244774 6174 244826
rect 6012 244772 6036 244774
rect 6092 244772 6116 244774
rect 6172 244772 6196 244774
rect 5956 244752 6252 244772
rect 5956 243740 6252 243760
rect 6012 243738 6036 243740
rect 6092 243738 6116 243740
rect 6172 243738 6196 243740
rect 6034 243686 6036 243738
rect 6098 243686 6110 243738
rect 6172 243686 6174 243738
rect 6012 243684 6036 243686
rect 6092 243684 6116 243686
rect 6172 243684 6196 243686
rect 5956 243664 6252 243684
rect 5956 242652 6252 242672
rect 6012 242650 6036 242652
rect 6092 242650 6116 242652
rect 6172 242650 6196 242652
rect 6034 242598 6036 242650
rect 6098 242598 6110 242650
rect 6172 242598 6174 242650
rect 6012 242596 6036 242598
rect 6092 242596 6116 242598
rect 6172 242596 6196 242598
rect 5956 242576 6252 242596
rect 5956 241564 6252 241584
rect 6012 241562 6036 241564
rect 6092 241562 6116 241564
rect 6172 241562 6196 241564
rect 6034 241510 6036 241562
rect 6098 241510 6110 241562
rect 6172 241510 6174 241562
rect 6012 241508 6036 241510
rect 6092 241508 6116 241510
rect 6172 241508 6196 241510
rect 5956 241488 6252 241508
rect 5956 240476 6252 240496
rect 6012 240474 6036 240476
rect 6092 240474 6116 240476
rect 6172 240474 6196 240476
rect 6034 240422 6036 240474
rect 6098 240422 6110 240474
rect 6172 240422 6174 240474
rect 6012 240420 6036 240422
rect 6092 240420 6116 240422
rect 6172 240420 6196 240422
rect 5956 240400 6252 240420
rect 5956 239388 6252 239408
rect 6012 239386 6036 239388
rect 6092 239386 6116 239388
rect 6172 239386 6196 239388
rect 6034 239334 6036 239386
rect 6098 239334 6110 239386
rect 6172 239334 6174 239386
rect 6012 239332 6036 239334
rect 6092 239332 6116 239334
rect 6172 239332 6196 239334
rect 5956 239312 6252 239332
rect 5956 238300 6252 238320
rect 6012 238298 6036 238300
rect 6092 238298 6116 238300
rect 6172 238298 6196 238300
rect 6034 238246 6036 238298
rect 6098 238246 6110 238298
rect 6172 238246 6174 238298
rect 6012 238244 6036 238246
rect 6092 238244 6116 238246
rect 6172 238244 6196 238246
rect 5956 238224 6252 238244
rect 5956 237212 6252 237232
rect 6012 237210 6036 237212
rect 6092 237210 6116 237212
rect 6172 237210 6196 237212
rect 6034 237158 6036 237210
rect 6098 237158 6110 237210
rect 6172 237158 6174 237210
rect 6012 237156 6036 237158
rect 6092 237156 6116 237158
rect 6172 237156 6196 237158
rect 5956 237136 6252 237156
rect 5956 236124 6252 236144
rect 6012 236122 6036 236124
rect 6092 236122 6116 236124
rect 6172 236122 6196 236124
rect 6034 236070 6036 236122
rect 6098 236070 6110 236122
rect 6172 236070 6174 236122
rect 6012 236068 6036 236070
rect 6092 236068 6116 236070
rect 6172 236068 6196 236070
rect 5956 236048 6252 236068
rect 5956 235036 6252 235056
rect 6012 235034 6036 235036
rect 6092 235034 6116 235036
rect 6172 235034 6196 235036
rect 6034 234982 6036 235034
rect 6098 234982 6110 235034
rect 6172 234982 6174 235034
rect 6012 234980 6036 234982
rect 6092 234980 6116 234982
rect 6172 234980 6196 234982
rect 5956 234960 6252 234980
rect 5956 233948 6252 233968
rect 6012 233946 6036 233948
rect 6092 233946 6116 233948
rect 6172 233946 6196 233948
rect 6034 233894 6036 233946
rect 6098 233894 6110 233946
rect 6172 233894 6174 233946
rect 6012 233892 6036 233894
rect 6092 233892 6116 233894
rect 6172 233892 6196 233894
rect 5956 233872 6252 233892
rect 5540 233640 5592 233646
rect 5540 233582 5592 233588
rect 5956 232860 6252 232880
rect 6012 232858 6036 232860
rect 6092 232858 6116 232860
rect 6172 232858 6196 232860
rect 6034 232806 6036 232858
rect 6098 232806 6110 232858
rect 6172 232806 6174 232858
rect 6012 232804 6036 232806
rect 6092 232804 6116 232806
rect 6172 232804 6196 232806
rect 5956 232784 6252 232804
rect 5956 231772 6252 231792
rect 6012 231770 6036 231772
rect 6092 231770 6116 231772
rect 6172 231770 6196 231772
rect 6034 231718 6036 231770
rect 6098 231718 6110 231770
rect 6172 231718 6174 231770
rect 6012 231716 6036 231718
rect 6092 231716 6116 231718
rect 6172 231716 6196 231718
rect 5956 231696 6252 231716
rect 5956 230684 6252 230704
rect 6012 230682 6036 230684
rect 6092 230682 6116 230684
rect 6172 230682 6196 230684
rect 6034 230630 6036 230682
rect 6098 230630 6110 230682
rect 6172 230630 6174 230682
rect 6012 230628 6036 230630
rect 6092 230628 6116 230630
rect 6172 230628 6196 230630
rect 5956 230608 6252 230628
rect 5956 229596 6252 229616
rect 6012 229594 6036 229596
rect 6092 229594 6116 229596
rect 6172 229594 6196 229596
rect 6034 229542 6036 229594
rect 6098 229542 6110 229594
rect 6172 229542 6174 229594
rect 6012 229540 6036 229542
rect 6092 229540 6116 229542
rect 6172 229540 6196 229542
rect 5956 229520 6252 229540
rect 5956 228508 6252 228528
rect 6012 228506 6036 228508
rect 6092 228506 6116 228508
rect 6172 228506 6196 228508
rect 6034 228454 6036 228506
rect 6098 228454 6110 228506
rect 6172 228454 6174 228506
rect 6012 228452 6036 228454
rect 6092 228452 6116 228454
rect 6172 228452 6196 228454
rect 5956 228432 6252 228452
rect 5956 227420 6252 227440
rect 6012 227418 6036 227420
rect 6092 227418 6116 227420
rect 6172 227418 6196 227420
rect 6034 227366 6036 227418
rect 6098 227366 6110 227418
rect 6172 227366 6174 227418
rect 6012 227364 6036 227366
rect 6092 227364 6116 227366
rect 6172 227364 6196 227366
rect 5956 227344 6252 227364
rect 5816 226432 5868 226438
rect 5816 226374 5868 226380
rect 5828 225486 5856 226374
rect 5956 226332 6252 226352
rect 6012 226330 6036 226332
rect 6092 226330 6116 226332
rect 6172 226330 6196 226332
rect 6034 226278 6036 226330
rect 6098 226278 6110 226330
rect 6172 226278 6174 226330
rect 6012 226276 6036 226278
rect 6092 226276 6116 226278
rect 6172 226276 6196 226278
rect 5956 226256 6252 226276
rect 6288 225554 6316 282503
rect 6366 249248 6422 249257
rect 6366 249183 6422 249192
rect 6380 239290 6408 249183
rect 6368 239284 6420 239290
rect 6368 239226 6420 239232
rect 6748 234258 6776 332574
rect 6826 332520 6882 332574
rect 7944 332574 8078 332602
rect 7944 332466 7972 332574
rect 8022 332520 8078 332574
rect 8300 332580 8352 332586
rect 8300 332522 8352 332528
rect 9310 332580 9366 333000
rect 9310 332528 9312 332580
rect 9364 332528 9366 332580
rect 7944 332438 8064 332466
rect 7622 330236 7918 330256
rect 7678 330234 7702 330236
rect 7758 330234 7782 330236
rect 7838 330234 7862 330236
rect 7700 330182 7702 330234
rect 7764 330182 7776 330234
rect 7838 330182 7840 330234
rect 7678 330180 7702 330182
rect 7758 330180 7782 330182
rect 7838 330180 7862 330182
rect 7622 330160 7918 330180
rect 7622 329148 7918 329168
rect 7678 329146 7702 329148
rect 7758 329146 7782 329148
rect 7838 329146 7862 329148
rect 7700 329094 7702 329146
rect 7764 329094 7776 329146
rect 7838 329094 7840 329146
rect 7678 329092 7702 329094
rect 7758 329092 7782 329094
rect 7838 329092 7862 329094
rect 7622 329072 7918 329092
rect 7622 328060 7918 328080
rect 7678 328058 7702 328060
rect 7758 328058 7782 328060
rect 7838 328058 7862 328060
rect 7700 328006 7702 328058
rect 7764 328006 7776 328058
rect 7838 328006 7840 328058
rect 7678 328004 7702 328006
rect 7758 328004 7782 328006
rect 7838 328004 7862 328006
rect 7622 327984 7918 328004
rect 7622 326972 7918 326992
rect 7678 326970 7702 326972
rect 7758 326970 7782 326972
rect 7838 326970 7862 326972
rect 7700 326918 7702 326970
rect 7764 326918 7776 326970
rect 7838 326918 7840 326970
rect 7678 326916 7702 326918
rect 7758 326916 7782 326918
rect 7838 326916 7862 326918
rect 7622 326896 7918 326916
rect 7622 325884 7918 325904
rect 7678 325882 7702 325884
rect 7758 325882 7782 325884
rect 7838 325882 7862 325884
rect 7700 325830 7702 325882
rect 7764 325830 7776 325882
rect 7838 325830 7840 325882
rect 7678 325828 7702 325830
rect 7758 325828 7782 325830
rect 7838 325828 7862 325830
rect 7622 325808 7918 325828
rect 7622 324796 7918 324816
rect 7678 324794 7702 324796
rect 7758 324794 7782 324796
rect 7838 324794 7862 324796
rect 7700 324742 7702 324794
rect 7764 324742 7776 324794
rect 7838 324742 7840 324794
rect 7678 324740 7702 324742
rect 7758 324740 7782 324742
rect 7838 324740 7862 324742
rect 7622 324720 7918 324740
rect 7622 323708 7918 323728
rect 7678 323706 7702 323708
rect 7758 323706 7782 323708
rect 7838 323706 7862 323708
rect 7700 323654 7702 323706
rect 7764 323654 7776 323706
rect 7838 323654 7840 323706
rect 7678 323652 7702 323654
rect 7758 323652 7782 323654
rect 7838 323652 7862 323654
rect 7622 323632 7918 323652
rect 7622 322620 7918 322640
rect 7678 322618 7702 322620
rect 7758 322618 7782 322620
rect 7838 322618 7862 322620
rect 7700 322566 7702 322618
rect 7764 322566 7776 322618
rect 7838 322566 7840 322618
rect 7678 322564 7702 322566
rect 7758 322564 7782 322566
rect 7838 322564 7862 322566
rect 7622 322544 7918 322564
rect 7622 321532 7918 321552
rect 7678 321530 7702 321532
rect 7758 321530 7782 321532
rect 7838 321530 7862 321532
rect 7700 321478 7702 321530
rect 7764 321478 7776 321530
rect 7838 321478 7840 321530
rect 7678 321476 7702 321478
rect 7758 321476 7782 321478
rect 7838 321476 7862 321478
rect 7622 321456 7918 321476
rect 7622 320444 7918 320464
rect 7678 320442 7702 320444
rect 7758 320442 7782 320444
rect 7838 320442 7862 320444
rect 7700 320390 7702 320442
rect 7764 320390 7776 320442
rect 7838 320390 7840 320442
rect 7678 320388 7702 320390
rect 7758 320388 7782 320390
rect 7838 320388 7862 320390
rect 7622 320368 7918 320388
rect 7622 319356 7918 319376
rect 7678 319354 7702 319356
rect 7758 319354 7782 319356
rect 7838 319354 7862 319356
rect 7700 319302 7702 319354
rect 7764 319302 7776 319354
rect 7838 319302 7840 319354
rect 7678 319300 7702 319302
rect 7758 319300 7782 319302
rect 7838 319300 7862 319302
rect 7622 319280 7918 319300
rect 7622 318268 7918 318288
rect 7678 318266 7702 318268
rect 7758 318266 7782 318268
rect 7838 318266 7862 318268
rect 7700 318214 7702 318266
rect 7764 318214 7776 318266
rect 7838 318214 7840 318266
rect 7678 318212 7702 318214
rect 7758 318212 7782 318214
rect 7838 318212 7862 318214
rect 7622 318192 7918 318212
rect 7622 317180 7918 317200
rect 7678 317178 7702 317180
rect 7758 317178 7782 317180
rect 7838 317178 7862 317180
rect 7700 317126 7702 317178
rect 7764 317126 7776 317178
rect 7838 317126 7840 317178
rect 7678 317124 7702 317126
rect 7758 317124 7782 317126
rect 7838 317124 7862 317126
rect 7622 317104 7918 317124
rect 7622 316092 7918 316112
rect 7678 316090 7702 316092
rect 7758 316090 7782 316092
rect 7838 316090 7862 316092
rect 7700 316038 7702 316090
rect 7764 316038 7776 316090
rect 7838 316038 7840 316090
rect 7678 316036 7702 316038
rect 7758 316036 7782 316038
rect 7838 316036 7862 316038
rect 7622 316016 7918 316036
rect 7286 315888 7342 315897
rect 7286 315823 7342 315832
rect 6828 239080 6880 239086
rect 6828 239022 6880 239028
rect 6736 234252 6788 234258
rect 6736 234194 6788 234200
rect 6748 233850 6776 234194
rect 6736 233844 6788 233850
rect 6736 233786 6788 233792
rect 6840 233782 6868 239022
rect 6920 234184 6972 234190
rect 6920 234126 6972 234132
rect 6828 233776 6880 233782
rect 6828 233718 6880 233724
rect 6932 233510 6960 234126
rect 6920 233504 6972 233510
rect 6920 233446 6972 233452
rect 7012 225888 7064 225894
rect 7012 225830 7064 225836
rect 6276 225548 6328 225554
rect 6276 225490 6328 225496
rect 5816 225480 5868 225486
rect 5816 225422 5868 225428
rect 5632 225344 5684 225350
rect 5632 225286 5684 225292
rect 5448 224460 5500 224466
rect 5448 224402 5500 224408
rect 5356 224392 5408 224398
rect 5356 224334 5408 224340
rect 5644 72078 5672 225286
rect 5828 225146 5856 225422
rect 5956 225244 6252 225264
rect 6012 225242 6036 225244
rect 6092 225242 6116 225244
rect 6172 225242 6196 225244
rect 6034 225190 6036 225242
rect 6098 225190 6110 225242
rect 6172 225190 6174 225242
rect 6012 225188 6036 225190
rect 6092 225188 6116 225190
rect 6172 225188 6196 225190
rect 5956 225168 6252 225188
rect 6288 225146 6316 225490
rect 5816 225140 5868 225146
rect 5816 225082 5868 225088
rect 6276 225140 6328 225146
rect 6276 225082 6328 225088
rect 6920 225004 6972 225010
rect 6920 224946 6972 224952
rect 6932 224602 6960 224946
rect 7024 224942 7052 225830
rect 7012 224936 7064 224942
rect 7012 224878 7064 224884
rect 7024 224602 7052 224878
rect 6920 224596 6972 224602
rect 6920 224538 6972 224544
rect 7012 224596 7064 224602
rect 7012 224538 7064 224544
rect 5816 224460 5868 224466
rect 5816 224402 5868 224408
rect 5828 224058 5856 224402
rect 6276 224392 6328 224398
rect 6276 224334 6328 224340
rect 5956 224156 6252 224176
rect 6012 224154 6036 224156
rect 6092 224154 6116 224156
rect 6172 224154 6196 224156
rect 6034 224102 6036 224154
rect 6098 224102 6110 224154
rect 6172 224102 6174 224154
rect 6012 224100 6036 224102
rect 6092 224100 6116 224102
rect 6172 224100 6196 224102
rect 5956 224080 6252 224100
rect 6288 224058 6316 224334
rect 6552 224256 6604 224262
rect 6552 224198 6604 224204
rect 5816 224052 5868 224058
rect 5816 223994 5868 224000
rect 6276 224052 6328 224058
rect 6276 223994 6328 224000
rect 5956 223068 6252 223088
rect 6012 223066 6036 223068
rect 6092 223066 6116 223068
rect 6172 223066 6196 223068
rect 6034 223014 6036 223066
rect 6098 223014 6110 223066
rect 6172 223014 6174 223066
rect 6012 223012 6036 223014
rect 6092 223012 6116 223014
rect 6172 223012 6196 223014
rect 5956 222992 6252 223012
rect 5956 221980 6252 222000
rect 6012 221978 6036 221980
rect 6092 221978 6116 221980
rect 6172 221978 6196 221980
rect 6034 221926 6036 221978
rect 6098 221926 6110 221978
rect 6172 221926 6174 221978
rect 6012 221924 6036 221926
rect 6092 221924 6116 221926
rect 6172 221924 6196 221926
rect 5956 221904 6252 221924
rect 5956 220892 6252 220912
rect 6012 220890 6036 220892
rect 6092 220890 6116 220892
rect 6172 220890 6196 220892
rect 6034 220838 6036 220890
rect 6098 220838 6110 220890
rect 6172 220838 6174 220890
rect 6012 220836 6036 220838
rect 6092 220836 6116 220838
rect 6172 220836 6196 220838
rect 5956 220816 6252 220836
rect 5956 219804 6252 219824
rect 6012 219802 6036 219804
rect 6092 219802 6116 219804
rect 6172 219802 6196 219804
rect 6034 219750 6036 219802
rect 6098 219750 6110 219802
rect 6172 219750 6174 219802
rect 6012 219748 6036 219750
rect 6092 219748 6116 219750
rect 6172 219748 6196 219750
rect 5956 219728 6252 219748
rect 5956 218716 6252 218736
rect 6012 218714 6036 218716
rect 6092 218714 6116 218716
rect 6172 218714 6196 218716
rect 6034 218662 6036 218714
rect 6098 218662 6110 218714
rect 6172 218662 6174 218714
rect 6012 218660 6036 218662
rect 6092 218660 6116 218662
rect 6172 218660 6196 218662
rect 5956 218640 6252 218660
rect 5956 217628 6252 217648
rect 6012 217626 6036 217628
rect 6092 217626 6116 217628
rect 6172 217626 6196 217628
rect 6034 217574 6036 217626
rect 6098 217574 6110 217626
rect 6172 217574 6174 217626
rect 6012 217572 6036 217574
rect 6092 217572 6116 217574
rect 6172 217572 6196 217574
rect 5956 217552 6252 217572
rect 5956 216540 6252 216560
rect 6012 216538 6036 216540
rect 6092 216538 6116 216540
rect 6172 216538 6196 216540
rect 6034 216486 6036 216538
rect 6098 216486 6110 216538
rect 6172 216486 6174 216538
rect 6012 216484 6036 216486
rect 6092 216484 6116 216486
rect 6172 216484 6196 216486
rect 5956 216464 6252 216484
rect 5956 215452 6252 215472
rect 6012 215450 6036 215452
rect 6092 215450 6116 215452
rect 6172 215450 6196 215452
rect 6034 215398 6036 215450
rect 6098 215398 6110 215450
rect 6172 215398 6174 215450
rect 6012 215396 6036 215398
rect 6092 215396 6116 215398
rect 6172 215396 6196 215398
rect 5956 215376 6252 215396
rect 5956 214364 6252 214384
rect 6012 214362 6036 214364
rect 6092 214362 6116 214364
rect 6172 214362 6196 214364
rect 6034 214310 6036 214362
rect 6098 214310 6110 214362
rect 6172 214310 6174 214362
rect 6012 214308 6036 214310
rect 6092 214308 6116 214310
rect 6172 214308 6196 214310
rect 5956 214288 6252 214308
rect 5956 213276 6252 213296
rect 6012 213274 6036 213276
rect 6092 213274 6116 213276
rect 6172 213274 6196 213276
rect 6034 213222 6036 213274
rect 6098 213222 6110 213274
rect 6172 213222 6174 213274
rect 6012 213220 6036 213222
rect 6092 213220 6116 213222
rect 6172 213220 6196 213222
rect 5956 213200 6252 213220
rect 5956 212188 6252 212208
rect 6012 212186 6036 212188
rect 6092 212186 6116 212188
rect 6172 212186 6196 212188
rect 6034 212134 6036 212186
rect 6098 212134 6110 212186
rect 6172 212134 6174 212186
rect 6012 212132 6036 212134
rect 6092 212132 6116 212134
rect 6172 212132 6196 212134
rect 5956 212112 6252 212132
rect 5956 211100 6252 211120
rect 6012 211098 6036 211100
rect 6092 211098 6116 211100
rect 6172 211098 6196 211100
rect 6034 211046 6036 211098
rect 6098 211046 6110 211098
rect 6172 211046 6174 211098
rect 6012 211044 6036 211046
rect 6092 211044 6116 211046
rect 6172 211044 6196 211046
rect 5956 211024 6252 211044
rect 5956 210012 6252 210032
rect 6012 210010 6036 210012
rect 6092 210010 6116 210012
rect 6172 210010 6196 210012
rect 6034 209958 6036 210010
rect 6098 209958 6110 210010
rect 6172 209958 6174 210010
rect 6012 209956 6036 209958
rect 6092 209956 6116 209958
rect 6172 209956 6196 209958
rect 5956 209936 6252 209956
rect 5956 208924 6252 208944
rect 6012 208922 6036 208924
rect 6092 208922 6116 208924
rect 6172 208922 6196 208924
rect 6034 208870 6036 208922
rect 6098 208870 6110 208922
rect 6172 208870 6174 208922
rect 6012 208868 6036 208870
rect 6092 208868 6116 208870
rect 6172 208868 6196 208870
rect 5956 208848 6252 208868
rect 5956 207836 6252 207856
rect 6012 207834 6036 207836
rect 6092 207834 6116 207836
rect 6172 207834 6196 207836
rect 6034 207782 6036 207834
rect 6098 207782 6110 207834
rect 6172 207782 6174 207834
rect 6012 207780 6036 207782
rect 6092 207780 6116 207782
rect 6172 207780 6196 207782
rect 5956 207760 6252 207780
rect 5956 206748 6252 206768
rect 6012 206746 6036 206748
rect 6092 206746 6116 206748
rect 6172 206746 6196 206748
rect 6034 206694 6036 206746
rect 6098 206694 6110 206746
rect 6172 206694 6174 206746
rect 6012 206692 6036 206694
rect 6092 206692 6116 206694
rect 6172 206692 6196 206694
rect 5956 206672 6252 206692
rect 5956 205660 6252 205680
rect 6012 205658 6036 205660
rect 6092 205658 6116 205660
rect 6172 205658 6196 205660
rect 6034 205606 6036 205658
rect 6098 205606 6110 205658
rect 6172 205606 6174 205658
rect 6012 205604 6036 205606
rect 6092 205604 6116 205606
rect 6172 205604 6196 205606
rect 5956 205584 6252 205604
rect 5956 204572 6252 204592
rect 6012 204570 6036 204572
rect 6092 204570 6116 204572
rect 6172 204570 6196 204572
rect 6034 204518 6036 204570
rect 6098 204518 6110 204570
rect 6172 204518 6174 204570
rect 6012 204516 6036 204518
rect 6092 204516 6116 204518
rect 6172 204516 6196 204518
rect 5956 204496 6252 204516
rect 5956 203484 6252 203504
rect 6012 203482 6036 203484
rect 6092 203482 6116 203484
rect 6172 203482 6196 203484
rect 6034 203430 6036 203482
rect 6098 203430 6110 203482
rect 6172 203430 6174 203482
rect 6012 203428 6036 203430
rect 6092 203428 6116 203430
rect 6172 203428 6196 203430
rect 5956 203408 6252 203428
rect 5956 202396 6252 202416
rect 6012 202394 6036 202396
rect 6092 202394 6116 202396
rect 6172 202394 6196 202396
rect 6034 202342 6036 202394
rect 6098 202342 6110 202394
rect 6172 202342 6174 202394
rect 6012 202340 6036 202342
rect 6092 202340 6116 202342
rect 6172 202340 6196 202342
rect 5956 202320 6252 202340
rect 5956 201308 6252 201328
rect 6012 201306 6036 201308
rect 6092 201306 6116 201308
rect 6172 201306 6196 201308
rect 6034 201254 6036 201306
rect 6098 201254 6110 201306
rect 6172 201254 6174 201306
rect 6012 201252 6036 201254
rect 6092 201252 6116 201254
rect 6172 201252 6196 201254
rect 5956 201232 6252 201252
rect 5956 200220 6252 200240
rect 6012 200218 6036 200220
rect 6092 200218 6116 200220
rect 6172 200218 6196 200220
rect 6034 200166 6036 200218
rect 6098 200166 6110 200218
rect 6172 200166 6174 200218
rect 6012 200164 6036 200166
rect 6092 200164 6116 200166
rect 6172 200164 6196 200166
rect 5956 200144 6252 200164
rect 5956 199132 6252 199152
rect 6012 199130 6036 199132
rect 6092 199130 6116 199132
rect 6172 199130 6196 199132
rect 6034 199078 6036 199130
rect 6098 199078 6110 199130
rect 6172 199078 6174 199130
rect 6012 199076 6036 199078
rect 6092 199076 6116 199078
rect 6172 199076 6196 199078
rect 5956 199056 6252 199076
rect 5956 198044 6252 198064
rect 6012 198042 6036 198044
rect 6092 198042 6116 198044
rect 6172 198042 6196 198044
rect 6034 197990 6036 198042
rect 6098 197990 6110 198042
rect 6172 197990 6174 198042
rect 6012 197988 6036 197990
rect 6092 197988 6116 197990
rect 6172 197988 6196 197990
rect 5956 197968 6252 197988
rect 5956 196956 6252 196976
rect 6012 196954 6036 196956
rect 6092 196954 6116 196956
rect 6172 196954 6196 196956
rect 6034 196902 6036 196954
rect 6098 196902 6110 196954
rect 6172 196902 6174 196954
rect 6012 196900 6036 196902
rect 6092 196900 6116 196902
rect 6172 196900 6196 196902
rect 5956 196880 6252 196900
rect 5956 195868 6252 195888
rect 6012 195866 6036 195868
rect 6092 195866 6116 195868
rect 6172 195866 6196 195868
rect 6034 195814 6036 195866
rect 6098 195814 6110 195866
rect 6172 195814 6174 195866
rect 6012 195812 6036 195814
rect 6092 195812 6116 195814
rect 6172 195812 6196 195814
rect 5956 195792 6252 195812
rect 5956 194780 6252 194800
rect 6012 194778 6036 194780
rect 6092 194778 6116 194780
rect 6172 194778 6196 194780
rect 6034 194726 6036 194778
rect 6098 194726 6110 194778
rect 6172 194726 6174 194778
rect 6012 194724 6036 194726
rect 6092 194724 6116 194726
rect 6172 194724 6196 194726
rect 5956 194704 6252 194724
rect 5956 193692 6252 193712
rect 6012 193690 6036 193692
rect 6092 193690 6116 193692
rect 6172 193690 6196 193692
rect 6034 193638 6036 193690
rect 6098 193638 6110 193690
rect 6172 193638 6174 193690
rect 6012 193636 6036 193638
rect 6092 193636 6116 193638
rect 6172 193636 6196 193638
rect 5956 193616 6252 193636
rect 5956 192604 6252 192624
rect 6012 192602 6036 192604
rect 6092 192602 6116 192604
rect 6172 192602 6196 192604
rect 6034 192550 6036 192602
rect 6098 192550 6110 192602
rect 6172 192550 6174 192602
rect 6012 192548 6036 192550
rect 6092 192548 6116 192550
rect 6172 192548 6196 192550
rect 5956 192528 6252 192548
rect 5956 191516 6252 191536
rect 6012 191514 6036 191516
rect 6092 191514 6116 191516
rect 6172 191514 6196 191516
rect 6034 191462 6036 191514
rect 6098 191462 6110 191514
rect 6172 191462 6174 191514
rect 6012 191460 6036 191462
rect 6092 191460 6116 191462
rect 6172 191460 6196 191462
rect 5956 191440 6252 191460
rect 5956 190428 6252 190448
rect 6012 190426 6036 190428
rect 6092 190426 6116 190428
rect 6172 190426 6196 190428
rect 6034 190374 6036 190426
rect 6098 190374 6110 190426
rect 6172 190374 6174 190426
rect 6012 190372 6036 190374
rect 6092 190372 6116 190374
rect 6172 190372 6196 190374
rect 5956 190352 6252 190372
rect 5956 189340 6252 189360
rect 6012 189338 6036 189340
rect 6092 189338 6116 189340
rect 6172 189338 6196 189340
rect 6034 189286 6036 189338
rect 6098 189286 6110 189338
rect 6172 189286 6174 189338
rect 6012 189284 6036 189286
rect 6092 189284 6116 189286
rect 6172 189284 6196 189286
rect 5956 189264 6252 189284
rect 5956 188252 6252 188272
rect 6012 188250 6036 188252
rect 6092 188250 6116 188252
rect 6172 188250 6196 188252
rect 6034 188198 6036 188250
rect 6098 188198 6110 188250
rect 6172 188198 6174 188250
rect 6012 188196 6036 188198
rect 6092 188196 6116 188198
rect 6172 188196 6196 188198
rect 5956 188176 6252 188196
rect 5956 187164 6252 187184
rect 6012 187162 6036 187164
rect 6092 187162 6116 187164
rect 6172 187162 6196 187164
rect 6034 187110 6036 187162
rect 6098 187110 6110 187162
rect 6172 187110 6174 187162
rect 6012 187108 6036 187110
rect 6092 187108 6116 187110
rect 6172 187108 6196 187110
rect 5956 187088 6252 187108
rect 5956 186076 6252 186096
rect 6012 186074 6036 186076
rect 6092 186074 6116 186076
rect 6172 186074 6196 186076
rect 6034 186022 6036 186074
rect 6098 186022 6110 186074
rect 6172 186022 6174 186074
rect 6012 186020 6036 186022
rect 6092 186020 6116 186022
rect 6172 186020 6196 186022
rect 5956 186000 6252 186020
rect 5956 184988 6252 185008
rect 6012 184986 6036 184988
rect 6092 184986 6116 184988
rect 6172 184986 6196 184988
rect 6034 184934 6036 184986
rect 6098 184934 6110 184986
rect 6172 184934 6174 184986
rect 6012 184932 6036 184934
rect 6092 184932 6116 184934
rect 6172 184932 6196 184934
rect 5956 184912 6252 184932
rect 5956 183900 6252 183920
rect 6012 183898 6036 183900
rect 6092 183898 6116 183900
rect 6172 183898 6196 183900
rect 6034 183846 6036 183898
rect 6098 183846 6110 183898
rect 6172 183846 6174 183898
rect 6012 183844 6036 183846
rect 6092 183844 6116 183846
rect 6172 183844 6196 183846
rect 5956 183824 6252 183844
rect 5956 182812 6252 182832
rect 6012 182810 6036 182812
rect 6092 182810 6116 182812
rect 6172 182810 6196 182812
rect 6034 182758 6036 182810
rect 6098 182758 6110 182810
rect 6172 182758 6174 182810
rect 6012 182756 6036 182758
rect 6092 182756 6116 182758
rect 6172 182756 6196 182758
rect 5956 182736 6252 182756
rect 5956 181724 6252 181744
rect 6012 181722 6036 181724
rect 6092 181722 6116 181724
rect 6172 181722 6196 181724
rect 6034 181670 6036 181722
rect 6098 181670 6110 181722
rect 6172 181670 6174 181722
rect 6012 181668 6036 181670
rect 6092 181668 6116 181670
rect 6172 181668 6196 181670
rect 5956 181648 6252 181668
rect 5956 180636 6252 180656
rect 6012 180634 6036 180636
rect 6092 180634 6116 180636
rect 6172 180634 6196 180636
rect 6034 180582 6036 180634
rect 6098 180582 6110 180634
rect 6172 180582 6174 180634
rect 6012 180580 6036 180582
rect 6092 180580 6116 180582
rect 6172 180580 6196 180582
rect 5956 180560 6252 180580
rect 5956 179548 6252 179568
rect 6012 179546 6036 179548
rect 6092 179546 6116 179548
rect 6172 179546 6196 179548
rect 6034 179494 6036 179546
rect 6098 179494 6110 179546
rect 6172 179494 6174 179546
rect 6012 179492 6036 179494
rect 6092 179492 6116 179494
rect 6172 179492 6196 179494
rect 5956 179472 6252 179492
rect 5956 178460 6252 178480
rect 6012 178458 6036 178460
rect 6092 178458 6116 178460
rect 6172 178458 6196 178460
rect 6034 178406 6036 178458
rect 6098 178406 6110 178458
rect 6172 178406 6174 178458
rect 6012 178404 6036 178406
rect 6092 178404 6116 178406
rect 6172 178404 6196 178406
rect 5956 178384 6252 178404
rect 5956 177372 6252 177392
rect 6012 177370 6036 177372
rect 6092 177370 6116 177372
rect 6172 177370 6196 177372
rect 6034 177318 6036 177370
rect 6098 177318 6110 177370
rect 6172 177318 6174 177370
rect 6012 177316 6036 177318
rect 6092 177316 6116 177318
rect 6172 177316 6196 177318
rect 5956 177296 6252 177316
rect 5956 176284 6252 176304
rect 6012 176282 6036 176284
rect 6092 176282 6116 176284
rect 6172 176282 6196 176284
rect 6034 176230 6036 176282
rect 6098 176230 6110 176282
rect 6172 176230 6174 176282
rect 6012 176228 6036 176230
rect 6092 176228 6116 176230
rect 6172 176228 6196 176230
rect 5956 176208 6252 176228
rect 5956 175196 6252 175216
rect 6012 175194 6036 175196
rect 6092 175194 6116 175196
rect 6172 175194 6196 175196
rect 6034 175142 6036 175194
rect 6098 175142 6110 175194
rect 6172 175142 6174 175194
rect 6012 175140 6036 175142
rect 6092 175140 6116 175142
rect 6172 175140 6196 175142
rect 5956 175120 6252 175140
rect 5956 174108 6252 174128
rect 6012 174106 6036 174108
rect 6092 174106 6116 174108
rect 6172 174106 6196 174108
rect 6034 174054 6036 174106
rect 6098 174054 6110 174106
rect 6172 174054 6174 174106
rect 6012 174052 6036 174054
rect 6092 174052 6116 174054
rect 6172 174052 6196 174054
rect 5956 174032 6252 174052
rect 5956 173020 6252 173040
rect 6012 173018 6036 173020
rect 6092 173018 6116 173020
rect 6172 173018 6196 173020
rect 6034 172966 6036 173018
rect 6098 172966 6110 173018
rect 6172 172966 6174 173018
rect 6012 172964 6036 172966
rect 6092 172964 6116 172966
rect 6172 172964 6196 172966
rect 5956 172944 6252 172964
rect 6564 172242 6592 224198
rect 7010 216200 7066 216209
rect 7010 216135 7066 216144
rect 6736 214056 6788 214062
rect 6736 213998 6788 214004
rect 6748 211750 6776 213998
rect 6736 211744 6788 211750
rect 6736 211686 6788 211692
rect 6642 182608 6698 182617
rect 6642 182543 6698 182552
rect 6656 172378 6684 182543
rect 6644 172372 6696 172378
rect 6644 172314 6696 172320
rect 6552 172236 6604 172242
rect 6552 172178 6604 172184
rect 5956 171932 6252 171952
rect 6012 171930 6036 171932
rect 6092 171930 6116 171932
rect 6172 171930 6196 171932
rect 6034 171878 6036 171930
rect 6098 171878 6110 171930
rect 6172 171878 6174 171930
rect 6012 171876 6036 171878
rect 6092 171876 6116 171878
rect 6172 171876 6196 171878
rect 5956 171856 6252 171876
rect 5956 170844 6252 170864
rect 6012 170842 6036 170844
rect 6092 170842 6116 170844
rect 6172 170842 6196 170844
rect 6034 170790 6036 170842
rect 6098 170790 6110 170842
rect 6172 170790 6174 170842
rect 6012 170788 6036 170790
rect 6092 170788 6116 170790
rect 6172 170788 6196 170790
rect 5956 170768 6252 170788
rect 5956 169756 6252 169776
rect 6012 169754 6036 169756
rect 6092 169754 6116 169756
rect 6172 169754 6196 169756
rect 6034 169702 6036 169754
rect 6098 169702 6110 169754
rect 6172 169702 6174 169754
rect 6012 169700 6036 169702
rect 6092 169700 6116 169702
rect 6172 169700 6196 169702
rect 5956 169680 6252 169700
rect 5956 168668 6252 168688
rect 6012 168666 6036 168668
rect 6092 168666 6116 168668
rect 6172 168666 6196 168668
rect 6034 168614 6036 168666
rect 6098 168614 6110 168666
rect 6172 168614 6174 168666
rect 6012 168612 6036 168614
rect 6092 168612 6116 168614
rect 6172 168612 6196 168614
rect 5956 168592 6252 168612
rect 5956 167580 6252 167600
rect 6012 167578 6036 167580
rect 6092 167578 6116 167580
rect 6172 167578 6196 167580
rect 6034 167526 6036 167578
rect 6098 167526 6110 167578
rect 6172 167526 6174 167578
rect 6012 167524 6036 167526
rect 6092 167524 6116 167526
rect 6172 167524 6196 167526
rect 5956 167504 6252 167524
rect 5956 166492 6252 166512
rect 6012 166490 6036 166492
rect 6092 166490 6116 166492
rect 6172 166490 6196 166492
rect 6034 166438 6036 166490
rect 6098 166438 6110 166490
rect 6172 166438 6174 166490
rect 6012 166436 6036 166438
rect 6092 166436 6116 166438
rect 6172 166436 6196 166438
rect 5956 166416 6252 166436
rect 5956 165404 6252 165424
rect 6012 165402 6036 165404
rect 6092 165402 6116 165404
rect 6172 165402 6196 165404
rect 6034 165350 6036 165402
rect 6098 165350 6110 165402
rect 6172 165350 6174 165402
rect 6012 165348 6036 165350
rect 6092 165348 6116 165350
rect 6172 165348 6196 165350
rect 5956 165328 6252 165348
rect 5956 164316 6252 164336
rect 6012 164314 6036 164316
rect 6092 164314 6116 164316
rect 6172 164314 6196 164316
rect 6034 164262 6036 164314
rect 6098 164262 6110 164314
rect 6172 164262 6174 164314
rect 6012 164260 6036 164262
rect 6092 164260 6116 164262
rect 6172 164260 6196 164262
rect 5956 164240 6252 164260
rect 5956 163228 6252 163248
rect 6012 163226 6036 163228
rect 6092 163226 6116 163228
rect 6172 163226 6196 163228
rect 6034 163174 6036 163226
rect 6098 163174 6110 163226
rect 6172 163174 6174 163226
rect 6012 163172 6036 163174
rect 6092 163172 6116 163174
rect 6172 163172 6196 163174
rect 5956 163152 6252 163172
rect 5956 162140 6252 162160
rect 6012 162138 6036 162140
rect 6092 162138 6116 162140
rect 6172 162138 6196 162140
rect 6034 162086 6036 162138
rect 6098 162086 6110 162138
rect 6172 162086 6174 162138
rect 6012 162084 6036 162086
rect 6092 162084 6116 162086
rect 6172 162084 6196 162086
rect 5956 162064 6252 162084
rect 5956 161052 6252 161072
rect 6012 161050 6036 161052
rect 6092 161050 6116 161052
rect 6172 161050 6196 161052
rect 6034 160998 6036 161050
rect 6098 160998 6110 161050
rect 6172 160998 6174 161050
rect 6012 160996 6036 160998
rect 6092 160996 6116 160998
rect 6172 160996 6196 160998
rect 5956 160976 6252 160996
rect 5956 159964 6252 159984
rect 6012 159962 6036 159964
rect 6092 159962 6116 159964
rect 6172 159962 6196 159964
rect 6034 159910 6036 159962
rect 6098 159910 6110 159962
rect 6172 159910 6174 159962
rect 6012 159908 6036 159910
rect 6092 159908 6116 159910
rect 6172 159908 6196 159910
rect 5956 159888 6252 159908
rect 5956 158876 6252 158896
rect 6012 158874 6036 158876
rect 6092 158874 6116 158876
rect 6172 158874 6196 158876
rect 6034 158822 6036 158874
rect 6098 158822 6110 158874
rect 6172 158822 6174 158874
rect 6012 158820 6036 158822
rect 6092 158820 6116 158822
rect 6172 158820 6196 158822
rect 5956 158800 6252 158820
rect 5956 157788 6252 157808
rect 6012 157786 6036 157788
rect 6092 157786 6116 157788
rect 6172 157786 6196 157788
rect 6034 157734 6036 157786
rect 6098 157734 6110 157786
rect 6172 157734 6174 157786
rect 6012 157732 6036 157734
rect 6092 157732 6116 157734
rect 6172 157732 6196 157734
rect 5956 157712 6252 157732
rect 5956 156700 6252 156720
rect 6012 156698 6036 156700
rect 6092 156698 6116 156700
rect 6172 156698 6196 156700
rect 6034 156646 6036 156698
rect 6098 156646 6110 156698
rect 6172 156646 6174 156698
rect 6012 156644 6036 156646
rect 6092 156644 6116 156646
rect 6172 156644 6196 156646
rect 5956 156624 6252 156644
rect 5956 155612 6252 155632
rect 6012 155610 6036 155612
rect 6092 155610 6116 155612
rect 6172 155610 6196 155612
rect 6034 155558 6036 155610
rect 6098 155558 6110 155610
rect 6172 155558 6174 155610
rect 6012 155556 6036 155558
rect 6092 155556 6116 155558
rect 6172 155556 6196 155558
rect 5956 155536 6252 155556
rect 5956 154524 6252 154544
rect 6012 154522 6036 154524
rect 6092 154522 6116 154524
rect 6172 154522 6196 154524
rect 6034 154470 6036 154522
rect 6098 154470 6110 154522
rect 6172 154470 6174 154522
rect 6012 154468 6036 154470
rect 6092 154468 6116 154470
rect 6172 154468 6196 154470
rect 5956 154448 6252 154468
rect 5956 153436 6252 153456
rect 6012 153434 6036 153436
rect 6092 153434 6116 153436
rect 6172 153434 6196 153436
rect 6034 153382 6036 153434
rect 6098 153382 6110 153434
rect 6172 153382 6174 153434
rect 6012 153380 6036 153382
rect 6092 153380 6116 153382
rect 6172 153380 6196 153382
rect 5956 153360 6252 153380
rect 5956 152348 6252 152368
rect 6012 152346 6036 152348
rect 6092 152346 6116 152348
rect 6172 152346 6196 152348
rect 6034 152294 6036 152346
rect 6098 152294 6110 152346
rect 6172 152294 6174 152346
rect 6012 152292 6036 152294
rect 6092 152292 6116 152294
rect 6172 152292 6196 152294
rect 5956 152272 6252 152292
rect 5956 151260 6252 151280
rect 6012 151258 6036 151260
rect 6092 151258 6116 151260
rect 6172 151258 6196 151260
rect 6034 151206 6036 151258
rect 6098 151206 6110 151258
rect 6172 151206 6174 151258
rect 6012 151204 6036 151206
rect 6092 151204 6116 151206
rect 6172 151204 6196 151206
rect 5956 151184 6252 151204
rect 5956 150172 6252 150192
rect 6012 150170 6036 150172
rect 6092 150170 6116 150172
rect 6172 150170 6196 150172
rect 6034 150118 6036 150170
rect 6098 150118 6110 150170
rect 6172 150118 6174 150170
rect 6012 150116 6036 150118
rect 6092 150116 6116 150118
rect 6172 150116 6196 150118
rect 5956 150096 6252 150116
rect 5956 149084 6252 149104
rect 6012 149082 6036 149084
rect 6092 149082 6116 149084
rect 6172 149082 6196 149084
rect 6034 149030 6036 149082
rect 6098 149030 6110 149082
rect 6172 149030 6174 149082
rect 6012 149028 6036 149030
rect 6092 149028 6116 149030
rect 6172 149028 6196 149030
rect 5956 149008 6252 149028
rect 5956 147996 6252 148016
rect 6012 147994 6036 147996
rect 6092 147994 6116 147996
rect 6172 147994 6196 147996
rect 6034 147942 6036 147994
rect 6098 147942 6110 147994
rect 6172 147942 6174 147994
rect 6012 147940 6036 147942
rect 6092 147940 6116 147942
rect 6172 147940 6196 147942
rect 5956 147920 6252 147940
rect 5956 146908 6252 146928
rect 6012 146906 6036 146908
rect 6092 146906 6116 146908
rect 6172 146906 6196 146908
rect 6034 146854 6036 146906
rect 6098 146854 6110 146906
rect 6172 146854 6174 146906
rect 6012 146852 6036 146854
rect 6092 146852 6116 146854
rect 6172 146852 6196 146854
rect 5956 146832 6252 146852
rect 5956 145820 6252 145840
rect 6012 145818 6036 145820
rect 6092 145818 6116 145820
rect 6172 145818 6196 145820
rect 6034 145766 6036 145818
rect 6098 145766 6110 145818
rect 6172 145766 6174 145818
rect 6012 145764 6036 145766
rect 6092 145764 6116 145766
rect 6172 145764 6196 145766
rect 5956 145744 6252 145764
rect 5956 144732 6252 144752
rect 6012 144730 6036 144732
rect 6092 144730 6116 144732
rect 6172 144730 6196 144732
rect 6034 144678 6036 144730
rect 6098 144678 6110 144730
rect 6172 144678 6174 144730
rect 6012 144676 6036 144678
rect 6092 144676 6116 144678
rect 6172 144676 6196 144678
rect 5956 144656 6252 144676
rect 5956 143644 6252 143664
rect 6012 143642 6036 143644
rect 6092 143642 6116 143644
rect 6172 143642 6196 143644
rect 6034 143590 6036 143642
rect 6098 143590 6110 143642
rect 6172 143590 6174 143642
rect 6012 143588 6036 143590
rect 6092 143588 6116 143590
rect 6172 143588 6196 143590
rect 5956 143568 6252 143588
rect 5956 142556 6252 142576
rect 6012 142554 6036 142556
rect 6092 142554 6116 142556
rect 6172 142554 6196 142556
rect 6034 142502 6036 142554
rect 6098 142502 6110 142554
rect 6172 142502 6174 142554
rect 6012 142500 6036 142502
rect 6092 142500 6116 142502
rect 6172 142500 6196 142502
rect 5956 142480 6252 142500
rect 5956 141468 6252 141488
rect 6012 141466 6036 141468
rect 6092 141466 6116 141468
rect 6172 141466 6196 141468
rect 6034 141414 6036 141466
rect 6098 141414 6110 141466
rect 6172 141414 6174 141466
rect 6012 141412 6036 141414
rect 6092 141412 6116 141414
rect 6172 141412 6196 141414
rect 5956 141392 6252 141412
rect 5956 140380 6252 140400
rect 6012 140378 6036 140380
rect 6092 140378 6116 140380
rect 6172 140378 6196 140380
rect 6034 140326 6036 140378
rect 6098 140326 6110 140378
rect 6172 140326 6174 140378
rect 6012 140324 6036 140326
rect 6092 140324 6116 140326
rect 6172 140324 6196 140326
rect 5956 140304 6252 140324
rect 5956 139292 6252 139312
rect 6012 139290 6036 139292
rect 6092 139290 6116 139292
rect 6172 139290 6196 139292
rect 6034 139238 6036 139290
rect 6098 139238 6110 139290
rect 6172 139238 6174 139290
rect 6012 139236 6036 139238
rect 6092 139236 6116 139238
rect 6172 139236 6196 139238
rect 5956 139216 6252 139236
rect 5956 138204 6252 138224
rect 6012 138202 6036 138204
rect 6092 138202 6116 138204
rect 6172 138202 6196 138204
rect 6034 138150 6036 138202
rect 6098 138150 6110 138202
rect 6172 138150 6174 138202
rect 6012 138148 6036 138150
rect 6092 138148 6116 138150
rect 6172 138148 6196 138150
rect 5956 138128 6252 138148
rect 5956 137116 6252 137136
rect 6012 137114 6036 137116
rect 6092 137114 6116 137116
rect 6172 137114 6196 137116
rect 6034 137062 6036 137114
rect 6098 137062 6110 137114
rect 6172 137062 6174 137114
rect 6012 137060 6036 137062
rect 6092 137060 6116 137062
rect 6172 137060 6196 137062
rect 5956 137040 6252 137060
rect 5956 136028 6252 136048
rect 6012 136026 6036 136028
rect 6092 136026 6116 136028
rect 6172 136026 6196 136028
rect 6034 135974 6036 136026
rect 6098 135974 6110 136026
rect 6172 135974 6174 136026
rect 6012 135972 6036 135974
rect 6092 135972 6116 135974
rect 6172 135972 6196 135974
rect 5956 135952 6252 135972
rect 5956 134940 6252 134960
rect 6012 134938 6036 134940
rect 6092 134938 6116 134940
rect 6172 134938 6196 134940
rect 6034 134886 6036 134938
rect 6098 134886 6110 134938
rect 6172 134886 6174 134938
rect 6012 134884 6036 134886
rect 6092 134884 6116 134886
rect 6172 134884 6196 134886
rect 5956 134864 6252 134884
rect 5956 133852 6252 133872
rect 6012 133850 6036 133852
rect 6092 133850 6116 133852
rect 6172 133850 6196 133852
rect 6034 133798 6036 133850
rect 6098 133798 6110 133850
rect 6172 133798 6174 133850
rect 6012 133796 6036 133798
rect 6092 133796 6116 133798
rect 6172 133796 6196 133798
rect 5956 133776 6252 133796
rect 5956 132764 6252 132784
rect 6012 132762 6036 132764
rect 6092 132762 6116 132764
rect 6172 132762 6196 132764
rect 6034 132710 6036 132762
rect 6098 132710 6110 132762
rect 6172 132710 6174 132762
rect 6012 132708 6036 132710
rect 6092 132708 6116 132710
rect 6172 132708 6196 132710
rect 5956 132688 6252 132708
rect 5956 131676 6252 131696
rect 6012 131674 6036 131676
rect 6092 131674 6116 131676
rect 6172 131674 6196 131676
rect 6034 131622 6036 131674
rect 6098 131622 6110 131674
rect 6172 131622 6174 131674
rect 6012 131620 6036 131622
rect 6092 131620 6116 131622
rect 6172 131620 6196 131622
rect 5956 131600 6252 131620
rect 5956 130588 6252 130608
rect 6012 130586 6036 130588
rect 6092 130586 6116 130588
rect 6172 130586 6196 130588
rect 6034 130534 6036 130586
rect 6098 130534 6110 130586
rect 6172 130534 6174 130586
rect 6012 130532 6036 130534
rect 6092 130532 6116 130534
rect 6172 130532 6196 130534
rect 5956 130512 6252 130532
rect 5956 129500 6252 129520
rect 6012 129498 6036 129500
rect 6092 129498 6116 129500
rect 6172 129498 6196 129500
rect 6034 129446 6036 129498
rect 6098 129446 6110 129498
rect 6172 129446 6174 129498
rect 6012 129444 6036 129446
rect 6092 129444 6116 129446
rect 6172 129444 6196 129446
rect 5956 129424 6252 129444
rect 5956 128412 6252 128432
rect 6012 128410 6036 128412
rect 6092 128410 6116 128412
rect 6172 128410 6196 128412
rect 6034 128358 6036 128410
rect 6098 128358 6110 128410
rect 6172 128358 6174 128410
rect 6012 128356 6036 128358
rect 6092 128356 6116 128358
rect 6172 128356 6196 128358
rect 5956 128336 6252 128356
rect 5956 127324 6252 127344
rect 6012 127322 6036 127324
rect 6092 127322 6116 127324
rect 6172 127322 6196 127324
rect 6034 127270 6036 127322
rect 6098 127270 6110 127322
rect 6172 127270 6174 127322
rect 6012 127268 6036 127270
rect 6092 127268 6116 127270
rect 6172 127268 6196 127270
rect 5956 127248 6252 127268
rect 5956 126236 6252 126256
rect 6012 126234 6036 126236
rect 6092 126234 6116 126236
rect 6172 126234 6196 126236
rect 6034 126182 6036 126234
rect 6098 126182 6110 126234
rect 6172 126182 6174 126234
rect 6012 126180 6036 126182
rect 6092 126180 6116 126182
rect 6172 126180 6196 126182
rect 5956 126160 6252 126180
rect 5956 125148 6252 125168
rect 6012 125146 6036 125148
rect 6092 125146 6116 125148
rect 6172 125146 6196 125148
rect 6034 125094 6036 125146
rect 6098 125094 6110 125146
rect 6172 125094 6174 125146
rect 6012 125092 6036 125094
rect 6092 125092 6116 125094
rect 6172 125092 6196 125094
rect 5956 125072 6252 125092
rect 5956 124060 6252 124080
rect 6012 124058 6036 124060
rect 6092 124058 6116 124060
rect 6172 124058 6196 124060
rect 6034 124006 6036 124058
rect 6098 124006 6110 124058
rect 6172 124006 6174 124058
rect 6012 124004 6036 124006
rect 6092 124004 6116 124006
rect 6172 124004 6196 124006
rect 5956 123984 6252 124004
rect 5956 122972 6252 122992
rect 6012 122970 6036 122972
rect 6092 122970 6116 122972
rect 6172 122970 6196 122972
rect 6034 122918 6036 122970
rect 6098 122918 6110 122970
rect 6172 122918 6174 122970
rect 6012 122916 6036 122918
rect 6092 122916 6116 122918
rect 6172 122916 6196 122918
rect 5956 122896 6252 122916
rect 5956 121884 6252 121904
rect 6012 121882 6036 121884
rect 6092 121882 6116 121884
rect 6172 121882 6196 121884
rect 6034 121830 6036 121882
rect 6098 121830 6110 121882
rect 6172 121830 6174 121882
rect 6012 121828 6036 121830
rect 6092 121828 6116 121830
rect 6172 121828 6196 121830
rect 5956 121808 6252 121828
rect 5956 120796 6252 120816
rect 6012 120794 6036 120796
rect 6092 120794 6116 120796
rect 6172 120794 6196 120796
rect 6034 120742 6036 120794
rect 6098 120742 6110 120794
rect 6172 120742 6174 120794
rect 6012 120740 6036 120742
rect 6092 120740 6116 120742
rect 6172 120740 6196 120742
rect 5956 120720 6252 120740
rect 5956 119708 6252 119728
rect 6012 119706 6036 119708
rect 6092 119706 6116 119708
rect 6172 119706 6196 119708
rect 6034 119654 6036 119706
rect 6098 119654 6110 119706
rect 6172 119654 6174 119706
rect 6012 119652 6036 119654
rect 6092 119652 6116 119654
rect 6172 119652 6196 119654
rect 5956 119632 6252 119652
rect 5956 118620 6252 118640
rect 6012 118618 6036 118620
rect 6092 118618 6116 118620
rect 6172 118618 6196 118620
rect 6034 118566 6036 118618
rect 6098 118566 6110 118618
rect 6172 118566 6174 118618
rect 6012 118564 6036 118566
rect 6092 118564 6116 118566
rect 6172 118564 6196 118566
rect 5956 118544 6252 118564
rect 5956 117532 6252 117552
rect 6012 117530 6036 117532
rect 6092 117530 6116 117532
rect 6172 117530 6196 117532
rect 6034 117478 6036 117530
rect 6098 117478 6110 117530
rect 6172 117478 6174 117530
rect 6012 117476 6036 117478
rect 6092 117476 6116 117478
rect 6172 117476 6196 117478
rect 5956 117456 6252 117476
rect 6748 116793 6776 211686
rect 7024 211002 7052 216135
rect 7300 214266 7328 315823
rect 8036 315178 8064 332438
rect 7380 315172 7432 315178
rect 7380 315114 7432 315120
rect 8024 315172 8076 315178
rect 8024 315114 8076 315120
rect 7392 242010 7420 315114
rect 7622 315004 7918 315024
rect 7678 315002 7702 315004
rect 7758 315002 7782 315004
rect 7838 315002 7862 315004
rect 7700 314950 7702 315002
rect 7764 314950 7776 315002
rect 7838 314950 7840 315002
rect 7678 314948 7702 314950
rect 7758 314948 7782 314950
rect 7838 314948 7862 314950
rect 7622 314928 7918 314948
rect 7622 313916 7918 313936
rect 7678 313914 7702 313916
rect 7758 313914 7782 313916
rect 7838 313914 7862 313916
rect 7700 313862 7702 313914
rect 7764 313862 7776 313914
rect 7838 313862 7840 313914
rect 7678 313860 7702 313862
rect 7758 313860 7782 313862
rect 7838 313860 7862 313862
rect 7622 313840 7918 313860
rect 7622 312828 7918 312848
rect 7678 312826 7702 312828
rect 7758 312826 7782 312828
rect 7838 312826 7862 312828
rect 7700 312774 7702 312826
rect 7764 312774 7776 312826
rect 7838 312774 7840 312826
rect 7678 312772 7702 312774
rect 7758 312772 7782 312774
rect 7838 312772 7862 312774
rect 7622 312752 7918 312772
rect 7622 311740 7918 311760
rect 7678 311738 7702 311740
rect 7758 311738 7782 311740
rect 7838 311738 7862 311740
rect 7700 311686 7702 311738
rect 7764 311686 7776 311738
rect 7838 311686 7840 311738
rect 7678 311684 7702 311686
rect 7758 311684 7782 311686
rect 7838 311684 7862 311686
rect 7622 311664 7918 311684
rect 7622 310652 7918 310672
rect 7678 310650 7702 310652
rect 7758 310650 7782 310652
rect 7838 310650 7862 310652
rect 7700 310598 7702 310650
rect 7764 310598 7776 310650
rect 7838 310598 7840 310650
rect 7678 310596 7702 310598
rect 7758 310596 7782 310598
rect 7838 310596 7862 310598
rect 7622 310576 7918 310596
rect 7622 309564 7918 309584
rect 7678 309562 7702 309564
rect 7758 309562 7782 309564
rect 7838 309562 7862 309564
rect 7700 309510 7702 309562
rect 7764 309510 7776 309562
rect 7838 309510 7840 309562
rect 7678 309508 7702 309510
rect 7758 309508 7782 309510
rect 7838 309508 7862 309510
rect 7622 309488 7918 309508
rect 7622 308476 7918 308496
rect 7678 308474 7702 308476
rect 7758 308474 7782 308476
rect 7838 308474 7862 308476
rect 7700 308422 7702 308474
rect 7764 308422 7776 308474
rect 7838 308422 7840 308474
rect 7678 308420 7702 308422
rect 7758 308420 7782 308422
rect 7838 308420 7862 308422
rect 7622 308400 7918 308420
rect 7622 307388 7918 307408
rect 7678 307386 7702 307388
rect 7758 307386 7782 307388
rect 7838 307386 7862 307388
rect 7700 307334 7702 307386
rect 7764 307334 7776 307386
rect 7838 307334 7840 307386
rect 7678 307332 7702 307334
rect 7758 307332 7782 307334
rect 7838 307332 7862 307334
rect 7622 307312 7918 307332
rect 7622 306300 7918 306320
rect 7678 306298 7702 306300
rect 7758 306298 7782 306300
rect 7838 306298 7862 306300
rect 7700 306246 7702 306298
rect 7764 306246 7776 306298
rect 7838 306246 7840 306298
rect 7678 306244 7702 306246
rect 7758 306244 7782 306246
rect 7838 306244 7862 306246
rect 7622 306224 7918 306244
rect 7622 305212 7918 305232
rect 7678 305210 7702 305212
rect 7758 305210 7782 305212
rect 7838 305210 7862 305212
rect 7700 305158 7702 305210
rect 7764 305158 7776 305210
rect 7838 305158 7840 305210
rect 7678 305156 7702 305158
rect 7758 305156 7782 305158
rect 7838 305156 7862 305158
rect 7622 305136 7918 305156
rect 7622 304124 7918 304144
rect 7678 304122 7702 304124
rect 7758 304122 7782 304124
rect 7838 304122 7862 304124
rect 7700 304070 7702 304122
rect 7764 304070 7776 304122
rect 7838 304070 7840 304122
rect 7678 304068 7702 304070
rect 7758 304068 7782 304070
rect 7838 304068 7862 304070
rect 7622 304048 7918 304068
rect 7622 303036 7918 303056
rect 7678 303034 7702 303036
rect 7758 303034 7782 303036
rect 7838 303034 7862 303036
rect 7700 302982 7702 303034
rect 7764 302982 7776 303034
rect 7838 302982 7840 303034
rect 7678 302980 7702 302982
rect 7758 302980 7782 302982
rect 7838 302980 7862 302982
rect 7622 302960 7918 302980
rect 7622 301948 7918 301968
rect 7678 301946 7702 301948
rect 7758 301946 7782 301948
rect 7838 301946 7862 301948
rect 7700 301894 7702 301946
rect 7764 301894 7776 301946
rect 7838 301894 7840 301946
rect 7678 301892 7702 301894
rect 7758 301892 7782 301894
rect 7838 301892 7862 301894
rect 7622 301872 7918 301892
rect 7622 300860 7918 300880
rect 7678 300858 7702 300860
rect 7758 300858 7782 300860
rect 7838 300858 7862 300860
rect 7700 300806 7702 300858
rect 7764 300806 7776 300858
rect 7838 300806 7840 300858
rect 7678 300804 7702 300806
rect 7758 300804 7782 300806
rect 7838 300804 7862 300806
rect 7622 300784 7918 300804
rect 7622 299772 7918 299792
rect 7678 299770 7702 299772
rect 7758 299770 7782 299772
rect 7838 299770 7862 299772
rect 7700 299718 7702 299770
rect 7764 299718 7776 299770
rect 7838 299718 7840 299770
rect 7678 299716 7702 299718
rect 7758 299716 7782 299718
rect 7838 299716 7862 299718
rect 7622 299696 7918 299716
rect 7622 298684 7918 298704
rect 7678 298682 7702 298684
rect 7758 298682 7782 298684
rect 7838 298682 7862 298684
rect 7700 298630 7702 298682
rect 7764 298630 7776 298682
rect 7838 298630 7840 298682
rect 7678 298628 7702 298630
rect 7758 298628 7782 298630
rect 7838 298628 7862 298630
rect 7622 298608 7918 298628
rect 7622 297596 7918 297616
rect 7678 297594 7702 297596
rect 7758 297594 7782 297596
rect 7838 297594 7862 297596
rect 7700 297542 7702 297594
rect 7764 297542 7776 297594
rect 7838 297542 7840 297594
rect 7678 297540 7702 297542
rect 7758 297540 7782 297542
rect 7838 297540 7862 297542
rect 7622 297520 7918 297540
rect 7622 296508 7918 296528
rect 7678 296506 7702 296508
rect 7758 296506 7782 296508
rect 7838 296506 7862 296508
rect 7700 296454 7702 296506
rect 7764 296454 7776 296506
rect 7838 296454 7840 296506
rect 7678 296452 7702 296454
rect 7758 296452 7782 296454
rect 7838 296452 7862 296454
rect 7622 296432 7918 296452
rect 7622 295420 7918 295440
rect 7678 295418 7702 295420
rect 7758 295418 7782 295420
rect 7838 295418 7862 295420
rect 7700 295366 7702 295418
rect 7764 295366 7776 295418
rect 7838 295366 7840 295418
rect 7678 295364 7702 295366
rect 7758 295364 7782 295366
rect 7838 295364 7862 295366
rect 7622 295344 7918 295364
rect 7622 294332 7918 294352
rect 7678 294330 7702 294332
rect 7758 294330 7782 294332
rect 7838 294330 7862 294332
rect 7700 294278 7702 294330
rect 7764 294278 7776 294330
rect 7838 294278 7840 294330
rect 7678 294276 7702 294278
rect 7758 294276 7782 294278
rect 7838 294276 7862 294278
rect 7622 294256 7918 294276
rect 7622 293244 7918 293264
rect 7678 293242 7702 293244
rect 7758 293242 7782 293244
rect 7838 293242 7862 293244
rect 7700 293190 7702 293242
rect 7764 293190 7776 293242
rect 7838 293190 7840 293242
rect 7678 293188 7702 293190
rect 7758 293188 7782 293190
rect 7838 293188 7862 293190
rect 7622 293168 7918 293188
rect 7622 292156 7918 292176
rect 7678 292154 7702 292156
rect 7758 292154 7782 292156
rect 7838 292154 7862 292156
rect 7700 292102 7702 292154
rect 7764 292102 7776 292154
rect 7838 292102 7840 292154
rect 7678 292100 7702 292102
rect 7758 292100 7782 292102
rect 7838 292100 7862 292102
rect 7622 292080 7918 292100
rect 7622 291068 7918 291088
rect 7678 291066 7702 291068
rect 7758 291066 7782 291068
rect 7838 291066 7862 291068
rect 7700 291014 7702 291066
rect 7764 291014 7776 291066
rect 7838 291014 7840 291066
rect 7678 291012 7702 291014
rect 7758 291012 7782 291014
rect 7838 291012 7862 291014
rect 7622 290992 7918 291012
rect 7622 289980 7918 290000
rect 7678 289978 7702 289980
rect 7758 289978 7782 289980
rect 7838 289978 7862 289980
rect 7700 289926 7702 289978
rect 7764 289926 7776 289978
rect 7838 289926 7840 289978
rect 7678 289924 7702 289926
rect 7758 289924 7782 289926
rect 7838 289924 7862 289926
rect 7622 289904 7918 289924
rect 7622 288892 7918 288912
rect 7678 288890 7702 288892
rect 7758 288890 7782 288892
rect 7838 288890 7862 288892
rect 7700 288838 7702 288890
rect 7764 288838 7776 288890
rect 7838 288838 7840 288890
rect 7678 288836 7702 288838
rect 7758 288836 7782 288838
rect 7838 288836 7862 288838
rect 7622 288816 7918 288836
rect 7622 287804 7918 287824
rect 7678 287802 7702 287804
rect 7758 287802 7782 287804
rect 7838 287802 7862 287804
rect 7700 287750 7702 287802
rect 7764 287750 7776 287802
rect 7838 287750 7840 287802
rect 7678 287748 7702 287750
rect 7758 287748 7782 287750
rect 7838 287748 7862 287750
rect 7622 287728 7918 287748
rect 7622 286716 7918 286736
rect 7678 286714 7702 286716
rect 7758 286714 7782 286716
rect 7838 286714 7862 286716
rect 7700 286662 7702 286714
rect 7764 286662 7776 286714
rect 7838 286662 7840 286714
rect 7678 286660 7702 286662
rect 7758 286660 7782 286662
rect 7838 286660 7862 286662
rect 7622 286640 7918 286660
rect 7622 285628 7918 285648
rect 7678 285626 7702 285628
rect 7758 285626 7782 285628
rect 7838 285626 7862 285628
rect 7700 285574 7702 285626
rect 7764 285574 7776 285626
rect 7838 285574 7840 285626
rect 7678 285572 7702 285574
rect 7758 285572 7782 285574
rect 7838 285572 7862 285574
rect 7622 285552 7918 285572
rect 7622 284540 7918 284560
rect 7678 284538 7702 284540
rect 7758 284538 7782 284540
rect 7838 284538 7862 284540
rect 7700 284486 7702 284538
rect 7764 284486 7776 284538
rect 7838 284486 7840 284538
rect 7678 284484 7702 284486
rect 7758 284484 7782 284486
rect 7838 284484 7862 284486
rect 7622 284464 7918 284484
rect 7622 283452 7918 283472
rect 7678 283450 7702 283452
rect 7758 283450 7782 283452
rect 7838 283450 7862 283452
rect 7700 283398 7702 283450
rect 7764 283398 7776 283450
rect 7838 283398 7840 283450
rect 7678 283396 7702 283398
rect 7758 283396 7782 283398
rect 7838 283396 7862 283398
rect 7622 283376 7918 283396
rect 7622 282364 7918 282384
rect 7678 282362 7702 282364
rect 7758 282362 7782 282364
rect 7838 282362 7862 282364
rect 7700 282310 7702 282362
rect 7764 282310 7776 282362
rect 7838 282310 7840 282362
rect 7678 282308 7702 282310
rect 7758 282308 7782 282310
rect 7838 282308 7862 282310
rect 7622 282288 7918 282308
rect 7622 281276 7918 281296
rect 7678 281274 7702 281276
rect 7758 281274 7782 281276
rect 7838 281274 7862 281276
rect 7700 281222 7702 281274
rect 7764 281222 7776 281274
rect 7838 281222 7840 281274
rect 7678 281220 7702 281222
rect 7758 281220 7782 281222
rect 7838 281220 7862 281222
rect 7622 281200 7918 281220
rect 7622 280188 7918 280208
rect 7678 280186 7702 280188
rect 7758 280186 7782 280188
rect 7838 280186 7862 280188
rect 7700 280134 7702 280186
rect 7764 280134 7776 280186
rect 7838 280134 7840 280186
rect 7678 280132 7702 280134
rect 7758 280132 7782 280134
rect 7838 280132 7862 280134
rect 7622 280112 7918 280132
rect 7622 279100 7918 279120
rect 7678 279098 7702 279100
rect 7758 279098 7782 279100
rect 7838 279098 7862 279100
rect 7700 279046 7702 279098
rect 7764 279046 7776 279098
rect 7838 279046 7840 279098
rect 7678 279044 7702 279046
rect 7758 279044 7782 279046
rect 7838 279044 7862 279046
rect 7622 279024 7918 279044
rect 7622 278012 7918 278032
rect 7678 278010 7702 278012
rect 7758 278010 7782 278012
rect 7838 278010 7862 278012
rect 7700 277958 7702 278010
rect 7764 277958 7776 278010
rect 7838 277958 7840 278010
rect 7678 277956 7702 277958
rect 7758 277956 7782 277958
rect 7838 277956 7862 277958
rect 7622 277936 7918 277956
rect 7622 276924 7918 276944
rect 7678 276922 7702 276924
rect 7758 276922 7782 276924
rect 7838 276922 7862 276924
rect 7700 276870 7702 276922
rect 7764 276870 7776 276922
rect 7838 276870 7840 276922
rect 7678 276868 7702 276870
rect 7758 276868 7782 276870
rect 7838 276868 7862 276870
rect 7622 276848 7918 276868
rect 7622 275836 7918 275856
rect 7678 275834 7702 275836
rect 7758 275834 7782 275836
rect 7838 275834 7862 275836
rect 7700 275782 7702 275834
rect 7764 275782 7776 275834
rect 7838 275782 7840 275834
rect 7678 275780 7702 275782
rect 7758 275780 7782 275782
rect 7838 275780 7862 275782
rect 7622 275760 7918 275780
rect 7622 274748 7918 274768
rect 7678 274746 7702 274748
rect 7758 274746 7782 274748
rect 7838 274746 7862 274748
rect 7700 274694 7702 274746
rect 7764 274694 7776 274746
rect 7838 274694 7840 274746
rect 7678 274692 7702 274694
rect 7758 274692 7782 274694
rect 7838 274692 7862 274694
rect 7622 274672 7918 274692
rect 7622 273660 7918 273680
rect 7678 273658 7702 273660
rect 7758 273658 7782 273660
rect 7838 273658 7862 273660
rect 7700 273606 7702 273658
rect 7764 273606 7776 273658
rect 7838 273606 7840 273658
rect 7678 273604 7702 273606
rect 7758 273604 7782 273606
rect 7838 273604 7862 273606
rect 7622 273584 7918 273604
rect 7622 272572 7918 272592
rect 7678 272570 7702 272572
rect 7758 272570 7782 272572
rect 7838 272570 7862 272572
rect 7700 272518 7702 272570
rect 7764 272518 7776 272570
rect 7838 272518 7840 272570
rect 7678 272516 7702 272518
rect 7758 272516 7782 272518
rect 7838 272516 7862 272518
rect 7622 272496 7918 272516
rect 7622 271484 7918 271504
rect 7678 271482 7702 271484
rect 7758 271482 7782 271484
rect 7838 271482 7862 271484
rect 7700 271430 7702 271482
rect 7764 271430 7776 271482
rect 7838 271430 7840 271482
rect 7678 271428 7702 271430
rect 7758 271428 7782 271430
rect 7838 271428 7862 271430
rect 7622 271408 7918 271428
rect 7622 270396 7918 270416
rect 7678 270394 7702 270396
rect 7758 270394 7782 270396
rect 7838 270394 7862 270396
rect 7700 270342 7702 270394
rect 7764 270342 7776 270394
rect 7838 270342 7840 270394
rect 7678 270340 7702 270342
rect 7758 270340 7782 270342
rect 7838 270340 7862 270342
rect 7622 270320 7918 270340
rect 7622 269308 7918 269328
rect 7678 269306 7702 269308
rect 7758 269306 7782 269308
rect 7838 269306 7862 269308
rect 7700 269254 7702 269306
rect 7764 269254 7776 269306
rect 7838 269254 7840 269306
rect 7678 269252 7702 269254
rect 7758 269252 7782 269254
rect 7838 269252 7862 269254
rect 7622 269232 7918 269252
rect 7622 268220 7918 268240
rect 7678 268218 7702 268220
rect 7758 268218 7782 268220
rect 7838 268218 7862 268220
rect 7700 268166 7702 268218
rect 7764 268166 7776 268218
rect 7838 268166 7840 268218
rect 7678 268164 7702 268166
rect 7758 268164 7782 268166
rect 7838 268164 7862 268166
rect 7622 268144 7918 268164
rect 7622 267132 7918 267152
rect 7678 267130 7702 267132
rect 7758 267130 7782 267132
rect 7838 267130 7862 267132
rect 7700 267078 7702 267130
rect 7764 267078 7776 267130
rect 7838 267078 7840 267130
rect 7678 267076 7702 267078
rect 7758 267076 7782 267078
rect 7838 267076 7862 267078
rect 7622 267056 7918 267076
rect 7622 266044 7918 266064
rect 7678 266042 7702 266044
rect 7758 266042 7782 266044
rect 7838 266042 7862 266044
rect 7700 265990 7702 266042
rect 7764 265990 7776 266042
rect 7838 265990 7840 266042
rect 7678 265988 7702 265990
rect 7758 265988 7782 265990
rect 7838 265988 7862 265990
rect 7622 265968 7918 265988
rect 7622 264956 7918 264976
rect 7678 264954 7702 264956
rect 7758 264954 7782 264956
rect 7838 264954 7862 264956
rect 7700 264902 7702 264954
rect 7764 264902 7776 264954
rect 7838 264902 7840 264954
rect 7678 264900 7702 264902
rect 7758 264900 7782 264902
rect 7838 264900 7862 264902
rect 7622 264880 7918 264900
rect 7622 263868 7918 263888
rect 7678 263866 7702 263868
rect 7758 263866 7782 263868
rect 7838 263866 7862 263868
rect 7700 263814 7702 263866
rect 7764 263814 7776 263866
rect 7838 263814 7840 263866
rect 7678 263812 7702 263814
rect 7758 263812 7782 263814
rect 7838 263812 7862 263814
rect 7622 263792 7918 263812
rect 7622 262780 7918 262800
rect 7678 262778 7702 262780
rect 7758 262778 7782 262780
rect 7838 262778 7862 262780
rect 7700 262726 7702 262778
rect 7764 262726 7776 262778
rect 7838 262726 7840 262778
rect 7678 262724 7702 262726
rect 7758 262724 7782 262726
rect 7838 262724 7862 262726
rect 7622 262704 7918 262724
rect 7622 261692 7918 261712
rect 7678 261690 7702 261692
rect 7758 261690 7782 261692
rect 7838 261690 7862 261692
rect 7700 261638 7702 261690
rect 7764 261638 7776 261690
rect 7838 261638 7840 261690
rect 7678 261636 7702 261638
rect 7758 261636 7782 261638
rect 7838 261636 7862 261638
rect 7622 261616 7918 261636
rect 7622 260604 7918 260624
rect 7678 260602 7702 260604
rect 7758 260602 7782 260604
rect 7838 260602 7862 260604
rect 7700 260550 7702 260602
rect 7764 260550 7776 260602
rect 7838 260550 7840 260602
rect 7678 260548 7702 260550
rect 7758 260548 7782 260550
rect 7838 260548 7862 260550
rect 7622 260528 7918 260548
rect 7622 259516 7918 259536
rect 7678 259514 7702 259516
rect 7758 259514 7782 259516
rect 7838 259514 7862 259516
rect 7700 259462 7702 259514
rect 7764 259462 7776 259514
rect 7838 259462 7840 259514
rect 7678 259460 7702 259462
rect 7758 259460 7782 259462
rect 7838 259460 7862 259462
rect 7622 259440 7918 259460
rect 7622 258428 7918 258448
rect 7678 258426 7702 258428
rect 7758 258426 7782 258428
rect 7838 258426 7862 258428
rect 7700 258374 7702 258426
rect 7764 258374 7776 258426
rect 7838 258374 7840 258426
rect 7678 258372 7702 258374
rect 7758 258372 7782 258374
rect 7838 258372 7862 258374
rect 7622 258352 7918 258372
rect 7622 257340 7918 257360
rect 7678 257338 7702 257340
rect 7758 257338 7782 257340
rect 7838 257338 7862 257340
rect 7700 257286 7702 257338
rect 7764 257286 7776 257338
rect 7838 257286 7840 257338
rect 7678 257284 7702 257286
rect 7758 257284 7782 257286
rect 7838 257284 7862 257286
rect 7622 257264 7918 257284
rect 7622 256252 7918 256272
rect 7678 256250 7702 256252
rect 7758 256250 7782 256252
rect 7838 256250 7862 256252
rect 7700 256198 7702 256250
rect 7764 256198 7776 256250
rect 7838 256198 7840 256250
rect 7678 256196 7702 256198
rect 7758 256196 7782 256198
rect 7838 256196 7862 256198
rect 7622 256176 7918 256196
rect 7622 255164 7918 255184
rect 7678 255162 7702 255164
rect 7758 255162 7782 255164
rect 7838 255162 7862 255164
rect 7700 255110 7702 255162
rect 7764 255110 7776 255162
rect 7838 255110 7840 255162
rect 7678 255108 7702 255110
rect 7758 255108 7782 255110
rect 7838 255108 7862 255110
rect 7622 255088 7918 255108
rect 7622 254076 7918 254096
rect 7678 254074 7702 254076
rect 7758 254074 7782 254076
rect 7838 254074 7862 254076
rect 7700 254022 7702 254074
rect 7764 254022 7776 254074
rect 7838 254022 7840 254074
rect 7678 254020 7702 254022
rect 7758 254020 7782 254022
rect 7838 254020 7862 254022
rect 7622 254000 7918 254020
rect 7622 252988 7918 253008
rect 7678 252986 7702 252988
rect 7758 252986 7782 252988
rect 7838 252986 7862 252988
rect 7700 252934 7702 252986
rect 7764 252934 7776 252986
rect 7838 252934 7840 252986
rect 7678 252932 7702 252934
rect 7758 252932 7782 252934
rect 7838 252932 7862 252934
rect 7622 252912 7918 252932
rect 7622 251900 7918 251920
rect 7678 251898 7702 251900
rect 7758 251898 7782 251900
rect 7838 251898 7862 251900
rect 7700 251846 7702 251898
rect 7764 251846 7776 251898
rect 7838 251846 7840 251898
rect 7678 251844 7702 251846
rect 7758 251844 7782 251846
rect 7838 251844 7862 251846
rect 7622 251824 7918 251844
rect 7622 250812 7918 250832
rect 7678 250810 7702 250812
rect 7758 250810 7782 250812
rect 7838 250810 7862 250812
rect 7700 250758 7702 250810
rect 7764 250758 7776 250810
rect 7838 250758 7840 250810
rect 7678 250756 7702 250758
rect 7758 250756 7782 250758
rect 7838 250756 7862 250758
rect 7622 250736 7918 250756
rect 7622 249724 7918 249744
rect 7678 249722 7702 249724
rect 7758 249722 7782 249724
rect 7838 249722 7862 249724
rect 7700 249670 7702 249722
rect 7764 249670 7776 249722
rect 7838 249670 7840 249722
rect 7678 249668 7702 249670
rect 7758 249668 7782 249670
rect 7838 249668 7862 249670
rect 7622 249648 7918 249668
rect 7622 248636 7918 248656
rect 7678 248634 7702 248636
rect 7758 248634 7782 248636
rect 7838 248634 7862 248636
rect 7700 248582 7702 248634
rect 7764 248582 7776 248634
rect 7838 248582 7840 248634
rect 7678 248580 7702 248582
rect 7758 248580 7782 248582
rect 7838 248580 7862 248582
rect 7622 248560 7918 248580
rect 7622 247548 7918 247568
rect 7678 247546 7702 247548
rect 7758 247546 7782 247548
rect 7838 247546 7862 247548
rect 7700 247494 7702 247546
rect 7764 247494 7776 247546
rect 7838 247494 7840 247546
rect 7678 247492 7702 247494
rect 7758 247492 7782 247494
rect 7838 247492 7862 247494
rect 7622 247472 7918 247492
rect 7622 246460 7918 246480
rect 7678 246458 7702 246460
rect 7758 246458 7782 246460
rect 7838 246458 7862 246460
rect 7700 246406 7702 246458
rect 7764 246406 7776 246458
rect 7838 246406 7840 246458
rect 7678 246404 7702 246406
rect 7758 246404 7782 246406
rect 7838 246404 7862 246406
rect 7622 246384 7918 246404
rect 7622 245372 7918 245392
rect 7678 245370 7702 245372
rect 7758 245370 7782 245372
rect 7838 245370 7862 245372
rect 7700 245318 7702 245370
rect 7764 245318 7776 245370
rect 7838 245318 7840 245370
rect 7678 245316 7702 245318
rect 7758 245316 7782 245318
rect 7838 245316 7862 245318
rect 7622 245296 7918 245316
rect 7622 244284 7918 244304
rect 7678 244282 7702 244284
rect 7758 244282 7782 244284
rect 7838 244282 7862 244284
rect 7700 244230 7702 244282
rect 7764 244230 7776 244282
rect 7838 244230 7840 244282
rect 7678 244228 7702 244230
rect 7758 244228 7782 244230
rect 7838 244228 7862 244230
rect 7622 244208 7918 244228
rect 7622 243196 7918 243216
rect 7678 243194 7702 243196
rect 7758 243194 7782 243196
rect 7838 243194 7862 243196
rect 7700 243142 7702 243194
rect 7764 243142 7776 243194
rect 7838 243142 7840 243194
rect 7678 243140 7702 243142
rect 7758 243140 7782 243142
rect 7838 243140 7862 243142
rect 7622 243120 7918 243140
rect 7622 242108 7918 242128
rect 7678 242106 7702 242108
rect 7758 242106 7782 242108
rect 7838 242106 7862 242108
rect 7700 242054 7702 242106
rect 7764 242054 7776 242106
rect 7838 242054 7840 242106
rect 7678 242052 7702 242054
rect 7758 242052 7782 242054
rect 7838 242052 7862 242054
rect 7622 242032 7918 242052
rect 7380 242004 7432 242010
rect 7380 241946 7432 241952
rect 7472 241868 7524 241874
rect 7472 241810 7524 241816
rect 7484 241126 7512 241810
rect 7472 241120 7524 241126
rect 7472 241062 7524 241068
rect 7484 234054 7512 241062
rect 7622 241020 7918 241040
rect 7678 241018 7702 241020
rect 7758 241018 7782 241020
rect 7838 241018 7862 241020
rect 7700 240966 7702 241018
rect 7764 240966 7776 241018
rect 7838 240966 7840 241018
rect 7678 240964 7702 240966
rect 7758 240964 7782 240966
rect 7838 240964 7862 240966
rect 7622 240944 7918 240964
rect 7622 239932 7918 239952
rect 7678 239930 7702 239932
rect 7758 239930 7782 239932
rect 7838 239930 7862 239932
rect 7700 239878 7702 239930
rect 7764 239878 7776 239930
rect 7838 239878 7840 239930
rect 7678 239876 7702 239878
rect 7758 239876 7782 239878
rect 7838 239876 7862 239878
rect 7622 239856 7918 239876
rect 7622 238844 7918 238864
rect 7678 238842 7702 238844
rect 7758 238842 7782 238844
rect 7838 238842 7862 238844
rect 7700 238790 7702 238842
rect 7764 238790 7776 238842
rect 7838 238790 7840 238842
rect 7678 238788 7702 238790
rect 7758 238788 7782 238790
rect 7838 238788 7862 238790
rect 7622 238768 7918 238788
rect 7622 237756 7918 237776
rect 7678 237754 7702 237756
rect 7758 237754 7782 237756
rect 7838 237754 7862 237756
rect 7700 237702 7702 237754
rect 7764 237702 7776 237754
rect 7838 237702 7840 237754
rect 7678 237700 7702 237702
rect 7758 237700 7782 237702
rect 7838 237700 7862 237702
rect 7622 237680 7918 237700
rect 7622 236668 7918 236688
rect 7678 236666 7702 236668
rect 7758 236666 7782 236668
rect 7838 236666 7862 236668
rect 7700 236614 7702 236666
rect 7764 236614 7776 236666
rect 7838 236614 7840 236666
rect 7678 236612 7702 236614
rect 7758 236612 7782 236614
rect 7838 236612 7862 236614
rect 7622 236592 7918 236612
rect 7622 235580 7918 235600
rect 7678 235578 7702 235580
rect 7758 235578 7782 235580
rect 7838 235578 7862 235580
rect 7700 235526 7702 235578
rect 7764 235526 7776 235578
rect 7838 235526 7840 235578
rect 7678 235524 7702 235526
rect 7758 235524 7782 235526
rect 7838 235524 7862 235526
rect 7622 235504 7918 235524
rect 7622 234492 7918 234512
rect 7678 234490 7702 234492
rect 7758 234490 7782 234492
rect 7838 234490 7862 234492
rect 7700 234438 7702 234490
rect 7764 234438 7776 234490
rect 7838 234438 7840 234490
rect 7678 234436 7702 234438
rect 7758 234436 7782 234438
rect 7838 234436 7862 234438
rect 7622 234416 7918 234436
rect 7472 234048 7524 234054
rect 7472 233990 7524 233996
rect 8208 234048 8260 234054
rect 8208 233990 8260 233996
rect 7622 233404 7918 233424
rect 7678 233402 7702 233404
rect 7758 233402 7782 233404
rect 7838 233402 7862 233404
rect 7700 233350 7702 233402
rect 7764 233350 7776 233402
rect 7838 233350 7840 233402
rect 7678 233348 7702 233350
rect 7758 233348 7782 233350
rect 7838 233348 7862 233350
rect 7622 233328 7918 233348
rect 7622 232316 7918 232336
rect 7678 232314 7702 232316
rect 7758 232314 7782 232316
rect 7838 232314 7862 232316
rect 7700 232262 7702 232314
rect 7764 232262 7776 232314
rect 7838 232262 7840 232314
rect 7678 232260 7702 232262
rect 7758 232260 7782 232262
rect 7838 232260 7862 232262
rect 7622 232240 7918 232260
rect 7622 231228 7918 231248
rect 7678 231226 7702 231228
rect 7758 231226 7782 231228
rect 7838 231226 7862 231228
rect 7700 231174 7702 231226
rect 7764 231174 7776 231226
rect 7838 231174 7840 231226
rect 7678 231172 7702 231174
rect 7758 231172 7782 231174
rect 7838 231172 7862 231174
rect 7622 231152 7918 231172
rect 7622 230140 7918 230160
rect 7678 230138 7702 230140
rect 7758 230138 7782 230140
rect 7838 230138 7862 230140
rect 7700 230086 7702 230138
rect 7764 230086 7776 230138
rect 7838 230086 7840 230138
rect 7678 230084 7702 230086
rect 7758 230084 7782 230086
rect 7838 230084 7862 230086
rect 7622 230064 7918 230084
rect 7622 229052 7918 229072
rect 7678 229050 7702 229052
rect 7758 229050 7782 229052
rect 7838 229050 7862 229052
rect 7700 228998 7702 229050
rect 7764 228998 7776 229050
rect 7838 228998 7840 229050
rect 7678 228996 7702 228998
rect 7758 228996 7782 228998
rect 7838 228996 7862 228998
rect 7622 228976 7918 228996
rect 7622 227964 7918 227984
rect 7678 227962 7702 227964
rect 7758 227962 7782 227964
rect 7838 227962 7862 227964
rect 7700 227910 7702 227962
rect 7764 227910 7776 227962
rect 7838 227910 7840 227962
rect 7678 227908 7702 227910
rect 7758 227908 7782 227910
rect 7838 227908 7862 227910
rect 7622 227888 7918 227908
rect 7622 226876 7918 226896
rect 7678 226874 7702 226876
rect 7758 226874 7782 226876
rect 7838 226874 7862 226876
rect 7700 226822 7702 226874
rect 7764 226822 7776 226874
rect 7838 226822 7840 226874
rect 7678 226820 7702 226822
rect 7758 226820 7782 226822
rect 7838 226820 7862 226822
rect 7622 226800 7918 226820
rect 7622 225788 7918 225808
rect 7678 225786 7702 225788
rect 7758 225786 7782 225788
rect 7838 225786 7862 225788
rect 7700 225734 7702 225786
rect 7764 225734 7776 225786
rect 7838 225734 7840 225786
rect 7678 225732 7702 225734
rect 7758 225732 7782 225734
rect 7838 225732 7862 225734
rect 7622 225712 7918 225732
rect 8024 224800 8076 224806
rect 8024 224742 8076 224748
rect 7622 224700 7918 224720
rect 7678 224698 7702 224700
rect 7758 224698 7782 224700
rect 7838 224698 7862 224700
rect 7700 224646 7702 224698
rect 7764 224646 7776 224698
rect 7838 224646 7840 224698
rect 7678 224644 7702 224646
rect 7758 224644 7782 224646
rect 7838 224644 7862 224646
rect 7622 224624 7918 224644
rect 7622 223612 7918 223632
rect 7678 223610 7702 223612
rect 7758 223610 7782 223612
rect 7838 223610 7862 223612
rect 7700 223558 7702 223610
rect 7764 223558 7776 223610
rect 7838 223558 7840 223610
rect 7678 223556 7702 223558
rect 7758 223556 7782 223558
rect 7838 223556 7862 223558
rect 7622 223536 7918 223556
rect 7622 222524 7918 222544
rect 7678 222522 7702 222524
rect 7758 222522 7782 222524
rect 7838 222522 7862 222524
rect 7700 222470 7702 222522
rect 7764 222470 7776 222522
rect 7838 222470 7840 222522
rect 7678 222468 7702 222470
rect 7758 222468 7782 222470
rect 7838 222468 7862 222470
rect 7622 222448 7918 222468
rect 7622 221436 7918 221456
rect 7678 221434 7702 221436
rect 7758 221434 7782 221436
rect 7838 221434 7862 221436
rect 7700 221382 7702 221434
rect 7764 221382 7776 221434
rect 7838 221382 7840 221434
rect 7678 221380 7702 221382
rect 7758 221380 7782 221382
rect 7838 221380 7862 221382
rect 7622 221360 7918 221380
rect 7622 220348 7918 220368
rect 7678 220346 7702 220348
rect 7758 220346 7782 220348
rect 7838 220346 7862 220348
rect 7700 220294 7702 220346
rect 7764 220294 7776 220346
rect 7838 220294 7840 220346
rect 7678 220292 7702 220294
rect 7758 220292 7782 220294
rect 7838 220292 7862 220294
rect 7622 220272 7918 220292
rect 7622 219260 7918 219280
rect 7678 219258 7702 219260
rect 7758 219258 7782 219260
rect 7838 219258 7862 219260
rect 7700 219206 7702 219258
rect 7764 219206 7776 219258
rect 7838 219206 7840 219258
rect 7678 219204 7702 219206
rect 7758 219204 7782 219206
rect 7838 219204 7862 219206
rect 7622 219184 7918 219204
rect 7622 218172 7918 218192
rect 7678 218170 7702 218172
rect 7758 218170 7782 218172
rect 7838 218170 7862 218172
rect 7700 218118 7702 218170
rect 7764 218118 7776 218170
rect 7838 218118 7840 218170
rect 7678 218116 7702 218118
rect 7758 218116 7782 218118
rect 7838 218116 7862 218118
rect 7622 218096 7918 218116
rect 7622 217084 7918 217104
rect 7678 217082 7702 217084
rect 7758 217082 7782 217084
rect 7838 217082 7862 217084
rect 7700 217030 7702 217082
rect 7764 217030 7776 217082
rect 7838 217030 7840 217082
rect 7678 217028 7702 217030
rect 7758 217028 7782 217030
rect 7838 217028 7862 217030
rect 7622 217008 7918 217028
rect 7622 215996 7918 216016
rect 7678 215994 7702 215996
rect 7758 215994 7782 215996
rect 7838 215994 7862 215996
rect 7700 215942 7702 215994
rect 7764 215942 7776 215994
rect 7838 215942 7840 215994
rect 7678 215940 7702 215942
rect 7758 215940 7782 215942
rect 7838 215940 7862 215942
rect 7622 215920 7918 215940
rect 7622 214908 7918 214928
rect 7678 214906 7702 214908
rect 7758 214906 7782 214908
rect 7838 214906 7862 214908
rect 7700 214854 7702 214906
rect 7764 214854 7776 214906
rect 7838 214854 7840 214906
rect 7678 214852 7702 214854
rect 7758 214852 7782 214854
rect 7838 214852 7862 214854
rect 7622 214832 7918 214852
rect 7288 214260 7340 214266
rect 7288 214202 7340 214208
rect 7622 213820 7918 213840
rect 7678 213818 7702 213820
rect 7758 213818 7782 213820
rect 7838 213818 7862 213820
rect 7700 213766 7702 213818
rect 7764 213766 7776 213818
rect 7838 213766 7840 213818
rect 7678 213764 7702 213766
rect 7758 213764 7782 213766
rect 7838 213764 7862 213766
rect 7622 213744 7918 213764
rect 7622 212732 7918 212752
rect 7678 212730 7702 212732
rect 7758 212730 7782 212732
rect 7838 212730 7862 212732
rect 7700 212678 7702 212730
rect 7764 212678 7776 212730
rect 7838 212678 7840 212730
rect 7678 212676 7702 212678
rect 7758 212676 7782 212678
rect 7838 212676 7862 212678
rect 7622 212656 7918 212676
rect 7622 211644 7918 211664
rect 7678 211642 7702 211644
rect 7758 211642 7782 211644
rect 7838 211642 7862 211644
rect 7700 211590 7702 211642
rect 7764 211590 7776 211642
rect 7838 211590 7840 211642
rect 7678 211588 7702 211590
rect 7758 211588 7782 211590
rect 7838 211588 7862 211590
rect 7622 211568 7918 211588
rect 7012 210996 7064 211002
rect 7012 210938 7064 210944
rect 7622 210556 7918 210576
rect 7678 210554 7702 210556
rect 7758 210554 7782 210556
rect 7838 210554 7862 210556
rect 7700 210502 7702 210554
rect 7764 210502 7776 210554
rect 7838 210502 7840 210554
rect 7678 210500 7702 210502
rect 7758 210500 7782 210502
rect 7838 210500 7862 210502
rect 7622 210480 7918 210500
rect 7622 209468 7918 209488
rect 7678 209466 7702 209468
rect 7758 209466 7782 209468
rect 7838 209466 7862 209468
rect 7700 209414 7702 209466
rect 7764 209414 7776 209466
rect 7838 209414 7840 209466
rect 7678 209412 7702 209414
rect 7758 209412 7782 209414
rect 7838 209412 7862 209414
rect 7622 209392 7918 209412
rect 7622 208380 7918 208400
rect 7678 208378 7702 208380
rect 7758 208378 7782 208380
rect 7838 208378 7862 208380
rect 7700 208326 7702 208378
rect 7764 208326 7776 208378
rect 7838 208326 7840 208378
rect 7678 208324 7702 208326
rect 7758 208324 7782 208326
rect 7838 208324 7862 208326
rect 7622 208304 7918 208324
rect 7622 207292 7918 207312
rect 7678 207290 7702 207292
rect 7758 207290 7782 207292
rect 7838 207290 7862 207292
rect 7700 207238 7702 207290
rect 7764 207238 7776 207290
rect 7838 207238 7840 207290
rect 7678 207236 7702 207238
rect 7758 207236 7782 207238
rect 7838 207236 7862 207238
rect 7622 207216 7918 207236
rect 7622 206204 7918 206224
rect 7678 206202 7702 206204
rect 7758 206202 7782 206204
rect 7838 206202 7862 206204
rect 7700 206150 7702 206202
rect 7764 206150 7776 206202
rect 7838 206150 7840 206202
rect 7678 206148 7702 206150
rect 7758 206148 7782 206150
rect 7838 206148 7862 206150
rect 7622 206128 7918 206148
rect 7622 205116 7918 205136
rect 7678 205114 7702 205116
rect 7758 205114 7782 205116
rect 7838 205114 7862 205116
rect 7700 205062 7702 205114
rect 7764 205062 7776 205114
rect 7838 205062 7840 205114
rect 7678 205060 7702 205062
rect 7758 205060 7782 205062
rect 7838 205060 7862 205062
rect 7622 205040 7918 205060
rect 7622 204028 7918 204048
rect 7678 204026 7702 204028
rect 7758 204026 7782 204028
rect 7838 204026 7862 204028
rect 7700 203974 7702 204026
rect 7764 203974 7776 204026
rect 7838 203974 7840 204026
rect 7678 203972 7702 203974
rect 7758 203972 7782 203974
rect 7838 203972 7862 203974
rect 7622 203952 7918 203972
rect 7622 202940 7918 202960
rect 7678 202938 7702 202940
rect 7758 202938 7782 202940
rect 7838 202938 7862 202940
rect 7700 202886 7702 202938
rect 7764 202886 7776 202938
rect 7838 202886 7840 202938
rect 7678 202884 7702 202886
rect 7758 202884 7782 202886
rect 7838 202884 7862 202886
rect 7622 202864 7918 202884
rect 7622 201852 7918 201872
rect 7678 201850 7702 201852
rect 7758 201850 7782 201852
rect 7838 201850 7862 201852
rect 7700 201798 7702 201850
rect 7764 201798 7776 201850
rect 7838 201798 7840 201850
rect 7678 201796 7702 201798
rect 7758 201796 7782 201798
rect 7838 201796 7862 201798
rect 7622 201776 7918 201796
rect 7622 200764 7918 200784
rect 7678 200762 7702 200764
rect 7758 200762 7782 200764
rect 7838 200762 7862 200764
rect 7700 200710 7702 200762
rect 7764 200710 7776 200762
rect 7838 200710 7840 200762
rect 7678 200708 7702 200710
rect 7758 200708 7782 200710
rect 7838 200708 7862 200710
rect 7622 200688 7918 200708
rect 7622 199676 7918 199696
rect 7678 199674 7702 199676
rect 7758 199674 7782 199676
rect 7838 199674 7862 199676
rect 7700 199622 7702 199674
rect 7764 199622 7776 199674
rect 7838 199622 7840 199674
rect 7678 199620 7702 199622
rect 7758 199620 7782 199622
rect 7838 199620 7862 199622
rect 7622 199600 7918 199620
rect 7622 198588 7918 198608
rect 7678 198586 7702 198588
rect 7758 198586 7782 198588
rect 7838 198586 7862 198588
rect 7700 198534 7702 198586
rect 7764 198534 7776 198586
rect 7838 198534 7840 198586
rect 7678 198532 7702 198534
rect 7758 198532 7782 198534
rect 7838 198532 7862 198534
rect 7622 198512 7918 198532
rect 7622 197500 7918 197520
rect 7678 197498 7702 197500
rect 7758 197498 7782 197500
rect 7838 197498 7862 197500
rect 7700 197446 7702 197498
rect 7764 197446 7776 197498
rect 7838 197446 7840 197498
rect 7678 197444 7702 197446
rect 7758 197444 7782 197446
rect 7838 197444 7862 197446
rect 7622 197424 7918 197444
rect 7622 196412 7918 196432
rect 7678 196410 7702 196412
rect 7758 196410 7782 196412
rect 7838 196410 7862 196412
rect 7700 196358 7702 196410
rect 7764 196358 7776 196410
rect 7838 196358 7840 196410
rect 7678 196356 7702 196358
rect 7758 196356 7782 196358
rect 7838 196356 7862 196358
rect 7622 196336 7918 196356
rect 7622 195324 7918 195344
rect 7678 195322 7702 195324
rect 7758 195322 7782 195324
rect 7838 195322 7862 195324
rect 7700 195270 7702 195322
rect 7764 195270 7776 195322
rect 7838 195270 7840 195322
rect 7678 195268 7702 195270
rect 7758 195268 7782 195270
rect 7838 195268 7862 195270
rect 7622 195248 7918 195268
rect 7622 194236 7918 194256
rect 7678 194234 7702 194236
rect 7758 194234 7782 194236
rect 7838 194234 7862 194236
rect 7700 194182 7702 194234
rect 7764 194182 7776 194234
rect 7838 194182 7840 194234
rect 7678 194180 7702 194182
rect 7758 194180 7782 194182
rect 7838 194180 7862 194182
rect 7622 194160 7918 194180
rect 7622 193148 7918 193168
rect 7678 193146 7702 193148
rect 7758 193146 7782 193148
rect 7838 193146 7862 193148
rect 7700 193094 7702 193146
rect 7764 193094 7776 193146
rect 7838 193094 7840 193146
rect 7678 193092 7702 193094
rect 7758 193092 7782 193094
rect 7838 193092 7862 193094
rect 7622 193072 7918 193092
rect 7622 192060 7918 192080
rect 7678 192058 7702 192060
rect 7758 192058 7782 192060
rect 7838 192058 7862 192060
rect 7700 192006 7702 192058
rect 7764 192006 7776 192058
rect 7838 192006 7840 192058
rect 7678 192004 7702 192006
rect 7758 192004 7782 192006
rect 7838 192004 7862 192006
rect 7622 191984 7918 192004
rect 7622 190972 7918 190992
rect 7678 190970 7702 190972
rect 7758 190970 7782 190972
rect 7838 190970 7862 190972
rect 7700 190918 7702 190970
rect 7764 190918 7776 190970
rect 7838 190918 7840 190970
rect 7678 190916 7702 190918
rect 7758 190916 7782 190918
rect 7838 190916 7862 190918
rect 7622 190896 7918 190916
rect 7622 189884 7918 189904
rect 7678 189882 7702 189884
rect 7758 189882 7782 189884
rect 7838 189882 7862 189884
rect 7700 189830 7702 189882
rect 7764 189830 7776 189882
rect 7838 189830 7840 189882
rect 7678 189828 7702 189830
rect 7758 189828 7782 189830
rect 7838 189828 7862 189830
rect 7622 189808 7918 189828
rect 7622 188796 7918 188816
rect 7678 188794 7702 188796
rect 7758 188794 7782 188796
rect 7838 188794 7862 188796
rect 7700 188742 7702 188794
rect 7764 188742 7776 188794
rect 7838 188742 7840 188794
rect 7678 188740 7702 188742
rect 7758 188740 7782 188742
rect 7838 188740 7862 188742
rect 7622 188720 7918 188740
rect 7622 187708 7918 187728
rect 7678 187706 7702 187708
rect 7758 187706 7782 187708
rect 7838 187706 7862 187708
rect 7700 187654 7702 187706
rect 7764 187654 7776 187706
rect 7838 187654 7840 187706
rect 7678 187652 7702 187654
rect 7758 187652 7782 187654
rect 7838 187652 7862 187654
rect 7622 187632 7918 187652
rect 7622 186620 7918 186640
rect 7678 186618 7702 186620
rect 7758 186618 7782 186620
rect 7838 186618 7862 186620
rect 7700 186566 7702 186618
rect 7764 186566 7776 186618
rect 7838 186566 7840 186618
rect 7678 186564 7702 186566
rect 7758 186564 7782 186566
rect 7838 186564 7862 186566
rect 7622 186544 7918 186564
rect 7622 185532 7918 185552
rect 7678 185530 7702 185532
rect 7758 185530 7782 185532
rect 7838 185530 7862 185532
rect 7700 185478 7702 185530
rect 7764 185478 7776 185530
rect 7838 185478 7840 185530
rect 7678 185476 7702 185478
rect 7758 185476 7782 185478
rect 7838 185476 7862 185478
rect 7622 185456 7918 185476
rect 7622 184444 7918 184464
rect 7678 184442 7702 184444
rect 7758 184442 7782 184444
rect 7838 184442 7862 184444
rect 7700 184390 7702 184442
rect 7764 184390 7776 184442
rect 7838 184390 7840 184442
rect 7678 184388 7702 184390
rect 7758 184388 7782 184390
rect 7838 184388 7862 184390
rect 7622 184368 7918 184388
rect 7622 183356 7918 183376
rect 7678 183354 7702 183356
rect 7758 183354 7782 183356
rect 7838 183354 7862 183356
rect 7700 183302 7702 183354
rect 7764 183302 7776 183354
rect 7838 183302 7840 183354
rect 7678 183300 7702 183302
rect 7758 183300 7782 183302
rect 7838 183300 7862 183302
rect 7622 183280 7918 183300
rect 7622 182268 7918 182288
rect 7678 182266 7702 182268
rect 7758 182266 7782 182268
rect 7838 182266 7862 182268
rect 7700 182214 7702 182266
rect 7764 182214 7776 182266
rect 7838 182214 7840 182266
rect 7678 182212 7702 182214
rect 7758 182212 7782 182214
rect 7838 182212 7862 182214
rect 7622 182192 7918 182212
rect 7622 181180 7918 181200
rect 7678 181178 7702 181180
rect 7758 181178 7782 181180
rect 7838 181178 7862 181180
rect 7700 181126 7702 181178
rect 7764 181126 7776 181178
rect 7838 181126 7840 181178
rect 7678 181124 7702 181126
rect 7758 181124 7782 181126
rect 7838 181124 7862 181126
rect 7622 181104 7918 181124
rect 7622 180092 7918 180112
rect 7678 180090 7702 180092
rect 7758 180090 7782 180092
rect 7838 180090 7862 180092
rect 7700 180038 7702 180090
rect 7764 180038 7776 180090
rect 7838 180038 7840 180090
rect 7678 180036 7702 180038
rect 7758 180036 7782 180038
rect 7838 180036 7862 180038
rect 7622 180016 7918 180036
rect 7622 179004 7918 179024
rect 7678 179002 7702 179004
rect 7758 179002 7782 179004
rect 7838 179002 7862 179004
rect 7700 178950 7702 179002
rect 7764 178950 7776 179002
rect 7838 178950 7840 179002
rect 7678 178948 7702 178950
rect 7758 178948 7782 178950
rect 7838 178948 7862 178950
rect 7622 178928 7918 178948
rect 7622 177916 7918 177936
rect 7678 177914 7702 177916
rect 7758 177914 7782 177916
rect 7838 177914 7862 177916
rect 7700 177862 7702 177914
rect 7764 177862 7776 177914
rect 7838 177862 7840 177914
rect 7678 177860 7702 177862
rect 7758 177860 7782 177862
rect 7838 177860 7862 177862
rect 7622 177840 7918 177860
rect 7622 176828 7918 176848
rect 7678 176826 7702 176828
rect 7758 176826 7782 176828
rect 7838 176826 7862 176828
rect 7700 176774 7702 176826
rect 7764 176774 7776 176826
rect 7838 176774 7840 176826
rect 7678 176772 7702 176774
rect 7758 176772 7782 176774
rect 7838 176772 7862 176774
rect 7622 176752 7918 176772
rect 7622 175740 7918 175760
rect 7678 175738 7702 175740
rect 7758 175738 7782 175740
rect 7838 175738 7862 175740
rect 7700 175686 7702 175738
rect 7764 175686 7776 175738
rect 7838 175686 7840 175738
rect 7678 175684 7702 175686
rect 7758 175684 7782 175686
rect 7838 175684 7862 175686
rect 7622 175664 7918 175684
rect 7622 174652 7918 174672
rect 7678 174650 7702 174652
rect 7758 174650 7782 174652
rect 7838 174650 7862 174652
rect 7700 174598 7702 174650
rect 7764 174598 7776 174650
rect 7838 174598 7840 174650
rect 7678 174596 7702 174598
rect 7758 174596 7782 174598
rect 7838 174596 7862 174598
rect 7622 174576 7918 174596
rect 7622 173564 7918 173584
rect 7678 173562 7702 173564
rect 7758 173562 7782 173564
rect 7838 173562 7862 173564
rect 7700 173510 7702 173562
rect 7764 173510 7776 173562
rect 7838 173510 7840 173562
rect 7678 173508 7702 173510
rect 7758 173508 7782 173510
rect 7838 173508 7862 173510
rect 7622 173488 7918 173508
rect 7622 172476 7918 172496
rect 7678 172474 7702 172476
rect 7758 172474 7782 172476
rect 7838 172474 7862 172476
rect 7700 172422 7702 172474
rect 7764 172422 7776 172474
rect 7838 172422 7840 172474
rect 7678 172420 7702 172422
rect 7758 172420 7782 172422
rect 7838 172420 7862 172422
rect 7622 172400 7918 172420
rect 6828 172236 6880 172242
rect 6828 172178 6880 172184
rect 7472 172236 7524 172242
rect 7472 172178 7524 172184
rect 6734 116784 6790 116793
rect 6734 116719 6790 116728
rect 5956 116444 6252 116464
rect 6012 116442 6036 116444
rect 6092 116442 6116 116444
rect 6172 116442 6196 116444
rect 6034 116390 6036 116442
rect 6098 116390 6110 116442
rect 6172 116390 6174 116442
rect 6012 116388 6036 116390
rect 6092 116388 6116 116390
rect 6172 116388 6196 116390
rect 5956 116368 6252 116388
rect 5956 115356 6252 115376
rect 6012 115354 6036 115356
rect 6092 115354 6116 115356
rect 6172 115354 6196 115356
rect 6034 115302 6036 115354
rect 6098 115302 6110 115354
rect 6172 115302 6174 115354
rect 6012 115300 6036 115302
rect 6092 115300 6116 115302
rect 6172 115300 6196 115302
rect 5956 115280 6252 115300
rect 5956 114268 6252 114288
rect 6012 114266 6036 114268
rect 6092 114266 6116 114268
rect 6172 114266 6196 114268
rect 6034 114214 6036 114266
rect 6098 114214 6110 114266
rect 6172 114214 6174 114266
rect 6012 114212 6036 114214
rect 6092 114212 6116 114214
rect 6172 114212 6196 114214
rect 5956 114192 6252 114212
rect 5956 113180 6252 113200
rect 6012 113178 6036 113180
rect 6092 113178 6116 113180
rect 6172 113178 6196 113180
rect 6034 113126 6036 113178
rect 6098 113126 6110 113178
rect 6172 113126 6174 113178
rect 6012 113124 6036 113126
rect 6092 113124 6116 113126
rect 6172 113124 6196 113126
rect 5956 113104 6252 113124
rect 5956 112092 6252 112112
rect 6012 112090 6036 112092
rect 6092 112090 6116 112092
rect 6172 112090 6196 112092
rect 6034 112038 6036 112090
rect 6098 112038 6110 112090
rect 6172 112038 6174 112090
rect 6012 112036 6036 112038
rect 6092 112036 6116 112038
rect 6172 112036 6196 112038
rect 5956 112016 6252 112036
rect 5956 111004 6252 111024
rect 6012 111002 6036 111004
rect 6092 111002 6116 111004
rect 6172 111002 6196 111004
rect 6034 110950 6036 111002
rect 6098 110950 6110 111002
rect 6172 110950 6174 111002
rect 6012 110948 6036 110950
rect 6092 110948 6116 110950
rect 6172 110948 6196 110950
rect 5956 110928 6252 110948
rect 5956 109916 6252 109936
rect 6012 109914 6036 109916
rect 6092 109914 6116 109916
rect 6172 109914 6196 109916
rect 6034 109862 6036 109914
rect 6098 109862 6110 109914
rect 6172 109862 6174 109914
rect 6012 109860 6036 109862
rect 6092 109860 6116 109862
rect 6172 109860 6196 109862
rect 5956 109840 6252 109860
rect 5956 108828 6252 108848
rect 6012 108826 6036 108828
rect 6092 108826 6116 108828
rect 6172 108826 6196 108828
rect 6034 108774 6036 108826
rect 6098 108774 6110 108826
rect 6172 108774 6174 108826
rect 6012 108772 6036 108774
rect 6092 108772 6116 108774
rect 6172 108772 6196 108774
rect 5956 108752 6252 108772
rect 5956 107740 6252 107760
rect 6012 107738 6036 107740
rect 6092 107738 6116 107740
rect 6172 107738 6196 107740
rect 6034 107686 6036 107738
rect 6098 107686 6110 107738
rect 6172 107686 6174 107738
rect 6012 107684 6036 107686
rect 6092 107684 6116 107686
rect 6172 107684 6196 107686
rect 5956 107664 6252 107684
rect 5956 106652 6252 106672
rect 6012 106650 6036 106652
rect 6092 106650 6116 106652
rect 6172 106650 6196 106652
rect 6034 106598 6036 106650
rect 6098 106598 6110 106650
rect 6172 106598 6174 106650
rect 6012 106596 6036 106598
rect 6092 106596 6116 106598
rect 6172 106596 6196 106598
rect 5956 106576 6252 106596
rect 5956 105564 6252 105584
rect 6012 105562 6036 105564
rect 6092 105562 6116 105564
rect 6172 105562 6196 105564
rect 6034 105510 6036 105562
rect 6098 105510 6110 105562
rect 6172 105510 6174 105562
rect 6012 105508 6036 105510
rect 6092 105508 6116 105510
rect 6172 105508 6196 105510
rect 5956 105488 6252 105508
rect 5956 104476 6252 104496
rect 6012 104474 6036 104476
rect 6092 104474 6116 104476
rect 6172 104474 6196 104476
rect 6034 104422 6036 104474
rect 6098 104422 6110 104474
rect 6172 104422 6174 104474
rect 6012 104420 6036 104422
rect 6092 104420 6116 104422
rect 6172 104420 6196 104422
rect 5956 104400 6252 104420
rect 5956 103388 6252 103408
rect 6012 103386 6036 103388
rect 6092 103386 6116 103388
rect 6172 103386 6196 103388
rect 6034 103334 6036 103386
rect 6098 103334 6110 103386
rect 6172 103334 6174 103386
rect 6012 103332 6036 103334
rect 6092 103332 6116 103334
rect 6172 103332 6196 103334
rect 5956 103312 6252 103332
rect 5956 102300 6252 102320
rect 6012 102298 6036 102300
rect 6092 102298 6116 102300
rect 6172 102298 6196 102300
rect 6034 102246 6036 102298
rect 6098 102246 6110 102298
rect 6172 102246 6174 102298
rect 6012 102244 6036 102246
rect 6092 102244 6116 102246
rect 6172 102244 6196 102246
rect 5956 102224 6252 102244
rect 5956 101212 6252 101232
rect 6012 101210 6036 101212
rect 6092 101210 6116 101212
rect 6172 101210 6196 101212
rect 6034 101158 6036 101210
rect 6098 101158 6110 101210
rect 6172 101158 6174 101210
rect 6012 101156 6036 101158
rect 6092 101156 6116 101158
rect 6172 101156 6196 101158
rect 5956 101136 6252 101156
rect 5956 100124 6252 100144
rect 6012 100122 6036 100124
rect 6092 100122 6116 100124
rect 6172 100122 6196 100124
rect 6034 100070 6036 100122
rect 6098 100070 6110 100122
rect 6172 100070 6174 100122
rect 6012 100068 6036 100070
rect 6092 100068 6116 100070
rect 6172 100068 6196 100070
rect 5956 100048 6252 100068
rect 5956 99036 6252 99056
rect 6012 99034 6036 99036
rect 6092 99034 6116 99036
rect 6172 99034 6196 99036
rect 6034 98982 6036 99034
rect 6098 98982 6110 99034
rect 6172 98982 6174 99034
rect 6012 98980 6036 98982
rect 6092 98980 6116 98982
rect 6172 98980 6196 98982
rect 5956 98960 6252 98980
rect 5956 97948 6252 97968
rect 6012 97946 6036 97948
rect 6092 97946 6116 97948
rect 6172 97946 6196 97948
rect 6034 97894 6036 97946
rect 6098 97894 6110 97946
rect 6172 97894 6174 97946
rect 6012 97892 6036 97894
rect 6092 97892 6116 97894
rect 6172 97892 6196 97894
rect 5956 97872 6252 97892
rect 5956 96860 6252 96880
rect 6012 96858 6036 96860
rect 6092 96858 6116 96860
rect 6172 96858 6196 96860
rect 6034 96806 6036 96858
rect 6098 96806 6110 96858
rect 6172 96806 6174 96858
rect 6012 96804 6036 96806
rect 6092 96804 6116 96806
rect 6172 96804 6196 96806
rect 5956 96784 6252 96804
rect 5956 95772 6252 95792
rect 6012 95770 6036 95772
rect 6092 95770 6116 95772
rect 6172 95770 6196 95772
rect 6034 95718 6036 95770
rect 6098 95718 6110 95770
rect 6172 95718 6174 95770
rect 6012 95716 6036 95718
rect 6092 95716 6116 95718
rect 6172 95716 6196 95718
rect 5956 95696 6252 95716
rect 5956 94684 6252 94704
rect 6012 94682 6036 94684
rect 6092 94682 6116 94684
rect 6172 94682 6196 94684
rect 6034 94630 6036 94682
rect 6098 94630 6110 94682
rect 6172 94630 6174 94682
rect 6012 94628 6036 94630
rect 6092 94628 6116 94630
rect 6172 94628 6196 94630
rect 5956 94608 6252 94628
rect 5956 93596 6252 93616
rect 6012 93594 6036 93596
rect 6092 93594 6116 93596
rect 6172 93594 6196 93596
rect 6034 93542 6036 93594
rect 6098 93542 6110 93594
rect 6172 93542 6174 93594
rect 6012 93540 6036 93542
rect 6092 93540 6116 93542
rect 6172 93540 6196 93542
rect 5956 93520 6252 93540
rect 5956 92508 6252 92528
rect 6012 92506 6036 92508
rect 6092 92506 6116 92508
rect 6172 92506 6196 92508
rect 6034 92454 6036 92506
rect 6098 92454 6110 92506
rect 6172 92454 6174 92506
rect 6012 92452 6036 92454
rect 6092 92452 6116 92454
rect 6172 92452 6196 92454
rect 5956 92432 6252 92452
rect 5956 91420 6252 91440
rect 6012 91418 6036 91420
rect 6092 91418 6116 91420
rect 6172 91418 6196 91420
rect 6034 91366 6036 91418
rect 6098 91366 6110 91418
rect 6172 91366 6174 91418
rect 6012 91364 6036 91366
rect 6092 91364 6116 91366
rect 6172 91364 6196 91366
rect 5956 91344 6252 91364
rect 5956 90332 6252 90352
rect 6012 90330 6036 90332
rect 6092 90330 6116 90332
rect 6172 90330 6196 90332
rect 6034 90278 6036 90330
rect 6098 90278 6110 90330
rect 6172 90278 6174 90330
rect 6012 90276 6036 90278
rect 6092 90276 6116 90278
rect 6172 90276 6196 90278
rect 5956 90256 6252 90276
rect 5956 89244 6252 89264
rect 6012 89242 6036 89244
rect 6092 89242 6116 89244
rect 6172 89242 6196 89244
rect 6034 89190 6036 89242
rect 6098 89190 6110 89242
rect 6172 89190 6174 89242
rect 6012 89188 6036 89190
rect 6092 89188 6116 89190
rect 6172 89188 6196 89190
rect 5956 89168 6252 89188
rect 5956 88156 6252 88176
rect 6012 88154 6036 88156
rect 6092 88154 6116 88156
rect 6172 88154 6196 88156
rect 6034 88102 6036 88154
rect 6098 88102 6110 88154
rect 6172 88102 6174 88154
rect 6012 88100 6036 88102
rect 6092 88100 6116 88102
rect 6172 88100 6196 88102
rect 5956 88080 6252 88100
rect 5956 87068 6252 87088
rect 6012 87066 6036 87068
rect 6092 87066 6116 87068
rect 6172 87066 6196 87068
rect 6034 87014 6036 87066
rect 6098 87014 6110 87066
rect 6172 87014 6174 87066
rect 6012 87012 6036 87014
rect 6092 87012 6116 87014
rect 6172 87012 6196 87014
rect 5956 86992 6252 87012
rect 5956 85980 6252 86000
rect 6012 85978 6036 85980
rect 6092 85978 6116 85980
rect 6172 85978 6196 85980
rect 6034 85926 6036 85978
rect 6098 85926 6110 85978
rect 6172 85926 6174 85978
rect 6012 85924 6036 85926
rect 6092 85924 6116 85926
rect 6172 85924 6196 85926
rect 5956 85904 6252 85924
rect 5956 84892 6252 84912
rect 6012 84890 6036 84892
rect 6092 84890 6116 84892
rect 6172 84890 6196 84892
rect 6034 84838 6036 84890
rect 6098 84838 6110 84890
rect 6172 84838 6174 84890
rect 6012 84836 6036 84838
rect 6092 84836 6116 84838
rect 6172 84836 6196 84838
rect 5956 84816 6252 84836
rect 5956 83804 6252 83824
rect 6012 83802 6036 83804
rect 6092 83802 6116 83804
rect 6172 83802 6196 83804
rect 6034 83750 6036 83802
rect 6098 83750 6110 83802
rect 6172 83750 6174 83802
rect 6012 83748 6036 83750
rect 6092 83748 6116 83750
rect 6172 83748 6196 83750
rect 5956 83728 6252 83748
rect 5956 82716 6252 82736
rect 6012 82714 6036 82716
rect 6092 82714 6116 82716
rect 6172 82714 6196 82716
rect 6034 82662 6036 82714
rect 6098 82662 6110 82714
rect 6172 82662 6174 82714
rect 6012 82660 6036 82662
rect 6092 82660 6116 82662
rect 6172 82660 6196 82662
rect 5956 82640 6252 82660
rect 5956 81628 6252 81648
rect 6012 81626 6036 81628
rect 6092 81626 6116 81628
rect 6172 81626 6196 81628
rect 6034 81574 6036 81626
rect 6098 81574 6110 81626
rect 6172 81574 6174 81626
rect 6012 81572 6036 81574
rect 6092 81572 6116 81574
rect 6172 81572 6196 81574
rect 5956 81552 6252 81572
rect 5956 80540 6252 80560
rect 6012 80538 6036 80540
rect 6092 80538 6116 80540
rect 6172 80538 6196 80540
rect 6034 80486 6036 80538
rect 6098 80486 6110 80538
rect 6172 80486 6174 80538
rect 6012 80484 6036 80486
rect 6092 80484 6116 80486
rect 6172 80484 6196 80486
rect 5956 80464 6252 80484
rect 5956 79452 6252 79472
rect 6012 79450 6036 79452
rect 6092 79450 6116 79452
rect 6172 79450 6196 79452
rect 6034 79398 6036 79450
rect 6098 79398 6110 79450
rect 6172 79398 6174 79450
rect 6012 79396 6036 79398
rect 6092 79396 6116 79398
rect 6172 79396 6196 79398
rect 5956 79376 6252 79396
rect 5956 78364 6252 78384
rect 6012 78362 6036 78364
rect 6092 78362 6116 78364
rect 6172 78362 6196 78364
rect 6034 78310 6036 78362
rect 6098 78310 6110 78362
rect 6172 78310 6174 78362
rect 6012 78308 6036 78310
rect 6092 78308 6116 78310
rect 6172 78308 6196 78310
rect 5956 78288 6252 78308
rect 5956 77276 6252 77296
rect 6012 77274 6036 77276
rect 6092 77274 6116 77276
rect 6172 77274 6196 77276
rect 6034 77222 6036 77274
rect 6098 77222 6110 77274
rect 6172 77222 6174 77274
rect 6012 77220 6036 77222
rect 6092 77220 6116 77222
rect 6172 77220 6196 77222
rect 5956 77200 6252 77220
rect 5956 76188 6252 76208
rect 6012 76186 6036 76188
rect 6092 76186 6116 76188
rect 6172 76186 6196 76188
rect 6034 76134 6036 76186
rect 6098 76134 6110 76186
rect 6172 76134 6174 76186
rect 6012 76132 6036 76134
rect 6092 76132 6116 76134
rect 6172 76132 6196 76134
rect 5956 76112 6252 76132
rect 5956 75100 6252 75120
rect 6012 75098 6036 75100
rect 6092 75098 6116 75100
rect 6172 75098 6196 75100
rect 6034 75046 6036 75098
rect 6098 75046 6110 75098
rect 6172 75046 6174 75098
rect 6012 75044 6036 75046
rect 6092 75044 6116 75046
rect 6172 75044 6196 75046
rect 5956 75024 6252 75044
rect 5956 74012 6252 74032
rect 6012 74010 6036 74012
rect 6092 74010 6116 74012
rect 6172 74010 6196 74012
rect 6034 73958 6036 74010
rect 6098 73958 6110 74010
rect 6172 73958 6174 74010
rect 6012 73956 6036 73958
rect 6092 73956 6116 73958
rect 6172 73956 6196 73958
rect 5956 73936 6252 73956
rect 5956 72924 6252 72944
rect 6012 72922 6036 72924
rect 6092 72922 6116 72924
rect 6172 72922 6196 72924
rect 6034 72870 6036 72922
rect 6098 72870 6110 72922
rect 6172 72870 6174 72922
rect 6012 72868 6036 72870
rect 6092 72868 6116 72870
rect 6172 72868 6196 72870
rect 5956 72848 6252 72868
rect 5632 72072 5684 72078
rect 5632 72014 5684 72020
rect 5644 71942 5672 72014
rect 5632 71936 5684 71942
rect 5632 71878 5684 71884
rect 6736 71936 6788 71942
rect 6736 71878 6788 71884
rect 5956 71836 6252 71856
rect 6012 71834 6036 71836
rect 6092 71834 6116 71836
rect 6172 71834 6196 71836
rect 6034 71782 6036 71834
rect 6098 71782 6110 71834
rect 6172 71782 6174 71834
rect 6012 71780 6036 71782
rect 6092 71780 6116 71782
rect 6172 71780 6196 71782
rect 5956 71760 6252 71780
rect 5956 70748 6252 70768
rect 6012 70746 6036 70748
rect 6092 70746 6116 70748
rect 6172 70746 6196 70748
rect 6034 70694 6036 70746
rect 6098 70694 6110 70746
rect 6172 70694 6174 70746
rect 6012 70692 6036 70694
rect 6092 70692 6116 70694
rect 6172 70692 6196 70694
rect 5956 70672 6252 70692
rect 5956 69660 6252 69680
rect 6012 69658 6036 69660
rect 6092 69658 6116 69660
rect 6172 69658 6196 69660
rect 6034 69606 6036 69658
rect 6098 69606 6110 69658
rect 6172 69606 6174 69658
rect 6012 69604 6036 69606
rect 6092 69604 6116 69606
rect 6172 69604 6196 69606
rect 5956 69584 6252 69604
rect 5956 68572 6252 68592
rect 6012 68570 6036 68572
rect 6092 68570 6116 68572
rect 6172 68570 6196 68572
rect 6034 68518 6036 68570
rect 6098 68518 6110 68570
rect 6172 68518 6174 68570
rect 6012 68516 6036 68518
rect 6092 68516 6116 68518
rect 6172 68516 6196 68518
rect 5956 68496 6252 68516
rect 5956 67484 6252 67504
rect 6012 67482 6036 67484
rect 6092 67482 6116 67484
rect 6172 67482 6196 67484
rect 6034 67430 6036 67482
rect 6098 67430 6110 67482
rect 6172 67430 6174 67482
rect 6012 67428 6036 67430
rect 6092 67428 6116 67430
rect 6172 67428 6196 67430
rect 5956 67408 6252 67428
rect 5956 66396 6252 66416
rect 6012 66394 6036 66396
rect 6092 66394 6116 66396
rect 6172 66394 6196 66396
rect 6034 66342 6036 66394
rect 6098 66342 6110 66394
rect 6172 66342 6174 66394
rect 6012 66340 6036 66342
rect 6092 66340 6116 66342
rect 6172 66340 6196 66342
rect 5956 66320 6252 66340
rect 5956 65308 6252 65328
rect 6012 65306 6036 65308
rect 6092 65306 6116 65308
rect 6172 65306 6196 65308
rect 6034 65254 6036 65306
rect 6098 65254 6110 65306
rect 6172 65254 6174 65306
rect 6012 65252 6036 65254
rect 6092 65252 6116 65254
rect 6172 65252 6196 65254
rect 5956 65232 6252 65252
rect 5956 64220 6252 64240
rect 6012 64218 6036 64220
rect 6092 64218 6116 64220
rect 6172 64218 6196 64220
rect 6034 64166 6036 64218
rect 6098 64166 6110 64218
rect 6172 64166 6174 64218
rect 6012 64164 6036 64166
rect 6092 64164 6116 64166
rect 6172 64164 6196 64166
rect 5956 64144 6252 64164
rect 5956 63132 6252 63152
rect 6012 63130 6036 63132
rect 6092 63130 6116 63132
rect 6172 63130 6196 63132
rect 6034 63078 6036 63130
rect 6098 63078 6110 63130
rect 6172 63078 6174 63130
rect 6012 63076 6036 63078
rect 6092 63076 6116 63078
rect 6172 63076 6196 63078
rect 5956 63056 6252 63076
rect 5956 62044 6252 62064
rect 6012 62042 6036 62044
rect 6092 62042 6116 62044
rect 6172 62042 6196 62044
rect 6034 61990 6036 62042
rect 6098 61990 6110 62042
rect 6172 61990 6174 62042
rect 6012 61988 6036 61990
rect 6092 61988 6116 61990
rect 6172 61988 6196 61990
rect 5956 61968 6252 61988
rect 5956 60956 6252 60976
rect 6012 60954 6036 60956
rect 6092 60954 6116 60956
rect 6172 60954 6196 60956
rect 6034 60902 6036 60954
rect 6098 60902 6110 60954
rect 6172 60902 6174 60954
rect 6012 60900 6036 60902
rect 6092 60900 6116 60902
rect 6172 60900 6196 60902
rect 5956 60880 6252 60900
rect 5956 59868 6252 59888
rect 6012 59866 6036 59868
rect 6092 59866 6116 59868
rect 6172 59866 6196 59868
rect 6034 59814 6036 59866
rect 6098 59814 6110 59866
rect 6172 59814 6174 59866
rect 6012 59812 6036 59814
rect 6092 59812 6116 59814
rect 6172 59812 6196 59814
rect 5956 59792 6252 59812
rect 5956 58780 6252 58800
rect 6012 58778 6036 58780
rect 6092 58778 6116 58780
rect 6172 58778 6196 58780
rect 6034 58726 6036 58778
rect 6098 58726 6110 58778
rect 6172 58726 6174 58778
rect 6012 58724 6036 58726
rect 6092 58724 6116 58726
rect 6172 58724 6196 58726
rect 5956 58704 6252 58724
rect 5956 57692 6252 57712
rect 6012 57690 6036 57692
rect 6092 57690 6116 57692
rect 6172 57690 6196 57692
rect 6034 57638 6036 57690
rect 6098 57638 6110 57690
rect 6172 57638 6174 57690
rect 6012 57636 6036 57638
rect 6092 57636 6116 57638
rect 6172 57636 6196 57638
rect 5956 57616 6252 57636
rect 5956 56604 6252 56624
rect 6012 56602 6036 56604
rect 6092 56602 6116 56604
rect 6172 56602 6196 56604
rect 6034 56550 6036 56602
rect 6098 56550 6110 56602
rect 6172 56550 6174 56602
rect 6012 56548 6036 56550
rect 6092 56548 6116 56550
rect 6172 56548 6196 56550
rect 5956 56528 6252 56548
rect 5956 55516 6252 55536
rect 6012 55514 6036 55516
rect 6092 55514 6116 55516
rect 6172 55514 6196 55516
rect 6034 55462 6036 55514
rect 6098 55462 6110 55514
rect 6172 55462 6174 55514
rect 6012 55460 6036 55462
rect 6092 55460 6116 55462
rect 6172 55460 6196 55462
rect 5956 55440 6252 55460
rect 5956 54428 6252 54448
rect 6012 54426 6036 54428
rect 6092 54426 6116 54428
rect 6172 54426 6196 54428
rect 6034 54374 6036 54426
rect 6098 54374 6110 54426
rect 6172 54374 6174 54426
rect 6012 54372 6036 54374
rect 6092 54372 6116 54374
rect 6172 54372 6196 54374
rect 5956 54352 6252 54372
rect 5956 53340 6252 53360
rect 6012 53338 6036 53340
rect 6092 53338 6116 53340
rect 6172 53338 6196 53340
rect 6034 53286 6036 53338
rect 6098 53286 6110 53338
rect 6172 53286 6174 53338
rect 6012 53284 6036 53286
rect 6092 53284 6116 53286
rect 6172 53284 6196 53286
rect 5956 53264 6252 53284
rect 5956 52252 6252 52272
rect 6012 52250 6036 52252
rect 6092 52250 6116 52252
rect 6172 52250 6196 52252
rect 6034 52198 6036 52250
rect 6098 52198 6110 52250
rect 6172 52198 6174 52250
rect 6012 52196 6036 52198
rect 6092 52196 6116 52198
rect 6172 52196 6196 52198
rect 5956 52176 6252 52196
rect 5956 51164 6252 51184
rect 6012 51162 6036 51164
rect 6092 51162 6116 51164
rect 6172 51162 6196 51164
rect 6034 51110 6036 51162
rect 6098 51110 6110 51162
rect 6172 51110 6174 51162
rect 6012 51108 6036 51110
rect 6092 51108 6116 51110
rect 6172 51108 6196 51110
rect 5956 51088 6252 51108
rect 6748 50862 6776 71878
rect 6736 50856 6788 50862
rect 6736 50798 6788 50804
rect 6840 50425 6868 172178
rect 7484 171834 7512 172178
rect 7472 171828 7524 171834
rect 7472 171770 7524 171776
rect 7622 171388 7918 171408
rect 7678 171386 7702 171388
rect 7758 171386 7782 171388
rect 7838 171386 7862 171388
rect 7700 171334 7702 171386
rect 7764 171334 7776 171386
rect 7838 171334 7840 171386
rect 7678 171332 7702 171334
rect 7758 171332 7782 171334
rect 7838 171332 7862 171334
rect 7622 171312 7918 171332
rect 7622 170300 7918 170320
rect 7678 170298 7702 170300
rect 7758 170298 7782 170300
rect 7838 170298 7862 170300
rect 7700 170246 7702 170298
rect 7764 170246 7776 170298
rect 7838 170246 7840 170298
rect 7678 170244 7702 170246
rect 7758 170244 7782 170246
rect 7838 170244 7862 170246
rect 7622 170224 7918 170244
rect 7622 169212 7918 169232
rect 7678 169210 7702 169212
rect 7758 169210 7782 169212
rect 7838 169210 7862 169212
rect 7700 169158 7702 169210
rect 7764 169158 7776 169210
rect 7838 169158 7840 169210
rect 7678 169156 7702 169158
rect 7758 169156 7782 169158
rect 7838 169156 7862 169158
rect 7622 169136 7918 169156
rect 7622 168124 7918 168144
rect 7678 168122 7702 168124
rect 7758 168122 7782 168124
rect 7838 168122 7862 168124
rect 7700 168070 7702 168122
rect 7764 168070 7776 168122
rect 7838 168070 7840 168122
rect 7678 168068 7702 168070
rect 7758 168068 7782 168070
rect 7838 168068 7862 168070
rect 7622 168048 7918 168068
rect 7622 167036 7918 167056
rect 7678 167034 7702 167036
rect 7758 167034 7782 167036
rect 7838 167034 7862 167036
rect 7700 166982 7702 167034
rect 7764 166982 7776 167034
rect 7838 166982 7840 167034
rect 7678 166980 7702 166982
rect 7758 166980 7782 166982
rect 7838 166980 7862 166982
rect 7622 166960 7918 166980
rect 7622 165948 7918 165968
rect 7678 165946 7702 165948
rect 7758 165946 7782 165948
rect 7838 165946 7862 165948
rect 7700 165894 7702 165946
rect 7764 165894 7776 165946
rect 7838 165894 7840 165946
rect 7678 165892 7702 165894
rect 7758 165892 7782 165894
rect 7838 165892 7862 165894
rect 7622 165872 7918 165892
rect 7622 164860 7918 164880
rect 7678 164858 7702 164860
rect 7758 164858 7782 164860
rect 7838 164858 7862 164860
rect 7700 164806 7702 164858
rect 7764 164806 7776 164858
rect 7838 164806 7840 164858
rect 7678 164804 7702 164806
rect 7758 164804 7782 164806
rect 7838 164804 7862 164806
rect 7622 164784 7918 164804
rect 7622 163772 7918 163792
rect 7678 163770 7702 163772
rect 7758 163770 7782 163772
rect 7838 163770 7862 163772
rect 7700 163718 7702 163770
rect 7764 163718 7776 163770
rect 7838 163718 7840 163770
rect 7678 163716 7702 163718
rect 7758 163716 7782 163718
rect 7838 163716 7862 163718
rect 7622 163696 7918 163716
rect 7622 162684 7918 162704
rect 7678 162682 7702 162684
rect 7758 162682 7782 162684
rect 7838 162682 7862 162684
rect 7700 162630 7702 162682
rect 7764 162630 7776 162682
rect 7838 162630 7840 162682
rect 7678 162628 7702 162630
rect 7758 162628 7782 162630
rect 7838 162628 7862 162630
rect 7622 162608 7918 162628
rect 7622 161596 7918 161616
rect 7678 161594 7702 161596
rect 7758 161594 7782 161596
rect 7838 161594 7862 161596
rect 7700 161542 7702 161594
rect 7764 161542 7776 161594
rect 7838 161542 7840 161594
rect 7678 161540 7702 161542
rect 7758 161540 7782 161542
rect 7838 161540 7862 161542
rect 7622 161520 7918 161540
rect 7622 160508 7918 160528
rect 7678 160506 7702 160508
rect 7758 160506 7782 160508
rect 7838 160506 7862 160508
rect 7700 160454 7702 160506
rect 7764 160454 7776 160506
rect 7838 160454 7840 160506
rect 7678 160452 7702 160454
rect 7758 160452 7782 160454
rect 7838 160452 7862 160454
rect 7622 160432 7918 160452
rect 7622 159420 7918 159440
rect 7678 159418 7702 159420
rect 7758 159418 7782 159420
rect 7838 159418 7862 159420
rect 7700 159366 7702 159418
rect 7764 159366 7776 159418
rect 7838 159366 7840 159418
rect 7678 159364 7702 159366
rect 7758 159364 7782 159366
rect 7838 159364 7862 159366
rect 7622 159344 7918 159364
rect 7622 158332 7918 158352
rect 7678 158330 7702 158332
rect 7758 158330 7782 158332
rect 7838 158330 7862 158332
rect 7700 158278 7702 158330
rect 7764 158278 7776 158330
rect 7838 158278 7840 158330
rect 7678 158276 7702 158278
rect 7758 158276 7782 158278
rect 7838 158276 7862 158278
rect 7622 158256 7918 158276
rect 8036 158166 8064 224742
rect 6920 158160 6972 158166
rect 6920 158102 6972 158108
rect 8024 158160 8076 158166
rect 8024 158102 8076 158108
rect 6826 50416 6882 50425
rect 6826 50351 6882 50360
rect 5956 50076 6252 50096
rect 6012 50074 6036 50076
rect 6092 50074 6116 50076
rect 6172 50074 6196 50076
rect 6034 50022 6036 50074
rect 6098 50022 6110 50074
rect 6172 50022 6174 50074
rect 6012 50020 6036 50022
rect 6092 50020 6116 50022
rect 6172 50020 6196 50022
rect 5956 50000 6252 50020
rect 5956 48988 6252 49008
rect 6012 48986 6036 48988
rect 6092 48986 6116 48988
rect 6172 48986 6196 48988
rect 6034 48934 6036 48986
rect 6098 48934 6110 48986
rect 6172 48934 6174 48986
rect 6012 48932 6036 48934
rect 6092 48932 6116 48934
rect 6172 48932 6196 48934
rect 5956 48912 6252 48932
rect 5956 47900 6252 47920
rect 6012 47898 6036 47900
rect 6092 47898 6116 47900
rect 6172 47898 6196 47900
rect 6034 47846 6036 47898
rect 6098 47846 6110 47898
rect 6172 47846 6174 47898
rect 6012 47844 6036 47846
rect 6092 47844 6116 47846
rect 6172 47844 6196 47846
rect 5956 47824 6252 47844
rect 5956 46812 6252 46832
rect 6012 46810 6036 46812
rect 6092 46810 6116 46812
rect 6172 46810 6196 46812
rect 6034 46758 6036 46810
rect 6098 46758 6110 46810
rect 6172 46758 6174 46810
rect 6012 46756 6036 46758
rect 6092 46756 6116 46758
rect 6172 46756 6196 46758
rect 5956 46736 6252 46756
rect 5956 45724 6252 45744
rect 6012 45722 6036 45724
rect 6092 45722 6116 45724
rect 6172 45722 6196 45724
rect 6034 45670 6036 45722
rect 6098 45670 6110 45722
rect 6172 45670 6174 45722
rect 6012 45668 6036 45670
rect 6092 45668 6116 45670
rect 6172 45668 6196 45670
rect 5956 45648 6252 45668
rect 5956 44636 6252 44656
rect 6012 44634 6036 44636
rect 6092 44634 6116 44636
rect 6172 44634 6196 44636
rect 6034 44582 6036 44634
rect 6098 44582 6110 44634
rect 6172 44582 6174 44634
rect 6012 44580 6036 44582
rect 6092 44580 6116 44582
rect 6172 44580 6196 44582
rect 5956 44560 6252 44580
rect 5956 43548 6252 43568
rect 6012 43546 6036 43548
rect 6092 43546 6116 43548
rect 6172 43546 6196 43548
rect 6034 43494 6036 43546
rect 6098 43494 6110 43546
rect 6172 43494 6174 43546
rect 6012 43492 6036 43494
rect 6092 43492 6116 43494
rect 6172 43492 6196 43494
rect 5956 43472 6252 43492
rect 5956 42460 6252 42480
rect 6012 42458 6036 42460
rect 6092 42458 6116 42460
rect 6172 42458 6196 42460
rect 6034 42406 6036 42458
rect 6098 42406 6110 42458
rect 6172 42406 6174 42458
rect 6012 42404 6036 42406
rect 6092 42404 6116 42406
rect 6172 42404 6196 42406
rect 5956 42384 6252 42404
rect 5956 41372 6252 41392
rect 6012 41370 6036 41372
rect 6092 41370 6116 41372
rect 6172 41370 6196 41372
rect 6034 41318 6036 41370
rect 6098 41318 6110 41370
rect 6172 41318 6174 41370
rect 6012 41316 6036 41318
rect 6092 41316 6116 41318
rect 6172 41316 6196 41318
rect 5956 41296 6252 41316
rect 5956 40284 6252 40304
rect 6012 40282 6036 40284
rect 6092 40282 6116 40284
rect 6172 40282 6196 40284
rect 6034 40230 6036 40282
rect 6098 40230 6110 40282
rect 6172 40230 6174 40282
rect 6012 40228 6036 40230
rect 6092 40228 6116 40230
rect 6172 40228 6196 40230
rect 5956 40208 6252 40228
rect 5956 39196 6252 39216
rect 6012 39194 6036 39196
rect 6092 39194 6116 39196
rect 6172 39194 6196 39196
rect 6034 39142 6036 39194
rect 6098 39142 6110 39194
rect 6172 39142 6174 39194
rect 6012 39140 6036 39142
rect 6092 39140 6116 39142
rect 6172 39140 6196 39142
rect 5956 39120 6252 39140
rect 5956 38108 6252 38128
rect 6012 38106 6036 38108
rect 6092 38106 6116 38108
rect 6172 38106 6196 38108
rect 6034 38054 6036 38106
rect 6098 38054 6110 38106
rect 6172 38054 6174 38106
rect 6012 38052 6036 38054
rect 6092 38052 6116 38054
rect 6172 38052 6196 38054
rect 5956 38032 6252 38052
rect 5956 37020 6252 37040
rect 6012 37018 6036 37020
rect 6092 37018 6116 37020
rect 6172 37018 6196 37020
rect 6034 36966 6036 37018
rect 6098 36966 6110 37018
rect 6172 36966 6174 37018
rect 6012 36964 6036 36966
rect 6092 36964 6116 36966
rect 6172 36964 6196 36966
rect 5956 36944 6252 36964
rect 5956 35932 6252 35952
rect 6012 35930 6036 35932
rect 6092 35930 6116 35932
rect 6172 35930 6196 35932
rect 6034 35878 6036 35930
rect 6098 35878 6110 35930
rect 6172 35878 6174 35930
rect 6012 35876 6036 35878
rect 6092 35876 6116 35878
rect 6172 35876 6196 35878
rect 5956 35856 6252 35876
rect 5956 34844 6252 34864
rect 6012 34842 6036 34844
rect 6092 34842 6116 34844
rect 6172 34842 6196 34844
rect 6034 34790 6036 34842
rect 6098 34790 6110 34842
rect 6172 34790 6174 34842
rect 6012 34788 6036 34790
rect 6092 34788 6116 34790
rect 6172 34788 6196 34790
rect 5956 34768 6252 34788
rect 5956 33756 6252 33776
rect 6012 33754 6036 33756
rect 6092 33754 6116 33756
rect 6172 33754 6196 33756
rect 6034 33702 6036 33754
rect 6098 33702 6110 33754
rect 6172 33702 6174 33754
rect 6012 33700 6036 33702
rect 6092 33700 6116 33702
rect 6172 33700 6196 33702
rect 5956 33680 6252 33700
rect 5956 32668 6252 32688
rect 6012 32666 6036 32668
rect 6092 32666 6116 32668
rect 6172 32666 6196 32668
rect 6034 32614 6036 32666
rect 6098 32614 6110 32666
rect 6172 32614 6174 32666
rect 6012 32612 6036 32614
rect 6092 32612 6116 32614
rect 6172 32612 6196 32614
rect 5956 32592 6252 32612
rect 5956 31580 6252 31600
rect 6012 31578 6036 31580
rect 6092 31578 6116 31580
rect 6172 31578 6196 31580
rect 6034 31526 6036 31578
rect 6098 31526 6110 31578
rect 6172 31526 6174 31578
rect 6012 31524 6036 31526
rect 6092 31524 6116 31526
rect 6172 31524 6196 31526
rect 5956 31504 6252 31524
rect 5956 30492 6252 30512
rect 6012 30490 6036 30492
rect 6092 30490 6116 30492
rect 6172 30490 6196 30492
rect 6034 30438 6036 30490
rect 6098 30438 6110 30490
rect 6172 30438 6174 30490
rect 6012 30436 6036 30438
rect 6092 30436 6116 30438
rect 6172 30436 6196 30438
rect 5956 30416 6252 30436
rect 5956 29404 6252 29424
rect 6012 29402 6036 29404
rect 6092 29402 6116 29404
rect 6172 29402 6196 29404
rect 6034 29350 6036 29402
rect 6098 29350 6110 29402
rect 6172 29350 6174 29402
rect 6012 29348 6036 29350
rect 6092 29348 6116 29350
rect 6172 29348 6196 29350
rect 5956 29328 6252 29348
rect 5956 28316 6252 28336
rect 6012 28314 6036 28316
rect 6092 28314 6116 28316
rect 6172 28314 6196 28316
rect 6034 28262 6036 28314
rect 6098 28262 6110 28314
rect 6172 28262 6174 28314
rect 6012 28260 6036 28262
rect 6092 28260 6116 28262
rect 6172 28260 6196 28262
rect 5956 28240 6252 28260
rect 5956 27228 6252 27248
rect 6012 27226 6036 27228
rect 6092 27226 6116 27228
rect 6172 27226 6196 27228
rect 6034 27174 6036 27226
rect 6098 27174 6110 27226
rect 6172 27174 6174 27226
rect 6012 27172 6036 27174
rect 6092 27172 6116 27174
rect 6172 27172 6196 27174
rect 5956 27152 6252 27172
rect 5956 26140 6252 26160
rect 6012 26138 6036 26140
rect 6092 26138 6116 26140
rect 6172 26138 6196 26140
rect 6034 26086 6036 26138
rect 6098 26086 6110 26138
rect 6172 26086 6174 26138
rect 6012 26084 6036 26086
rect 6092 26084 6116 26086
rect 6172 26084 6196 26086
rect 5956 26064 6252 26084
rect 5956 25052 6252 25072
rect 6012 25050 6036 25052
rect 6092 25050 6116 25052
rect 6172 25050 6196 25052
rect 6034 24998 6036 25050
rect 6098 24998 6110 25050
rect 6172 24998 6174 25050
rect 6012 24996 6036 24998
rect 6092 24996 6116 24998
rect 6172 24996 6196 24998
rect 5956 24976 6252 24996
rect 5956 23964 6252 23984
rect 6012 23962 6036 23964
rect 6092 23962 6116 23964
rect 6172 23962 6196 23964
rect 6034 23910 6036 23962
rect 6098 23910 6110 23962
rect 6172 23910 6174 23962
rect 6012 23908 6036 23910
rect 6092 23908 6116 23910
rect 6172 23908 6196 23910
rect 5956 23888 6252 23908
rect 5956 22876 6252 22896
rect 6012 22874 6036 22876
rect 6092 22874 6116 22876
rect 6172 22874 6196 22876
rect 6034 22822 6036 22874
rect 6098 22822 6110 22874
rect 6172 22822 6174 22874
rect 6012 22820 6036 22822
rect 6092 22820 6116 22822
rect 6172 22820 6196 22822
rect 5956 22800 6252 22820
rect 5956 21788 6252 21808
rect 6012 21786 6036 21788
rect 6092 21786 6116 21788
rect 6172 21786 6196 21788
rect 6034 21734 6036 21786
rect 6098 21734 6110 21786
rect 6172 21734 6174 21786
rect 6012 21732 6036 21734
rect 6092 21732 6116 21734
rect 6172 21732 6196 21734
rect 5956 21712 6252 21732
rect 5956 20700 6252 20720
rect 6012 20698 6036 20700
rect 6092 20698 6116 20700
rect 6172 20698 6196 20700
rect 6034 20646 6036 20698
rect 6098 20646 6110 20698
rect 6172 20646 6174 20698
rect 6012 20644 6036 20646
rect 6092 20644 6116 20646
rect 6172 20644 6196 20646
rect 5956 20624 6252 20644
rect 5956 19612 6252 19632
rect 6012 19610 6036 19612
rect 6092 19610 6116 19612
rect 6172 19610 6196 19612
rect 6034 19558 6036 19610
rect 6098 19558 6110 19610
rect 6172 19558 6174 19610
rect 6012 19556 6036 19558
rect 6092 19556 6116 19558
rect 6172 19556 6196 19558
rect 5956 19536 6252 19556
rect 5956 18524 6252 18544
rect 6012 18522 6036 18524
rect 6092 18522 6116 18524
rect 6172 18522 6196 18524
rect 6034 18470 6036 18522
rect 6098 18470 6110 18522
rect 6172 18470 6174 18522
rect 6012 18468 6036 18470
rect 6092 18468 6116 18470
rect 6172 18468 6196 18470
rect 5956 18448 6252 18468
rect 5956 17436 6252 17456
rect 6012 17434 6036 17436
rect 6092 17434 6116 17436
rect 6172 17434 6196 17436
rect 6034 17382 6036 17434
rect 6098 17382 6110 17434
rect 6172 17382 6174 17434
rect 6012 17380 6036 17382
rect 6092 17380 6116 17382
rect 6172 17380 6196 17382
rect 5956 17360 6252 17380
rect 4802 17232 4858 17241
rect 4802 17167 4858 17176
rect 4289 16892 4585 16912
rect 4345 16890 4369 16892
rect 4425 16890 4449 16892
rect 4505 16890 4529 16892
rect 4367 16838 4369 16890
rect 4431 16838 4443 16890
rect 4505 16838 4507 16890
rect 4345 16836 4369 16838
rect 4425 16836 4449 16838
rect 4505 16836 4529 16838
rect 4289 16816 4585 16836
rect 5956 16348 6252 16368
rect 6012 16346 6036 16348
rect 6092 16346 6116 16348
rect 6172 16346 6196 16348
rect 6034 16294 6036 16346
rect 6098 16294 6110 16346
rect 6172 16294 6174 16346
rect 6012 16292 6036 16294
rect 6092 16292 6116 16294
rect 6172 16292 6196 16294
rect 5956 16272 6252 16292
rect 4289 15804 4585 15824
rect 4345 15802 4369 15804
rect 4425 15802 4449 15804
rect 4505 15802 4529 15804
rect 4367 15750 4369 15802
rect 4431 15750 4443 15802
rect 4505 15750 4507 15802
rect 4345 15748 4369 15750
rect 4425 15748 4449 15750
rect 4505 15748 4529 15750
rect 4289 15728 4585 15748
rect 5956 15260 6252 15280
rect 6012 15258 6036 15260
rect 6092 15258 6116 15260
rect 6172 15258 6196 15260
rect 6034 15206 6036 15258
rect 6098 15206 6110 15258
rect 6172 15206 6174 15258
rect 6012 15204 6036 15206
rect 6092 15204 6116 15206
rect 6172 15204 6196 15206
rect 5956 15184 6252 15204
rect 4289 14716 4585 14736
rect 4345 14714 4369 14716
rect 4425 14714 4449 14716
rect 4505 14714 4529 14716
rect 4367 14662 4369 14714
rect 4431 14662 4443 14714
rect 4505 14662 4507 14714
rect 4345 14660 4369 14662
rect 4425 14660 4449 14662
rect 4505 14660 4529 14662
rect 4289 14640 4585 14660
rect 5956 14172 6252 14192
rect 6012 14170 6036 14172
rect 6092 14170 6116 14172
rect 6172 14170 6196 14172
rect 6034 14118 6036 14170
rect 6098 14118 6110 14170
rect 6172 14118 6174 14170
rect 6012 14116 6036 14118
rect 6092 14116 6116 14118
rect 6172 14116 6196 14118
rect 5956 14096 6252 14116
rect 4289 13628 4585 13648
rect 4345 13626 4369 13628
rect 4425 13626 4449 13628
rect 4505 13626 4529 13628
rect 4367 13574 4369 13626
rect 4431 13574 4443 13626
rect 4505 13574 4507 13626
rect 4345 13572 4369 13574
rect 4425 13572 4449 13574
rect 4505 13572 4529 13574
rect 4289 13552 4585 13572
rect 5956 13084 6252 13104
rect 6012 13082 6036 13084
rect 6092 13082 6116 13084
rect 6172 13082 6196 13084
rect 6034 13030 6036 13082
rect 6098 13030 6110 13082
rect 6172 13030 6174 13082
rect 6012 13028 6036 13030
rect 6092 13028 6116 13030
rect 6172 13028 6196 13030
rect 5956 13008 6252 13028
rect 4289 12540 4585 12560
rect 4345 12538 4369 12540
rect 4425 12538 4449 12540
rect 4505 12538 4529 12540
rect 4367 12486 4369 12538
rect 4431 12486 4443 12538
rect 4505 12486 4507 12538
rect 4345 12484 4369 12486
rect 4425 12484 4449 12486
rect 4505 12484 4529 12486
rect 4289 12464 4585 12484
rect 5956 11996 6252 12016
rect 6012 11994 6036 11996
rect 6092 11994 6116 11996
rect 6172 11994 6196 11996
rect 6034 11942 6036 11994
rect 6098 11942 6110 11994
rect 6172 11942 6174 11994
rect 6012 11940 6036 11942
rect 6092 11940 6116 11942
rect 6172 11940 6196 11942
rect 5956 11920 6252 11940
rect 4289 11452 4585 11472
rect 4345 11450 4369 11452
rect 4425 11450 4449 11452
rect 4505 11450 4529 11452
rect 4367 11398 4369 11450
rect 4431 11398 4443 11450
rect 4505 11398 4507 11450
rect 4345 11396 4369 11398
rect 4425 11396 4449 11398
rect 4505 11396 4529 11398
rect 4289 11376 4585 11396
rect 5956 10908 6252 10928
rect 6012 10906 6036 10908
rect 6092 10906 6116 10908
rect 6172 10906 6196 10908
rect 6034 10854 6036 10906
rect 6098 10854 6110 10906
rect 6172 10854 6174 10906
rect 6012 10852 6036 10854
rect 6092 10852 6116 10854
rect 6172 10852 6196 10854
rect 5956 10832 6252 10852
rect 4289 10364 4585 10384
rect 4345 10362 4369 10364
rect 4425 10362 4449 10364
rect 4505 10362 4529 10364
rect 4367 10310 4369 10362
rect 4431 10310 4443 10362
rect 4505 10310 4507 10362
rect 4345 10308 4369 10310
rect 4425 10308 4449 10310
rect 4505 10308 4529 10310
rect 4289 10288 4585 10308
rect 5956 9820 6252 9840
rect 6012 9818 6036 9820
rect 6092 9818 6116 9820
rect 6172 9818 6196 9820
rect 6034 9766 6036 9818
rect 6098 9766 6110 9818
rect 6172 9766 6174 9818
rect 6012 9764 6036 9766
rect 6092 9764 6116 9766
rect 6172 9764 6196 9766
rect 5956 9744 6252 9764
rect 4289 9276 4585 9296
rect 4345 9274 4369 9276
rect 4425 9274 4449 9276
rect 4505 9274 4529 9276
rect 4367 9222 4369 9274
rect 4431 9222 4443 9274
rect 4505 9222 4507 9274
rect 4345 9220 4369 9222
rect 4425 9220 4449 9222
rect 4505 9220 4529 9222
rect 4289 9200 4585 9220
rect 5956 8732 6252 8752
rect 6012 8730 6036 8732
rect 6092 8730 6116 8732
rect 6172 8730 6196 8732
rect 6034 8678 6036 8730
rect 6098 8678 6110 8730
rect 6172 8678 6174 8730
rect 6012 8676 6036 8678
rect 6092 8676 6116 8678
rect 6172 8676 6196 8678
rect 5956 8656 6252 8676
rect 4289 8188 4585 8208
rect 4345 8186 4369 8188
rect 4425 8186 4449 8188
rect 4505 8186 4529 8188
rect 4367 8134 4369 8186
rect 4431 8134 4443 8186
rect 4505 8134 4507 8186
rect 4345 8132 4369 8134
rect 4425 8132 4449 8134
rect 4505 8132 4529 8134
rect 4289 8112 4585 8132
rect 5956 7644 6252 7664
rect 6012 7642 6036 7644
rect 6092 7642 6116 7644
rect 6172 7642 6196 7644
rect 6034 7590 6036 7642
rect 6098 7590 6110 7642
rect 6172 7590 6174 7642
rect 6012 7588 6036 7590
rect 6092 7588 6116 7590
rect 6172 7588 6196 7590
rect 5956 7568 6252 7588
rect 4289 7100 4585 7120
rect 4345 7098 4369 7100
rect 4425 7098 4449 7100
rect 4505 7098 4529 7100
rect 4367 7046 4369 7098
rect 4431 7046 4443 7098
rect 4505 7046 4507 7098
rect 4345 7044 4369 7046
rect 4425 7044 4449 7046
rect 4505 7044 4529 7046
rect 4289 7024 4585 7044
rect 5956 6556 6252 6576
rect 6012 6554 6036 6556
rect 6092 6554 6116 6556
rect 6172 6554 6196 6556
rect 6034 6502 6036 6554
rect 6098 6502 6110 6554
rect 6172 6502 6174 6554
rect 6012 6500 6036 6502
rect 6092 6500 6116 6502
rect 6172 6500 6196 6502
rect 5956 6480 6252 6500
rect 4289 6012 4585 6032
rect 4345 6010 4369 6012
rect 4425 6010 4449 6012
rect 4505 6010 4529 6012
rect 4367 5958 4369 6010
rect 4431 5958 4443 6010
rect 4505 5958 4507 6010
rect 4345 5956 4369 5958
rect 4425 5956 4449 5958
rect 4505 5956 4529 5958
rect 4289 5936 4585 5956
rect 5956 5468 6252 5488
rect 6012 5466 6036 5468
rect 6092 5466 6116 5468
rect 6172 5466 6196 5468
rect 6034 5414 6036 5466
rect 6098 5414 6110 5466
rect 6172 5414 6174 5466
rect 6012 5412 6036 5414
rect 6092 5412 6116 5414
rect 6172 5412 6196 5414
rect 5956 5392 6252 5412
rect 4289 4924 4585 4944
rect 4345 4922 4369 4924
rect 4425 4922 4449 4924
rect 4505 4922 4529 4924
rect 4367 4870 4369 4922
rect 4431 4870 4443 4922
rect 4505 4870 4507 4922
rect 4345 4868 4369 4870
rect 4425 4868 4449 4870
rect 4505 4868 4529 4870
rect 4289 4848 4585 4868
rect 5956 4380 6252 4400
rect 6012 4378 6036 4380
rect 6092 4378 6116 4380
rect 6172 4378 6196 4380
rect 6034 4326 6036 4378
rect 6098 4326 6110 4378
rect 6172 4326 6174 4378
rect 6012 4324 6036 4326
rect 6092 4324 6116 4326
rect 6172 4324 6196 4326
rect 5956 4304 6252 4324
rect 6932 4154 6960 158102
rect 7622 157244 7918 157264
rect 7678 157242 7702 157244
rect 7758 157242 7782 157244
rect 7838 157242 7862 157244
rect 7700 157190 7702 157242
rect 7764 157190 7776 157242
rect 7838 157190 7840 157242
rect 7678 157188 7702 157190
rect 7758 157188 7782 157190
rect 7838 157188 7862 157190
rect 7622 157168 7918 157188
rect 7622 156156 7918 156176
rect 7678 156154 7702 156156
rect 7758 156154 7782 156156
rect 7838 156154 7862 156156
rect 7700 156102 7702 156154
rect 7764 156102 7776 156154
rect 7838 156102 7840 156154
rect 7678 156100 7702 156102
rect 7758 156100 7782 156102
rect 7838 156100 7862 156102
rect 7622 156080 7918 156100
rect 7622 155068 7918 155088
rect 7678 155066 7702 155068
rect 7758 155066 7782 155068
rect 7838 155066 7862 155068
rect 7700 155014 7702 155066
rect 7764 155014 7776 155066
rect 7838 155014 7840 155066
rect 7678 155012 7702 155014
rect 7758 155012 7782 155014
rect 7838 155012 7862 155014
rect 7622 154992 7918 155012
rect 7622 153980 7918 154000
rect 7678 153978 7702 153980
rect 7758 153978 7782 153980
rect 7838 153978 7862 153980
rect 7700 153926 7702 153978
rect 7764 153926 7776 153978
rect 7838 153926 7840 153978
rect 7678 153924 7702 153926
rect 7758 153924 7782 153926
rect 7838 153924 7862 153926
rect 7622 153904 7918 153924
rect 7622 152892 7918 152912
rect 7678 152890 7702 152892
rect 7758 152890 7782 152892
rect 7838 152890 7862 152892
rect 7700 152838 7702 152890
rect 7764 152838 7776 152890
rect 7838 152838 7840 152890
rect 7678 152836 7702 152838
rect 7758 152836 7782 152838
rect 7838 152836 7862 152838
rect 7622 152816 7918 152836
rect 7622 151804 7918 151824
rect 7678 151802 7702 151804
rect 7758 151802 7782 151804
rect 7838 151802 7862 151804
rect 7700 151750 7702 151802
rect 7764 151750 7776 151802
rect 7838 151750 7840 151802
rect 7678 151748 7702 151750
rect 7758 151748 7782 151750
rect 7838 151748 7862 151750
rect 7622 151728 7918 151748
rect 7622 150716 7918 150736
rect 7678 150714 7702 150716
rect 7758 150714 7782 150716
rect 7838 150714 7862 150716
rect 7700 150662 7702 150714
rect 7764 150662 7776 150714
rect 7838 150662 7840 150714
rect 7678 150660 7702 150662
rect 7758 150660 7782 150662
rect 7838 150660 7862 150662
rect 7622 150640 7918 150660
rect 7622 149628 7918 149648
rect 7678 149626 7702 149628
rect 7758 149626 7782 149628
rect 7838 149626 7862 149628
rect 7700 149574 7702 149626
rect 7764 149574 7776 149626
rect 7838 149574 7840 149626
rect 7678 149572 7702 149574
rect 7758 149572 7782 149574
rect 7838 149572 7862 149574
rect 7622 149552 7918 149572
rect 7622 148540 7918 148560
rect 7678 148538 7702 148540
rect 7758 148538 7782 148540
rect 7838 148538 7862 148540
rect 7700 148486 7702 148538
rect 7764 148486 7776 148538
rect 7838 148486 7840 148538
rect 7678 148484 7702 148486
rect 7758 148484 7782 148486
rect 7838 148484 7862 148486
rect 7622 148464 7918 148484
rect 7622 147452 7918 147472
rect 7678 147450 7702 147452
rect 7758 147450 7782 147452
rect 7838 147450 7862 147452
rect 7700 147398 7702 147450
rect 7764 147398 7776 147450
rect 7838 147398 7840 147450
rect 7678 147396 7702 147398
rect 7758 147396 7782 147398
rect 7838 147396 7862 147398
rect 7622 147376 7918 147396
rect 7622 146364 7918 146384
rect 7678 146362 7702 146364
rect 7758 146362 7782 146364
rect 7838 146362 7862 146364
rect 7700 146310 7702 146362
rect 7764 146310 7776 146362
rect 7838 146310 7840 146362
rect 7678 146308 7702 146310
rect 7758 146308 7782 146310
rect 7838 146308 7862 146310
rect 7622 146288 7918 146308
rect 7622 145276 7918 145296
rect 7678 145274 7702 145276
rect 7758 145274 7782 145276
rect 7838 145274 7862 145276
rect 7700 145222 7702 145274
rect 7764 145222 7776 145274
rect 7838 145222 7840 145274
rect 7678 145220 7702 145222
rect 7758 145220 7782 145222
rect 7838 145220 7862 145222
rect 7622 145200 7918 145220
rect 7622 144188 7918 144208
rect 7678 144186 7702 144188
rect 7758 144186 7782 144188
rect 7838 144186 7862 144188
rect 7700 144134 7702 144186
rect 7764 144134 7776 144186
rect 7838 144134 7840 144186
rect 7678 144132 7702 144134
rect 7758 144132 7782 144134
rect 7838 144132 7862 144134
rect 7622 144112 7918 144132
rect 7622 143100 7918 143120
rect 7678 143098 7702 143100
rect 7758 143098 7782 143100
rect 7838 143098 7862 143100
rect 7700 143046 7702 143098
rect 7764 143046 7776 143098
rect 7838 143046 7840 143098
rect 7678 143044 7702 143046
rect 7758 143044 7782 143046
rect 7838 143044 7862 143046
rect 7622 143024 7918 143044
rect 7622 142012 7918 142032
rect 7678 142010 7702 142012
rect 7758 142010 7782 142012
rect 7838 142010 7862 142012
rect 7700 141958 7702 142010
rect 7764 141958 7776 142010
rect 7838 141958 7840 142010
rect 7678 141956 7702 141958
rect 7758 141956 7782 141958
rect 7838 141956 7862 141958
rect 7622 141936 7918 141956
rect 7622 140924 7918 140944
rect 7678 140922 7702 140924
rect 7758 140922 7782 140924
rect 7838 140922 7862 140924
rect 7700 140870 7702 140922
rect 7764 140870 7776 140922
rect 7838 140870 7840 140922
rect 7678 140868 7702 140870
rect 7758 140868 7782 140870
rect 7838 140868 7862 140870
rect 7622 140848 7918 140868
rect 7622 139836 7918 139856
rect 7678 139834 7702 139836
rect 7758 139834 7782 139836
rect 7838 139834 7862 139836
rect 7700 139782 7702 139834
rect 7764 139782 7776 139834
rect 7838 139782 7840 139834
rect 7678 139780 7702 139782
rect 7758 139780 7782 139782
rect 7838 139780 7862 139782
rect 7622 139760 7918 139780
rect 7622 138748 7918 138768
rect 7678 138746 7702 138748
rect 7758 138746 7782 138748
rect 7838 138746 7862 138748
rect 7700 138694 7702 138746
rect 7764 138694 7776 138746
rect 7838 138694 7840 138746
rect 7678 138692 7702 138694
rect 7758 138692 7782 138694
rect 7838 138692 7862 138694
rect 7622 138672 7918 138692
rect 7622 137660 7918 137680
rect 7678 137658 7702 137660
rect 7758 137658 7782 137660
rect 7838 137658 7862 137660
rect 7700 137606 7702 137658
rect 7764 137606 7776 137658
rect 7838 137606 7840 137658
rect 7678 137604 7702 137606
rect 7758 137604 7782 137606
rect 7838 137604 7862 137606
rect 7622 137584 7918 137604
rect 7622 136572 7918 136592
rect 7678 136570 7702 136572
rect 7758 136570 7782 136572
rect 7838 136570 7862 136572
rect 7700 136518 7702 136570
rect 7764 136518 7776 136570
rect 7838 136518 7840 136570
rect 7678 136516 7702 136518
rect 7758 136516 7782 136518
rect 7838 136516 7862 136518
rect 7622 136496 7918 136516
rect 7622 135484 7918 135504
rect 7678 135482 7702 135484
rect 7758 135482 7782 135484
rect 7838 135482 7862 135484
rect 7700 135430 7702 135482
rect 7764 135430 7776 135482
rect 7838 135430 7840 135482
rect 7678 135428 7702 135430
rect 7758 135428 7782 135430
rect 7838 135428 7862 135430
rect 7622 135408 7918 135428
rect 7622 134396 7918 134416
rect 7678 134394 7702 134396
rect 7758 134394 7782 134396
rect 7838 134394 7862 134396
rect 7700 134342 7702 134394
rect 7764 134342 7776 134394
rect 7838 134342 7840 134394
rect 7678 134340 7702 134342
rect 7758 134340 7782 134342
rect 7838 134340 7862 134342
rect 7622 134320 7918 134340
rect 7622 133308 7918 133328
rect 7678 133306 7702 133308
rect 7758 133306 7782 133308
rect 7838 133306 7862 133308
rect 7700 133254 7702 133306
rect 7764 133254 7776 133306
rect 7838 133254 7840 133306
rect 7678 133252 7702 133254
rect 7758 133252 7782 133254
rect 7838 133252 7862 133254
rect 7622 133232 7918 133252
rect 7622 132220 7918 132240
rect 7678 132218 7702 132220
rect 7758 132218 7782 132220
rect 7838 132218 7862 132220
rect 7700 132166 7702 132218
rect 7764 132166 7776 132218
rect 7838 132166 7840 132218
rect 7678 132164 7702 132166
rect 7758 132164 7782 132166
rect 7838 132164 7862 132166
rect 7622 132144 7918 132164
rect 7622 131132 7918 131152
rect 7678 131130 7702 131132
rect 7758 131130 7782 131132
rect 7838 131130 7862 131132
rect 7700 131078 7702 131130
rect 7764 131078 7776 131130
rect 7838 131078 7840 131130
rect 7678 131076 7702 131078
rect 7758 131076 7782 131078
rect 7838 131076 7862 131078
rect 7622 131056 7918 131076
rect 7622 130044 7918 130064
rect 7678 130042 7702 130044
rect 7758 130042 7782 130044
rect 7838 130042 7862 130044
rect 7700 129990 7702 130042
rect 7764 129990 7776 130042
rect 7838 129990 7840 130042
rect 7678 129988 7702 129990
rect 7758 129988 7782 129990
rect 7838 129988 7862 129990
rect 7622 129968 7918 129988
rect 7622 128956 7918 128976
rect 7678 128954 7702 128956
rect 7758 128954 7782 128956
rect 7838 128954 7862 128956
rect 7700 128902 7702 128954
rect 7764 128902 7776 128954
rect 7838 128902 7840 128954
rect 7678 128900 7702 128902
rect 7758 128900 7782 128902
rect 7838 128900 7862 128902
rect 7622 128880 7918 128900
rect 7622 127868 7918 127888
rect 7678 127866 7702 127868
rect 7758 127866 7782 127868
rect 7838 127866 7862 127868
rect 7700 127814 7702 127866
rect 7764 127814 7776 127866
rect 7838 127814 7840 127866
rect 7678 127812 7702 127814
rect 7758 127812 7782 127814
rect 7838 127812 7862 127814
rect 7622 127792 7918 127812
rect 7622 126780 7918 126800
rect 7678 126778 7702 126780
rect 7758 126778 7782 126780
rect 7838 126778 7862 126780
rect 7700 126726 7702 126778
rect 7764 126726 7776 126778
rect 7838 126726 7840 126778
rect 7678 126724 7702 126726
rect 7758 126724 7782 126726
rect 7838 126724 7862 126726
rect 7622 126704 7918 126724
rect 7622 125692 7918 125712
rect 7678 125690 7702 125692
rect 7758 125690 7782 125692
rect 7838 125690 7862 125692
rect 7700 125638 7702 125690
rect 7764 125638 7776 125690
rect 7838 125638 7840 125690
rect 7678 125636 7702 125638
rect 7758 125636 7782 125638
rect 7838 125636 7862 125638
rect 7622 125616 7918 125636
rect 7622 124604 7918 124624
rect 7678 124602 7702 124604
rect 7758 124602 7782 124604
rect 7838 124602 7862 124604
rect 7700 124550 7702 124602
rect 7764 124550 7776 124602
rect 7838 124550 7840 124602
rect 7678 124548 7702 124550
rect 7758 124548 7782 124550
rect 7838 124548 7862 124550
rect 7622 124528 7918 124548
rect 7622 123516 7918 123536
rect 7678 123514 7702 123516
rect 7758 123514 7782 123516
rect 7838 123514 7862 123516
rect 7700 123462 7702 123514
rect 7764 123462 7776 123514
rect 7838 123462 7840 123514
rect 7678 123460 7702 123462
rect 7758 123460 7782 123462
rect 7838 123460 7862 123462
rect 7622 123440 7918 123460
rect 7622 122428 7918 122448
rect 7678 122426 7702 122428
rect 7758 122426 7782 122428
rect 7838 122426 7862 122428
rect 7700 122374 7702 122426
rect 7764 122374 7776 122426
rect 7838 122374 7840 122426
rect 7678 122372 7702 122374
rect 7758 122372 7782 122374
rect 7838 122372 7862 122374
rect 7622 122352 7918 122372
rect 7622 121340 7918 121360
rect 7678 121338 7702 121340
rect 7758 121338 7782 121340
rect 7838 121338 7862 121340
rect 7700 121286 7702 121338
rect 7764 121286 7776 121338
rect 7838 121286 7840 121338
rect 7678 121284 7702 121286
rect 7758 121284 7782 121286
rect 7838 121284 7862 121286
rect 7622 121264 7918 121284
rect 7622 120252 7918 120272
rect 7678 120250 7702 120252
rect 7758 120250 7782 120252
rect 7838 120250 7862 120252
rect 7700 120198 7702 120250
rect 7764 120198 7776 120250
rect 7838 120198 7840 120250
rect 7678 120196 7702 120198
rect 7758 120196 7782 120198
rect 7838 120196 7862 120198
rect 7622 120176 7918 120196
rect 7622 119164 7918 119184
rect 7678 119162 7702 119164
rect 7758 119162 7782 119164
rect 7838 119162 7862 119164
rect 7700 119110 7702 119162
rect 7764 119110 7776 119162
rect 7838 119110 7840 119162
rect 7678 119108 7702 119110
rect 7758 119108 7782 119110
rect 7838 119108 7862 119110
rect 7622 119088 7918 119108
rect 7622 118076 7918 118096
rect 7678 118074 7702 118076
rect 7758 118074 7782 118076
rect 7838 118074 7862 118076
rect 7700 118022 7702 118074
rect 7764 118022 7776 118074
rect 7838 118022 7840 118074
rect 7678 118020 7702 118022
rect 7758 118020 7782 118022
rect 7838 118020 7862 118022
rect 7622 118000 7918 118020
rect 7622 116988 7918 117008
rect 7678 116986 7702 116988
rect 7758 116986 7782 116988
rect 7838 116986 7862 116988
rect 7700 116934 7702 116986
rect 7764 116934 7776 116986
rect 7838 116934 7840 116986
rect 7678 116932 7702 116934
rect 7758 116932 7782 116934
rect 7838 116932 7862 116934
rect 7622 116912 7918 116932
rect 7622 115900 7918 115920
rect 7678 115898 7702 115900
rect 7758 115898 7782 115900
rect 7838 115898 7862 115900
rect 7700 115846 7702 115898
rect 7764 115846 7776 115898
rect 7838 115846 7840 115898
rect 7678 115844 7702 115846
rect 7758 115844 7782 115846
rect 7838 115844 7862 115846
rect 7622 115824 7918 115844
rect 7622 114812 7918 114832
rect 7678 114810 7702 114812
rect 7758 114810 7782 114812
rect 7838 114810 7862 114812
rect 7700 114758 7702 114810
rect 7764 114758 7776 114810
rect 7838 114758 7840 114810
rect 7678 114756 7702 114758
rect 7758 114756 7782 114758
rect 7838 114756 7862 114758
rect 7622 114736 7918 114756
rect 7622 113724 7918 113744
rect 7678 113722 7702 113724
rect 7758 113722 7782 113724
rect 7838 113722 7862 113724
rect 7700 113670 7702 113722
rect 7764 113670 7776 113722
rect 7838 113670 7840 113722
rect 7678 113668 7702 113670
rect 7758 113668 7782 113670
rect 7838 113668 7862 113670
rect 7622 113648 7918 113668
rect 7622 112636 7918 112656
rect 7678 112634 7702 112636
rect 7758 112634 7782 112636
rect 7838 112634 7862 112636
rect 7700 112582 7702 112634
rect 7764 112582 7776 112634
rect 7838 112582 7840 112634
rect 7678 112580 7702 112582
rect 7758 112580 7782 112582
rect 7838 112580 7862 112582
rect 7622 112560 7918 112580
rect 7622 111548 7918 111568
rect 7678 111546 7702 111548
rect 7758 111546 7782 111548
rect 7838 111546 7862 111548
rect 7700 111494 7702 111546
rect 7764 111494 7776 111546
rect 7838 111494 7840 111546
rect 7678 111492 7702 111494
rect 7758 111492 7782 111494
rect 7838 111492 7862 111494
rect 7622 111472 7918 111492
rect 7622 110460 7918 110480
rect 7678 110458 7702 110460
rect 7758 110458 7782 110460
rect 7838 110458 7862 110460
rect 7700 110406 7702 110458
rect 7764 110406 7776 110458
rect 7838 110406 7840 110458
rect 7678 110404 7702 110406
rect 7758 110404 7782 110406
rect 7838 110404 7862 110406
rect 7622 110384 7918 110404
rect 7622 109372 7918 109392
rect 7678 109370 7702 109372
rect 7758 109370 7782 109372
rect 7838 109370 7862 109372
rect 7700 109318 7702 109370
rect 7764 109318 7776 109370
rect 7838 109318 7840 109370
rect 7678 109316 7702 109318
rect 7758 109316 7782 109318
rect 7838 109316 7862 109318
rect 7622 109296 7918 109316
rect 7622 108284 7918 108304
rect 7678 108282 7702 108284
rect 7758 108282 7782 108284
rect 7838 108282 7862 108284
rect 7700 108230 7702 108282
rect 7764 108230 7776 108282
rect 7838 108230 7840 108282
rect 7678 108228 7702 108230
rect 7758 108228 7782 108230
rect 7838 108228 7862 108230
rect 7622 108208 7918 108228
rect 7622 107196 7918 107216
rect 7678 107194 7702 107196
rect 7758 107194 7782 107196
rect 7838 107194 7862 107196
rect 7700 107142 7702 107194
rect 7764 107142 7776 107194
rect 7838 107142 7840 107194
rect 7678 107140 7702 107142
rect 7758 107140 7782 107142
rect 7838 107140 7862 107142
rect 7622 107120 7918 107140
rect 7622 106108 7918 106128
rect 7678 106106 7702 106108
rect 7758 106106 7782 106108
rect 7838 106106 7862 106108
rect 7700 106054 7702 106106
rect 7764 106054 7776 106106
rect 7838 106054 7840 106106
rect 7678 106052 7702 106054
rect 7758 106052 7782 106054
rect 7838 106052 7862 106054
rect 7622 106032 7918 106052
rect 7622 105020 7918 105040
rect 7678 105018 7702 105020
rect 7758 105018 7782 105020
rect 7838 105018 7862 105020
rect 7700 104966 7702 105018
rect 7764 104966 7776 105018
rect 7838 104966 7840 105018
rect 7678 104964 7702 104966
rect 7758 104964 7782 104966
rect 7838 104964 7862 104966
rect 7622 104944 7918 104964
rect 7622 103932 7918 103952
rect 7678 103930 7702 103932
rect 7758 103930 7782 103932
rect 7838 103930 7862 103932
rect 7700 103878 7702 103930
rect 7764 103878 7776 103930
rect 7838 103878 7840 103930
rect 7678 103876 7702 103878
rect 7758 103876 7782 103878
rect 7838 103876 7862 103878
rect 7622 103856 7918 103876
rect 7622 102844 7918 102864
rect 7678 102842 7702 102844
rect 7758 102842 7782 102844
rect 7838 102842 7862 102844
rect 7700 102790 7702 102842
rect 7764 102790 7776 102842
rect 7838 102790 7840 102842
rect 7678 102788 7702 102790
rect 7758 102788 7782 102790
rect 7838 102788 7862 102790
rect 7622 102768 7918 102788
rect 7622 101756 7918 101776
rect 7678 101754 7702 101756
rect 7758 101754 7782 101756
rect 7838 101754 7862 101756
rect 7700 101702 7702 101754
rect 7764 101702 7776 101754
rect 7838 101702 7840 101754
rect 7678 101700 7702 101702
rect 7758 101700 7782 101702
rect 7838 101700 7862 101702
rect 7622 101680 7918 101700
rect 7622 100668 7918 100688
rect 7678 100666 7702 100668
rect 7758 100666 7782 100668
rect 7838 100666 7862 100668
rect 7700 100614 7702 100666
rect 7764 100614 7776 100666
rect 7838 100614 7840 100666
rect 7678 100612 7702 100614
rect 7758 100612 7782 100614
rect 7838 100612 7862 100614
rect 7622 100592 7918 100612
rect 7622 99580 7918 99600
rect 7678 99578 7702 99580
rect 7758 99578 7782 99580
rect 7838 99578 7862 99580
rect 7700 99526 7702 99578
rect 7764 99526 7776 99578
rect 7838 99526 7840 99578
rect 7678 99524 7702 99526
rect 7758 99524 7782 99526
rect 7838 99524 7862 99526
rect 7622 99504 7918 99524
rect 7622 98492 7918 98512
rect 7678 98490 7702 98492
rect 7758 98490 7782 98492
rect 7838 98490 7862 98492
rect 7700 98438 7702 98490
rect 7764 98438 7776 98490
rect 7838 98438 7840 98490
rect 7678 98436 7702 98438
rect 7758 98436 7782 98438
rect 7838 98436 7862 98438
rect 7622 98416 7918 98436
rect 7622 97404 7918 97424
rect 7678 97402 7702 97404
rect 7758 97402 7782 97404
rect 7838 97402 7862 97404
rect 7700 97350 7702 97402
rect 7764 97350 7776 97402
rect 7838 97350 7840 97402
rect 7678 97348 7702 97350
rect 7758 97348 7782 97350
rect 7838 97348 7862 97350
rect 7622 97328 7918 97348
rect 7622 96316 7918 96336
rect 7678 96314 7702 96316
rect 7758 96314 7782 96316
rect 7838 96314 7862 96316
rect 7700 96262 7702 96314
rect 7764 96262 7776 96314
rect 7838 96262 7840 96314
rect 7678 96260 7702 96262
rect 7758 96260 7782 96262
rect 7838 96260 7862 96262
rect 7622 96240 7918 96260
rect 7622 95228 7918 95248
rect 7678 95226 7702 95228
rect 7758 95226 7782 95228
rect 7838 95226 7862 95228
rect 7700 95174 7702 95226
rect 7764 95174 7776 95226
rect 7838 95174 7840 95226
rect 7678 95172 7702 95174
rect 7758 95172 7782 95174
rect 7838 95172 7862 95174
rect 7622 95152 7918 95172
rect 7622 94140 7918 94160
rect 7678 94138 7702 94140
rect 7758 94138 7782 94140
rect 7838 94138 7862 94140
rect 7700 94086 7702 94138
rect 7764 94086 7776 94138
rect 7838 94086 7840 94138
rect 7678 94084 7702 94086
rect 7758 94084 7782 94086
rect 7838 94084 7862 94086
rect 7622 94064 7918 94084
rect 7622 93052 7918 93072
rect 7678 93050 7702 93052
rect 7758 93050 7782 93052
rect 7838 93050 7862 93052
rect 7700 92998 7702 93050
rect 7764 92998 7776 93050
rect 7838 92998 7840 93050
rect 7678 92996 7702 92998
rect 7758 92996 7782 92998
rect 7838 92996 7862 92998
rect 7622 92976 7918 92996
rect 7622 91964 7918 91984
rect 7678 91962 7702 91964
rect 7758 91962 7782 91964
rect 7838 91962 7862 91964
rect 7700 91910 7702 91962
rect 7764 91910 7776 91962
rect 7838 91910 7840 91962
rect 7678 91908 7702 91910
rect 7758 91908 7782 91910
rect 7838 91908 7862 91910
rect 7622 91888 7918 91908
rect 7622 90876 7918 90896
rect 7678 90874 7702 90876
rect 7758 90874 7782 90876
rect 7838 90874 7862 90876
rect 7700 90822 7702 90874
rect 7764 90822 7776 90874
rect 7838 90822 7840 90874
rect 7678 90820 7702 90822
rect 7758 90820 7782 90822
rect 7838 90820 7862 90822
rect 7622 90800 7918 90820
rect 7622 89788 7918 89808
rect 7678 89786 7702 89788
rect 7758 89786 7782 89788
rect 7838 89786 7862 89788
rect 7700 89734 7702 89786
rect 7764 89734 7776 89786
rect 7838 89734 7840 89786
rect 7678 89732 7702 89734
rect 7758 89732 7782 89734
rect 7838 89732 7862 89734
rect 7622 89712 7918 89732
rect 7622 88700 7918 88720
rect 7678 88698 7702 88700
rect 7758 88698 7782 88700
rect 7838 88698 7862 88700
rect 7700 88646 7702 88698
rect 7764 88646 7776 88698
rect 7838 88646 7840 88698
rect 7678 88644 7702 88646
rect 7758 88644 7782 88646
rect 7838 88644 7862 88646
rect 7622 88624 7918 88644
rect 7622 87612 7918 87632
rect 7678 87610 7702 87612
rect 7758 87610 7782 87612
rect 7838 87610 7862 87612
rect 7700 87558 7702 87610
rect 7764 87558 7776 87610
rect 7838 87558 7840 87610
rect 7678 87556 7702 87558
rect 7758 87556 7782 87558
rect 7838 87556 7862 87558
rect 7622 87536 7918 87556
rect 7622 86524 7918 86544
rect 7678 86522 7702 86524
rect 7758 86522 7782 86524
rect 7838 86522 7862 86524
rect 7700 86470 7702 86522
rect 7764 86470 7776 86522
rect 7838 86470 7840 86522
rect 7678 86468 7702 86470
rect 7758 86468 7782 86470
rect 7838 86468 7862 86470
rect 7622 86448 7918 86468
rect 7622 85436 7918 85456
rect 7678 85434 7702 85436
rect 7758 85434 7782 85436
rect 7838 85434 7862 85436
rect 7700 85382 7702 85434
rect 7764 85382 7776 85434
rect 7838 85382 7840 85434
rect 7678 85380 7702 85382
rect 7758 85380 7782 85382
rect 7838 85380 7862 85382
rect 7622 85360 7918 85380
rect 7622 84348 7918 84368
rect 7678 84346 7702 84348
rect 7758 84346 7782 84348
rect 7838 84346 7862 84348
rect 7700 84294 7702 84346
rect 7764 84294 7776 84346
rect 7838 84294 7840 84346
rect 7678 84292 7702 84294
rect 7758 84292 7782 84294
rect 7838 84292 7862 84294
rect 7622 84272 7918 84292
rect 8220 83745 8248 233990
rect 8312 225010 8340 332522
rect 9310 332520 9366 332528
rect 9324 332491 9352 332520
rect 8300 225004 8352 225010
rect 8300 224946 8352 224952
rect 8206 83736 8262 83745
rect 8206 83671 8262 83680
rect 7622 83260 7918 83280
rect 7678 83258 7702 83260
rect 7758 83258 7782 83260
rect 7838 83258 7862 83260
rect 7700 83206 7702 83258
rect 7764 83206 7776 83258
rect 7838 83206 7840 83258
rect 7678 83204 7702 83206
rect 7758 83204 7782 83206
rect 7838 83204 7862 83206
rect 7622 83184 7918 83204
rect 7622 82172 7918 82192
rect 7678 82170 7702 82172
rect 7758 82170 7782 82172
rect 7838 82170 7862 82172
rect 7700 82118 7702 82170
rect 7764 82118 7776 82170
rect 7838 82118 7840 82170
rect 7678 82116 7702 82118
rect 7758 82116 7782 82118
rect 7838 82116 7862 82118
rect 7622 82096 7918 82116
rect 7622 81084 7918 81104
rect 7678 81082 7702 81084
rect 7758 81082 7782 81084
rect 7838 81082 7862 81084
rect 7700 81030 7702 81082
rect 7764 81030 7776 81082
rect 7838 81030 7840 81082
rect 7678 81028 7702 81030
rect 7758 81028 7782 81030
rect 7838 81028 7862 81030
rect 7622 81008 7918 81028
rect 7622 79996 7918 80016
rect 7678 79994 7702 79996
rect 7758 79994 7782 79996
rect 7838 79994 7862 79996
rect 7700 79942 7702 79994
rect 7764 79942 7776 79994
rect 7838 79942 7840 79994
rect 7678 79940 7702 79942
rect 7758 79940 7782 79942
rect 7838 79940 7862 79942
rect 7622 79920 7918 79940
rect 7622 78908 7918 78928
rect 7678 78906 7702 78908
rect 7758 78906 7782 78908
rect 7838 78906 7862 78908
rect 7700 78854 7702 78906
rect 7764 78854 7776 78906
rect 7838 78854 7840 78906
rect 7678 78852 7702 78854
rect 7758 78852 7782 78854
rect 7838 78852 7862 78854
rect 7622 78832 7918 78852
rect 7622 77820 7918 77840
rect 7678 77818 7702 77820
rect 7758 77818 7782 77820
rect 7838 77818 7862 77820
rect 7700 77766 7702 77818
rect 7764 77766 7776 77818
rect 7838 77766 7840 77818
rect 7678 77764 7702 77766
rect 7758 77764 7782 77766
rect 7838 77764 7862 77766
rect 7622 77744 7918 77764
rect 7622 76732 7918 76752
rect 7678 76730 7702 76732
rect 7758 76730 7782 76732
rect 7838 76730 7862 76732
rect 7700 76678 7702 76730
rect 7764 76678 7776 76730
rect 7838 76678 7840 76730
rect 7678 76676 7702 76678
rect 7758 76676 7782 76678
rect 7838 76676 7862 76678
rect 7622 76656 7918 76676
rect 7622 75644 7918 75664
rect 7678 75642 7702 75644
rect 7758 75642 7782 75644
rect 7838 75642 7862 75644
rect 7700 75590 7702 75642
rect 7764 75590 7776 75642
rect 7838 75590 7840 75642
rect 7678 75588 7702 75590
rect 7758 75588 7782 75590
rect 7838 75588 7862 75590
rect 7622 75568 7918 75588
rect 7622 74556 7918 74576
rect 7678 74554 7702 74556
rect 7758 74554 7782 74556
rect 7838 74554 7862 74556
rect 7700 74502 7702 74554
rect 7764 74502 7776 74554
rect 7838 74502 7840 74554
rect 7678 74500 7702 74502
rect 7758 74500 7782 74502
rect 7838 74500 7862 74502
rect 7622 74480 7918 74500
rect 7622 73468 7918 73488
rect 7678 73466 7702 73468
rect 7758 73466 7782 73468
rect 7838 73466 7862 73468
rect 7700 73414 7702 73466
rect 7764 73414 7776 73466
rect 7838 73414 7840 73466
rect 7678 73412 7702 73414
rect 7758 73412 7782 73414
rect 7838 73412 7862 73414
rect 7622 73392 7918 73412
rect 7622 72380 7918 72400
rect 7678 72378 7702 72380
rect 7758 72378 7782 72380
rect 7838 72378 7862 72380
rect 7700 72326 7702 72378
rect 7764 72326 7776 72378
rect 7838 72326 7840 72378
rect 7678 72324 7702 72326
rect 7758 72324 7782 72326
rect 7838 72324 7862 72326
rect 7622 72304 7918 72324
rect 7622 71292 7918 71312
rect 7678 71290 7702 71292
rect 7758 71290 7782 71292
rect 7838 71290 7862 71292
rect 7700 71238 7702 71290
rect 7764 71238 7776 71290
rect 7838 71238 7840 71290
rect 7678 71236 7702 71238
rect 7758 71236 7782 71238
rect 7838 71236 7862 71238
rect 7622 71216 7918 71236
rect 7622 70204 7918 70224
rect 7678 70202 7702 70204
rect 7758 70202 7782 70204
rect 7838 70202 7862 70204
rect 7700 70150 7702 70202
rect 7764 70150 7776 70202
rect 7838 70150 7840 70202
rect 7678 70148 7702 70150
rect 7758 70148 7782 70150
rect 7838 70148 7862 70150
rect 7622 70128 7918 70148
rect 7622 69116 7918 69136
rect 7678 69114 7702 69116
rect 7758 69114 7782 69116
rect 7838 69114 7862 69116
rect 7700 69062 7702 69114
rect 7764 69062 7776 69114
rect 7838 69062 7840 69114
rect 7678 69060 7702 69062
rect 7758 69060 7782 69062
rect 7838 69060 7862 69062
rect 7622 69040 7918 69060
rect 7622 68028 7918 68048
rect 7678 68026 7702 68028
rect 7758 68026 7782 68028
rect 7838 68026 7862 68028
rect 7700 67974 7702 68026
rect 7764 67974 7776 68026
rect 7838 67974 7840 68026
rect 7678 67972 7702 67974
rect 7758 67972 7782 67974
rect 7838 67972 7862 67974
rect 7622 67952 7918 67972
rect 7622 66940 7918 66960
rect 7678 66938 7702 66940
rect 7758 66938 7782 66940
rect 7838 66938 7862 66940
rect 7700 66886 7702 66938
rect 7764 66886 7776 66938
rect 7838 66886 7840 66938
rect 7678 66884 7702 66886
rect 7758 66884 7782 66886
rect 7838 66884 7862 66886
rect 7622 66864 7918 66884
rect 7622 65852 7918 65872
rect 7678 65850 7702 65852
rect 7758 65850 7782 65852
rect 7838 65850 7862 65852
rect 7700 65798 7702 65850
rect 7764 65798 7776 65850
rect 7838 65798 7840 65850
rect 7678 65796 7702 65798
rect 7758 65796 7782 65798
rect 7838 65796 7862 65798
rect 7622 65776 7918 65796
rect 7622 64764 7918 64784
rect 7678 64762 7702 64764
rect 7758 64762 7782 64764
rect 7838 64762 7862 64764
rect 7700 64710 7702 64762
rect 7764 64710 7776 64762
rect 7838 64710 7840 64762
rect 7678 64708 7702 64710
rect 7758 64708 7782 64710
rect 7838 64708 7862 64710
rect 7622 64688 7918 64708
rect 7622 63676 7918 63696
rect 7678 63674 7702 63676
rect 7758 63674 7782 63676
rect 7838 63674 7862 63676
rect 7700 63622 7702 63674
rect 7764 63622 7776 63674
rect 7838 63622 7840 63674
rect 7678 63620 7702 63622
rect 7758 63620 7782 63622
rect 7838 63620 7862 63622
rect 7622 63600 7918 63620
rect 7622 62588 7918 62608
rect 7678 62586 7702 62588
rect 7758 62586 7782 62588
rect 7838 62586 7862 62588
rect 7700 62534 7702 62586
rect 7764 62534 7776 62586
rect 7838 62534 7840 62586
rect 7678 62532 7702 62534
rect 7758 62532 7782 62534
rect 7838 62532 7862 62534
rect 7622 62512 7918 62532
rect 7622 61500 7918 61520
rect 7678 61498 7702 61500
rect 7758 61498 7782 61500
rect 7838 61498 7862 61500
rect 7700 61446 7702 61498
rect 7764 61446 7776 61498
rect 7838 61446 7840 61498
rect 7678 61444 7702 61446
rect 7758 61444 7782 61446
rect 7838 61444 7862 61446
rect 7622 61424 7918 61444
rect 7622 60412 7918 60432
rect 7678 60410 7702 60412
rect 7758 60410 7782 60412
rect 7838 60410 7862 60412
rect 7700 60358 7702 60410
rect 7764 60358 7776 60410
rect 7838 60358 7840 60410
rect 7678 60356 7702 60358
rect 7758 60356 7782 60358
rect 7838 60356 7862 60358
rect 7622 60336 7918 60356
rect 7622 59324 7918 59344
rect 7678 59322 7702 59324
rect 7758 59322 7782 59324
rect 7838 59322 7862 59324
rect 7700 59270 7702 59322
rect 7764 59270 7776 59322
rect 7838 59270 7840 59322
rect 7678 59268 7702 59270
rect 7758 59268 7782 59270
rect 7838 59268 7862 59270
rect 7622 59248 7918 59268
rect 7622 58236 7918 58256
rect 7678 58234 7702 58236
rect 7758 58234 7782 58236
rect 7838 58234 7862 58236
rect 7700 58182 7702 58234
rect 7764 58182 7776 58234
rect 7838 58182 7840 58234
rect 7678 58180 7702 58182
rect 7758 58180 7782 58182
rect 7838 58180 7862 58182
rect 7622 58160 7918 58180
rect 7622 57148 7918 57168
rect 7678 57146 7702 57148
rect 7758 57146 7782 57148
rect 7838 57146 7862 57148
rect 7700 57094 7702 57146
rect 7764 57094 7776 57146
rect 7838 57094 7840 57146
rect 7678 57092 7702 57094
rect 7758 57092 7782 57094
rect 7838 57092 7862 57094
rect 7622 57072 7918 57092
rect 7622 56060 7918 56080
rect 7678 56058 7702 56060
rect 7758 56058 7782 56060
rect 7838 56058 7862 56060
rect 7700 56006 7702 56058
rect 7764 56006 7776 56058
rect 7838 56006 7840 56058
rect 7678 56004 7702 56006
rect 7758 56004 7782 56006
rect 7838 56004 7862 56006
rect 7622 55984 7918 56004
rect 7622 54972 7918 54992
rect 7678 54970 7702 54972
rect 7758 54970 7782 54972
rect 7838 54970 7862 54972
rect 7700 54918 7702 54970
rect 7764 54918 7776 54970
rect 7838 54918 7840 54970
rect 7678 54916 7702 54918
rect 7758 54916 7782 54918
rect 7838 54916 7862 54918
rect 7622 54896 7918 54916
rect 7622 53884 7918 53904
rect 7678 53882 7702 53884
rect 7758 53882 7782 53884
rect 7838 53882 7862 53884
rect 7700 53830 7702 53882
rect 7764 53830 7776 53882
rect 7838 53830 7840 53882
rect 7678 53828 7702 53830
rect 7758 53828 7782 53830
rect 7838 53828 7862 53830
rect 7622 53808 7918 53828
rect 7622 52796 7918 52816
rect 7678 52794 7702 52796
rect 7758 52794 7782 52796
rect 7838 52794 7862 52796
rect 7700 52742 7702 52794
rect 7764 52742 7776 52794
rect 7838 52742 7840 52794
rect 7678 52740 7702 52742
rect 7758 52740 7782 52742
rect 7838 52740 7862 52742
rect 7622 52720 7918 52740
rect 7622 51708 7918 51728
rect 7678 51706 7702 51708
rect 7758 51706 7782 51708
rect 7838 51706 7862 51708
rect 7700 51654 7702 51706
rect 7764 51654 7776 51706
rect 7838 51654 7840 51706
rect 7678 51652 7702 51654
rect 7758 51652 7782 51654
rect 7838 51652 7862 51654
rect 7622 51632 7918 51652
rect 8208 50992 8260 50998
rect 8208 50934 8260 50940
rect 7622 50620 7918 50640
rect 7678 50618 7702 50620
rect 7758 50618 7782 50620
rect 7838 50618 7862 50620
rect 7700 50566 7702 50618
rect 7764 50566 7776 50618
rect 7838 50566 7840 50618
rect 7678 50564 7702 50566
rect 7758 50564 7782 50566
rect 7838 50564 7862 50566
rect 7622 50544 7918 50564
rect 7622 49532 7918 49552
rect 7678 49530 7702 49532
rect 7758 49530 7782 49532
rect 7838 49530 7862 49532
rect 7700 49478 7702 49530
rect 7764 49478 7776 49530
rect 7838 49478 7840 49530
rect 7678 49476 7702 49478
rect 7758 49476 7782 49478
rect 7838 49476 7862 49478
rect 7622 49456 7918 49476
rect 7622 48444 7918 48464
rect 7678 48442 7702 48444
rect 7758 48442 7782 48444
rect 7838 48442 7862 48444
rect 7700 48390 7702 48442
rect 7764 48390 7776 48442
rect 7838 48390 7840 48442
rect 7678 48388 7702 48390
rect 7758 48388 7782 48390
rect 7838 48388 7862 48390
rect 7622 48368 7918 48388
rect 7622 47356 7918 47376
rect 7678 47354 7702 47356
rect 7758 47354 7782 47356
rect 7838 47354 7862 47356
rect 7700 47302 7702 47354
rect 7764 47302 7776 47354
rect 7838 47302 7840 47354
rect 7678 47300 7702 47302
rect 7758 47300 7782 47302
rect 7838 47300 7862 47302
rect 7622 47280 7918 47300
rect 7622 46268 7918 46288
rect 7678 46266 7702 46268
rect 7758 46266 7782 46268
rect 7838 46266 7862 46268
rect 7700 46214 7702 46266
rect 7764 46214 7776 46266
rect 7838 46214 7840 46266
rect 7678 46212 7702 46214
rect 7758 46212 7782 46214
rect 7838 46212 7862 46214
rect 7622 46192 7918 46212
rect 7622 45180 7918 45200
rect 7678 45178 7702 45180
rect 7758 45178 7782 45180
rect 7838 45178 7862 45180
rect 7700 45126 7702 45178
rect 7764 45126 7776 45178
rect 7838 45126 7840 45178
rect 7678 45124 7702 45126
rect 7758 45124 7782 45126
rect 7838 45124 7862 45126
rect 7622 45104 7918 45124
rect 7622 44092 7918 44112
rect 7678 44090 7702 44092
rect 7758 44090 7782 44092
rect 7838 44090 7862 44092
rect 7700 44038 7702 44090
rect 7764 44038 7776 44090
rect 7838 44038 7840 44090
rect 7678 44036 7702 44038
rect 7758 44036 7782 44038
rect 7838 44036 7862 44038
rect 7622 44016 7918 44036
rect 7622 43004 7918 43024
rect 7678 43002 7702 43004
rect 7758 43002 7782 43004
rect 7838 43002 7862 43004
rect 7700 42950 7702 43002
rect 7764 42950 7776 43002
rect 7838 42950 7840 43002
rect 7678 42948 7702 42950
rect 7758 42948 7782 42950
rect 7838 42948 7862 42950
rect 7622 42928 7918 42948
rect 7622 41916 7918 41936
rect 7678 41914 7702 41916
rect 7758 41914 7782 41916
rect 7838 41914 7862 41916
rect 7700 41862 7702 41914
rect 7764 41862 7776 41914
rect 7838 41862 7840 41914
rect 7678 41860 7702 41862
rect 7758 41860 7782 41862
rect 7838 41860 7862 41862
rect 7622 41840 7918 41860
rect 7622 40828 7918 40848
rect 7678 40826 7702 40828
rect 7758 40826 7782 40828
rect 7838 40826 7862 40828
rect 7700 40774 7702 40826
rect 7764 40774 7776 40826
rect 7838 40774 7840 40826
rect 7678 40772 7702 40774
rect 7758 40772 7782 40774
rect 7838 40772 7862 40774
rect 7622 40752 7918 40772
rect 7622 39740 7918 39760
rect 7678 39738 7702 39740
rect 7758 39738 7782 39740
rect 7838 39738 7862 39740
rect 7700 39686 7702 39738
rect 7764 39686 7776 39738
rect 7838 39686 7840 39738
rect 7678 39684 7702 39686
rect 7758 39684 7782 39686
rect 7838 39684 7862 39686
rect 7622 39664 7918 39684
rect 7622 38652 7918 38672
rect 7678 38650 7702 38652
rect 7758 38650 7782 38652
rect 7838 38650 7862 38652
rect 7700 38598 7702 38650
rect 7764 38598 7776 38650
rect 7838 38598 7840 38650
rect 7678 38596 7702 38598
rect 7758 38596 7782 38598
rect 7838 38596 7862 38598
rect 7622 38576 7918 38596
rect 7622 37564 7918 37584
rect 7678 37562 7702 37564
rect 7758 37562 7782 37564
rect 7838 37562 7862 37564
rect 7700 37510 7702 37562
rect 7764 37510 7776 37562
rect 7838 37510 7840 37562
rect 7678 37508 7702 37510
rect 7758 37508 7782 37510
rect 7838 37508 7862 37510
rect 7622 37488 7918 37508
rect 7622 36476 7918 36496
rect 7678 36474 7702 36476
rect 7758 36474 7782 36476
rect 7838 36474 7862 36476
rect 7700 36422 7702 36474
rect 7764 36422 7776 36474
rect 7838 36422 7840 36474
rect 7678 36420 7702 36422
rect 7758 36420 7782 36422
rect 7838 36420 7862 36422
rect 7622 36400 7918 36420
rect 7622 35388 7918 35408
rect 7678 35386 7702 35388
rect 7758 35386 7782 35388
rect 7838 35386 7862 35388
rect 7700 35334 7702 35386
rect 7764 35334 7776 35386
rect 7838 35334 7840 35386
rect 7678 35332 7702 35334
rect 7758 35332 7782 35334
rect 7838 35332 7862 35334
rect 7622 35312 7918 35332
rect 7622 34300 7918 34320
rect 7678 34298 7702 34300
rect 7758 34298 7782 34300
rect 7838 34298 7862 34300
rect 7700 34246 7702 34298
rect 7764 34246 7776 34298
rect 7838 34246 7840 34298
rect 7678 34244 7702 34246
rect 7758 34244 7782 34246
rect 7838 34244 7862 34246
rect 7622 34224 7918 34244
rect 7622 33212 7918 33232
rect 7678 33210 7702 33212
rect 7758 33210 7782 33212
rect 7838 33210 7862 33212
rect 7700 33158 7702 33210
rect 7764 33158 7776 33210
rect 7838 33158 7840 33210
rect 7678 33156 7702 33158
rect 7758 33156 7782 33158
rect 7838 33156 7862 33158
rect 7622 33136 7918 33156
rect 7622 32124 7918 32144
rect 7678 32122 7702 32124
rect 7758 32122 7782 32124
rect 7838 32122 7862 32124
rect 7700 32070 7702 32122
rect 7764 32070 7776 32122
rect 7838 32070 7840 32122
rect 7678 32068 7702 32070
rect 7758 32068 7782 32070
rect 7838 32068 7862 32070
rect 7622 32048 7918 32068
rect 7622 31036 7918 31056
rect 7678 31034 7702 31036
rect 7758 31034 7782 31036
rect 7838 31034 7862 31036
rect 7700 30982 7702 31034
rect 7764 30982 7776 31034
rect 7838 30982 7840 31034
rect 7678 30980 7702 30982
rect 7758 30980 7782 30982
rect 7838 30980 7862 30982
rect 7622 30960 7918 30980
rect 7622 29948 7918 29968
rect 7678 29946 7702 29948
rect 7758 29946 7782 29948
rect 7838 29946 7862 29948
rect 7700 29894 7702 29946
rect 7764 29894 7776 29946
rect 7838 29894 7840 29946
rect 7678 29892 7702 29894
rect 7758 29892 7782 29894
rect 7838 29892 7862 29894
rect 7622 29872 7918 29892
rect 7622 28860 7918 28880
rect 7678 28858 7702 28860
rect 7758 28858 7782 28860
rect 7838 28858 7862 28860
rect 7700 28806 7702 28858
rect 7764 28806 7776 28858
rect 7838 28806 7840 28858
rect 7678 28804 7702 28806
rect 7758 28804 7782 28806
rect 7838 28804 7862 28806
rect 7622 28784 7918 28804
rect 7622 27772 7918 27792
rect 7678 27770 7702 27772
rect 7758 27770 7782 27772
rect 7838 27770 7862 27772
rect 7700 27718 7702 27770
rect 7764 27718 7776 27770
rect 7838 27718 7840 27770
rect 7678 27716 7702 27718
rect 7758 27716 7782 27718
rect 7838 27716 7862 27718
rect 7622 27696 7918 27716
rect 7622 26684 7918 26704
rect 7678 26682 7702 26684
rect 7758 26682 7782 26684
rect 7838 26682 7862 26684
rect 7700 26630 7702 26682
rect 7764 26630 7776 26682
rect 7838 26630 7840 26682
rect 7678 26628 7702 26630
rect 7758 26628 7782 26630
rect 7838 26628 7862 26630
rect 7622 26608 7918 26628
rect 7622 25596 7918 25616
rect 7678 25594 7702 25596
rect 7758 25594 7782 25596
rect 7838 25594 7862 25596
rect 7700 25542 7702 25594
rect 7764 25542 7776 25594
rect 7838 25542 7840 25594
rect 7678 25540 7702 25542
rect 7758 25540 7782 25542
rect 7838 25540 7862 25542
rect 7622 25520 7918 25540
rect 7622 24508 7918 24528
rect 7678 24506 7702 24508
rect 7758 24506 7782 24508
rect 7838 24506 7862 24508
rect 7700 24454 7702 24506
rect 7764 24454 7776 24506
rect 7838 24454 7840 24506
rect 7678 24452 7702 24454
rect 7758 24452 7782 24454
rect 7838 24452 7862 24454
rect 7622 24432 7918 24452
rect 7622 23420 7918 23440
rect 7678 23418 7702 23420
rect 7758 23418 7782 23420
rect 7838 23418 7862 23420
rect 7700 23366 7702 23418
rect 7764 23366 7776 23418
rect 7838 23366 7840 23418
rect 7678 23364 7702 23366
rect 7758 23364 7782 23366
rect 7838 23364 7862 23366
rect 7622 23344 7918 23364
rect 7622 22332 7918 22352
rect 7678 22330 7702 22332
rect 7758 22330 7782 22332
rect 7838 22330 7862 22332
rect 7700 22278 7702 22330
rect 7764 22278 7776 22330
rect 7838 22278 7840 22330
rect 7678 22276 7702 22278
rect 7758 22276 7782 22278
rect 7838 22276 7862 22278
rect 7622 22256 7918 22276
rect 7622 21244 7918 21264
rect 7678 21242 7702 21244
rect 7758 21242 7782 21244
rect 7838 21242 7862 21244
rect 7700 21190 7702 21242
rect 7764 21190 7776 21242
rect 7838 21190 7840 21242
rect 7678 21188 7702 21190
rect 7758 21188 7782 21190
rect 7838 21188 7862 21190
rect 7622 21168 7918 21188
rect 7622 20156 7918 20176
rect 7678 20154 7702 20156
rect 7758 20154 7782 20156
rect 7838 20154 7862 20156
rect 7700 20102 7702 20154
rect 7764 20102 7776 20154
rect 7838 20102 7840 20154
rect 7678 20100 7702 20102
rect 7758 20100 7782 20102
rect 7838 20100 7862 20102
rect 7622 20080 7918 20100
rect 7622 19068 7918 19088
rect 7678 19066 7702 19068
rect 7758 19066 7782 19068
rect 7838 19066 7862 19068
rect 7700 19014 7702 19066
rect 7764 19014 7776 19066
rect 7838 19014 7840 19066
rect 7678 19012 7702 19014
rect 7758 19012 7782 19014
rect 7838 19012 7862 19014
rect 7622 18992 7918 19012
rect 7622 17980 7918 18000
rect 7678 17978 7702 17980
rect 7758 17978 7782 17980
rect 7838 17978 7862 17980
rect 7700 17926 7702 17978
rect 7764 17926 7776 17978
rect 7838 17926 7840 17978
rect 7678 17924 7702 17926
rect 7758 17924 7782 17926
rect 7838 17924 7862 17926
rect 7622 17904 7918 17924
rect 7622 16892 7918 16912
rect 7678 16890 7702 16892
rect 7758 16890 7782 16892
rect 7838 16890 7862 16892
rect 7700 16838 7702 16890
rect 7764 16838 7776 16890
rect 7838 16838 7840 16890
rect 7678 16836 7702 16838
rect 7758 16836 7782 16838
rect 7838 16836 7862 16838
rect 7622 16816 7918 16836
rect 7622 15804 7918 15824
rect 7678 15802 7702 15804
rect 7758 15802 7782 15804
rect 7838 15802 7862 15804
rect 7700 15750 7702 15802
rect 7764 15750 7776 15802
rect 7838 15750 7840 15802
rect 7678 15748 7702 15750
rect 7758 15748 7782 15750
rect 7838 15748 7862 15750
rect 7622 15728 7918 15748
rect 7622 14716 7918 14736
rect 7678 14714 7702 14716
rect 7758 14714 7782 14716
rect 7838 14714 7862 14716
rect 7700 14662 7702 14714
rect 7764 14662 7776 14714
rect 7838 14662 7840 14714
rect 7678 14660 7702 14662
rect 7758 14660 7782 14662
rect 7838 14660 7862 14662
rect 7622 14640 7918 14660
rect 7622 13628 7918 13648
rect 7678 13626 7702 13628
rect 7758 13626 7782 13628
rect 7838 13626 7862 13628
rect 7700 13574 7702 13626
rect 7764 13574 7776 13626
rect 7838 13574 7840 13626
rect 7678 13572 7702 13574
rect 7758 13572 7782 13574
rect 7838 13572 7862 13574
rect 7622 13552 7918 13572
rect 7622 12540 7918 12560
rect 7678 12538 7702 12540
rect 7758 12538 7782 12540
rect 7838 12538 7862 12540
rect 7700 12486 7702 12538
rect 7764 12486 7776 12538
rect 7838 12486 7840 12538
rect 7678 12484 7702 12486
rect 7758 12484 7782 12486
rect 7838 12484 7862 12486
rect 7622 12464 7918 12484
rect 7622 11452 7918 11472
rect 7678 11450 7702 11452
rect 7758 11450 7782 11452
rect 7838 11450 7862 11452
rect 7700 11398 7702 11450
rect 7764 11398 7776 11450
rect 7838 11398 7840 11450
rect 7678 11396 7702 11398
rect 7758 11396 7782 11398
rect 7838 11396 7862 11398
rect 7622 11376 7918 11396
rect 7622 10364 7918 10384
rect 7678 10362 7702 10364
rect 7758 10362 7782 10364
rect 7838 10362 7862 10364
rect 7700 10310 7702 10362
rect 7764 10310 7776 10362
rect 7838 10310 7840 10362
rect 7678 10308 7702 10310
rect 7758 10308 7782 10310
rect 7838 10308 7862 10310
rect 7622 10288 7918 10308
rect 7622 9276 7918 9296
rect 7678 9274 7702 9276
rect 7758 9274 7782 9276
rect 7838 9274 7862 9276
rect 7700 9222 7702 9274
rect 7764 9222 7776 9274
rect 7838 9222 7840 9274
rect 7678 9220 7702 9222
rect 7758 9220 7782 9222
rect 7838 9220 7862 9222
rect 7622 9200 7918 9220
rect 7622 8188 7918 8208
rect 7678 8186 7702 8188
rect 7758 8186 7782 8188
rect 7838 8186 7862 8188
rect 7700 8134 7702 8186
rect 7764 8134 7776 8186
rect 7838 8134 7840 8186
rect 7678 8132 7702 8134
rect 7758 8132 7782 8134
rect 7838 8132 7862 8134
rect 7622 8112 7918 8132
rect 7622 7100 7918 7120
rect 7678 7098 7702 7100
rect 7758 7098 7782 7100
rect 7838 7098 7862 7100
rect 7700 7046 7702 7098
rect 7764 7046 7776 7098
rect 7838 7046 7840 7098
rect 7678 7044 7702 7046
rect 7758 7044 7782 7046
rect 7838 7044 7862 7046
rect 7622 7024 7918 7044
rect 7622 6012 7918 6032
rect 7678 6010 7702 6012
rect 7758 6010 7782 6012
rect 7838 6010 7862 6012
rect 7700 5958 7702 6010
rect 7764 5958 7776 6010
rect 7838 5958 7840 6010
rect 7678 5956 7702 5958
rect 7758 5956 7782 5958
rect 7838 5956 7862 5958
rect 7622 5936 7918 5956
rect 7622 4924 7918 4944
rect 7678 4922 7702 4924
rect 7758 4922 7782 4924
rect 7838 4922 7862 4924
rect 7700 4870 7702 4922
rect 7764 4870 7776 4922
rect 7838 4870 7840 4922
rect 7678 4868 7702 4870
rect 7758 4868 7782 4870
rect 7838 4868 7862 4870
rect 7622 4848 7918 4868
rect 6840 4126 6960 4154
rect 4289 3836 4585 3856
rect 4345 3834 4369 3836
rect 4425 3834 4449 3836
rect 4505 3834 4529 3836
rect 4367 3782 4369 3834
rect 4431 3782 4443 3834
rect 4505 3782 4507 3834
rect 4345 3780 4369 3782
rect 4425 3780 4449 3782
rect 4505 3780 4529 3782
rect 4289 3760 4585 3780
rect 5956 3292 6252 3312
rect 6012 3290 6036 3292
rect 6092 3290 6116 3292
rect 6172 3290 6196 3292
rect 6034 3238 6036 3290
rect 6098 3238 6110 3290
rect 6172 3238 6174 3290
rect 6012 3236 6036 3238
rect 6092 3236 6116 3238
rect 6172 3236 6196 3238
rect 5956 3216 6252 3236
rect 4289 2748 4585 2768
rect 4345 2746 4369 2748
rect 4425 2746 4449 2748
rect 4505 2746 4529 2748
rect 4367 2694 4369 2746
rect 4431 2694 4443 2746
rect 4505 2694 4507 2746
rect 4345 2692 4369 2694
rect 4425 2692 4449 2694
rect 4505 2692 4529 2694
rect 4289 2672 4585 2692
rect 5956 2204 6252 2224
rect 6012 2202 6036 2204
rect 6092 2202 6116 2204
rect 6172 2202 6196 2204
rect 6034 2150 6036 2202
rect 6098 2150 6110 2202
rect 6172 2150 6174 2202
rect 6012 2148 6036 2150
rect 6092 2148 6116 2150
rect 6172 2148 6196 2150
rect 5956 2128 6252 2148
rect 2870 54 3004 82
rect 938 0 994 54
rect 2870 0 2926 54
rect 4894 0 4950 480
rect 6840 82 6868 4126
rect 7622 3836 7918 3856
rect 7678 3834 7702 3836
rect 7758 3834 7782 3836
rect 7838 3834 7862 3836
rect 7700 3782 7702 3834
rect 7764 3782 7776 3834
rect 7838 3782 7840 3834
rect 7678 3780 7702 3782
rect 7758 3780 7782 3782
rect 7838 3780 7862 3782
rect 7622 3760 7918 3780
rect 7622 2748 7918 2768
rect 7678 2746 7702 2748
rect 7758 2746 7782 2748
rect 7838 2746 7862 2748
rect 7700 2694 7702 2746
rect 7764 2694 7776 2746
rect 7838 2694 7840 2746
rect 7678 2692 7702 2694
rect 7758 2692 7782 2694
rect 7838 2692 7862 2694
rect 7622 2672 7918 2692
rect 6918 82 6974 480
rect 8220 134 8248 50934
rect 6840 54 6974 82
rect 8208 128 8260 134
rect 8208 70 8260 76
rect 8942 128 8998 480
rect 8942 76 8944 128
rect 8996 76 8998 128
rect 6918 0 6974 54
rect 8942 0 8998 76
<< via2 >>
rect 2622 330778 2678 330780
rect 2702 330778 2758 330780
rect 2782 330778 2838 330780
rect 2862 330778 2918 330780
rect 2622 330726 2648 330778
rect 2648 330726 2678 330778
rect 2702 330726 2712 330778
rect 2712 330726 2758 330778
rect 2782 330726 2828 330778
rect 2828 330726 2838 330778
rect 2862 330726 2892 330778
rect 2892 330726 2918 330778
rect 2622 330724 2678 330726
rect 2702 330724 2758 330726
rect 2782 330724 2838 330726
rect 2862 330724 2918 330726
rect 2622 329690 2678 329692
rect 2702 329690 2758 329692
rect 2782 329690 2838 329692
rect 2862 329690 2918 329692
rect 2622 329638 2648 329690
rect 2648 329638 2678 329690
rect 2702 329638 2712 329690
rect 2712 329638 2758 329690
rect 2782 329638 2828 329690
rect 2828 329638 2838 329690
rect 2862 329638 2892 329690
rect 2892 329638 2918 329690
rect 2622 329636 2678 329638
rect 2702 329636 2758 329638
rect 2782 329636 2838 329638
rect 2862 329636 2918 329638
rect 2622 328602 2678 328604
rect 2702 328602 2758 328604
rect 2782 328602 2838 328604
rect 2862 328602 2918 328604
rect 2622 328550 2648 328602
rect 2648 328550 2678 328602
rect 2702 328550 2712 328602
rect 2712 328550 2758 328602
rect 2782 328550 2828 328602
rect 2828 328550 2838 328602
rect 2862 328550 2892 328602
rect 2892 328550 2918 328602
rect 2622 328548 2678 328550
rect 2702 328548 2758 328550
rect 2782 328548 2838 328550
rect 2862 328548 2918 328550
rect 2622 327514 2678 327516
rect 2702 327514 2758 327516
rect 2782 327514 2838 327516
rect 2862 327514 2918 327516
rect 2622 327462 2648 327514
rect 2648 327462 2678 327514
rect 2702 327462 2712 327514
rect 2712 327462 2758 327514
rect 2782 327462 2828 327514
rect 2828 327462 2838 327514
rect 2862 327462 2892 327514
rect 2892 327462 2918 327514
rect 2622 327460 2678 327462
rect 2702 327460 2758 327462
rect 2782 327460 2838 327462
rect 2862 327460 2918 327462
rect 2622 326426 2678 326428
rect 2702 326426 2758 326428
rect 2782 326426 2838 326428
rect 2862 326426 2918 326428
rect 2622 326374 2648 326426
rect 2648 326374 2678 326426
rect 2702 326374 2712 326426
rect 2712 326374 2758 326426
rect 2782 326374 2828 326426
rect 2828 326374 2838 326426
rect 2862 326374 2892 326426
rect 2892 326374 2918 326426
rect 2622 326372 2678 326374
rect 2702 326372 2758 326374
rect 2782 326372 2838 326374
rect 2862 326372 2918 326374
rect 2622 325338 2678 325340
rect 2702 325338 2758 325340
rect 2782 325338 2838 325340
rect 2862 325338 2918 325340
rect 2622 325286 2648 325338
rect 2648 325286 2678 325338
rect 2702 325286 2712 325338
rect 2712 325286 2758 325338
rect 2782 325286 2828 325338
rect 2828 325286 2838 325338
rect 2862 325286 2892 325338
rect 2892 325286 2918 325338
rect 2622 325284 2678 325286
rect 2702 325284 2758 325286
rect 2782 325284 2838 325286
rect 2862 325284 2918 325286
rect 2622 324250 2678 324252
rect 2702 324250 2758 324252
rect 2782 324250 2838 324252
rect 2862 324250 2918 324252
rect 2622 324198 2648 324250
rect 2648 324198 2678 324250
rect 2702 324198 2712 324250
rect 2712 324198 2758 324250
rect 2782 324198 2828 324250
rect 2828 324198 2838 324250
rect 2862 324198 2892 324250
rect 2892 324198 2918 324250
rect 2622 324196 2678 324198
rect 2702 324196 2758 324198
rect 2782 324196 2838 324198
rect 2862 324196 2918 324198
rect 2622 323162 2678 323164
rect 2702 323162 2758 323164
rect 2782 323162 2838 323164
rect 2862 323162 2918 323164
rect 2622 323110 2648 323162
rect 2648 323110 2678 323162
rect 2702 323110 2712 323162
rect 2712 323110 2758 323162
rect 2782 323110 2828 323162
rect 2828 323110 2838 323162
rect 2862 323110 2892 323162
rect 2892 323110 2918 323162
rect 2622 323108 2678 323110
rect 2702 323108 2758 323110
rect 2782 323108 2838 323110
rect 2862 323108 2918 323110
rect 2622 322074 2678 322076
rect 2702 322074 2758 322076
rect 2782 322074 2838 322076
rect 2862 322074 2918 322076
rect 2622 322022 2648 322074
rect 2648 322022 2678 322074
rect 2702 322022 2712 322074
rect 2712 322022 2758 322074
rect 2782 322022 2828 322074
rect 2828 322022 2838 322074
rect 2862 322022 2892 322074
rect 2892 322022 2918 322074
rect 2622 322020 2678 322022
rect 2702 322020 2758 322022
rect 2782 322020 2838 322022
rect 2862 322020 2918 322022
rect 2622 320986 2678 320988
rect 2702 320986 2758 320988
rect 2782 320986 2838 320988
rect 2862 320986 2918 320988
rect 2622 320934 2648 320986
rect 2648 320934 2678 320986
rect 2702 320934 2712 320986
rect 2712 320934 2758 320986
rect 2782 320934 2828 320986
rect 2828 320934 2838 320986
rect 2862 320934 2892 320986
rect 2892 320934 2918 320986
rect 2622 320932 2678 320934
rect 2702 320932 2758 320934
rect 2782 320932 2838 320934
rect 2862 320932 2918 320934
rect 2622 319898 2678 319900
rect 2702 319898 2758 319900
rect 2782 319898 2838 319900
rect 2862 319898 2918 319900
rect 2622 319846 2648 319898
rect 2648 319846 2678 319898
rect 2702 319846 2712 319898
rect 2712 319846 2758 319898
rect 2782 319846 2828 319898
rect 2828 319846 2838 319898
rect 2862 319846 2892 319898
rect 2892 319846 2918 319898
rect 2622 319844 2678 319846
rect 2702 319844 2758 319846
rect 2782 319844 2838 319846
rect 2862 319844 2918 319846
rect 2622 318810 2678 318812
rect 2702 318810 2758 318812
rect 2782 318810 2838 318812
rect 2862 318810 2918 318812
rect 2622 318758 2648 318810
rect 2648 318758 2678 318810
rect 2702 318758 2712 318810
rect 2712 318758 2758 318810
rect 2782 318758 2828 318810
rect 2828 318758 2838 318810
rect 2862 318758 2892 318810
rect 2892 318758 2918 318810
rect 2622 318756 2678 318758
rect 2702 318756 2758 318758
rect 2782 318756 2838 318758
rect 2862 318756 2918 318758
rect 2622 317722 2678 317724
rect 2702 317722 2758 317724
rect 2782 317722 2838 317724
rect 2862 317722 2918 317724
rect 2622 317670 2648 317722
rect 2648 317670 2678 317722
rect 2702 317670 2712 317722
rect 2712 317670 2758 317722
rect 2782 317670 2828 317722
rect 2828 317670 2838 317722
rect 2862 317670 2892 317722
rect 2892 317670 2918 317722
rect 2622 317668 2678 317670
rect 2702 317668 2758 317670
rect 2782 317668 2838 317670
rect 2862 317668 2918 317670
rect 2622 316634 2678 316636
rect 2702 316634 2758 316636
rect 2782 316634 2838 316636
rect 2862 316634 2918 316636
rect 2622 316582 2648 316634
rect 2648 316582 2678 316634
rect 2702 316582 2712 316634
rect 2712 316582 2758 316634
rect 2782 316582 2828 316634
rect 2828 316582 2838 316634
rect 2862 316582 2892 316634
rect 2892 316582 2918 316634
rect 2622 316580 2678 316582
rect 2702 316580 2758 316582
rect 2782 316580 2838 316582
rect 2862 316580 2918 316582
rect 2622 315546 2678 315548
rect 2702 315546 2758 315548
rect 2782 315546 2838 315548
rect 2862 315546 2918 315548
rect 2622 315494 2648 315546
rect 2648 315494 2678 315546
rect 2702 315494 2712 315546
rect 2712 315494 2758 315546
rect 2782 315494 2828 315546
rect 2828 315494 2838 315546
rect 2862 315494 2892 315546
rect 2892 315494 2918 315546
rect 2622 315492 2678 315494
rect 2702 315492 2758 315494
rect 2782 315492 2838 315494
rect 2862 315492 2918 315494
rect 2622 314458 2678 314460
rect 2702 314458 2758 314460
rect 2782 314458 2838 314460
rect 2862 314458 2918 314460
rect 2622 314406 2648 314458
rect 2648 314406 2678 314458
rect 2702 314406 2712 314458
rect 2712 314406 2758 314458
rect 2782 314406 2828 314458
rect 2828 314406 2838 314458
rect 2862 314406 2892 314458
rect 2892 314406 2918 314458
rect 2622 314404 2678 314406
rect 2702 314404 2758 314406
rect 2782 314404 2838 314406
rect 2862 314404 2918 314406
rect 2622 313370 2678 313372
rect 2702 313370 2758 313372
rect 2782 313370 2838 313372
rect 2862 313370 2918 313372
rect 2622 313318 2648 313370
rect 2648 313318 2678 313370
rect 2702 313318 2712 313370
rect 2712 313318 2758 313370
rect 2782 313318 2828 313370
rect 2828 313318 2838 313370
rect 2862 313318 2892 313370
rect 2892 313318 2918 313370
rect 2622 313316 2678 313318
rect 2702 313316 2758 313318
rect 2782 313316 2838 313318
rect 2862 313316 2918 313318
rect 2622 312282 2678 312284
rect 2702 312282 2758 312284
rect 2782 312282 2838 312284
rect 2862 312282 2918 312284
rect 2622 312230 2648 312282
rect 2648 312230 2678 312282
rect 2702 312230 2712 312282
rect 2712 312230 2758 312282
rect 2782 312230 2828 312282
rect 2828 312230 2838 312282
rect 2862 312230 2892 312282
rect 2892 312230 2918 312282
rect 2622 312228 2678 312230
rect 2702 312228 2758 312230
rect 2782 312228 2838 312230
rect 2862 312228 2918 312230
rect 2622 311194 2678 311196
rect 2702 311194 2758 311196
rect 2782 311194 2838 311196
rect 2862 311194 2918 311196
rect 2622 311142 2648 311194
rect 2648 311142 2678 311194
rect 2702 311142 2712 311194
rect 2712 311142 2758 311194
rect 2782 311142 2828 311194
rect 2828 311142 2838 311194
rect 2862 311142 2892 311194
rect 2892 311142 2918 311194
rect 2622 311140 2678 311142
rect 2702 311140 2758 311142
rect 2782 311140 2838 311142
rect 2862 311140 2918 311142
rect 2622 310106 2678 310108
rect 2702 310106 2758 310108
rect 2782 310106 2838 310108
rect 2862 310106 2918 310108
rect 2622 310054 2648 310106
rect 2648 310054 2678 310106
rect 2702 310054 2712 310106
rect 2712 310054 2758 310106
rect 2782 310054 2828 310106
rect 2828 310054 2838 310106
rect 2862 310054 2892 310106
rect 2892 310054 2918 310106
rect 2622 310052 2678 310054
rect 2702 310052 2758 310054
rect 2782 310052 2838 310054
rect 2862 310052 2918 310054
rect 2622 309018 2678 309020
rect 2702 309018 2758 309020
rect 2782 309018 2838 309020
rect 2862 309018 2918 309020
rect 2622 308966 2648 309018
rect 2648 308966 2678 309018
rect 2702 308966 2712 309018
rect 2712 308966 2758 309018
rect 2782 308966 2828 309018
rect 2828 308966 2838 309018
rect 2862 308966 2892 309018
rect 2892 308966 2918 309018
rect 2622 308964 2678 308966
rect 2702 308964 2758 308966
rect 2782 308964 2838 308966
rect 2862 308964 2918 308966
rect 2226 308624 2282 308680
rect 2622 307930 2678 307932
rect 2702 307930 2758 307932
rect 2782 307930 2838 307932
rect 2862 307930 2918 307932
rect 2622 307878 2648 307930
rect 2648 307878 2678 307930
rect 2702 307878 2712 307930
rect 2712 307878 2758 307930
rect 2782 307878 2828 307930
rect 2828 307878 2838 307930
rect 2862 307878 2892 307930
rect 2892 307878 2918 307930
rect 2622 307876 2678 307878
rect 2702 307876 2758 307878
rect 2782 307876 2838 307878
rect 2862 307876 2918 307878
rect 2622 306842 2678 306844
rect 2702 306842 2758 306844
rect 2782 306842 2838 306844
rect 2862 306842 2918 306844
rect 2622 306790 2648 306842
rect 2648 306790 2678 306842
rect 2702 306790 2712 306842
rect 2712 306790 2758 306842
rect 2782 306790 2828 306842
rect 2828 306790 2838 306842
rect 2862 306790 2892 306842
rect 2892 306790 2918 306842
rect 2622 306788 2678 306790
rect 2702 306788 2758 306790
rect 2782 306788 2838 306790
rect 2862 306788 2918 306790
rect 2622 305754 2678 305756
rect 2702 305754 2758 305756
rect 2782 305754 2838 305756
rect 2862 305754 2918 305756
rect 2622 305702 2648 305754
rect 2648 305702 2678 305754
rect 2702 305702 2712 305754
rect 2712 305702 2758 305754
rect 2782 305702 2828 305754
rect 2828 305702 2838 305754
rect 2862 305702 2892 305754
rect 2892 305702 2918 305754
rect 2622 305700 2678 305702
rect 2702 305700 2758 305702
rect 2782 305700 2838 305702
rect 2862 305700 2918 305702
rect 2622 304666 2678 304668
rect 2702 304666 2758 304668
rect 2782 304666 2838 304668
rect 2862 304666 2918 304668
rect 2622 304614 2648 304666
rect 2648 304614 2678 304666
rect 2702 304614 2712 304666
rect 2712 304614 2758 304666
rect 2782 304614 2828 304666
rect 2828 304614 2838 304666
rect 2862 304614 2892 304666
rect 2892 304614 2918 304666
rect 2622 304612 2678 304614
rect 2702 304612 2758 304614
rect 2782 304612 2838 304614
rect 2862 304612 2918 304614
rect 2622 303578 2678 303580
rect 2702 303578 2758 303580
rect 2782 303578 2838 303580
rect 2862 303578 2918 303580
rect 2622 303526 2648 303578
rect 2648 303526 2678 303578
rect 2702 303526 2712 303578
rect 2712 303526 2758 303578
rect 2782 303526 2828 303578
rect 2828 303526 2838 303578
rect 2862 303526 2892 303578
rect 2892 303526 2918 303578
rect 2622 303524 2678 303526
rect 2702 303524 2758 303526
rect 2782 303524 2838 303526
rect 2862 303524 2918 303526
rect 2622 302490 2678 302492
rect 2702 302490 2758 302492
rect 2782 302490 2838 302492
rect 2862 302490 2918 302492
rect 2622 302438 2648 302490
rect 2648 302438 2678 302490
rect 2702 302438 2712 302490
rect 2712 302438 2758 302490
rect 2782 302438 2828 302490
rect 2828 302438 2838 302490
rect 2862 302438 2892 302490
rect 2892 302438 2918 302490
rect 2622 302436 2678 302438
rect 2702 302436 2758 302438
rect 2782 302436 2838 302438
rect 2862 302436 2918 302438
rect 2622 301402 2678 301404
rect 2702 301402 2758 301404
rect 2782 301402 2838 301404
rect 2862 301402 2918 301404
rect 2622 301350 2648 301402
rect 2648 301350 2678 301402
rect 2702 301350 2712 301402
rect 2712 301350 2758 301402
rect 2782 301350 2828 301402
rect 2828 301350 2838 301402
rect 2862 301350 2892 301402
rect 2892 301350 2918 301402
rect 2622 301348 2678 301350
rect 2702 301348 2758 301350
rect 2782 301348 2838 301350
rect 2862 301348 2918 301350
rect 2622 300314 2678 300316
rect 2702 300314 2758 300316
rect 2782 300314 2838 300316
rect 2862 300314 2918 300316
rect 2622 300262 2648 300314
rect 2648 300262 2678 300314
rect 2702 300262 2712 300314
rect 2712 300262 2758 300314
rect 2782 300262 2828 300314
rect 2828 300262 2838 300314
rect 2862 300262 2892 300314
rect 2892 300262 2918 300314
rect 2622 300260 2678 300262
rect 2702 300260 2758 300262
rect 2782 300260 2838 300262
rect 2862 300260 2918 300262
rect 2622 299226 2678 299228
rect 2702 299226 2758 299228
rect 2782 299226 2838 299228
rect 2862 299226 2918 299228
rect 2622 299174 2648 299226
rect 2648 299174 2678 299226
rect 2702 299174 2712 299226
rect 2712 299174 2758 299226
rect 2782 299174 2828 299226
rect 2828 299174 2838 299226
rect 2862 299174 2892 299226
rect 2892 299174 2918 299226
rect 2622 299172 2678 299174
rect 2702 299172 2758 299174
rect 2782 299172 2838 299174
rect 2862 299172 2918 299174
rect 2622 298138 2678 298140
rect 2702 298138 2758 298140
rect 2782 298138 2838 298140
rect 2862 298138 2918 298140
rect 2622 298086 2648 298138
rect 2648 298086 2678 298138
rect 2702 298086 2712 298138
rect 2712 298086 2758 298138
rect 2782 298086 2828 298138
rect 2828 298086 2838 298138
rect 2862 298086 2892 298138
rect 2892 298086 2918 298138
rect 2622 298084 2678 298086
rect 2702 298084 2758 298086
rect 2782 298084 2838 298086
rect 2862 298084 2918 298086
rect 2622 297050 2678 297052
rect 2702 297050 2758 297052
rect 2782 297050 2838 297052
rect 2862 297050 2918 297052
rect 2622 296998 2648 297050
rect 2648 296998 2678 297050
rect 2702 296998 2712 297050
rect 2712 296998 2758 297050
rect 2782 296998 2828 297050
rect 2828 296998 2838 297050
rect 2862 296998 2892 297050
rect 2892 296998 2918 297050
rect 2622 296996 2678 296998
rect 2702 296996 2758 296998
rect 2782 296996 2838 296998
rect 2862 296996 2918 296998
rect 2622 295962 2678 295964
rect 2702 295962 2758 295964
rect 2782 295962 2838 295964
rect 2862 295962 2918 295964
rect 2622 295910 2648 295962
rect 2648 295910 2678 295962
rect 2702 295910 2712 295962
rect 2712 295910 2758 295962
rect 2782 295910 2828 295962
rect 2828 295910 2838 295962
rect 2862 295910 2892 295962
rect 2892 295910 2918 295962
rect 2622 295908 2678 295910
rect 2702 295908 2758 295910
rect 2782 295908 2838 295910
rect 2862 295908 2918 295910
rect 2622 294874 2678 294876
rect 2702 294874 2758 294876
rect 2782 294874 2838 294876
rect 2862 294874 2918 294876
rect 2622 294822 2648 294874
rect 2648 294822 2678 294874
rect 2702 294822 2712 294874
rect 2712 294822 2758 294874
rect 2782 294822 2828 294874
rect 2828 294822 2838 294874
rect 2862 294822 2892 294874
rect 2892 294822 2918 294874
rect 2622 294820 2678 294822
rect 2702 294820 2758 294822
rect 2782 294820 2838 294822
rect 2862 294820 2918 294822
rect 2622 293786 2678 293788
rect 2702 293786 2758 293788
rect 2782 293786 2838 293788
rect 2862 293786 2918 293788
rect 2622 293734 2648 293786
rect 2648 293734 2678 293786
rect 2702 293734 2712 293786
rect 2712 293734 2758 293786
rect 2782 293734 2828 293786
rect 2828 293734 2838 293786
rect 2862 293734 2892 293786
rect 2892 293734 2918 293786
rect 2622 293732 2678 293734
rect 2702 293732 2758 293734
rect 2782 293732 2838 293734
rect 2862 293732 2918 293734
rect 2622 292698 2678 292700
rect 2702 292698 2758 292700
rect 2782 292698 2838 292700
rect 2862 292698 2918 292700
rect 2622 292646 2648 292698
rect 2648 292646 2678 292698
rect 2702 292646 2712 292698
rect 2712 292646 2758 292698
rect 2782 292646 2828 292698
rect 2828 292646 2838 292698
rect 2862 292646 2892 292698
rect 2892 292646 2918 292698
rect 2622 292644 2678 292646
rect 2702 292644 2758 292646
rect 2782 292644 2838 292646
rect 2862 292644 2918 292646
rect 2622 291610 2678 291612
rect 2702 291610 2758 291612
rect 2782 291610 2838 291612
rect 2862 291610 2918 291612
rect 2622 291558 2648 291610
rect 2648 291558 2678 291610
rect 2702 291558 2712 291610
rect 2712 291558 2758 291610
rect 2782 291558 2828 291610
rect 2828 291558 2838 291610
rect 2862 291558 2892 291610
rect 2892 291558 2918 291610
rect 2622 291556 2678 291558
rect 2702 291556 2758 291558
rect 2782 291556 2838 291558
rect 2862 291556 2918 291558
rect 2622 290522 2678 290524
rect 2702 290522 2758 290524
rect 2782 290522 2838 290524
rect 2862 290522 2918 290524
rect 2622 290470 2648 290522
rect 2648 290470 2678 290522
rect 2702 290470 2712 290522
rect 2712 290470 2758 290522
rect 2782 290470 2828 290522
rect 2828 290470 2838 290522
rect 2862 290470 2892 290522
rect 2892 290470 2918 290522
rect 2622 290468 2678 290470
rect 2702 290468 2758 290470
rect 2782 290468 2838 290470
rect 2862 290468 2918 290470
rect 2622 289434 2678 289436
rect 2702 289434 2758 289436
rect 2782 289434 2838 289436
rect 2862 289434 2918 289436
rect 2622 289382 2648 289434
rect 2648 289382 2678 289434
rect 2702 289382 2712 289434
rect 2712 289382 2758 289434
rect 2782 289382 2828 289434
rect 2828 289382 2838 289434
rect 2862 289382 2892 289434
rect 2892 289382 2918 289434
rect 2622 289380 2678 289382
rect 2702 289380 2758 289382
rect 2782 289380 2838 289382
rect 2862 289380 2918 289382
rect 2622 288346 2678 288348
rect 2702 288346 2758 288348
rect 2782 288346 2838 288348
rect 2862 288346 2918 288348
rect 2622 288294 2648 288346
rect 2648 288294 2678 288346
rect 2702 288294 2712 288346
rect 2712 288294 2758 288346
rect 2782 288294 2828 288346
rect 2828 288294 2838 288346
rect 2862 288294 2892 288346
rect 2892 288294 2918 288346
rect 2622 288292 2678 288294
rect 2702 288292 2758 288294
rect 2782 288292 2838 288294
rect 2862 288292 2918 288294
rect 2622 287258 2678 287260
rect 2702 287258 2758 287260
rect 2782 287258 2838 287260
rect 2862 287258 2918 287260
rect 2622 287206 2648 287258
rect 2648 287206 2678 287258
rect 2702 287206 2712 287258
rect 2712 287206 2758 287258
rect 2782 287206 2828 287258
rect 2828 287206 2838 287258
rect 2862 287206 2892 287258
rect 2892 287206 2918 287258
rect 2622 287204 2678 287206
rect 2702 287204 2758 287206
rect 2782 287204 2838 287206
rect 2862 287204 2918 287206
rect 2622 286170 2678 286172
rect 2702 286170 2758 286172
rect 2782 286170 2838 286172
rect 2862 286170 2918 286172
rect 2622 286118 2648 286170
rect 2648 286118 2678 286170
rect 2702 286118 2712 286170
rect 2712 286118 2758 286170
rect 2782 286118 2828 286170
rect 2828 286118 2838 286170
rect 2862 286118 2892 286170
rect 2892 286118 2918 286170
rect 2622 286116 2678 286118
rect 2702 286116 2758 286118
rect 2782 286116 2838 286118
rect 2862 286116 2918 286118
rect 2622 285082 2678 285084
rect 2702 285082 2758 285084
rect 2782 285082 2838 285084
rect 2862 285082 2918 285084
rect 2622 285030 2648 285082
rect 2648 285030 2678 285082
rect 2702 285030 2712 285082
rect 2712 285030 2758 285082
rect 2782 285030 2828 285082
rect 2828 285030 2838 285082
rect 2862 285030 2892 285082
rect 2892 285030 2918 285082
rect 2622 285028 2678 285030
rect 2702 285028 2758 285030
rect 2782 285028 2838 285030
rect 2862 285028 2918 285030
rect 2622 283994 2678 283996
rect 2702 283994 2758 283996
rect 2782 283994 2838 283996
rect 2862 283994 2918 283996
rect 2622 283942 2648 283994
rect 2648 283942 2678 283994
rect 2702 283942 2712 283994
rect 2712 283942 2758 283994
rect 2782 283942 2828 283994
rect 2828 283942 2838 283994
rect 2862 283942 2892 283994
rect 2892 283942 2918 283994
rect 2622 283940 2678 283942
rect 2702 283940 2758 283942
rect 2782 283940 2838 283942
rect 2862 283940 2918 283942
rect 2622 282906 2678 282908
rect 2702 282906 2758 282908
rect 2782 282906 2838 282908
rect 2862 282906 2918 282908
rect 2622 282854 2648 282906
rect 2648 282854 2678 282906
rect 2702 282854 2712 282906
rect 2712 282854 2758 282906
rect 2782 282854 2828 282906
rect 2828 282854 2838 282906
rect 2862 282854 2892 282906
rect 2892 282854 2918 282906
rect 2622 282852 2678 282854
rect 2702 282852 2758 282854
rect 2782 282852 2838 282854
rect 2862 282852 2918 282854
rect 2622 281818 2678 281820
rect 2702 281818 2758 281820
rect 2782 281818 2838 281820
rect 2862 281818 2918 281820
rect 2622 281766 2648 281818
rect 2648 281766 2678 281818
rect 2702 281766 2712 281818
rect 2712 281766 2758 281818
rect 2782 281766 2828 281818
rect 2828 281766 2838 281818
rect 2862 281766 2892 281818
rect 2892 281766 2918 281818
rect 2622 281764 2678 281766
rect 2702 281764 2758 281766
rect 2782 281764 2838 281766
rect 2862 281764 2918 281766
rect 2622 280730 2678 280732
rect 2702 280730 2758 280732
rect 2782 280730 2838 280732
rect 2862 280730 2918 280732
rect 2622 280678 2648 280730
rect 2648 280678 2678 280730
rect 2702 280678 2712 280730
rect 2712 280678 2758 280730
rect 2782 280678 2828 280730
rect 2828 280678 2838 280730
rect 2862 280678 2892 280730
rect 2892 280678 2918 280730
rect 2622 280676 2678 280678
rect 2702 280676 2758 280678
rect 2782 280676 2838 280678
rect 2862 280676 2918 280678
rect 2622 279642 2678 279644
rect 2702 279642 2758 279644
rect 2782 279642 2838 279644
rect 2862 279642 2918 279644
rect 2622 279590 2648 279642
rect 2648 279590 2678 279642
rect 2702 279590 2712 279642
rect 2712 279590 2758 279642
rect 2782 279590 2828 279642
rect 2828 279590 2838 279642
rect 2862 279590 2892 279642
rect 2892 279590 2918 279642
rect 2622 279588 2678 279590
rect 2702 279588 2758 279590
rect 2782 279588 2838 279590
rect 2862 279588 2918 279590
rect 2622 278554 2678 278556
rect 2702 278554 2758 278556
rect 2782 278554 2838 278556
rect 2862 278554 2918 278556
rect 2622 278502 2648 278554
rect 2648 278502 2678 278554
rect 2702 278502 2712 278554
rect 2712 278502 2758 278554
rect 2782 278502 2828 278554
rect 2828 278502 2838 278554
rect 2862 278502 2892 278554
rect 2892 278502 2918 278554
rect 2622 278500 2678 278502
rect 2702 278500 2758 278502
rect 2782 278500 2838 278502
rect 2862 278500 2918 278502
rect 2622 277466 2678 277468
rect 2702 277466 2758 277468
rect 2782 277466 2838 277468
rect 2862 277466 2918 277468
rect 2622 277414 2648 277466
rect 2648 277414 2678 277466
rect 2702 277414 2712 277466
rect 2712 277414 2758 277466
rect 2782 277414 2828 277466
rect 2828 277414 2838 277466
rect 2862 277414 2892 277466
rect 2892 277414 2918 277466
rect 2622 277412 2678 277414
rect 2702 277412 2758 277414
rect 2782 277412 2838 277414
rect 2862 277412 2918 277414
rect 2622 276378 2678 276380
rect 2702 276378 2758 276380
rect 2782 276378 2838 276380
rect 2862 276378 2918 276380
rect 2622 276326 2648 276378
rect 2648 276326 2678 276378
rect 2702 276326 2712 276378
rect 2712 276326 2758 276378
rect 2782 276326 2828 276378
rect 2828 276326 2838 276378
rect 2862 276326 2892 276378
rect 2892 276326 2918 276378
rect 2622 276324 2678 276326
rect 2702 276324 2758 276326
rect 2782 276324 2838 276326
rect 2862 276324 2918 276326
rect 2622 275290 2678 275292
rect 2702 275290 2758 275292
rect 2782 275290 2838 275292
rect 2862 275290 2918 275292
rect 2622 275238 2648 275290
rect 2648 275238 2678 275290
rect 2702 275238 2712 275290
rect 2712 275238 2758 275290
rect 2782 275238 2828 275290
rect 2828 275238 2838 275290
rect 2862 275238 2892 275290
rect 2892 275238 2918 275290
rect 2622 275236 2678 275238
rect 2702 275236 2758 275238
rect 2782 275236 2838 275238
rect 2862 275236 2918 275238
rect 2622 274202 2678 274204
rect 2702 274202 2758 274204
rect 2782 274202 2838 274204
rect 2862 274202 2918 274204
rect 2622 274150 2648 274202
rect 2648 274150 2678 274202
rect 2702 274150 2712 274202
rect 2712 274150 2758 274202
rect 2782 274150 2828 274202
rect 2828 274150 2838 274202
rect 2862 274150 2892 274202
rect 2892 274150 2918 274202
rect 2622 274148 2678 274150
rect 2702 274148 2758 274150
rect 2782 274148 2838 274150
rect 2862 274148 2918 274150
rect 2622 273114 2678 273116
rect 2702 273114 2758 273116
rect 2782 273114 2838 273116
rect 2862 273114 2918 273116
rect 2622 273062 2648 273114
rect 2648 273062 2678 273114
rect 2702 273062 2712 273114
rect 2712 273062 2758 273114
rect 2782 273062 2828 273114
rect 2828 273062 2838 273114
rect 2862 273062 2892 273114
rect 2892 273062 2918 273114
rect 2622 273060 2678 273062
rect 2702 273060 2758 273062
rect 2782 273060 2838 273062
rect 2862 273060 2918 273062
rect 2622 272026 2678 272028
rect 2702 272026 2758 272028
rect 2782 272026 2838 272028
rect 2862 272026 2918 272028
rect 2622 271974 2648 272026
rect 2648 271974 2678 272026
rect 2702 271974 2712 272026
rect 2712 271974 2758 272026
rect 2782 271974 2828 272026
rect 2828 271974 2838 272026
rect 2862 271974 2892 272026
rect 2892 271974 2918 272026
rect 2622 271972 2678 271974
rect 2702 271972 2758 271974
rect 2782 271972 2838 271974
rect 2862 271972 2918 271974
rect 2622 270938 2678 270940
rect 2702 270938 2758 270940
rect 2782 270938 2838 270940
rect 2862 270938 2918 270940
rect 2622 270886 2648 270938
rect 2648 270886 2678 270938
rect 2702 270886 2712 270938
rect 2712 270886 2758 270938
rect 2782 270886 2828 270938
rect 2828 270886 2838 270938
rect 2862 270886 2892 270938
rect 2892 270886 2918 270938
rect 2622 270884 2678 270886
rect 2702 270884 2758 270886
rect 2782 270884 2838 270886
rect 2862 270884 2918 270886
rect 2622 269850 2678 269852
rect 2702 269850 2758 269852
rect 2782 269850 2838 269852
rect 2862 269850 2918 269852
rect 2622 269798 2648 269850
rect 2648 269798 2678 269850
rect 2702 269798 2712 269850
rect 2712 269798 2758 269850
rect 2782 269798 2828 269850
rect 2828 269798 2838 269850
rect 2862 269798 2892 269850
rect 2892 269798 2918 269850
rect 2622 269796 2678 269798
rect 2702 269796 2758 269798
rect 2782 269796 2838 269798
rect 2862 269796 2918 269798
rect 2622 268762 2678 268764
rect 2702 268762 2758 268764
rect 2782 268762 2838 268764
rect 2862 268762 2918 268764
rect 2622 268710 2648 268762
rect 2648 268710 2678 268762
rect 2702 268710 2712 268762
rect 2712 268710 2758 268762
rect 2782 268710 2828 268762
rect 2828 268710 2838 268762
rect 2862 268710 2892 268762
rect 2892 268710 2918 268762
rect 2622 268708 2678 268710
rect 2702 268708 2758 268710
rect 2782 268708 2838 268710
rect 2862 268708 2918 268710
rect 2622 267674 2678 267676
rect 2702 267674 2758 267676
rect 2782 267674 2838 267676
rect 2862 267674 2918 267676
rect 2622 267622 2648 267674
rect 2648 267622 2678 267674
rect 2702 267622 2712 267674
rect 2712 267622 2758 267674
rect 2782 267622 2828 267674
rect 2828 267622 2838 267674
rect 2862 267622 2892 267674
rect 2892 267622 2918 267674
rect 2622 267620 2678 267622
rect 2702 267620 2758 267622
rect 2782 267620 2838 267622
rect 2862 267620 2918 267622
rect 2622 266586 2678 266588
rect 2702 266586 2758 266588
rect 2782 266586 2838 266588
rect 2862 266586 2918 266588
rect 2622 266534 2648 266586
rect 2648 266534 2678 266586
rect 2702 266534 2712 266586
rect 2712 266534 2758 266586
rect 2782 266534 2828 266586
rect 2828 266534 2838 266586
rect 2862 266534 2892 266586
rect 2892 266534 2918 266586
rect 2622 266532 2678 266534
rect 2702 266532 2758 266534
rect 2782 266532 2838 266534
rect 2862 266532 2918 266534
rect 2622 265498 2678 265500
rect 2702 265498 2758 265500
rect 2782 265498 2838 265500
rect 2862 265498 2918 265500
rect 2622 265446 2648 265498
rect 2648 265446 2678 265498
rect 2702 265446 2712 265498
rect 2712 265446 2758 265498
rect 2782 265446 2828 265498
rect 2828 265446 2838 265498
rect 2862 265446 2892 265498
rect 2892 265446 2918 265498
rect 2622 265444 2678 265446
rect 2702 265444 2758 265446
rect 2782 265444 2838 265446
rect 2862 265444 2918 265446
rect 2622 264410 2678 264412
rect 2702 264410 2758 264412
rect 2782 264410 2838 264412
rect 2862 264410 2918 264412
rect 2622 264358 2648 264410
rect 2648 264358 2678 264410
rect 2702 264358 2712 264410
rect 2712 264358 2758 264410
rect 2782 264358 2828 264410
rect 2828 264358 2838 264410
rect 2862 264358 2892 264410
rect 2892 264358 2918 264410
rect 2622 264356 2678 264358
rect 2702 264356 2758 264358
rect 2782 264356 2838 264358
rect 2862 264356 2918 264358
rect 2622 263322 2678 263324
rect 2702 263322 2758 263324
rect 2782 263322 2838 263324
rect 2862 263322 2918 263324
rect 2622 263270 2648 263322
rect 2648 263270 2678 263322
rect 2702 263270 2712 263322
rect 2712 263270 2758 263322
rect 2782 263270 2828 263322
rect 2828 263270 2838 263322
rect 2862 263270 2892 263322
rect 2892 263270 2918 263322
rect 2622 263268 2678 263270
rect 2702 263268 2758 263270
rect 2782 263268 2838 263270
rect 2862 263268 2918 263270
rect 2622 262234 2678 262236
rect 2702 262234 2758 262236
rect 2782 262234 2838 262236
rect 2862 262234 2918 262236
rect 2622 262182 2648 262234
rect 2648 262182 2678 262234
rect 2702 262182 2712 262234
rect 2712 262182 2758 262234
rect 2782 262182 2828 262234
rect 2828 262182 2838 262234
rect 2862 262182 2892 262234
rect 2892 262182 2918 262234
rect 2622 262180 2678 262182
rect 2702 262180 2758 262182
rect 2782 262180 2838 262182
rect 2862 262180 2918 262182
rect 2502 261296 2558 261352
rect 2622 261146 2678 261148
rect 2702 261146 2758 261148
rect 2782 261146 2838 261148
rect 2862 261146 2918 261148
rect 2622 261094 2648 261146
rect 2648 261094 2678 261146
rect 2702 261094 2712 261146
rect 2712 261094 2758 261146
rect 2782 261094 2828 261146
rect 2828 261094 2838 261146
rect 2862 261094 2892 261146
rect 2892 261094 2918 261146
rect 2622 261092 2678 261094
rect 2702 261092 2758 261094
rect 2782 261092 2838 261094
rect 2862 261092 2918 261094
rect 2622 260058 2678 260060
rect 2702 260058 2758 260060
rect 2782 260058 2838 260060
rect 2862 260058 2918 260060
rect 2622 260006 2648 260058
rect 2648 260006 2678 260058
rect 2702 260006 2712 260058
rect 2712 260006 2758 260058
rect 2782 260006 2828 260058
rect 2828 260006 2838 260058
rect 2862 260006 2892 260058
rect 2892 260006 2918 260058
rect 2622 260004 2678 260006
rect 2702 260004 2758 260006
rect 2782 260004 2838 260006
rect 2862 260004 2918 260006
rect 2622 258970 2678 258972
rect 2702 258970 2758 258972
rect 2782 258970 2838 258972
rect 2862 258970 2918 258972
rect 2622 258918 2648 258970
rect 2648 258918 2678 258970
rect 2702 258918 2712 258970
rect 2712 258918 2758 258970
rect 2782 258918 2828 258970
rect 2828 258918 2838 258970
rect 2862 258918 2892 258970
rect 2892 258918 2918 258970
rect 2622 258916 2678 258918
rect 2702 258916 2758 258918
rect 2782 258916 2838 258918
rect 2862 258916 2918 258918
rect 2622 257882 2678 257884
rect 2702 257882 2758 257884
rect 2782 257882 2838 257884
rect 2862 257882 2918 257884
rect 2622 257830 2648 257882
rect 2648 257830 2678 257882
rect 2702 257830 2712 257882
rect 2712 257830 2758 257882
rect 2782 257830 2828 257882
rect 2828 257830 2838 257882
rect 2862 257830 2892 257882
rect 2892 257830 2918 257882
rect 2622 257828 2678 257830
rect 2702 257828 2758 257830
rect 2782 257828 2838 257830
rect 2862 257828 2918 257830
rect 2622 256794 2678 256796
rect 2702 256794 2758 256796
rect 2782 256794 2838 256796
rect 2862 256794 2918 256796
rect 2622 256742 2648 256794
rect 2648 256742 2678 256794
rect 2702 256742 2712 256794
rect 2712 256742 2758 256794
rect 2782 256742 2828 256794
rect 2828 256742 2838 256794
rect 2862 256742 2892 256794
rect 2892 256742 2918 256794
rect 2622 256740 2678 256742
rect 2702 256740 2758 256742
rect 2782 256740 2838 256742
rect 2862 256740 2918 256742
rect 2622 255706 2678 255708
rect 2702 255706 2758 255708
rect 2782 255706 2838 255708
rect 2862 255706 2918 255708
rect 2622 255654 2648 255706
rect 2648 255654 2678 255706
rect 2702 255654 2712 255706
rect 2712 255654 2758 255706
rect 2782 255654 2828 255706
rect 2828 255654 2838 255706
rect 2862 255654 2892 255706
rect 2892 255654 2918 255706
rect 2622 255652 2678 255654
rect 2702 255652 2758 255654
rect 2782 255652 2838 255654
rect 2862 255652 2918 255654
rect 2622 254618 2678 254620
rect 2702 254618 2758 254620
rect 2782 254618 2838 254620
rect 2862 254618 2918 254620
rect 2622 254566 2648 254618
rect 2648 254566 2678 254618
rect 2702 254566 2712 254618
rect 2712 254566 2758 254618
rect 2782 254566 2828 254618
rect 2828 254566 2838 254618
rect 2862 254566 2892 254618
rect 2892 254566 2918 254618
rect 2622 254564 2678 254566
rect 2702 254564 2758 254566
rect 2782 254564 2838 254566
rect 2862 254564 2918 254566
rect 2622 253530 2678 253532
rect 2702 253530 2758 253532
rect 2782 253530 2838 253532
rect 2862 253530 2918 253532
rect 2622 253478 2648 253530
rect 2648 253478 2678 253530
rect 2702 253478 2712 253530
rect 2712 253478 2758 253530
rect 2782 253478 2828 253530
rect 2828 253478 2838 253530
rect 2862 253478 2892 253530
rect 2892 253478 2918 253530
rect 2622 253476 2678 253478
rect 2702 253476 2758 253478
rect 2782 253476 2838 253478
rect 2862 253476 2918 253478
rect 2622 252442 2678 252444
rect 2702 252442 2758 252444
rect 2782 252442 2838 252444
rect 2862 252442 2918 252444
rect 2622 252390 2648 252442
rect 2648 252390 2678 252442
rect 2702 252390 2712 252442
rect 2712 252390 2758 252442
rect 2782 252390 2828 252442
rect 2828 252390 2838 252442
rect 2862 252390 2892 252442
rect 2892 252390 2918 252442
rect 2622 252388 2678 252390
rect 2702 252388 2758 252390
rect 2782 252388 2838 252390
rect 2862 252388 2918 252390
rect 2622 251354 2678 251356
rect 2702 251354 2758 251356
rect 2782 251354 2838 251356
rect 2862 251354 2918 251356
rect 2622 251302 2648 251354
rect 2648 251302 2678 251354
rect 2702 251302 2712 251354
rect 2712 251302 2758 251354
rect 2782 251302 2828 251354
rect 2828 251302 2838 251354
rect 2862 251302 2892 251354
rect 2892 251302 2918 251354
rect 2622 251300 2678 251302
rect 2702 251300 2758 251302
rect 2782 251300 2838 251302
rect 2862 251300 2918 251302
rect 2622 250266 2678 250268
rect 2702 250266 2758 250268
rect 2782 250266 2838 250268
rect 2862 250266 2918 250268
rect 2622 250214 2648 250266
rect 2648 250214 2678 250266
rect 2702 250214 2712 250266
rect 2712 250214 2758 250266
rect 2782 250214 2828 250266
rect 2828 250214 2838 250266
rect 2862 250214 2892 250266
rect 2892 250214 2918 250266
rect 2622 250212 2678 250214
rect 2702 250212 2758 250214
rect 2782 250212 2838 250214
rect 2862 250212 2918 250214
rect 2622 249178 2678 249180
rect 2702 249178 2758 249180
rect 2782 249178 2838 249180
rect 2862 249178 2918 249180
rect 2622 249126 2648 249178
rect 2648 249126 2678 249178
rect 2702 249126 2712 249178
rect 2712 249126 2758 249178
rect 2782 249126 2828 249178
rect 2828 249126 2838 249178
rect 2862 249126 2892 249178
rect 2892 249126 2918 249178
rect 2622 249124 2678 249126
rect 2702 249124 2758 249126
rect 2782 249124 2838 249126
rect 2862 249124 2918 249126
rect 2622 248090 2678 248092
rect 2702 248090 2758 248092
rect 2782 248090 2838 248092
rect 2862 248090 2918 248092
rect 2622 248038 2648 248090
rect 2648 248038 2678 248090
rect 2702 248038 2712 248090
rect 2712 248038 2758 248090
rect 2782 248038 2828 248090
rect 2828 248038 2838 248090
rect 2862 248038 2892 248090
rect 2892 248038 2918 248090
rect 2622 248036 2678 248038
rect 2702 248036 2758 248038
rect 2782 248036 2838 248038
rect 2862 248036 2918 248038
rect 2622 247002 2678 247004
rect 2702 247002 2758 247004
rect 2782 247002 2838 247004
rect 2862 247002 2918 247004
rect 2622 246950 2648 247002
rect 2648 246950 2678 247002
rect 2702 246950 2712 247002
rect 2712 246950 2758 247002
rect 2782 246950 2828 247002
rect 2828 246950 2838 247002
rect 2862 246950 2892 247002
rect 2892 246950 2918 247002
rect 2622 246948 2678 246950
rect 2702 246948 2758 246950
rect 2782 246948 2838 246950
rect 2862 246948 2918 246950
rect 2622 245914 2678 245916
rect 2702 245914 2758 245916
rect 2782 245914 2838 245916
rect 2862 245914 2918 245916
rect 2622 245862 2648 245914
rect 2648 245862 2678 245914
rect 2702 245862 2712 245914
rect 2712 245862 2758 245914
rect 2782 245862 2828 245914
rect 2828 245862 2838 245914
rect 2862 245862 2892 245914
rect 2892 245862 2918 245914
rect 2622 245860 2678 245862
rect 2702 245860 2758 245862
rect 2782 245860 2838 245862
rect 2862 245860 2918 245862
rect 2622 244826 2678 244828
rect 2702 244826 2758 244828
rect 2782 244826 2838 244828
rect 2862 244826 2918 244828
rect 2622 244774 2648 244826
rect 2648 244774 2678 244826
rect 2702 244774 2712 244826
rect 2712 244774 2758 244826
rect 2782 244774 2828 244826
rect 2828 244774 2838 244826
rect 2862 244774 2892 244826
rect 2892 244774 2918 244826
rect 2622 244772 2678 244774
rect 2702 244772 2758 244774
rect 2782 244772 2838 244774
rect 2862 244772 2918 244774
rect 2622 243738 2678 243740
rect 2702 243738 2758 243740
rect 2782 243738 2838 243740
rect 2862 243738 2918 243740
rect 2622 243686 2648 243738
rect 2648 243686 2678 243738
rect 2702 243686 2712 243738
rect 2712 243686 2758 243738
rect 2782 243686 2828 243738
rect 2828 243686 2838 243738
rect 2862 243686 2892 243738
rect 2892 243686 2918 243738
rect 2622 243684 2678 243686
rect 2702 243684 2758 243686
rect 2782 243684 2838 243686
rect 2862 243684 2918 243686
rect 2622 242650 2678 242652
rect 2702 242650 2758 242652
rect 2782 242650 2838 242652
rect 2862 242650 2918 242652
rect 2622 242598 2648 242650
rect 2648 242598 2678 242650
rect 2702 242598 2712 242650
rect 2712 242598 2758 242650
rect 2782 242598 2828 242650
rect 2828 242598 2838 242650
rect 2862 242598 2892 242650
rect 2892 242598 2918 242650
rect 2622 242596 2678 242598
rect 2702 242596 2758 242598
rect 2782 242596 2838 242598
rect 2862 242596 2918 242598
rect 2622 241562 2678 241564
rect 2702 241562 2758 241564
rect 2782 241562 2838 241564
rect 2862 241562 2918 241564
rect 2622 241510 2648 241562
rect 2648 241510 2678 241562
rect 2702 241510 2712 241562
rect 2712 241510 2758 241562
rect 2782 241510 2828 241562
rect 2828 241510 2838 241562
rect 2862 241510 2892 241562
rect 2892 241510 2918 241562
rect 2622 241508 2678 241510
rect 2702 241508 2758 241510
rect 2782 241508 2838 241510
rect 2862 241508 2918 241510
rect 2622 240474 2678 240476
rect 2702 240474 2758 240476
rect 2782 240474 2838 240476
rect 2862 240474 2918 240476
rect 2622 240422 2648 240474
rect 2648 240422 2678 240474
rect 2702 240422 2712 240474
rect 2712 240422 2758 240474
rect 2782 240422 2828 240474
rect 2828 240422 2838 240474
rect 2862 240422 2892 240474
rect 2892 240422 2918 240474
rect 2622 240420 2678 240422
rect 2702 240420 2758 240422
rect 2782 240420 2838 240422
rect 2862 240420 2918 240422
rect 2622 239386 2678 239388
rect 2702 239386 2758 239388
rect 2782 239386 2838 239388
rect 2862 239386 2918 239388
rect 2622 239334 2648 239386
rect 2648 239334 2678 239386
rect 2702 239334 2712 239386
rect 2712 239334 2758 239386
rect 2782 239334 2828 239386
rect 2828 239334 2838 239386
rect 2862 239334 2892 239386
rect 2892 239334 2918 239386
rect 2622 239332 2678 239334
rect 2702 239332 2758 239334
rect 2782 239332 2838 239334
rect 2862 239332 2918 239334
rect 2622 238298 2678 238300
rect 2702 238298 2758 238300
rect 2782 238298 2838 238300
rect 2862 238298 2918 238300
rect 2622 238246 2648 238298
rect 2648 238246 2678 238298
rect 2702 238246 2712 238298
rect 2712 238246 2758 238298
rect 2782 238246 2828 238298
rect 2828 238246 2838 238298
rect 2862 238246 2892 238298
rect 2892 238246 2918 238298
rect 2622 238244 2678 238246
rect 2702 238244 2758 238246
rect 2782 238244 2838 238246
rect 2862 238244 2918 238246
rect 2622 237210 2678 237212
rect 2702 237210 2758 237212
rect 2782 237210 2838 237212
rect 2862 237210 2918 237212
rect 2622 237158 2648 237210
rect 2648 237158 2678 237210
rect 2702 237158 2712 237210
rect 2712 237158 2758 237210
rect 2782 237158 2828 237210
rect 2828 237158 2838 237210
rect 2862 237158 2892 237210
rect 2892 237158 2918 237210
rect 2622 237156 2678 237158
rect 2702 237156 2758 237158
rect 2782 237156 2838 237158
rect 2862 237156 2918 237158
rect 2622 236122 2678 236124
rect 2702 236122 2758 236124
rect 2782 236122 2838 236124
rect 2862 236122 2918 236124
rect 2622 236070 2648 236122
rect 2648 236070 2678 236122
rect 2702 236070 2712 236122
rect 2712 236070 2758 236122
rect 2782 236070 2828 236122
rect 2828 236070 2838 236122
rect 2862 236070 2892 236122
rect 2892 236070 2918 236122
rect 2622 236068 2678 236070
rect 2702 236068 2758 236070
rect 2782 236068 2838 236070
rect 2862 236068 2918 236070
rect 2622 235034 2678 235036
rect 2702 235034 2758 235036
rect 2782 235034 2838 235036
rect 2862 235034 2918 235036
rect 2622 234982 2648 235034
rect 2648 234982 2678 235034
rect 2702 234982 2712 235034
rect 2712 234982 2758 235034
rect 2782 234982 2828 235034
rect 2828 234982 2838 235034
rect 2862 234982 2892 235034
rect 2892 234982 2918 235034
rect 2622 234980 2678 234982
rect 2702 234980 2758 234982
rect 2782 234980 2838 234982
rect 2862 234980 2918 234982
rect 2622 233946 2678 233948
rect 2702 233946 2758 233948
rect 2782 233946 2838 233948
rect 2862 233946 2918 233948
rect 2622 233894 2648 233946
rect 2648 233894 2678 233946
rect 2702 233894 2712 233946
rect 2712 233894 2758 233946
rect 2782 233894 2828 233946
rect 2828 233894 2838 233946
rect 2862 233894 2892 233946
rect 2892 233894 2918 233946
rect 2622 233892 2678 233894
rect 2702 233892 2758 233894
rect 2782 233892 2838 233894
rect 2862 233892 2918 233894
rect 2622 232858 2678 232860
rect 2702 232858 2758 232860
rect 2782 232858 2838 232860
rect 2862 232858 2918 232860
rect 2622 232806 2648 232858
rect 2648 232806 2678 232858
rect 2702 232806 2712 232858
rect 2712 232806 2758 232858
rect 2782 232806 2828 232858
rect 2828 232806 2838 232858
rect 2862 232806 2892 232858
rect 2892 232806 2918 232858
rect 2622 232804 2678 232806
rect 2702 232804 2758 232806
rect 2782 232804 2838 232806
rect 2862 232804 2918 232806
rect 2622 231770 2678 231772
rect 2702 231770 2758 231772
rect 2782 231770 2838 231772
rect 2862 231770 2918 231772
rect 2622 231718 2648 231770
rect 2648 231718 2678 231770
rect 2702 231718 2712 231770
rect 2712 231718 2758 231770
rect 2782 231718 2828 231770
rect 2828 231718 2838 231770
rect 2862 231718 2892 231770
rect 2892 231718 2918 231770
rect 2622 231716 2678 231718
rect 2702 231716 2758 231718
rect 2782 231716 2838 231718
rect 2862 231716 2918 231718
rect 2622 230682 2678 230684
rect 2702 230682 2758 230684
rect 2782 230682 2838 230684
rect 2862 230682 2918 230684
rect 2622 230630 2648 230682
rect 2648 230630 2678 230682
rect 2702 230630 2712 230682
rect 2712 230630 2758 230682
rect 2782 230630 2828 230682
rect 2828 230630 2838 230682
rect 2862 230630 2892 230682
rect 2892 230630 2918 230682
rect 2622 230628 2678 230630
rect 2702 230628 2758 230630
rect 2782 230628 2838 230630
rect 2862 230628 2918 230630
rect 2622 229594 2678 229596
rect 2702 229594 2758 229596
rect 2782 229594 2838 229596
rect 2862 229594 2918 229596
rect 2622 229542 2648 229594
rect 2648 229542 2678 229594
rect 2702 229542 2712 229594
rect 2712 229542 2758 229594
rect 2782 229542 2828 229594
rect 2828 229542 2838 229594
rect 2862 229542 2892 229594
rect 2892 229542 2918 229594
rect 2622 229540 2678 229542
rect 2702 229540 2758 229542
rect 2782 229540 2838 229542
rect 2862 229540 2918 229542
rect 2622 228506 2678 228508
rect 2702 228506 2758 228508
rect 2782 228506 2838 228508
rect 2862 228506 2918 228508
rect 2622 228454 2648 228506
rect 2648 228454 2678 228506
rect 2702 228454 2712 228506
rect 2712 228454 2758 228506
rect 2782 228454 2828 228506
rect 2828 228454 2838 228506
rect 2862 228454 2892 228506
rect 2892 228454 2918 228506
rect 2622 228452 2678 228454
rect 2702 228452 2758 228454
rect 2782 228452 2838 228454
rect 2862 228452 2918 228454
rect 2622 227418 2678 227420
rect 2702 227418 2758 227420
rect 2782 227418 2838 227420
rect 2862 227418 2918 227420
rect 2622 227366 2648 227418
rect 2648 227366 2678 227418
rect 2702 227366 2712 227418
rect 2712 227366 2758 227418
rect 2782 227366 2828 227418
rect 2828 227366 2838 227418
rect 2862 227366 2892 227418
rect 2892 227366 2918 227418
rect 2622 227364 2678 227366
rect 2702 227364 2758 227366
rect 2782 227364 2838 227366
rect 2862 227364 2918 227366
rect 2622 226330 2678 226332
rect 2702 226330 2758 226332
rect 2782 226330 2838 226332
rect 2862 226330 2918 226332
rect 2622 226278 2648 226330
rect 2648 226278 2678 226330
rect 2702 226278 2712 226330
rect 2712 226278 2758 226330
rect 2782 226278 2828 226330
rect 2828 226278 2838 226330
rect 2862 226278 2892 226330
rect 2892 226278 2918 226330
rect 2622 226276 2678 226278
rect 2702 226276 2758 226278
rect 2782 226276 2838 226278
rect 2862 226276 2918 226278
rect 2622 225242 2678 225244
rect 2702 225242 2758 225244
rect 2782 225242 2838 225244
rect 2862 225242 2918 225244
rect 2622 225190 2648 225242
rect 2648 225190 2678 225242
rect 2702 225190 2712 225242
rect 2712 225190 2758 225242
rect 2782 225190 2828 225242
rect 2828 225190 2838 225242
rect 2862 225190 2892 225242
rect 2892 225190 2918 225242
rect 2622 225188 2678 225190
rect 2702 225188 2758 225190
rect 2782 225188 2838 225190
rect 2862 225188 2918 225190
rect 2622 224154 2678 224156
rect 2702 224154 2758 224156
rect 2782 224154 2838 224156
rect 2862 224154 2918 224156
rect 2622 224102 2648 224154
rect 2648 224102 2678 224154
rect 2702 224102 2712 224154
rect 2712 224102 2758 224154
rect 2782 224102 2828 224154
rect 2828 224102 2838 224154
rect 2862 224102 2892 224154
rect 2892 224102 2918 224154
rect 2622 224100 2678 224102
rect 2702 224100 2758 224102
rect 2782 224100 2838 224102
rect 2862 224100 2918 224102
rect 2622 223066 2678 223068
rect 2702 223066 2758 223068
rect 2782 223066 2838 223068
rect 2862 223066 2918 223068
rect 2622 223014 2648 223066
rect 2648 223014 2678 223066
rect 2702 223014 2712 223066
rect 2712 223014 2758 223066
rect 2782 223014 2828 223066
rect 2828 223014 2838 223066
rect 2862 223014 2892 223066
rect 2892 223014 2918 223066
rect 2622 223012 2678 223014
rect 2702 223012 2758 223014
rect 2782 223012 2838 223014
rect 2862 223012 2918 223014
rect 2622 221978 2678 221980
rect 2702 221978 2758 221980
rect 2782 221978 2838 221980
rect 2862 221978 2918 221980
rect 2622 221926 2648 221978
rect 2648 221926 2678 221978
rect 2702 221926 2712 221978
rect 2712 221926 2758 221978
rect 2782 221926 2828 221978
rect 2828 221926 2838 221978
rect 2862 221926 2892 221978
rect 2892 221926 2918 221978
rect 2622 221924 2678 221926
rect 2702 221924 2758 221926
rect 2782 221924 2838 221926
rect 2862 221924 2918 221926
rect 110 213968 166 214024
rect 18 118768 74 118824
rect 110 71168 166 71224
rect 2622 220890 2678 220892
rect 2702 220890 2758 220892
rect 2782 220890 2838 220892
rect 2862 220890 2918 220892
rect 2622 220838 2648 220890
rect 2648 220838 2678 220890
rect 2702 220838 2712 220890
rect 2712 220838 2758 220890
rect 2782 220838 2828 220890
rect 2828 220838 2838 220890
rect 2862 220838 2892 220890
rect 2892 220838 2918 220890
rect 2622 220836 2678 220838
rect 2702 220836 2758 220838
rect 2782 220836 2838 220838
rect 2862 220836 2918 220838
rect 2622 219802 2678 219804
rect 2702 219802 2758 219804
rect 2782 219802 2838 219804
rect 2862 219802 2918 219804
rect 2622 219750 2648 219802
rect 2648 219750 2678 219802
rect 2702 219750 2712 219802
rect 2712 219750 2758 219802
rect 2782 219750 2828 219802
rect 2828 219750 2838 219802
rect 2862 219750 2892 219802
rect 2892 219750 2918 219802
rect 2622 219748 2678 219750
rect 2702 219748 2758 219750
rect 2782 219748 2838 219750
rect 2862 219748 2918 219750
rect 2622 218714 2678 218716
rect 2702 218714 2758 218716
rect 2782 218714 2838 218716
rect 2862 218714 2918 218716
rect 2622 218662 2648 218714
rect 2648 218662 2678 218714
rect 2702 218662 2712 218714
rect 2712 218662 2758 218714
rect 2782 218662 2828 218714
rect 2828 218662 2838 218714
rect 2862 218662 2892 218714
rect 2892 218662 2918 218714
rect 2622 218660 2678 218662
rect 2702 218660 2758 218662
rect 2782 218660 2838 218662
rect 2862 218660 2918 218662
rect 2622 217626 2678 217628
rect 2702 217626 2758 217628
rect 2782 217626 2838 217628
rect 2862 217626 2918 217628
rect 2622 217574 2648 217626
rect 2648 217574 2678 217626
rect 2702 217574 2712 217626
rect 2712 217574 2758 217626
rect 2782 217574 2828 217626
rect 2828 217574 2838 217626
rect 2862 217574 2892 217626
rect 2892 217574 2918 217626
rect 2622 217572 2678 217574
rect 2702 217572 2758 217574
rect 2782 217572 2838 217574
rect 2862 217572 2918 217574
rect 2622 216538 2678 216540
rect 2702 216538 2758 216540
rect 2782 216538 2838 216540
rect 2862 216538 2918 216540
rect 2622 216486 2648 216538
rect 2648 216486 2678 216538
rect 2702 216486 2712 216538
rect 2712 216486 2758 216538
rect 2782 216486 2828 216538
rect 2828 216486 2838 216538
rect 2862 216486 2892 216538
rect 2892 216486 2918 216538
rect 2622 216484 2678 216486
rect 2702 216484 2758 216486
rect 2782 216484 2838 216486
rect 2862 216484 2918 216486
rect 2622 215450 2678 215452
rect 2702 215450 2758 215452
rect 2782 215450 2838 215452
rect 2862 215450 2918 215452
rect 2622 215398 2648 215450
rect 2648 215398 2678 215450
rect 2702 215398 2712 215450
rect 2712 215398 2758 215450
rect 2782 215398 2828 215450
rect 2828 215398 2838 215450
rect 2862 215398 2892 215450
rect 2892 215398 2918 215450
rect 2622 215396 2678 215398
rect 2702 215396 2758 215398
rect 2782 215396 2838 215398
rect 2862 215396 2918 215398
rect 2622 214362 2678 214364
rect 2702 214362 2758 214364
rect 2782 214362 2838 214364
rect 2862 214362 2918 214364
rect 2622 214310 2648 214362
rect 2648 214310 2678 214362
rect 2702 214310 2712 214362
rect 2712 214310 2758 214362
rect 2782 214310 2828 214362
rect 2828 214310 2838 214362
rect 2862 214310 2892 214362
rect 2892 214310 2918 214362
rect 2622 214308 2678 214310
rect 2702 214308 2758 214310
rect 2782 214308 2838 214310
rect 2862 214308 2918 214310
rect 2622 213274 2678 213276
rect 2702 213274 2758 213276
rect 2782 213274 2838 213276
rect 2862 213274 2918 213276
rect 2622 213222 2648 213274
rect 2648 213222 2678 213274
rect 2702 213222 2712 213274
rect 2712 213222 2758 213274
rect 2782 213222 2828 213274
rect 2828 213222 2838 213274
rect 2862 213222 2892 213274
rect 2892 213222 2918 213274
rect 2622 213220 2678 213222
rect 2702 213220 2758 213222
rect 2782 213220 2838 213222
rect 2862 213220 2918 213222
rect 2622 212186 2678 212188
rect 2702 212186 2758 212188
rect 2782 212186 2838 212188
rect 2862 212186 2918 212188
rect 2622 212134 2648 212186
rect 2648 212134 2678 212186
rect 2702 212134 2712 212186
rect 2712 212134 2758 212186
rect 2782 212134 2828 212186
rect 2828 212134 2838 212186
rect 2862 212134 2892 212186
rect 2892 212134 2918 212186
rect 2622 212132 2678 212134
rect 2702 212132 2758 212134
rect 2782 212132 2838 212134
rect 2862 212132 2918 212134
rect 2622 211098 2678 211100
rect 2702 211098 2758 211100
rect 2782 211098 2838 211100
rect 2862 211098 2918 211100
rect 2622 211046 2648 211098
rect 2648 211046 2678 211098
rect 2702 211046 2712 211098
rect 2712 211046 2758 211098
rect 2782 211046 2828 211098
rect 2828 211046 2838 211098
rect 2862 211046 2892 211098
rect 2892 211046 2918 211098
rect 2622 211044 2678 211046
rect 2702 211044 2758 211046
rect 2782 211044 2838 211046
rect 2862 211044 2918 211046
rect 2622 210010 2678 210012
rect 2702 210010 2758 210012
rect 2782 210010 2838 210012
rect 2862 210010 2918 210012
rect 2622 209958 2648 210010
rect 2648 209958 2678 210010
rect 2702 209958 2712 210010
rect 2712 209958 2758 210010
rect 2782 209958 2828 210010
rect 2828 209958 2838 210010
rect 2862 209958 2892 210010
rect 2892 209958 2918 210010
rect 2622 209956 2678 209958
rect 2702 209956 2758 209958
rect 2782 209956 2838 209958
rect 2862 209956 2918 209958
rect 2622 208922 2678 208924
rect 2702 208922 2758 208924
rect 2782 208922 2838 208924
rect 2862 208922 2918 208924
rect 2622 208870 2648 208922
rect 2648 208870 2678 208922
rect 2702 208870 2712 208922
rect 2712 208870 2758 208922
rect 2782 208870 2828 208922
rect 2828 208870 2838 208922
rect 2862 208870 2892 208922
rect 2892 208870 2918 208922
rect 2622 208868 2678 208870
rect 2702 208868 2758 208870
rect 2782 208868 2838 208870
rect 2862 208868 2918 208870
rect 2622 207834 2678 207836
rect 2702 207834 2758 207836
rect 2782 207834 2838 207836
rect 2862 207834 2918 207836
rect 2622 207782 2648 207834
rect 2648 207782 2678 207834
rect 2702 207782 2712 207834
rect 2712 207782 2758 207834
rect 2782 207782 2828 207834
rect 2828 207782 2838 207834
rect 2862 207782 2892 207834
rect 2892 207782 2918 207834
rect 2622 207780 2678 207782
rect 2702 207780 2758 207782
rect 2782 207780 2838 207782
rect 2862 207780 2918 207782
rect 2622 206746 2678 206748
rect 2702 206746 2758 206748
rect 2782 206746 2838 206748
rect 2862 206746 2918 206748
rect 2622 206694 2648 206746
rect 2648 206694 2678 206746
rect 2702 206694 2712 206746
rect 2712 206694 2758 206746
rect 2782 206694 2828 206746
rect 2828 206694 2838 206746
rect 2862 206694 2892 206746
rect 2892 206694 2918 206746
rect 2622 206692 2678 206694
rect 2702 206692 2758 206694
rect 2782 206692 2838 206694
rect 2862 206692 2918 206694
rect 2622 205658 2678 205660
rect 2702 205658 2758 205660
rect 2782 205658 2838 205660
rect 2862 205658 2918 205660
rect 2622 205606 2648 205658
rect 2648 205606 2678 205658
rect 2702 205606 2712 205658
rect 2712 205606 2758 205658
rect 2782 205606 2828 205658
rect 2828 205606 2838 205658
rect 2862 205606 2892 205658
rect 2892 205606 2918 205658
rect 2622 205604 2678 205606
rect 2702 205604 2758 205606
rect 2782 205604 2838 205606
rect 2862 205604 2918 205606
rect 2622 204570 2678 204572
rect 2702 204570 2758 204572
rect 2782 204570 2838 204572
rect 2862 204570 2918 204572
rect 2622 204518 2648 204570
rect 2648 204518 2678 204570
rect 2702 204518 2712 204570
rect 2712 204518 2758 204570
rect 2782 204518 2828 204570
rect 2828 204518 2838 204570
rect 2862 204518 2892 204570
rect 2892 204518 2918 204570
rect 2622 204516 2678 204518
rect 2702 204516 2758 204518
rect 2782 204516 2838 204518
rect 2862 204516 2918 204518
rect 2622 203482 2678 203484
rect 2702 203482 2758 203484
rect 2782 203482 2838 203484
rect 2862 203482 2918 203484
rect 2622 203430 2648 203482
rect 2648 203430 2678 203482
rect 2702 203430 2712 203482
rect 2712 203430 2758 203482
rect 2782 203430 2828 203482
rect 2828 203430 2838 203482
rect 2862 203430 2892 203482
rect 2892 203430 2918 203482
rect 2622 203428 2678 203430
rect 2702 203428 2758 203430
rect 2782 203428 2838 203430
rect 2862 203428 2918 203430
rect 2622 202394 2678 202396
rect 2702 202394 2758 202396
rect 2782 202394 2838 202396
rect 2862 202394 2918 202396
rect 2622 202342 2648 202394
rect 2648 202342 2678 202394
rect 2702 202342 2712 202394
rect 2712 202342 2758 202394
rect 2782 202342 2828 202394
rect 2828 202342 2838 202394
rect 2862 202342 2892 202394
rect 2892 202342 2918 202394
rect 2622 202340 2678 202342
rect 2702 202340 2758 202342
rect 2782 202340 2838 202342
rect 2862 202340 2918 202342
rect 2622 201306 2678 201308
rect 2702 201306 2758 201308
rect 2782 201306 2838 201308
rect 2862 201306 2918 201308
rect 2622 201254 2648 201306
rect 2648 201254 2678 201306
rect 2702 201254 2712 201306
rect 2712 201254 2758 201306
rect 2782 201254 2828 201306
rect 2828 201254 2838 201306
rect 2862 201254 2892 201306
rect 2892 201254 2918 201306
rect 2622 201252 2678 201254
rect 2702 201252 2758 201254
rect 2782 201252 2838 201254
rect 2862 201252 2918 201254
rect 2622 200218 2678 200220
rect 2702 200218 2758 200220
rect 2782 200218 2838 200220
rect 2862 200218 2918 200220
rect 2622 200166 2648 200218
rect 2648 200166 2678 200218
rect 2702 200166 2712 200218
rect 2712 200166 2758 200218
rect 2782 200166 2828 200218
rect 2828 200166 2838 200218
rect 2862 200166 2892 200218
rect 2892 200166 2918 200218
rect 2622 200164 2678 200166
rect 2702 200164 2758 200166
rect 2782 200164 2838 200166
rect 2862 200164 2918 200166
rect 2622 199130 2678 199132
rect 2702 199130 2758 199132
rect 2782 199130 2838 199132
rect 2862 199130 2918 199132
rect 2622 199078 2648 199130
rect 2648 199078 2678 199130
rect 2702 199078 2712 199130
rect 2712 199078 2758 199130
rect 2782 199078 2828 199130
rect 2828 199078 2838 199130
rect 2862 199078 2892 199130
rect 2892 199078 2918 199130
rect 2622 199076 2678 199078
rect 2702 199076 2758 199078
rect 2782 199076 2838 199078
rect 2862 199076 2918 199078
rect 2622 198042 2678 198044
rect 2702 198042 2758 198044
rect 2782 198042 2838 198044
rect 2862 198042 2918 198044
rect 2622 197990 2648 198042
rect 2648 197990 2678 198042
rect 2702 197990 2712 198042
rect 2712 197990 2758 198042
rect 2782 197990 2828 198042
rect 2828 197990 2838 198042
rect 2862 197990 2892 198042
rect 2892 197990 2918 198042
rect 2622 197988 2678 197990
rect 2702 197988 2758 197990
rect 2782 197988 2838 197990
rect 2862 197988 2918 197990
rect 2622 196954 2678 196956
rect 2702 196954 2758 196956
rect 2782 196954 2838 196956
rect 2862 196954 2918 196956
rect 2622 196902 2648 196954
rect 2648 196902 2678 196954
rect 2702 196902 2712 196954
rect 2712 196902 2758 196954
rect 2782 196902 2828 196954
rect 2828 196902 2838 196954
rect 2862 196902 2892 196954
rect 2892 196902 2918 196954
rect 2622 196900 2678 196902
rect 2702 196900 2758 196902
rect 2782 196900 2838 196902
rect 2862 196900 2918 196902
rect 2622 195866 2678 195868
rect 2702 195866 2758 195868
rect 2782 195866 2838 195868
rect 2862 195866 2918 195868
rect 2622 195814 2648 195866
rect 2648 195814 2678 195866
rect 2702 195814 2712 195866
rect 2712 195814 2758 195866
rect 2782 195814 2828 195866
rect 2828 195814 2838 195866
rect 2862 195814 2892 195866
rect 2892 195814 2918 195866
rect 2622 195812 2678 195814
rect 2702 195812 2758 195814
rect 2782 195812 2838 195814
rect 2862 195812 2918 195814
rect 2622 194778 2678 194780
rect 2702 194778 2758 194780
rect 2782 194778 2838 194780
rect 2862 194778 2918 194780
rect 2622 194726 2648 194778
rect 2648 194726 2678 194778
rect 2702 194726 2712 194778
rect 2712 194726 2758 194778
rect 2782 194726 2828 194778
rect 2828 194726 2838 194778
rect 2862 194726 2892 194778
rect 2892 194726 2918 194778
rect 2622 194724 2678 194726
rect 2702 194724 2758 194726
rect 2782 194724 2838 194726
rect 2862 194724 2918 194726
rect 2622 193690 2678 193692
rect 2702 193690 2758 193692
rect 2782 193690 2838 193692
rect 2862 193690 2918 193692
rect 2622 193638 2648 193690
rect 2648 193638 2678 193690
rect 2702 193638 2712 193690
rect 2712 193638 2758 193690
rect 2782 193638 2828 193690
rect 2828 193638 2838 193690
rect 2862 193638 2892 193690
rect 2892 193638 2918 193690
rect 2622 193636 2678 193638
rect 2702 193636 2758 193638
rect 2782 193636 2838 193638
rect 2862 193636 2918 193638
rect 2622 192602 2678 192604
rect 2702 192602 2758 192604
rect 2782 192602 2838 192604
rect 2862 192602 2918 192604
rect 2622 192550 2648 192602
rect 2648 192550 2678 192602
rect 2702 192550 2712 192602
rect 2712 192550 2758 192602
rect 2782 192550 2828 192602
rect 2828 192550 2838 192602
rect 2862 192550 2892 192602
rect 2892 192550 2918 192602
rect 2622 192548 2678 192550
rect 2702 192548 2758 192550
rect 2782 192548 2838 192550
rect 2862 192548 2918 192550
rect 2622 191514 2678 191516
rect 2702 191514 2758 191516
rect 2782 191514 2838 191516
rect 2862 191514 2918 191516
rect 2622 191462 2648 191514
rect 2648 191462 2678 191514
rect 2702 191462 2712 191514
rect 2712 191462 2758 191514
rect 2782 191462 2828 191514
rect 2828 191462 2838 191514
rect 2862 191462 2892 191514
rect 2892 191462 2918 191514
rect 2622 191460 2678 191462
rect 2702 191460 2758 191462
rect 2782 191460 2838 191462
rect 2862 191460 2918 191462
rect 2622 190426 2678 190428
rect 2702 190426 2758 190428
rect 2782 190426 2838 190428
rect 2862 190426 2918 190428
rect 2622 190374 2648 190426
rect 2648 190374 2678 190426
rect 2702 190374 2712 190426
rect 2712 190374 2758 190426
rect 2782 190374 2828 190426
rect 2828 190374 2838 190426
rect 2862 190374 2892 190426
rect 2892 190374 2918 190426
rect 2622 190372 2678 190374
rect 2702 190372 2758 190374
rect 2782 190372 2838 190374
rect 2862 190372 2918 190374
rect 2622 189338 2678 189340
rect 2702 189338 2758 189340
rect 2782 189338 2838 189340
rect 2862 189338 2918 189340
rect 2622 189286 2648 189338
rect 2648 189286 2678 189338
rect 2702 189286 2712 189338
rect 2712 189286 2758 189338
rect 2782 189286 2828 189338
rect 2828 189286 2838 189338
rect 2862 189286 2892 189338
rect 2892 189286 2918 189338
rect 2622 189284 2678 189286
rect 2702 189284 2758 189286
rect 2782 189284 2838 189286
rect 2862 189284 2918 189286
rect 2622 188250 2678 188252
rect 2702 188250 2758 188252
rect 2782 188250 2838 188252
rect 2862 188250 2918 188252
rect 2622 188198 2648 188250
rect 2648 188198 2678 188250
rect 2702 188198 2712 188250
rect 2712 188198 2758 188250
rect 2782 188198 2828 188250
rect 2828 188198 2838 188250
rect 2862 188198 2892 188250
rect 2892 188198 2918 188250
rect 2622 188196 2678 188198
rect 2702 188196 2758 188198
rect 2782 188196 2838 188198
rect 2862 188196 2918 188198
rect 2622 187162 2678 187164
rect 2702 187162 2758 187164
rect 2782 187162 2838 187164
rect 2862 187162 2918 187164
rect 2622 187110 2648 187162
rect 2648 187110 2678 187162
rect 2702 187110 2712 187162
rect 2712 187110 2758 187162
rect 2782 187110 2828 187162
rect 2828 187110 2838 187162
rect 2862 187110 2892 187162
rect 2892 187110 2918 187162
rect 2622 187108 2678 187110
rect 2702 187108 2758 187110
rect 2782 187108 2838 187110
rect 2862 187108 2918 187110
rect 2622 186074 2678 186076
rect 2702 186074 2758 186076
rect 2782 186074 2838 186076
rect 2862 186074 2918 186076
rect 2622 186022 2648 186074
rect 2648 186022 2678 186074
rect 2702 186022 2712 186074
rect 2712 186022 2758 186074
rect 2782 186022 2828 186074
rect 2828 186022 2838 186074
rect 2862 186022 2892 186074
rect 2892 186022 2918 186074
rect 2622 186020 2678 186022
rect 2702 186020 2758 186022
rect 2782 186020 2838 186022
rect 2862 186020 2918 186022
rect 2622 184986 2678 184988
rect 2702 184986 2758 184988
rect 2782 184986 2838 184988
rect 2862 184986 2918 184988
rect 2622 184934 2648 184986
rect 2648 184934 2678 184986
rect 2702 184934 2712 184986
rect 2712 184934 2758 184986
rect 2782 184934 2828 184986
rect 2828 184934 2838 184986
rect 2862 184934 2892 184986
rect 2892 184934 2918 184986
rect 2622 184932 2678 184934
rect 2702 184932 2758 184934
rect 2782 184932 2838 184934
rect 2862 184932 2918 184934
rect 2622 183898 2678 183900
rect 2702 183898 2758 183900
rect 2782 183898 2838 183900
rect 2862 183898 2918 183900
rect 2622 183846 2648 183898
rect 2648 183846 2678 183898
rect 2702 183846 2712 183898
rect 2712 183846 2758 183898
rect 2782 183846 2828 183898
rect 2828 183846 2838 183898
rect 2862 183846 2892 183898
rect 2892 183846 2918 183898
rect 2622 183844 2678 183846
rect 2702 183844 2758 183846
rect 2782 183844 2838 183846
rect 2862 183844 2918 183846
rect 2622 182810 2678 182812
rect 2702 182810 2758 182812
rect 2782 182810 2838 182812
rect 2862 182810 2918 182812
rect 2622 182758 2648 182810
rect 2648 182758 2678 182810
rect 2702 182758 2712 182810
rect 2712 182758 2758 182810
rect 2782 182758 2828 182810
rect 2828 182758 2838 182810
rect 2862 182758 2892 182810
rect 2892 182758 2918 182810
rect 2622 182756 2678 182758
rect 2702 182756 2758 182758
rect 2782 182756 2838 182758
rect 2862 182756 2918 182758
rect 2622 181722 2678 181724
rect 2702 181722 2758 181724
rect 2782 181722 2838 181724
rect 2862 181722 2918 181724
rect 2622 181670 2648 181722
rect 2648 181670 2678 181722
rect 2702 181670 2712 181722
rect 2712 181670 2758 181722
rect 2782 181670 2828 181722
rect 2828 181670 2838 181722
rect 2862 181670 2892 181722
rect 2892 181670 2918 181722
rect 2622 181668 2678 181670
rect 2702 181668 2758 181670
rect 2782 181668 2838 181670
rect 2862 181668 2918 181670
rect 2622 180634 2678 180636
rect 2702 180634 2758 180636
rect 2782 180634 2838 180636
rect 2862 180634 2918 180636
rect 2622 180582 2648 180634
rect 2648 180582 2678 180634
rect 2702 180582 2712 180634
rect 2712 180582 2758 180634
rect 2782 180582 2828 180634
rect 2828 180582 2838 180634
rect 2862 180582 2892 180634
rect 2892 180582 2918 180634
rect 2622 180580 2678 180582
rect 2702 180580 2758 180582
rect 2782 180580 2838 180582
rect 2862 180580 2918 180582
rect 2622 179546 2678 179548
rect 2702 179546 2758 179548
rect 2782 179546 2838 179548
rect 2862 179546 2918 179548
rect 2622 179494 2648 179546
rect 2648 179494 2678 179546
rect 2702 179494 2712 179546
rect 2712 179494 2758 179546
rect 2782 179494 2828 179546
rect 2828 179494 2838 179546
rect 2862 179494 2892 179546
rect 2892 179494 2918 179546
rect 2622 179492 2678 179494
rect 2702 179492 2758 179494
rect 2782 179492 2838 179494
rect 2862 179492 2918 179494
rect 2622 178458 2678 178460
rect 2702 178458 2758 178460
rect 2782 178458 2838 178460
rect 2862 178458 2918 178460
rect 2622 178406 2648 178458
rect 2648 178406 2678 178458
rect 2702 178406 2712 178458
rect 2712 178406 2758 178458
rect 2782 178406 2828 178458
rect 2828 178406 2838 178458
rect 2862 178406 2892 178458
rect 2892 178406 2918 178458
rect 2622 178404 2678 178406
rect 2702 178404 2758 178406
rect 2782 178404 2838 178406
rect 2862 178404 2918 178406
rect 2622 177370 2678 177372
rect 2702 177370 2758 177372
rect 2782 177370 2838 177372
rect 2862 177370 2918 177372
rect 2622 177318 2648 177370
rect 2648 177318 2678 177370
rect 2702 177318 2712 177370
rect 2712 177318 2758 177370
rect 2782 177318 2828 177370
rect 2828 177318 2838 177370
rect 2862 177318 2892 177370
rect 2892 177318 2918 177370
rect 2622 177316 2678 177318
rect 2702 177316 2758 177318
rect 2782 177316 2838 177318
rect 2862 177316 2918 177318
rect 2622 176282 2678 176284
rect 2702 176282 2758 176284
rect 2782 176282 2838 176284
rect 2862 176282 2918 176284
rect 2622 176230 2648 176282
rect 2648 176230 2678 176282
rect 2702 176230 2712 176282
rect 2712 176230 2758 176282
rect 2782 176230 2828 176282
rect 2828 176230 2838 176282
rect 2862 176230 2892 176282
rect 2892 176230 2918 176282
rect 2622 176228 2678 176230
rect 2702 176228 2758 176230
rect 2782 176228 2838 176230
rect 2862 176228 2918 176230
rect 2622 175194 2678 175196
rect 2702 175194 2758 175196
rect 2782 175194 2838 175196
rect 2862 175194 2918 175196
rect 2622 175142 2648 175194
rect 2648 175142 2678 175194
rect 2702 175142 2712 175194
rect 2712 175142 2758 175194
rect 2782 175142 2828 175194
rect 2828 175142 2838 175194
rect 2862 175142 2892 175194
rect 2892 175142 2918 175194
rect 2622 175140 2678 175142
rect 2702 175140 2758 175142
rect 2782 175140 2838 175142
rect 2862 175140 2918 175142
rect 2622 174106 2678 174108
rect 2702 174106 2758 174108
rect 2782 174106 2838 174108
rect 2862 174106 2918 174108
rect 2622 174054 2648 174106
rect 2648 174054 2678 174106
rect 2702 174054 2712 174106
rect 2712 174054 2758 174106
rect 2782 174054 2828 174106
rect 2828 174054 2838 174106
rect 2862 174054 2892 174106
rect 2892 174054 2918 174106
rect 2622 174052 2678 174054
rect 2702 174052 2758 174054
rect 2782 174052 2838 174054
rect 2862 174052 2918 174054
rect 2622 173018 2678 173020
rect 2702 173018 2758 173020
rect 2782 173018 2838 173020
rect 2862 173018 2918 173020
rect 2622 172966 2648 173018
rect 2648 172966 2678 173018
rect 2702 172966 2712 173018
rect 2712 172966 2758 173018
rect 2782 172966 2828 173018
rect 2828 172966 2838 173018
rect 2862 172966 2892 173018
rect 2892 172966 2918 173018
rect 2622 172964 2678 172966
rect 2702 172964 2758 172966
rect 2782 172964 2838 172966
rect 2862 172964 2918 172966
rect 2622 171930 2678 171932
rect 2702 171930 2758 171932
rect 2782 171930 2838 171932
rect 2862 171930 2918 171932
rect 2622 171878 2648 171930
rect 2648 171878 2678 171930
rect 2702 171878 2712 171930
rect 2712 171878 2758 171930
rect 2782 171878 2828 171930
rect 2828 171878 2838 171930
rect 2862 171878 2892 171930
rect 2892 171878 2918 171930
rect 2622 171876 2678 171878
rect 2702 171876 2758 171878
rect 2782 171876 2838 171878
rect 2862 171876 2918 171878
rect 2622 170842 2678 170844
rect 2702 170842 2758 170844
rect 2782 170842 2838 170844
rect 2862 170842 2918 170844
rect 2622 170790 2648 170842
rect 2648 170790 2678 170842
rect 2702 170790 2712 170842
rect 2712 170790 2758 170842
rect 2782 170790 2828 170842
rect 2828 170790 2838 170842
rect 2862 170790 2892 170842
rect 2892 170790 2918 170842
rect 2622 170788 2678 170790
rect 2702 170788 2758 170790
rect 2782 170788 2838 170790
rect 2862 170788 2918 170790
rect 2622 169754 2678 169756
rect 2702 169754 2758 169756
rect 2782 169754 2838 169756
rect 2862 169754 2918 169756
rect 2622 169702 2648 169754
rect 2648 169702 2678 169754
rect 2702 169702 2712 169754
rect 2712 169702 2758 169754
rect 2782 169702 2828 169754
rect 2828 169702 2838 169754
rect 2862 169702 2892 169754
rect 2892 169702 2918 169754
rect 2622 169700 2678 169702
rect 2702 169700 2758 169702
rect 2782 169700 2838 169702
rect 2862 169700 2918 169702
rect 2622 168666 2678 168668
rect 2702 168666 2758 168668
rect 2782 168666 2838 168668
rect 2862 168666 2918 168668
rect 2622 168614 2648 168666
rect 2648 168614 2678 168666
rect 2702 168614 2712 168666
rect 2712 168614 2758 168666
rect 2782 168614 2828 168666
rect 2828 168614 2838 168666
rect 2862 168614 2892 168666
rect 2892 168614 2918 168666
rect 2622 168612 2678 168614
rect 2702 168612 2758 168614
rect 2782 168612 2838 168614
rect 2862 168612 2918 168614
rect 2622 167578 2678 167580
rect 2702 167578 2758 167580
rect 2782 167578 2838 167580
rect 2862 167578 2918 167580
rect 2622 167526 2648 167578
rect 2648 167526 2678 167578
rect 2702 167526 2712 167578
rect 2712 167526 2758 167578
rect 2782 167526 2828 167578
rect 2828 167526 2838 167578
rect 2862 167526 2892 167578
rect 2892 167526 2918 167578
rect 2622 167524 2678 167526
rect 2702 167524 2758 167526
rect 2782 167524 2838 167526
rect 2862 167524 2918 167526
rect 2622 166490 2678 166492
rect 2702 166490 2758 166492
rect 2782 166490 2838 166492
rect 2862 166490 2918 166492
rect 2622 166438 2648 166490
rect 2648 166438 2678 166490
rect 2702 166438 2712 166490
rect 2712 166438 2758 166490
rect 2782 166438 2828 166490
rect 2828 166438 2838 166490
rect 2862 166438 2892 166490
rect 2892 166438 2918 166490
rect 2622 166436 2678 166438
rect 2702 166436 2758 166438
rect 2782 166436 2838 166438
rect 2862 166436 2918 166438
rect 2622 165402 2678 165404
rect 2702 165402 2758 165404
rect 2782 165402 2838 165404
rect 2862 165402 2918 165404
rect 2622 165350 2648 165402
rect 2648 165350 2678 165402
rect 2702 165350 2712 165402
rect 2712 165350 2758 165402
rect 2782 165350 2828 165402
rect 2828 165350 2838 165402
rect 2862 165350 2892 165402
rect 2892 165350 2918 165402
rect 2622 165348 2678 165350
rect 2702 165348 2758 165350
rect 2782 165348 2838 165350
rect 2862 165348 2918 165350
rect 2622 164314 2678 164316
rect 2702 164314 2758 164316
rect 2782 164314 2838 164316
rect 2862 164314 2918 164316
rect 2622 164262 2648 164314
rect 2648 164262 2678 164314
rect 2702 164262 2712 164314
rect 2712 164262 2758 164314
rect 2782 164262 2828 164314
rect 2828 164262 2838 164314
rect 2862 164262 2892 164314
rect 2892 164262 2918 164314
rect 2622 164260 2678 164262
rect 2702 164260 2758 164262
rect 2782 164260 2838 164262
rect 2862 164260 2918 164262
rect 2622 163226 2678 163228
rect 2702 163226 2758 163228
rect 2782 163226 2838 163228
rect 2862 163226 2918 163228
rect 2622 163174 2648 163226
rect 2648 163174 2678 163226
rect 2702 163174 2712 163226
rect 2712 163174 2758 163226
rect 2782 163174 2828 163226
rect 2828 163174 2838 163226
rect 2862 163174 2892 163226
rect 2892 163174 2918 163226
rect 2622 163172 2678 163174
rect 2702 163172 2758 163174
rect 2782 163172 2838 163174
rect 2862 163172 2918 163174
rect 2622 162138 2678 162140
rect 2702 162138 2758 162140
rect 2782 162138 2838 162140
rect 2862 162138 2918 162140
rect 2622 162086 2648 162138
rect 2648 162086 2678 162138
rect 2702 162086 2712 162138
rect 2712 162086 2758 162138
rect 2782 162086 2828 162138
rect 2828 162086 2838 162138
rect 2862 162086 2892 162138
rect 2892 162086 2918 162138
rect 2622 162084 2678 162086
rect 2702 162084 2758 162086
rect 2782 162084 2838 162086
rect 2862 162084 2918 162086
rect 2622 161050 2678 161052
rect 2702 161050 2758 161052
rect 2782 161050 2838 161052
rect 2862 161050 2918 161052
rect 2622 160998 2648 161050
rect 2648 160998 2678 161050
rect 2702 160998 2712 161050
rect 2712 160998 2758 161050
rect 2782 160998 2828 161050
rect 2828 160998 2838 161050
rect 2862 160998 2892 161050
rect 2892 160998 2918 161050
rect 2622 160996 2678 160998
rect 2702 160996 2758 160998
rect 2782 160996 2838 160998
rect 2862 160996 2918 160998
rect 2622 159962 2678 159964
rect 2702 159962 2758 159964
rect 2782 159962 2838 159964
rect 2862 159962 2918 159964
rect 2622 159910 2648 159962
rect 2648 159910 2678 159962
rect 2702 159910 2712 159962
rect 2712 159910 2758 159962
rect 2782 159910 2828 159962
rect 2828 159910 2838 159962
rect 2862 159910 2892 159962
rect 2892 159910 2918 159962
rect 2622 159908 2678 159910
rect 2702 159908 2758 159910
rect 2782 159908 2838 159910
rect 2862 159908 2918 159910
rect 2622 158874 2678 158876
rect 2702 158874 2758 158876
rect 2782 158874 2838 158876
rect 2862 158874 2918 158876
rect 2622 158822 2648 158874
rect 2648 158822 2678 158874
rect 2702 158822 2712 158874
rect 2712 158822 2758 158874
rect 2782 158822 2828 158874
rect 2828 158822 2838 158874
rect 2862 158822 2892 158874
rect 2892 158822 2918 158874
rect 2622 158820 2678 158822
rect 2702 158820 2758 158822
rect 2782 158820 2838 158822
rect 2862 158820 2918 158822
rect 2622 157786 2678 157788
rect 2702 157786 2758 157788
rect 2782 157786 2838 157788
rect 2862 157786 2918 157788
rect 2622 157734 2648 157786
rect 2648 157734 2678 157786
rect 2702 157734 2712 157786
rect 2712 157734 2758 157786
rect 2782 157734 2828 157786
rect 2828 157734 2838 157786
rect 2862 157734 2892 157786
rect 2892 157734 2918 157786
rect 2622 157732 2678 157734
rect 2702 157732 2758 157734
rect 2782 157732 2838 157734
rect 2862 157732 2918 157734
rect 2622 156698 2678 156700
rect 2702 156698 2758 156700
rect 2782 156698 2838 156700
rect 2862 156698 2918 156700
rect 2622 156646 2648 156698
rect 2648 156646 2678 156698
rect 2702 156646 2712 156698
rect 2712 156646 2758 156698
rect 2782 156646 2828 156698
rect 2828 156646 2838 156698
rect 2862 156646 2892 156698
rect 2892 156646 2918 156698
rect 2622 156644 2678 156646
rect 2702 156644 2758 156646
rect 2782 156644 2838 156646
rect 2862 156644 2918 156646
rect 2622 155610 2678 155612
rect 2702 155610 2758 155612
rect 2782 155610 2838 155612
rect 2862 155610 2918 155612
rect 2622 155558 2648 155610
rect 2648 155558 2678 155610
rect 2702 155558 2712 155610
rect 2712 155558 2758 155610
rect 2782 155558 2828 155610
rect 2828 155558 2838 155610
rect 2862 155558 2892 155610
rect 2892 155558 2918 155610
rect 2622 155556 2678 155558
rect 2702 155556 2758 155558
rect 2782 155556 2838 155558
rect 2862 155556 2918 155558
rect 2622 154522 2678 154524
rect 2702 154522 2758 154524
rect 2782 154522 2838 154524
rect 2862 154522 2918 154524
rect 2622 154470 2648 154522
rect 2648 154470 2678 154522
rect 2702 154470 2712 154522
rect 2712 154470 2758 154522
rect 2782 154470 2828 154522
rect 2828 154470 2838 154522
rect 2862 154470 2892 154522
rect 2892 154470 2918 154522
rect 2622 154468 2678 154470
rect 2702 154468 2758 154470
rect 2782 154468 2838 154470
rect 2862 154468 2918 154470
rect 2622 153434 2678 153436
rect 2702 153434 2758 153436
rect 2782 153434 2838 153436
rect 2862 153434 2918 153436
rect 2622 153382 2648 153434
rect 2648 153382 2678 153434
rect 2702 153382 2712 153434
rect 2712 153382 2758 153434
rect 2782 153382 2828 153434
rect 2828 153382 2838 153434
rect 2862 153382 2892 153434
rect 2892 153382 2918 153434
rect 2622 153380 2678 153382
rect 2702 153380 2758 153382
rect 2782 153380 2838 153382
rect 2862 153380 2918 153382
rect 2622 152346 2678 152348
rect 2702 152346 2758 152348
rect 2782 152346 2838 152348
rect 2862 152346 2918 152348
rect 2622 152294 2648 152346
rect 2648 152294 2678 152346
rect 2702 152294 2712 152346
rect 2712 152294 2758 152346
rect 2782 152294 2828 152346
rect 2828 152294 2838 152346
rect 2862 152294 2892 152346
rect 2892 152294 2918 152346
rect 2622 152292 2678 152294
rect 2702 152292 2758 152294
rect 2782 152292 2838 152294
rect 2862 152292 2918 152294
rect 2622 151258 2678 151260
rect 2702 151258 2758 151260
rect 2782 151258 2838 151260
rect 2862 151258 2918 151260
rect 2622 151206 2648 151258
rect 2648 151206 2678 151258
rect 2702 151206 2712 151258
rect 2712 151206 2758 151258
rect 2782 151206 2828 151258
rect 2828 151206 2838 151258
rect 2862 151206 2892 151258
rect 2892 151206 2918 151258
rect 2622 151204 2678 151206
rect 2702 151204 2758 151206
rect 2782 151204 2838 151206
rect 2862 151204 2918 151206
rect 2622 150170 2678 150172
rect 2702 150170 2758 150172
rect 2782 150170 2838 150172
rect 2862 150170 2918 150172
rect 2622 150118 2648 150170
rect 2648 150118 2678 150170
rect 2702 150118 2712 150170
rect 2712 150118 2758 150170
rect 2782 150118 2828 150170
rect 2828 150118 2838 150170
rect 2862 150118 2892 150170
rect 2892 150118 2918 150170
rect 2622 150116 2678 150118
rect 2702 150116 2758 150118
rect 2782 150116 2838 150118
rect 2862 150116 2918 150118
rect 2622 149082 2678 149084
rect 2702 149082 2758 149084
rect 2782 149082 2838 149084
rect 2862 149082 2918 149084
rect 2622 149030 2648 149082
rect 2648 149030 2678 149082
rect 2702 149030 2712 149082
rect 2712 149030 2758 149082
rect 2782 149030 2828 149082
rect 2828 149030 2838 149082
rect 2862 149030 2892 149082
rect 2892 149030 2918 149082
rect 2622 149028 2678 149030
rect 2702 149028 2758 149030
rect 2782 149028 2838 149030
rect 2862 149028 2918 149030
rect 2622 147994 2678 147996
rect 2702 147994 2758 147996
rect 2782 147994 2838 147996
rect 2862 147994 2918 147996
rect 2622 147942 2648 147994
rect 2648 147942 2678 147994
rect 2702 147942 2712 147994
rect 2712 147942 2758 147994
rect 2782 147942 2828 147994
rect 2828 147942 2838 147994
rect 2862 147942 2892 147994
rect 2892 147942 2918 147994
rect 2622 147940 2678 147942
rect 2702 147940 2758 147942
rect 2782 147940 2838 147942
rect 2862 147940 2918 147942
rect 2622 146906 2678 146908
rect 2702 146906 2758 146908
rect 2782 146906 2838 146908
rect 2862 146906 2918 146908
rect 2622 146854 2648 146906
rect 2648 146854 2678 146906
rect 2702 146854 2712 146906
rect 2712 146854 2758 146906
rect 2782 146854 2828 146906
rect 2828 146854 2838 146906
rect 2862 146854 2892 146906
rect 2892 146854 2918 146906
rect 2622 146852 2678 146854
rect 2702 146852 2758 146854
rect 2782 146852 2838 146854
rect 2862 146852 2918 146854
rect 2622 145818 2678 145820
rect 2702 145818 2758 145820
rect 2782 145818 2838 145820
rect 2862 145818 2918 145820
rect 2622 145766 2648 145818
rect 2648 145766 2678 145818
rect 2702 145766 2712 145818
rect 2712 145766 2758 145818
rect 2782 145766 2828 145818
rect 2828 145766 2838 145818
rect 2862 145766 2892 145818
rect 2892 145766 2918 145818
rect 2622 145764 2678 145766
rect 2702 145764 2758 145766
rect 2782 145764 2838 145766
rect 2862 145764 2918 145766
rect 2622 144730 2678 144732
rect 2702 144730 2758 144732
rect 2782 144730 2838 144732
rect 2862 144730 2918 144732
rect 2622 144678 2648 144730
rect 2648 144678 2678 144730
rect 2702 144678 2712 144730
rect 2712 144678 2758 144730
rect 2782 144678 2828 144730
rect 2828 144678 2838 144730
rect 2862 144678 2892 144730
rect 2892 144678 2918 144730
rect 2622 144676 2678 144678
rect 2702 144676 2758 144678
rect 2782 144676 2838 144678
rect 2862 144676 2918 144678
rect 2622 143642 2678 143644
rect 2702 143642 2758 143644
rect 2782 143642 2838 143644
rect 2862 143642 2918 143644
rect 2622 143590 2648 143642
rect 2648 143590 2678 143642
rect 2702 143590 2712 143642
rect 2712 143590 2758 143642
rect 2782 143590 2828 143642
rect 2828 143590 2838 143642
rect 2862 143590 2892 143642
rect 2892 143590 2918 143642
rect 2622 143588 2678 143590
rect 2702 143588 2758 143590
rect 2782 143588 2838 143590
rect 2862 143588 2918 143590
rect 2622 142554 2678 142556
rect 2702 142554 2758 142556
rect 2782 142554 2838 142556
rect 2862 142554 2918 142556
rect 2622 142502 2648 142554
rect 2648 142502 2678 142554
rect 2702 142502 2712 142554
rect 2712 142502 2758 142554
rect 2782 142502 2828 142554
rect 2828 142502 2838 142554
rect 2862 142502 2892 142554
rect 2892 142502 2918 142554
rect 2622 142500 2678 142502
rect 2702 142500 2758 142502
rect 2782 142500 2838 142502
rect 2862 142500 2918 142502
rect 2622 141466 2678 141468
rect 2702 141466 2758 141468
rect 2782 141466 2838 141468
rect 2862 141466 2918 141468
rect 2622 141414 2648 141466
rect 2648 141414 2678 141466
rect 2702 141414 2712 141466
rect 2712 141414 2758 141466
rect 2782 141414 2828 141466
rect 2828 141414 2838 141466
rect 2862 141414 2892 141466
rect 2892 141414 2918 141466
rect 2622 141412 2678 141414
rect 2702 141412 2758 141414
rect 2782 141412 2838 141414
rect 2862 141412 2918 141414
rect 2622 140378 2678 140380
rect 2702 140378 2758 140380
rect 2782 140378 2838 140380
rect 2862 140378 2918 140380
rect 2622 140326 2648 140378
rect 2648 140326 2678 140378
rect 2702 140326 2712 140378
rect 2712 140326 2758 140378
rect 2782 140326 2828 140378
rect 2828 140326 2838 140378
rect 2862 140326 2892 140378
rect 2892 140326 2918 140378
rect 2622 140324 2678 140326
rect 2702 140324 2758 140326
rect 2782 140324 2838 140326
rect 2862 140324 2918 140326
rect 2622 139290 2678 139292
rect 2702 139290 2758 139292
rect 2782 139290 2838 139292
rect 2862 139290 2918 139292
rect 2622 139238 2648 139290
rect 2648 139238 2678 139290
rect 2702 139238 2712 139290
rect 2712 139238 2758 139290
rect 2782 139238 2828 139290
rect 2828 139238 2838 139290
rect 2862 139238 2892 139290
rect 2892 139238 2918 139290
rect 2622 139236 2678 139238
rect 2702 139236 2758 139238
rect 2782 139236 2838 139238
rect 2862 139236 2918 139238
rect 2622 138202 2678 138204
rect 2702 138202 2758 138204
rect 2782 138202 2838 138204
rect 2862 138202 2918 138204
rect 2622 138150 2648 138202
rect 2648 138150 2678 138202
rect 2702 138150 2712 138202
rect 2712 138150 2758 138202
rect 2782 138150 2828 138202
rect 2828 138150 2838 138202
rect 2862 138150 2892 138202
rect 2892 138150 2918 138202
rect 2622 138148 2678 138150
rect 2702 138148 2758 138150
rect 2782 138148 2838 138150
rect 2862 138148 2918 138150
rect 2622 137114 2678 137116
rect 2702 137114 2758 137116
rect 2782 137114 2838 137116
rect 2862 137114 2918 137116
rect 2622 137062 2648 137114
rect 2648 137062 2678 137114
rect 2702 137062 2712 137114
rect 2712 137062 2758 137114
rect 2782 137062 2828 137114
rect 2828 137062 2838 137114
rect 2862 137062 2892 137114
rect 2892 137062 2918 137114
rect 2622 137060 2678 137062
rect 2702 137060 2758 137062
rect 2782 137060 2838 137062
rect 2862 137060 2918 137062
rect 2622 136026 2678 136028
rect 2702 136026 2758 136028
rect 2782 136026 2838 136028
rect 2862 136026 2918 136028
rect 2622 135974 2648 136026
rect 2648 135974 2678 136026
rect 2702 135974 2712 136026
rect 2712 135974 2758 136026
rect 2782 135974 2828 136026
rect 2828 135974 2838 136026
rect 2862 135974 2892 136026
rect 2892 135974 2918 136026
rect 2622 135972 2678 135974
rect 2702 135972 2758 135974
rect 2782 135972 2838 135974
rect 2862 135972 2918 135974
rect 2622 134938 2678 134940
rect 2702 134938 2758 134940
rect 2782 134938 2838 134940
rect 2862 134938 2918 134940
rect 2622 134886 2648 134938
rect 2648 134886 2678 134938
rect 2702 134886 2712 134938
rect 2712 134886 2758 134938
rect 2782 134886 2828 134938
rect 2828 134886 2838 134938
rect 2862 134886 2892 134938
rect 2892 134886 2918 134938
rect 2622 134884 2678 134886
rect 2702 134884 2758 134886
rect 2782 134884 2838 134886
rect 2862 134884 2918 134886
rect 2622 133850 2678 133852
rect 2702 133850 2758 133852
rect 2782 133850 2838 133852
rect 2862 133850 2918 133852
rect 2622 133798 2648 133850
rect 2648 133798 2678 133850
rect 2702 133798 2712 133850
rect 2712 133798 2758 133850
rect 2782 133798 2828 133850
rect 2828 133798 2838 133850
rect 2862 133798 2892 133850
rect 2892 133798 2918 133850
rect 2622 133796 2678 133798
rect 2702 133796 2758 133798
rect 2782 133796 2838 133798
rect 2862 133796 2918 133798
rect 2622 132762 2678 132764
rect 2702 132762 2758 132764
rect 2782 132762 2838 132764
rect 2862 132762 2918 132764
rect 2622 132710 2648 132762
rect 2648 132710 2678 132762
rect 2702 132710 2712 132762
rect 2712 132710 2758 132762
rect 2782 132710 2828 132762
rect 2828 132710 2838 132762
rect 2862 132710 2892 132762
rect 2892 132710 2918 132762
rect 2622 132708 2678 132710
rect 2702 132708 2758 132710
rect 2782 132708 2838 132710
rect 2862 132708 2918 132710
rect 2622 131674 2678 131676
rect 2702 131674 2758 131676
rect 2782 131674 2838 131676
rect 2862 131674 2918 131676
rect 2622 131622 2648 131674
rect 2648 131622 2678 131674
rect 2702 131622 2712 131674
rect 2712 131622 2758 131674
rect 2782 131622 2828 131674
rect 2828 131622 2838 131674
rect 2862 131622 2892 131674
rect 2892 131622 2918 131674
rect 2622 131620 2678 131622
rect 2702 131620 2758 131622
rect 2782 131620 2838 131622
rect 2862 131620 2918 131622
rect 2622 130586 2678 130588
rect 2702 130586 2758 130588
rect 2782 130586 2838 130588
rect 2862 130586 2918 130588
rect 2622 130534 2648 130586
rect 2648 130534 2678 130586
rect 2702 130534 2712 130586
rect 2712 130534 2758 130586
rect 2782 130534 2828 130586
rect 2828 130534 2838 130586
rect 2862 130534 2892 130586
rect 2892 130534 2918 130586
rect 2622 130532 2678 130534
rect 2702 130532 2758 130534
rect 2782 130532 2838 130534
rect 2862 130532 2918 130534
rect 2622 129498 2678 129500
rect 2702 129498 2758 129500
rect 2782 129498 2838 129500
rect 2862 129498 2918 129500
rect 2622 129446 2648 129498
rect 2648 129446 2678 129498
rect 2702 129446 2712 129498
rect 2712 129446 2758 129498
rect 2782 129446 2828 129498
rect 2828 129446 2838 129498
rect 2862 129446 2892 129498
rect 2892 129446 2918 129498
rect 2622 129444 2678 129446
rect 2702 129444 2758 129446
rect 2782 129444 2838 129446
rect 2862 129444 2918 129446
rect 2622 128410 2678 128412
rect 2702 128410 2758 128412
rect 2782 128410 2838 128412
rect 2862 128410 2918 128412
rect 2622 128358 2648 128410
rect 2648 128358 2678 128410
rect 2702 128358 2712 128410
rect 2712 128358 2758 128410
rect 2782 128358 2828 128410
rect 2828 128358 2838 128410
rect 2862 128358 2892 128410
rect 2892 128358 2918 128410
rect 2622 128356 2678 128358
rect 2702 128356 2758 128358
rect 2782 128356 2838 128358
rect 2862 128356 2918 128358
rect 2622 127322 2678 127324
rect 2702 127322 2758 127324
rect 2782 127322 2838 127324
rect 2862 127322 2918 127324
rect 2622 127270 2648 127322
rect 2648 127270 2678 127322
rect 2702 127270 2712 127322
rect 2712 127270 2758 127322
rect 2782 127270 2828 127322
rect 2828 127270 2838 127322
rect 2862 127270 2892 127322
rect 2892 127270 2918 127322
rect 2622 127268 2678 127270
rect 2702 127268 2758 127270
rect 2782 127268 2838 127270
rect 2862 127268 2918 127270
rect 2622 126234 2678 126236
rect 2702 126234 2758 126236
rect 2782 126234 2838 126236
rect 2862 126234 2918 126236
rect 2622 126182 2648 126234
rect 2648 126182 2678 126234
rect 2702 126182 2712 126234
rect 2712 126182 2758 126234
rect 2782 126182 2828 126234
rect 2828 126182 2838 126234
rect 2862 126182 2892 126234
rect 2892 126182 2918 126234
rect 2622 126180 2678 126182
rect 2702 126180 2758 126182
rect 2782 126180 2838 126182
rect 2862 126180 2918 126182
rect 2622 125146 2678 125148
rect 2702 125146 2758 125148
rect 2782 125146 2838 125148
rect 2862 125146 2918 125148
rect 2622 125094 2648 125146
rect 2648 125094 2678 125146
rect 2702 125094 2712 125146
rect 2712 125094 2758 125146
rect 2782 125094 2828 125146
rect 2828 125094 2838 125146
rect 2862 125094 2892 125146
rect 2892 125094 2918 125146
rect 2622 125092 2678 125094
rect 2702 125092 2758 125094
rect 2782 125092 2838 125094
rect 2862 125092 2918 125094
rect 2622 124058 2678 124060
rect 2702 124058 2758 124060
rect 2782 124058 2838 124060
rect 2862 124058 2918 124060
rect 2622 124006 2648 124058
rect 2648 124006 2678 124058
rect 2702 124006 2712 124058
rect 2712 124006 2758 124058
rect 2782 124006 2828 124058
rect 2828 124006 2838 124058
rect 2862 124006 2892 124058
rect 2892 124006 2918 124058
rect 2622 124004 2678 124006
rect 2702 124004 2758 124006
rect 2782 124004 2838 124006
rect 2862 124004 2918 124006
rect 2622 122970 2678 122972
rect 2702 122970 2758 122972
rect 2782 122970 2838 122972
rect 2862 122970 2918 122972
rect 2622 122918 2648 122970
rect 2648 122918 2678 122970
rect 2702 122918 2712 122970
rect 2712 122918 2758 122970
rect 2782 122918 2828 122970
rect 2828 122918 2838 122970
rect 2862 122918 2892 122970
rect 2892 122918 2918 122970
rect 2622 122916 2678 122918
rect 2702 122916 2758 122918
rect 2782 122916 2838 122918
rect 2862 122916 2918 122918
rect 2622 121882 2678 121884
rect 2702 121882 2758 121884
rect 2782 121882 2838 121884
rect 2862 121882 2918 121884
rect 2622 121830 2648 121882
rect 2648 121830 2678 121882
rect 2702 121830 2712 121882
rect 2712 121830 2758 121882
rect 2782 121830 2828 121882
rect 2828 121830 2838 121882
rect 2862 121830 2892 121882
rect 2892 121830 2918 121882
rect 2622 121828 2678 121830
rect 2702 121828 2758 121830
rect 2782 121828 2838 121830
rect 2862 121828 2918 121830
rect 2622 120794 2678 120796
rect 2702 120794 2758 120796
rect 2782 120794 2838 120796
rect 2862 120794 2918 120796
rect 2622 120742 2648 120794
rect 2648 120742 2678 120794
rect 2702 120742 2712 120794
rect 2712 120742 2758 120794
rect 2782 120742 2828 120794
rect 2828 120742 2838 120794
rect 2862 120742 2892 120794
rect 2892 120742 2918 120794
rect 2622 120740 2678 120742
rect 2702 120740 2758 120742
rect 2782 120740 2838 120742
rect 2862 120740 2918 120742
rect 2622 119706 2678 119708
rect 2702 119706 2758 119708
rect 2782 119706 2838 119708
rect 2862 119706 2918 119708
rect 2622 119654 2648 119706
rect 2648 119654 2678 119706
rect 2702 119654 2712 119706
rect 2712 119654 2758 119706
rect 2782 119654 2828 119706
rect 2828 119654 2838 119706
rect 2862 119654 2892 119706
rect 2892 119654 2918 119706
rect 2622 119652 2678 119654
rect 2702 119652 2758 119654
rect 2782 119652 2838 119654
rect 2862 119652 2918 119654
rect 2622 118618 2678 118620
rect 2702 118618 2758 118620
rect 2782 118618 2838 118620
rect 2862 118618 2918 118620
rect 2622 118566 2648 118618
rect 2648 118566 2678 118618
rect 2702 118566 2712 118618
rect 2712 118566 2758 118618
rect 2782 118566 2828 118618
rect 2828 118566 2838 118618
rect 2862 118566 2892 118618
rect 2892 118566 2918 118618
rect 2622 118564 2678 118566
rect 2702 118564 2758 118566
rect 2782 118564 2838 118566
rect 2862 118564 2918 118566
rect 2622 117530 2678 117532
rect 2702 117530 2758 117532
rect 2782 117530 2838 117532
rect 2862 117530 2918 117532
rect 2622 117478 2648 117530
rect 2648 117478 2678 117530
rect 2702 117478 2712 117530
rect 2712 117478 2758 117530
rect 2782 117478 2828 117530
rect 2828 117478 2838 117530
rect 2862 117478 2892 117530
rect 2892 117478 2918 117530
rect 2622 117476 2678 117478
rect 2702 117476 2758 117478
rect 2782 117476 2838 117478
rect 2862 117476 2918 117478
rect 2622 116442 2678 116444
rect 2702 116442 2758 116444
rect 2782 116442 2838 116444
rect 2862 116442 2918 116444
rect 2622 116390 2648 116442
rect 2648 116390 2678 116442
rect 2702 116390 2712 116442
rect 2712 116390 2758 116442
rect 2782 116390 2828 116442
rect 2828 116390 2838 116442
rect 2862 116390 2892 116442
rect 2892 116390 2918 116442
rect 2622 116388 2678 116390
rect 2702 116388 2758 116390
rect 2782 116388 2838 116390
rect 2862 116388 2918 116390
rect 2622 115354 2678 115356
rect 2702 115354 2758 115356
rect 2782 115354 2838 115356
rect 2862 115354 2918 115356
rect 2622 115302 2648 115354
rect 2648 115302 2678 115354
rect 2702 115302 2712 115354
rect 2712 115302 2758 115354
rect 2782 115302 2828 115354
rect 2828 115302 2838 115354
rect 2862 115302 2892 115354
rect 2892 115302 2918 115354
rect 2622 115300 2678 115302
rect 2702 115300 2758 115302
rect 2782 115300 2838 115302
rect 2862 115300 2918 115302
rect 2622 114266 2678 114268
rect 2702 114266 2758 114268
rect 2782 114266 2838 114268
rect 2862 114266 2918 114268
rect 2622 114214 2648 114266
rect 2648 114214 2678 114266
rect 2702 114214 2712 114266
rect 2712 114214 2758 114266
rect 2782 114214 2828 114266
rect 2828 114214 2838 114266
rect 2862 114214 2892 114266
rect 2892 114214 2918 114266
rect 2622 114212 2678 114214
rect 2702 114212 2758 114214
rect 2782 114212 2838 114214
rect 2862 114212 2918 114214
rect 2622 113178 2678 113180
rect 2702 113178 2758 113180
rect 2782 113178 2838 113180
rect 2862 113178 2918 113180
rect 2622 113126 2648 113178
rect 2648 113126 2678 113178
rect 2702 113126 2712 113178
rect 2712 113126 2758 113178
rect 2782 113126 2828 113178
rect 2828 113126 2838 113178
rect 2862 113126 2892 113178
rect 2892 113126 2918 113178
rect 2622 113124 2678 113126
rect 2702 113124 2758 113126
rect 2782 113124 2838 113126
rect 2862 113124 2918 113126
rect 2622 112090 2678 112092
rect 2702 112090 2758 112092
rect 2782 112090 2838 112092
rect 2862 112090 2918 112092
rect 2622 112038 2648 112090
rect 2648 112038 2678 112090
rect 2702 112038 2712 112090
rect 2712 112038 2758 112090
rect 2782 112038 2828 112090
rect 2828 112038 2838 112090
rect 2862 112038 2892 112090
rect 2892 112038 2918 112090
rect 2622 112036 2678 112038
rect 2702 112036 2758 112038
rect 2782 112036 2838 112038
rect 2862 112036 2918 112038
rect 2622 111002 2678 111004
rect 2702 111002 2758 111004
rect 2782 111002 2838 111004
rect 2862 111002 2918 111004
rect 2622 110950 2648 111002
rect 2648 110950 2678 111002
rect 2702 110950 2712 111002
rect 2712 110950 2758 111002
rect 2782 110950 2828 111002
rect 2828 110950 2838 111002
rect 2862 110950 2892 111002
rect 2892 110950 2918 111002
rect 2622 110948 2678 110950
rect 2702 110948 2758 110950
rect 2782 110948 2838 110950
rect 2862 110948 2918 110950
rect 2622 109914 2678 109916
rect 2702 109914 2758 109916
rect 2782 109914 2838 109916
rect 2862 109914 2918 109916
rect 2622 109862 2648 109914
rect 2648 109862 2678 109914
rect 2702 109862 2712 109914
rect 2712 109862 2758 109914
rect 2782 109862 2828 109914
rect 2828 109862 2838 109914
rect 2862 109862 2892 109914
rect 2892 109862 2918 109914
rect 2622 109860 2678 109862
rect 2702 109860 2758 109862
rect 2782 109860 2838 109862
rect 2862 109860 2918 109862
rect 2622 108826 2678 108828
rect 2702 108826 2758 108828
rect 2782 108826 2838 108828
rect 2862 108826 2918 108828
rect 2622 108774 2648 108826
rect 2648 108774 2678 108826
rect 2702 108774 2712 108826
rect 2712 108774 2758 108826
rect 2782 108774 2828 108826
rect 2828 108774 2838 108826
rect 2862 108774 2892 108826
rect 2892 108774 2918 108826
rect 2622 108772 2678 108774
rect 2702 108772 2758 108774
rect 2782 108772 2838 108774
rect 2862 108772 2918 108774
rect 2622 107738 2678 107740
rect 2702 107738 2758 107740
rect 2782 107738 2838 107740
rect 2862 107738 2918 107740
rect 2622 107686 2648 107738
rect 2648 107686 2678 107738
rect 2702 107686 2712 107738
rect 2712 107686 2758 107738
rect 2782 107686 2828 107738
rect 2828 107686 2838 107738
rect 2862 107686 2892 107738
rect 2892 107686 2918 107738
rect 2622 107684 2678 107686
rect 2702 107684 2758 107686
rect 2782 107684 2838 107686
rect 2862 107684 2918 107686
rect 2622 106650 2678 106652
rect 2702 106650 2758 106652
rect 2782 106650 2838 106652
rect 2862 106650 2918 106652
rect 2622 106598 2648 106650
rect 2648 106598 2678 106650
rect 2702 106598 2712 106650
rect 2712 106598 2758 106650
rect 2782 106598 2828 106650
rect 2828 106598 2838 106650
rect 2862 106598 2892 106650
rect 2892 106598 2918 106650
rect 2622 106596 2678 106598
rect 2702 106596 2758 106598
rect 2782 106596 2838 106598
rect 2862 106596 2918 106598
rect 2622 105562 2678 105564
rect 2702 105562 2758 105564
rect 2782 105562 2838 105564
rect 2862 105562 2918 105564
rect 2622 105510 2648 105562
rect 2648 105510 2678 105562
rect 2702 105510 2712 105562
rect 2712 105510 2758 105562
rect 2782 105510 2828 105562
rect 2828 105510 2838 105562
rect 2862 105510 2892 105562
rect 2892 105510 2918 105562
rect 2622 105508 2678 105510
rect 2702 105508 2758 105510
rect 2782 105508 2838 105510
rect 2862 105508 2918 105510
rect 2622 104474 2678 104476
rect 2702 104474 2758 104476
rect 2782 104474 2838 104476
rect 2862 104474 2918 104476
rect 2622 104422 2648 104474
rect 2648 104422 2678 104474
rect 2702 104422 2712 104474
rect 2712 104422 2758 104474
rect 2782 104422 2828 104474
rect 2828 104422 2838 104474
rect 2862 104422 2892 104474
rect 2892 104422 2918 104474
rect 2622 104420 2678 104422
rect 2702 104420 2758 104422
rect 2782 104420 2838 104422
rect 2862 104420 2918 104422
rect 2622 103386 2678 103388
rect 2702 103386 2758 103388
rect 2782 103386 2838 103388
rect 2862 103386 2918 103388
rect 2622 103334 2648 103386
rect 2648 103334 2678 103386
rect 2702 103334 2712 103386
rect 2712 103334 2758 103386
rect 2782 103334 2828 103386
rect 2828 103334 2838 103386
rect 2862 103334 2892 103386
rect 2892 103334 2918 103386
rect 2622 103332 2678 103334
rect 2702 103332 2758 103334
rect 2782 103332 2838 103334
rect 2862 103332 2918 103334
rect 2622 102298 2678 102300
rect 2702 102298 2758 102300
rect 2782 102298 2838 102300
rect 2862 102298 2918 102300
rect 2622 102246 2648 102298
rect 2648 102246 2678 102298
rect 2702 102246 2712 102298
rect 2712 102246 2758 102298
rect 2782 102246 2828 102298
rect 2828 102246 2838 102298
rect 2862 102246 2892 102298
rect 2892 102246 2918 102298
rect 2622 102244 2678 102246
rect 2702 102244 2758 102246
rect 2782 102244 2838 102246
rect 2862 102244 2918 102246
rect 2622 101210 2678 101212
rect 2702 101210 2758 101212
rect 2782 101210 2838 101212
rect 2862 101210 2918 101212
rect 2622 101158 2648 101210
rect 2648 101158 2678 101210
rect 2702 101158 2712 101210
rect 2712 101158 2758 101210
rect 2782 101158 2828 101210
rect 2828 101158 2838 101210
rect 2862 101158 2892 101210
rect 2892 101158 2918 101210
rect 2622 101156 2678 101158
rect 2702 101156 2758 101158
rect 2782 101156 2838 101158
rect 2862 101156 2918 101158
rect 2622 100122 2678 100124
rect 2702 100122 2758 100124
rect 2782 100122 2838 100124
rect 2862 100122 2918 100124
rect 2622 100070 2648 100122
rect 2648 100070 2678 100122
rect 2702 100070 2712 100122
rect 2712 100070 2758 100122
rect 2782 100070 2828 100122
rect 2828 100070 2838 100122
rect 2862 100070 2892 100122
rect 2892 100070 2918 100122
rect 2622 100068 2678 100070
rect 2702 100068 2758 100070
rect 2782 100068 2838 100070
rect 2862 100068 2918 100070
rect 2622 99034 2678 99036
rect 2702 99034 2758 99036
rect 2782 99034 2838 99036
rect 2862 99034 2918 99036
rect 2622 98982 2648 99034
rect 2648 98982 2678 99034
rect 2702 98982 2712 99034
rect 2712 98982 2758 99034
rect 2782 98982 2828 99034
rect 2828 98982 2838 99034
rect 2862 98982 2892 99034
rect 2892 98982 2918 99034
rect 2622 98980 2678 98982
rect 2702 98980 2758 98982
rect 2782 98980 2838 98982
rect 2862 98980 2918 98982
rect 2622 97946 2678 97948
rect 2702 97946 2758 97948
rect 2782 97946 2838 97948
rect 2862 97946 2918 97948
rect 2622 97894 2648 97946
rect 2648 97894 2678 97946
rect 2702 97894 2712 97946
rect 2712 97894 2758 97946
rect 2782 97894 2828 97946
rect 2828 97894 2838 97946
rect 2862 97894 2892 97946
rect 2892 97894 2918 97946
rect 2622 97892 2678 97894
rect 2702 97892 2758 97894
rect 2782 97892 2838 97894
rect 2862 97892 2918 97894
rect 2622 96858 2678 96860
rect 2702 96858 2758 96860
rect 2782 96858 2838 96860
rect 2862 96858 2918 96860
rect 2622 96806 2648 96858
rect 2648 96806 2678 96858
rect 2702 96806 2712 96858
rect 2712 96806 2758 96858
rect 2782 96806 2828 96858
rect 2828 96806 2838 96858
rect 2862 96806 2892 96858
rect 2892 96806 2918 96858
rect 2622 96804 2678 96806
rect 2702 96804 2758 96806
rect 2782 96804 2838 96806
rect 2862 96804 2918 96806
rect 2622 95770 2678 95772
rect 2702 95770 2758 95772
rect 2782 95770 2838 95772
rect 2862 95770 2918 95772
rect 2622 95718 2648 95770
rect 2648 95718 2678 95770
rect 2702 95718 2712 95770
rect 2712 95718 2758 95770
rect 2782 95718 2828 95770
rect 2828 95718 2838 95770
rect 2862 95718 2892 95770
rect 2892 95718 2918 95770
rect 2622 95716 2678 95718
rect 2702 95716 2758 95718
rect 2782 95716 2838 95718
rect 2862 95716 2918 95718
rect 2622 94682 2678 94684
rect 2702 94682 2758 94684
rect 2782 94682 2838 94684
rect 2862 94682 2918 94684
rect 2622 94630 2648 94682
rect 2648 94630 2678 94682
rect 2702 94630 2712 94682
rect 2712 94630 2758 94682
rect 2782 94630 2828 94682
rect 2828 94630 2838 94682
rect 2862 94630 2892 94682
rect 2892 94630 2918 94682
rect 2622 94628 2678 94630
rect 2702 94628 2758 94630
rect 2782 94628 2838 94630
rect 2862 94628 2918 94630
rect 2622 93594 2678 93596
rect 2702 93594 2758 93596
rect 2782 93594 2838 93596
rect 2862 93594 2918 93596
rect 2622 93542 2648 93594
rect 2648 93542 2678 93594
rect 2702 93542 2712 93594
rect 2712 93542 2758 93594
rect 2782 93542 2828 93594
rect 2828 93542 2838 93594
rect 2862 93542 2892 93594
rect 2892 93542 2918 93594
rect 2622 93540 2678 93542
rect 2702 93540 2758 93542
rect 2782 93540 2838 93542
rect 2862 93540 2918 93542
rect 2622 92506 2678 92508
rect 2702 92506 2758 92508
rect 2782 92506 2838 92508
rect 2862 92506 2918 92508
rect 2622 92454 2648 92506
rect 2648 92454 2678 92506
rect 2702 92454 2712 92506
rect 2712 92454 2758 92506
rect 2782 92454 2828 92506
rect 2828 92454 2838 92506
rect 2862 92454 2892 92506
rect 2892 92454 2918 92506
rect 2622 92452 2678 92454
rect 2702 92452 2758 92454
rect 2782 92452 2838 92454
rect 2862 92452 2918 92454
rect 2622 91418 2678 91420
rect 2702 91418 2758 91420
rect 2782 91418 2838 91420
rect 2862 91418 2918 91420
rect 2622 91366 2648 91418
rect 2648 91366 2678 91418
rect 2702 91366 2712 91418
rect 2712 91366 2758 91418
rect 2782 91366 2828 91418
rect 2828 91366 2838 91418
rect 2862 91366 2892 91418
rect 2892 91366 2918 91418
rect 2622 91364 2678 91366
rect 2702 91364 2758 91366
rect 2782 91364 2838 91366
rect 2862 91364 2918 91366
rect 2622 90330 2678 90332
rect 2702 90330 2758 90332
rect 2782 90330 2838 90332
rect 2862 90330 2918 90332
rect 2622 90278 2648 90330
rect 2648 90278 2678 90330
rect 2702 90278 2712 90330
rect 2712 90278 2758 90330
rect 2782 90278 2828 90330
rect 2828 90278 2838 90330
rect 2862 90278 2892 90330
rect 2892 90278 2918 90330
rect 2622 90276 2678 90278
rect 2702 90276 2758 90278
rect 2782 90276 2838 90278
rect 2862 90276 2918 90278
rect 2622 89242 2678 89244
rect 2702 89242 2758 89244
rect 2782 89242 2838 89244
rect 2862 89242 2918 89244
rect 2622 89190 2648 89242
rect 2648 89190 2678 89242
rect 2702 89190 2712 89242
rect 2712 89190 2758 89242
rect 2782 89190 2828 89242
rect 2828 89190 2838 89242
rect 2862 89190 2892 89242
rect 2892 89190 2918 89242
rect 2622 89188 2678 89190
rect 2702 89188 2758 89190
rect 2782 89188 2838 89190
rect 2862 89188 2918 89190
rect 2622 88154 2678 88156
rect 2702 88154 2758 88156
rect 2782 88154 2838 88156
rect 2862 88154 2918 88156
rect 2622 88102 2648 88154
rect 2648 88102 2678 88154
rect 2702 88102 2712 88154
rect 2712 88102 2758 88154
rect 2782 88102 2828 88154
rect 2828 88102 2838 88154
rect 2862 88102 2892 88154
rect 2892 88102 2918 88154
rect 2622 88100 2678 88102
rect 2702 88100 2758 88102
rect 2782 88100 2838 88102
rect 2862 88100 2918 88102
rect 2622 87066 2678 87068
rect 2702 87066 2758 87068
rect 2782 87066 2838 87068
rect 2862 87066 2918 87068
rect 2622 87014 2648 87066
rect 2648 87014 2678 87066
rect 2702 87014 2712 87066
rect 2712 87014 2758 87066
rect 2782 87014 2828 87066
rect 2828 87014 2838 87066
rect 2862 87014 2892 87066
rect 2892 87014 2918 87066
rect 2622 87012 2678 87014
rect 2702 87012 2758 87014
rect 2782 87012 2838 87014
rect 2862 87012 2918 87014
rect 2622 85978 2678 85980
rect 2702 85978 2758 85980
rect 2782 85978 2838 85980
rect 2862 85978 2918 85980
rect 2622 85926 2648 85978
rect 2648 85926 2678 85978
rect 2702 85926 2712 85978
rect 2712 85926 2758 85978
rect 2782 85926 2828 85978
rect 2828 85926 2838 85978
rect 2862 85926 2892 85978
rect 2892 85926 2918 85978
rect 2622 85924 2678 85926
rect 2702 85924 2758 85926
rect 2782 85924 2838 85926
rect 2862 85924 2918 85926
rect 2622 84890 2678 84892
rect 2702 84890 2758 84892
rect 2782 84890 2838 84892
rect 2862 84890 2918 84892
rect 2622 84838 2648 84890
rect 2648 84838 2678 84890
rect 2702 84838 2712 84890
rect 2712 84838 2758 84890
rect 2782 84838 2828 84890
rect 2828 84838 2838 84890
rect 2862 84838 2892 84890
rect 2892 84838 2918 84890
rect 2622 84836 2678 84838
rect 2702 84836 2758 84838
rect 2782 84836 2838 84838
rect 2862 84836 2918 84838
rect 2622 83802 2678 83804
rect 2702 83802 2758 83804
rect 2782 83802 2838 83804
rect 2862 83802 2918 83804
rect 2622 83750 2648 83802
rect 2648 83750 2678 83802
rect 2702 83750 2712 83802
rect 2712 83750 2758 83802
rect 2782 83750 2828 83802
rect 2828 83750 2838 83802
rect 2862 83750 2892 83802
rect 2892 83750 2918 83802
rect 2622 83748 2678 83750
rect 2702 83748 2758 83750
rect 2782 83748 2838 83750
rect 2862 83748 2918 83750
rect 2622 82714 2678 82716
rect 2702 82714 2758 82716
rect 2782 82714 2838 82716
rect 2862 82714 2918 82716
rect 2622 82662 2648 82714
rect 2648 82662 2678 82714
rect 2702 82662 2712 82714
rect 2712 82662 2758 82714
rect 2782 82662 2828 82714
rect 2828 82662 2838 82714
rect 2862 82662 2892 82714
rect 2892 82662 2918 82714
rect 2622 82660 2678 82662
rect 2702 82660 2758 82662
rect 2782 82660 2838 82662
rect 2862 82660 2918 82662
rect 2622 81626 2678 81628
rect 2702 81626 2758 81628
rect 2782 81626 2838 81628
rect 2862 81626 2918 81628
rect 2622 81574 2648 81626
rect 2648 81574 2678 81626
rect 2702 81574 2712 81626
rect 2712 81574 2758 81626
rect 2782 81574 2828 81626
rect 2828 81574 2838 81626
rect 2862 81574 2892 81626
rect 2892 81574 2918 81626
rect 2622 81572 2678 81574
rect 2702 81572 2758 81574
rect 2782 81572 2838 81574
rect 2862 81572 2918 81574
rect 2622 80538 2678 80540
rect 2702 80538 2758 80540
rect 2782 80538 2838 80540
rect 2862 80538 2918 80540
rect 2622 80486 2648 80538
rect 2648 80486 2678 80538
rect 2702 80486 2712 80538
rect 2712 80486 2758 80538
rect 2782 80486 2828 80538
rect 2828 80486 2838 80538
rect 2862 80486 2892 80538
rect 2892 80486 2918 80538
rect 2622 80484 2678 80486
rect 2702 80484 2758 80486
rect 2782 80484 2838 80486
rect 2862 80484 2918 80486
rect 2622 79450 2678 79452
rect 2702 79450 2758 79452
rect 2782 79450 2838 79452
rect 2862 79450 2918 79452
rect 2622 79398 2648 79450
rect 2648 79398 2678 79450
rect 2702 79398 2712 79450
rect 2712 79398 2758 79450
rect 2782 79398 2828 79450
rect 2828 79398 2838 79450
rect 2862 79398 2892 79450
rect 2892 79398 2918 79450
rect 2622 79396 2678 79398
rect 2702 79396 2758 79398
rect 2782 79396 2838 79398
rect 2862 79396 2918 79398
rect 2622 78362 2678 78364
rect 2702 78362 2758 78364
rect 2782 78362 2838 78364
rect 2862 78362 2918 78364
rect 2622 78310 2648 78362
rect 2648 78310 2678 78362
rect 2702 78310 2712 78362
rect 2712 78310 2758 78362
rect 2782 78310 2828 78362
rect 2828 78310 2838 78362
rect 2862 78310 2892 78362
rect 2892 78310 2918 78362
rect 2622 78308 2678 78310
rect 2702 78308 2758 78310
rect 2782 78308 2838 78310
rect 2862 78308 2918 78310
rect 2622 77274 2678 77276
rect 2702 77274 2758 77276
rect 2782 77274 2838 77276
rect 2862 77274 2918 77276
rect 2622 77222 2648 77274
rect 2648 77222 2678 77274
rect 2702 77222 2712 77274
rect 2712 77222 2758 77274
rect 2782 77222 2828 77274
rect 2828 77222 2838 77274
rect 2862 77222 2892 77274
rect 2892 77222 2918 77274
rect 2622 77220 2678 77222
rect 2702 77220 2758 77222
rect 2782 77220 2838 77222
rect 2862 77220 2918 77222
rect 2622 76186 2678 76188
rect 2702 76186 2758 76188
rect 2782 76186 2838 76188
rect 2862 76186 2918 76188
rect 2622 76134 2648 76186
rect 2648 76134 2678 76186
rect 2702 76134 2712 76186
rect 2712 76134 2758 76186
rect 2782 76134 2828 76186
rect 2828 76134 2838 76186
rect 2862 76134 2892 76186
rect 2892 76134 2918 76186
rect 2622 76132 2678 76134
rect 2702 76132 2758 76134
rect 2782 76132 2838 76134
rect 2862 76132 2918 76134
rect 2622 75098 2678 75100
rect 2702 75098 2758 75100
rect 2782 75098 2838 75100
rect 2862 75098 2918 75100
rect 2622 75046 2648 75098
rect 2648 75046 2678 75098
rect 2702 75046 2712 75098
rect 2712 75046 2758 75098
rect 2782 75046 2828 75098
rect 2828 75046 2838 75098
rect 2862 75046 2892 75098
rect 2892 75046 2918 75098
rect 2622 75044 2678 75046
rect 2702 75044 2758 75046
rect 2782 75044 2838 75046
rect 2862 75044 2918 75046
rect 2622 74010 2678 74012
rect 2702 74010 2758 74012
rect 2782 74010 2838 74012
rect 2862 74010 2918 74012
rect 2622 73958 2648 74010
rect 2648 73958 2678 74010
rect 2702 73958 2712 74010
rect 2712 73958 2758 74010
rect 2782 73958 2828 74010
rect 2828 73958 2838 74010
rect 2862 73958 2892 74010
rect 2892 73958 2918 74010
rect 2622 73956 2678 73958
rect 2702 73956 2758 73958
rect 2782 73956 2838 73958
rect 2862 73956 2918 73958
rect 2622 72922 2678 72924
rect 2702 72922 2758 72924
rect 2782 72922 2838 72924
rect 2862 72922 2918 72924
rect 2622 72870 2648 72922
rect 2648 72870 2678 72922
rect 2702 72870 2712 72922
rect 2712 72870 2758 72922
rect 2782 72870 2828 72922
rect 2828 72870 2838 72922
rect 2862 72870 2892 72922
rect 2892 72870 2918 72922
rect 2622 72868 2678 72870
rect 2702 72868 2758 72870
rect 2782 72868 2838 72870
rect 2862 72868 2918 72870
rect 2622 71834 2678 71836
rect 2702 71834 2758 71836
rect 2782 71834 2838 71836
rect 2862 71834 2918 71836
rect 2622 71782 2648 71834
rect 2648 71782 2678 71834
rect 2702 71782 2712 71834
rect 2712 71782 2758 71834
rect 2782 71782 2828 71834
rect 2828 71782 2838 71834
rect 2862 71782 2892 71834
rect 2892 71782 2918 71834
rect 2622 71780 2678 71782
rect 2702 71780 2758 71782
rect 2782 71780 2838 71782
rect 2862 71780 2918 71782
rect 2622 70746 2678 70748
rect 2702 70746 2758 70748
rect 2782 70746 2838 70748
rect 2862 70746 2918 70748
rect 2622 70694 2648 70746
rect 2648 70694 2678 70746
rect 2702 70694 2712 70746
rect 2712 70694 2758 70746
rect 2782 70694 2828 70746
rect 2828 70694 2838 70746
rect 2862 70694 2892 70746
rect 2892 70694 2918 70746
rect 2622 70692 2678 70694
rect 2702 70692 2758 70694
rect 2782 70692 2838 70694
rect 2862 70692 2918 70694
rect 2622 69658 2678 69660
rect 2702 69658 2758 69660
rect 2782 69658 2838 69660
rect 2862 69658 2918 69660
rect 2622 69606 2648 69658
rect 2648 69606 2678 69658
rect 2702 69606 2712 69658
rect 2712 69606 2758 69658
rect 2782 69606 2828 69658
rect 2828 69606 2838 69658
rect 2862 69606 2892 69658
rect 2892 69606 2918 69658
rect 2622 69604 2678 69606
rect 2702 69604 2758 69606
rect 2782 69604 2838 69606
rect 2862 69604 2918 69606
rect 2622 68570 2678 68572
rect 2702 68570 2758 68572
rect 2782 68570 2838 68572
rect 2862 68570 2918 68572
rect 2622 68518 2648 68570
rect 2648 68518 2678 68570
rect 2702 68518 2712 68570
rect 2712 68518 2758 68570
rect 2782 68518 2828 68570
rect 2828 68518 2838 68570
rect 2862 68518 2892 68570
rect 2892 68518 2918 68570
rect 2622 68516 2678 68518
rect 2702 68516 2758 68518
rect 2782 68516 2838 68518
rect 2862 68516 2918 68518
rect 2622 67482 2678 67484
rect 2702 67482 2758 67484
rect 2782 67482 2838 67484
rect 2862 67482 2918 67484
rect 2622 67430 2648 67482
rect 2648 67430 2678 67482
rect 2702 67430 2712 67482
rect 2712 67430 2758 67482
rect 2782 67430 2828 67482
rect 2828 67430 2838 67482
rect 2862 67430 2892 67482
rect 2892 67430 2918 67482
rect 2622 67428 2678 67430
rect 2702 67428 2758 67430
rect 2782 67428 2838 67430
rect 2862 67428 2918 67430
rect 2622 66394 2678 66396
rect 2702 66394 2758 66396
rect 2782 66394 2838 66396
rect 2862 66394 2918 66396
rect 2622 66342 2648 66394
rect 2648 66342 2678 66394
rect 2702 66342 2712 66394
rect 2712 66342 2758 66394
rect 2782 66342 2828 66394
rect 2828 66342 2838 66394
rect 2862 66342 2892 66394
rect 2892 66342 2918 66394
rect 2622 66340 2678 66342
rect 2702 66340 2758 66342
rect 2782 66340 2838 66342
rect 2862 66340 2918 66342
rect 2622 65306 2678 65308
rect 2702 65306 2758 65308
rect 2782 65306 2838 65308
rect 2862 65306 2918 65308
rect 2622 65254 2648 65306
rect 2648 65254 2678 65306
rect 2702 65254 2712 65306
rect 2712 65254 2758 65306
rect 2782 65254 2828 65306
rect 2828 65254 2838 65306
rect 2862 65254 2892 65306
rect 2892 65254 2918 65306
rect 2622 65252 2678 65254
rect 2702 65252 2758 65254
rect 2782 65252 2838 65254
rect 2862 65252 2918 65254
rect 2622 64218 2678 64220
rect 2702 64218 2758 64220
rect 2782 64218 2838 64220
rect 2862 64218 2918 64220
rect 2622 64166 2648 64218
rect 2648 64166 2678 64218
rect 2702 64166 2712 64218
rect 2712 64166 2758 64218
rect 2782 64166 2828 64218
rect 2828 64166 2838 64218
rect 2862 64166 2892 64218
rect 2892 64166 2918 64218
rect 2622 64164 2678 64166
rect 2702 64164 2758 64166
rect 2782 64164 2838 64166
rect 2862 64164 2918 64166
rect 2622 63130 2678 63132
rect 2702 63130 2758 63132
rect 2782 63130 2838 63132
rect 2862 63130 2918 63132
rect 2622 63078 2648 63130
rect 2648 63078 2678 63130
rect 2702 63078 2712 63130
rect 2712 63078 2758 63130
rect 2782 63078 2828 63130
rect 2828 63078 2838 63130
rect 2862 63078 2892 63130
rect 2892 63078 2918 63130
rect 2622 63076 2678 63078
rect 2702 63076 2758 63078
rect 2782 63076 2838 63078
rect 2862 63076 2918 63078
rect 2622 62042 2678 62044
rect 2702 62042 2758 62044
rect 2782 62042 2838 62044
rect 2862 62042 2918 62044
rect 2622 61990 2648 62042
rect 2648 61990 2678 62042
rect 2702 61990 2712 62042
rect 2712 61990 2758 62042
rect 2782 61990 2828 62042
rect 2828 61990 2838 62042
rect 2862 61990 2892 62042
rect 2892 61990 2918 62042
rect 2622 61988 2678 61990
rect 2702 61988 2758 61990
rect 2782 61988 2838 61990
rect 2862 61988 2918 61990
rect 2622 60954 2678 60956
rect 2702 60954 2758 60956
rect 2782 60954 2838 60956
rect 2862 60954 2918 60956
rect 2622 60902 2648 60954
rect 2648 60902 2678 60954
rect 2702 60902 2712 60954
rect 2712 60902 2758 60954
rect 2782 60902 2828 60954
rect 2828 60902 2838 60954
rect 2862 60902 2892 60954
rect 2892 60902 2918 60954
rect 2622 60900 2678 60902
rect 2702 60900 2758 60902
rect 2782 60900 2838 60902
rect 2862 60900 2918 60902
rect 2622 59866 2678 59868
rect 2702 59866 2758 59868
rect 2782 59866 2838 59868
rect 2862 59866 2918 59868
rect 2622 59814 2648 59866
rect 2648 59814 2678 59866
rect 2702 59814 2712 59866
rect 2712 59814 2758 59866
rect 2782 59814 2828 59866
rect 2828 59814 2838 59866
rect 2862 59814 2892 59866
rect 2892 59814 2918 59866
rect 2622 59812 2678 59814
rect 2702 59812 2758 59814
rect 2782 59812 2838 59814
rect 2862 59812 2918 59814
rect 2622 58778 2678 58780
rect 2702 58778 2758 58780
rect 2782 58778 2838 58780
rect 2862 58778 2918 58780
rect 2622 58726 2648 58778
rect 2648 58726 2678 58778
rect 2702 58726 2712 58778
rect 2712 58726 2758 58778
rect 2782 58726 2828 58778
rect 2828 58726 2838 58778
rect 2862 58726 2892 58778
rect 2892 58726 2918 58778
rect 2622 58724 2678 58726
rect 2702 58724 2758 58726
rect 2782 58724 2838 58726
rect 2862 58724 2918 58726
rect 2622 57690 2678 57692
rect 2702 57690 2758 57692
rect 2782 57690 2838 57692
rect 2862 57690 2918 57692
rect 2622 57638 2648 57690
rect 2648 57638 2678 57690
rect 2702 57638 2712 57690
rect 2712 57638 2758 57690
rect 2782 57638 2828 57690
rect 2828 57638 2838 57690
rect 2862 57638 2892 57690
rect 2892 57638 2918 57690
rect 2622 57636 2678 57638
rect 2702 57636 2758 57638
rect 2782 57636 2838 57638
rect 2862 57636 2918 57638
rect 2622 56602 2678 56604
rect 2702 56602 2758 56604
rect 2782 56602 2838 56604
rect 2862 56602 2918 56604
rect 2622 56550 2648 56602
rect 2648 56550 2678 56602
rect 2702 56550 2712 56602
rect 2712 56550 2758 56602
rect 2782 56550 2828 56602
rect 2828 56550 2838 56602
rect 2862 56550 2892 56602
rect 2892 56550 2918 56602
rect 2622 56548 2678 56550
rect 2702 56548 2758 56550
rect 2782 56548 2838 56550
rect 2862 56548 2918 56550
rect 2622 55514 2678 55516
rect 2702 55514 2758 55516
rect 2782 55514 2838 55516
rect 2862 55514 2918 55516
rect 2622 55462 2648 55514
rect 2648 55462 2678 55514
rect 2702 55462 2712 55514
rect 2712 55462 2758 55514
rect 2782 55462 2828 55514
rect 2828 55462 2838 55514
rect 2862 55462 2892 55514
rect 2892 55462 2918 55514
rect 2622 55460 2678 55462
rect 2702 55460 2758 55462
rect 2782 55460 2838 55462
rect 2862 55460 2918 55462
rect 2622 54426 2678 54428
rect 2702 54426 2758 54428
rect 2782 54426 2838 54428
rect 2862 54426 2918 54428
rect 2622 54374 2648 54426
rect 2648 54374 2678 54426
rect 2702 54374 2712 54426
rect 2712 54374 2758 54426
rect 2782 54374 2828 54426
rect 2828 54374 2838 54426
rect 2862 54374 2892 54426
rect 2892 54374 2918 54426
rect 2622 54372 2678 54374
rect 2702 54372 2758 54374
rect 2782 54372 2838 54374
rect 2862 54372 2918 54374
rect 2622 53338 2678 53340
rect 2702 53338 2758 53340
rect 2782 53338 2838 53340
rect 2862 53338 2918 53340
rect 2622 53286 2648 53338
rect 2648 53286 2678 53338
rect 2702 53286 2712 53338
rect 2712 53286 2758 53338
rect 2782 53286 2828 53338
rect 2828 53286 2838 53338
rect 2862 53286 2892 53338
rect 2892 53286 2918 53338
rect 2622 53284 2678 53286
rect 2702 53284 2758 53286
rect 2782 53284 2838 53286
rect 2862 53284 2918 53286
rect 2622 52250 2678 52252
rect 2702 52250 2758 52252
rect 2782 52250 2838 52252
rect 2862 52250 2918 52252
rect 2622 52198 2648 52250
rect 2648 52198 2678 52250
rect 2702 52198 2712 52250
rect 2712 52198 2758 52250
rect 2782 52198 2828 52250
rect 2828 52198 2838 52250
rect 2862 52198 2892 52250
rect 2892 52198 2918 52250
rect 2622 52196 2678 52198
rect 2702 52196 2758 52198
rect 2782 52196 2838 52198
rect 2862 52196 2918 52198
rect 2622 51162 2678 51164
rect 2702 51162 2758 51164
rect 2782 51162 2838 51164
rect 2862 51162 2918 51164
rect 2622 51110 2648 51162
rect 2648 51110 2678 51162
rect 2702 51110 2712 51162
rect 2712 51110 2758 51162
rect 2782 51110 2828 51162
rect 2828 51110 2838 51162
rect 2862 51110 2892 51162
rect 2892 51110 2918 51162
rect 2622 51108 2678 51110
rect 2702 51108 2758 51110
rect 2782 51108 2838 51110
rect 2862 51108 2918 51110
rect 2622 50074 2678 50076
rect 2702 50074 2758 50076
rect 2782 50074 2838 50076
rect 2862 50074 2918 50076
rect 2622 50022 2648 50074
rect 2648 50022 2678 50074
rect 2702 50022 2712 50074
rect 2712 50022 2758 50074
rect 2782 50022 2828 50074
rect 2828 50022 2838 50074
rect 2862 50022 2892 50074
rect 2892 50022 2918 50074
rect 2622 50020 2678 50022
rect 2702 50020 2758 50022
rect 2782 50020 2838 50022
rect 2862 50020 2918 50022
rect 2622 48986 2678 48988
rect 2702 48986 2758 48988
rect 2782 48986 2838 48988
rect 2862 48986 2918 48988
rect 2622 48934 2648 48986
rect 2648 48934 2678 48986
rect 2702 48934 2712 48986
rect 2712 48934 2758 48986
rect 2782 48934 2828 48986
rect 2828 48934 2838 48986
rect 2862 48934 2892 48986
rect 2892 48934 2918 48986
rect 2622 48932 2678 48934
rect 2702 48932 2758 48934
rect 2782 48932 2838 48934
rect 2862 48932 2918 48934
rect 2622 47898 2678 47900
rect 2702 47898 2758 47900
rect 2782 47898 2838 47900
rect 2862 47898 2918 47900
rect 2622 47846 2648 47898
rect 2648 47846 2678 47898
rect 2702 47846 2712 47898
rect 2712 47846 2758 47898
rect 2782 47846 2828 47898
rect 2828 47846 2838 47898
rect 2862 47846 2892 47898
rect 2892 47846 2918 47898
rect 2622 47844 2678 47846
rect 2702 47844 2758 47846
rect 2782 47844 2838 47846
rect 2862 47844 2918 47846
rect 2622 46810 2678 46812
rect 2702 46810 2758 46812
rect 2782 46810 2838 46812
rect 2862 46810 2918 46812
rect 2622 46758 2648 46810
rect 2648 46758 2678 46810
rect 2702 46758 2712 46810
rect 2712 46758 2758 46810
rect 2782 46758 2828 46810
rect 2828 46758 2838 46810
rect 2862 46758 2892 46810
rect 2892 46758 2918 46810
rect 2622 46756 2678 46758
rect 2702 46756 2758 46758
rect 2782 46756 2838 46758
rect 2862 46756 2918 46758
rect 2622 45722 2678 45724
rect 2702 45722 2758 45724
rect 2782 45722 2838 45724
rect 2862 45722 2918 45724
rect 2622 45670 2648 45722
rect 2648 45670 2678 45722
rect 2702 45670 2712 45722
rect 2712 45670 2758 45722
rect 2782 45670 2828 45722
rect 2828 45670 2838 45722
rect 2862 45670 2892 45722
rect 2892 45670 2918 45722
rect 2622 45668 2678 45670
rect 2702 45668 2758 45670
rect 2782 45668 2838 45670
rect 2862 45668 2918 45670
rect 2622 44634 2678 44636
rect 2702 44634 2758 44636
rect 2782 44634 2838 44636
rect 2862 44634 2918 44636
rect 2622 44582 2648 44634
rect 2648 44582 2678 44634
rect 2702 44582 2712 44634
rect 2712 44582 2758 44634
rect 2782 44582 2828 44634
rect 2828 44582 2838 44634
rect 2862 44582 2892 44634
rect 2892 44582 2918 44634
rect 2622 44580 2678 44582
rect 2702 44580 2758 44582
rect 2782 44580 2838 44582
rect 2862 44580 2918 44582
rect 2622 43546 2678 43548
rect 2702 43546 2758 43548
rect 2782 43546 2838 43548
rect 2862 43546 2918 43548
rect 2622 43494 2648 43546
rect 2648 43494 2678 43546
rect 2702 43494 2712 43546
rect 2712 43494 2758 43546
rect 2782 43494 2828 43546
rect 2828 43494 2838 43546
rect 2862 43494 2892 43546
rect 2892 43494 2918 43546
rect 2622 43492 2678 43494
rect 2702 43492 2758 43494
rect 2782 43492 2838 43494
rect 2862 43492 2918 43494
rect 2622 42458 2678 42460
rect 2702 42458 2758 42460
rect 2782 42458 2838 42460
rect 2862 42458 2918 42460
rect 2622 42406 2648 42458
rect 2648 42406 2678 42458
rect 2702 42406 2712 42458
rect 2712 42406 2758 42458
rect 2782 42406 2828 42458
rect 2828 42406 2838 42458
rect 2862 42406 2892 42458
rect 2892 42406 2918 42458
rect 2622 42404 2678 42406
rect 2702 42404 2758 42406
rect 2782 42404 2838 42406
rect 2862 42404 2918 42406
rect 2622 41370 2678 41372
rect 2702 41370 2758 41372
rect 2782 41370 2838 41372
rect 2862 41370 2918 41372
rect 2622 41318 2648 41370
rect 2648 41318 2678 41370
rect 2702 41318 2712 41370
rect 2712 41318 2758 41370
rect 2782 41318 2828 41370
rect 2828 41318 2838 41370
rect 2862 41318 2892 41370
rect 2892 41318 2918 41370
rect 2622 41316 2678 41318
rect 2702 41316 2758 41318
rect 2782 41316 2838 41318
rect 2862 41316 2918 41318
rect 2622 40282 2678 40284
rect 2702 40282 2758 40284
rect 2782 40282 2838 40284
rect 2862 40282 2918 40284
rect 2622 40230 2648 40282
rect 2648 40230 2678 40282
rect 2702 40230 2712 40282
rect 2712 40230 2758 40282
rect 2782 40230 2828 40282
rect 2828 40230 2838 40282
rect 2862 40230 2892 40282
rect 2892 40230 2918 40282
rect 2622 40228 2678 40230
rect 2702 40228 2758 40230
rect 2782 40228 2838 40230
rect 2862 40228 2918 40230
rect 2622 39194 2678 39196
rect 2702 39194 2758 39196
rect 2782 39194 2838 39196
rect 2862 39194 2918 39196
rect 2622 39142 2648 39194
rect 2648 39142 2678 39194
rect 2702 39142 2712 39194
rect 2712 39142 2758 39194
rect 2782 39142 2828 39194
rect 2828 39142 2838 39194
rect 2862 39142 2892 39194
rect 2892 39142 2918 39194
rect 2622 39140 2678 39142
rect 2702 39140 2758 39142
rect 2782 39140 2838 39142
rect 2862 39140 2918 39142
rect 2622 38106 2678 38108
rect 2702 38106 2758 38108
rect 2782 38106 2838 38108
rect 2862 38106 2918 38108
rect 2622 38054 2648 38106
rect 2648 38054 2678 38106
rect 2702 38054 2712 38106
rect 2712 38054 2758 38106
rect 2782 38054 2828 38106
rect 2828 38054 2838 38106
rect 2862 38054 2892 38106
rect 2892 38054 2918 38106
rect 2622 38052 2678 38054
rect 2702 38052 2758 38054
rect 2782 38052 2838 38054
rect 2862 38052 2918 38054
rect 2622 37018 2678 37020
rect 2702 37018 2758 37020
rect 2782 37018 2838 37020
rect 2862 37018 2918 37020
rect 2622 36966 2648 37018
rect 2648 36966 2678 37018
rect 2702 36966 2712 37018
rect 2712 36966 2758 37018
rect 2782 36966 2828 37018
rect 2828 36966 2838 37018
rect 2862 36966 2892 37018
rect 2892 36966 2918 37018
rect 2622 36964 2678 36966
rect 2702 36964 2758 36966
rect 2782 36964 2838 36966
rect 2862 36964 2918 36966
rect 2622 35930 2678 35932
rect 2702 35930 2758 35932
rect 2782 35930 2838 35932
rect 2862 35930 2918 35932
rect 2622 35878 2648 35930
rect 2648 35878 2678 35930
rect 2702 35878 2712 35930
rect 2712 35878 2758 35930
rect 2782 35878 2828 35930
rect 2828 35878 2838 35930
rect 2862 35878 2892 35930
rect 2892 35878 2918 35930
rect 2622 35876 2678 35878
rect 2702 35876 2758 35878
rect 2782 35876 2838 35878
rect 2862 35876 2918 35878
rect 2622 34842 2678 34844
rect 2702 34842 2758 34844
rect 2782 34842 2838 34844
rect 2862 34842 2918 34844
rect 2622 34790 2648 34842
rect 2648 34790 2678 34842
rect 2702 34790 2712 34842
rect 2712 34790 2758 34842
rect 2782 34790 2828 34842
rect 2828 34790 2838 34842
rect 2862 34790 2892 34842
rect 2892 34790 2918 34842
rect 2622 34788 2678 34790
rect 2702 34788 2758 34790
rect 2782 34788 2838 34790
rect 2862 34788 2918 34790
rect 2622 33754 2678 33756
rect 2702 33754 2758 33756
rect 2782 33754 2838 33756
rect 2862 33754 2918 33756
rect 2622 33702 2648 33754
rect 2648 33702 2678 33754
rect 2702 33702 2712 33754
rect 2712 33702 2758 33754
rect 2782 33702 2828 33754
rect 2828 33702 2838 33754
rect 2862 33702 2892 33754
rect 2892 33702 2918 33754
rect 2622 33700 2678 33702
rect 2702 33700 2758 33702
rect 2782 33700 2838 33702
rect 2862 33700 2918 33702
rect 2622 32666 2678 32668
rect 2702 32666 2758 32668
rect 2782 32666 2838 32668
rect 2862 32666 2918 32668
rect 2622 32614 2648 32666
rect 2648 32614 2678 32666
rect 2702 32614 2712 32666
rect 2712 32614 2758 32666
rect 2782 32614 2828 32666
rect 2828 32614 2838 32666
rect 2862 32614 2892 32666
rect 2892 32614 2918 32666
rect 2622 32612 2678 32614
rect 2702 32612 2758 32614
rect 2782 32612 2838 32614
rect 2862 32612 2918 32614
rect 2622 31578 2678 31580
rect 2702 31578 2758 31580
rect 2782 31578 2838 31580
rect 2862 31578 2918 31580
rect 2622 31526 2648 31578
rect 2648 31526 2678 31578
rect 2702 31526 2712 31578
rect 2712 31526 2758 31578
rect 2782 31526 2828 31578
rect 2828 31526 2838 31578
rect 2862 31526 2892 31578
rect 2892 31526 2918 31578
rect 2622 31524 2678 31526
rect 2702 31524 2758 31526
rect 2782 31524 2838 31526
rect 2862 31524 2918 31526
rect 2622 30490 2678 30492
rect 2702 30490 2758 30492
rect 2782 30490 2838 30492
rect 2862 30490 2918 30492
rect 2622 30438 2648 30490
rect 2648 30438 2678 30490
rect 2702 30438 2712 30490
rect 2712 30438 2758 30490
rect 2782 30438 2828 30490
rect 2828 30438 2838 30490
rect 2862 30438 2892 30490
rect 2892 30438 2918 30490
rect 2622 30436 2678 30438
rect 2702 30436 2758 30438
rect 2782 30436 2838 30438
rect 2862 30436 2918 30438
rect 2622 29402 2678 29404
rect 2702 29402 2758 29404
rect 2782 29402 2838 29404
rect 2862 29402 2918 29404
rect 2622 29350 2648 29402
rect 2648 29350 2678 29402
rect 2702 29350 2712 29402
rect 2712 29350 2758 29402
rect 2782 29350 2828 29402
rect 2828 29350 2838 29402
rect 2862 29350 2892 29402
rect 2892 29350 2918 29402
rect 2622 29348 2678 29350
rect 2702 29348 2758 29350
rect 2782 29348 2838 29350
rect 2862 29348 2918 29350
rect 2622 28314 2678 28316
rect 2702 28314 2758 28316
rect 2782 28314 2838 28316
rect 2862 28314 2918 28316
rect 2622 28262 2648 28314
rect 2648 28262 2678 28314
rect 2702 28262 2712 28314
rect 2712 28262 2758 28314
rect 2782 28262 2828 28314
rect 2828 28262 2838 28314
rect 2862 28262 2892 28314
rect 2892 28262 2918 28314
rect 2622 28260 2678 28262
rect 2702 28260 2758 28262
rect 2782 28260 2838 28262
rect 2862 28260 2918 28262
rect 2622 27226 2678 27228
rect 2702 27226 2758 27228
rect 2782 27226 2838 27228
rect 2862 27226 2918 27228
rect 2622 27174 2648 27226
rect 2648 27174 2678 27226
rect 2702 27174 2712 27226
rect 2712 27174 2758 27226
rect 2782 27174 2828 27226
rect 2828 27174 2838 27226
rect 2862 27174 2892 27226
rect 2892 27174 2918 27226
rect 2622 27172 2678 27174
rect 2702 27172 2758 27174
rect 2782 27172 2838 27174
rect 2862 27172 2918 27174
rect 2622 26138 2678 26140
rect 2702 26138 2758 26140
rect 2782 26138 2838 26140
rect 2862 26138 2918 26140
rect 2622 26086 2648 26138
rect 2648 26086 2678 26138
rect 2702 26086 2712 26138
rect 2712 26086 2758 26138
rect 2782 26086 2828 26138
rect 2828 26086 2838 26138
rect 2862 26086 2892 26138
rect 2892 26086 2918 26138
rect 2622 26084 2678 26086
rect 2702 26084 2758 26086
rect 2782 26084 2838 26086
rect 2862 26084 2918 26086
rect 2622 25050 2678 25052
rect 2702 25050 2758 25052
rect 2782 25050 2838 25052
rect 2862 25050 2918 25052
rect 2622 24998 2648 25050
rect 2648 24998 2678 25050
rect 2702 24998 2712 25050
rect 2712 24998 2758 25050
rect 2782 24998 2828 25050
rect 2828 24998 2838 25050
rect 2862 24998 2892 25050
rect 2892 24998 2918 25050
rect 2622 24996 2678 24998
rect 2702 24996 2758 24998
rect 2782 24996 2838 24998
rect 2862 24996 2918 24998
rect 2622 23962 2678 23964
rect 2702 23962 2758 23964
rect 2782 23962 2838 23964
rect 2862 23962 2918 23964
rect 2622 23910 2648 23962
rect 2648 23910 2678 23962
rect 2702 23910 2712 23962
rect 2712 23910 2758 23962
rect 2782 23910 2828 23962
rect 2828 23910 2838 23962
rect 2862 23910 2892 23962
rect 2892 23910 2918 23962
rect 2622 23908 2678 23910
rect 2702 23908 2758 23910
rect 2782 23908 2838 23910
rect 2862 23908 2918 23910
rect 2622 22874 2678 22876
rect 2702 22874 2758 22876
rect 2782 22874 2838 22876
rect 2862 22874 2918 22876
rect 2622 22822 2648 22874
rect 2648 22822 2678 22874
rect 2702 22822 2712 22874
rect 2712 22822 2758 22874
rect 2782 22822 2828 22874
rect 2828 22822 2838 22874
rect 2862 22822 2892 22874
rect 2892 22822 2918 22874
rect 2622 22820 2678 22822
rect 2702 22820 2758 22822
rect 2782 22820 2838 22822
rect 2862 22820 2918 22822
rect 2622 21786 2678 21788
rect 2702 21786 2758 21788
rect 2782 21786 2838 21788
rect 2862 21786 2918 21788
rect 2622 21734 2648 21786
rect 2648 21734 2678 21786
rect 2702 21734 2712 21786
rect 2712 21734 2758 21786
rect 2782 21734 2828 21786
rect 2828 21734 2838 21786
rect 2862 21734 2892 21786
rect 2892 21734 2918 21786
rect 2622 21732 2678 21734
rect 2702 21732 2758 21734
rect 2782 21732 2838 21734
rect 2862 21732 2918 21734
rect 2622 20698 2678 20700
rect 2702 20698 2758 20700
rect 2782 20698 2838 20700
rect 2862 20698 2918 20700
rect 2622 20646 2648 20698
rect 2648 20646 2678 20698
rect 2702 20646 2712 20698
rect 2712 20646 2758 20698
rect 2782 20646 2828 20698
rect 2828 20646 2838 20698
rect 2862 20646 2892 20698
rect 2892 20646 2918 20698
rect 2622 20644 2678 20646
rect 2702 20644 2758 20646
rect 2782 20644 2838 20646
rect 2862 20644 2918 20646
rect 2622 19610 2678 19612
rect 2702 19610 2758 19612
rect 2782 19610 2838 19612
rect 2862 19610 2918 19612
rect 2622 19558 2648 19610
rect 2648 19558 2678 19610
rect 2702 19558 2712 19610
rect 2712 19558 2758 19610
rect 2782 19558 2828 19610
rect 2828 19558 2838 19610
rect 2862 19558 2892 19610
rect 2892 19558 2918 19610
rect 2622 19556 2678 19558
rect 2702 19556 2758 19558
rect 2782 19556 2838 19558
rect 2862 19556 2918 19558
rect 2622 18522 2678 18524
rect 2702 18522 2758 18524
rect 2782 18522 2838 18524
rect 2862 18522 2918 18524
rect 2622 18470 2648 18522
rect 2648 18470 2678 18522
rect 2702 18470 2712 18522
rect 2712 18470 2758 18522
rect 2782 18470 2828 18522
rect 2828 18470 2838 18522
rect 2862 18470 2892 18522
rect 2892 18470 2918 18522
rect 2622 18468 2678 18470
rect 2702 18468 2758 18470
rect 2782 18468 2838 18470
rect 2862 18468 2918 18470
rect 2622 17434 2678 17436
rect 2702 17434 2758 17436
rect 2782 17434 2838 17436
rect 2862 17434 2918 17436
rect 2622 17382 2648 17434
rect 2648 17382 2678 17434
rect 2702 17382 2712 17434
rect 2712 17382 2758 17434
rect 2782 17382 2828 17434
rect 2828 17382 2838 17434
rect 2862 17382 2892 17434
rect 2892 17382 2918 17434
rect 2622 17380 2678 17382
rect 2702 17380 2758 17382
rect 2782 17380 2838 17382
rect 2862 17380 2918 17382
rect 2622 16346 2678 16348
rect 2702 16346 2758 16348
rect 2782 16346 2838 16348
rect 2862 16346 2918 16348
rect 2622 16294 2648 16346
rect 2648 16294 2678 16346
rect 2702 16294 2712 16346
rect 2712 16294 2758 16346
rect 2782 16294 2828 16346
rect 2828 16294 2838 16346
rect 2862 16294 2892 16346
rect 2892 16294 2918 16346
rect 2622 16292 2678 16294
rect 2702 16292 2758 16294
rect 2782 16292 2838 16294
rect 2862 16292 2918 16294
rect 2622 15258 2678 15260
rect 2702 15258 2758 15260
rect 2782 15258 2838 15260
rect 2862 15258 2918 15260
rect 2622 15206 2648 15258
rect 2648 15206 2678 15258
rect 2702 15206 2712 15258
rect 2712 15206 2758 15258
rect 2782 15206 2828 15258
rect 2828 15206 2838 15258
rect 2862 15206 2892 15258
rect 2892 15206 2918 15258
rect 2622 15204 2678 15206
rect 2702 15204 2758 15206
rect 2782 15204 2838 15206
rect 2862 15204 2918 15206
rect 2622 14170 2678 14172
rect 2702 14170 2758 14172
rect 2782 14170 2838 14172
rect 2862 14170 2918 14172
rect 2622 14118 2648 14170
rect 2648 14118 2678 14170
rect 2702 14118 2712 14170
rect 2712 14118 2758 14170
rect 2782 14118 2828 14170
rect 2828 14118 2838 14170
rect 2862 14118 2892 14170
rect 2892 14118 2918 14170
rect 2622 14116 2678 14118
rect 2702 14116 2758 14118
rect 2782 14116 2838 14118
rect 2862 14116 2918 14118
rect 2622 13082 2678 13084
rect 2702 13082 2758 13084
rect 2782 13082 2838 13084
rect 2862 13082 2918 13084
rect 2622 13030 2648 13082
rect 2648 13030 2678 13082
rect 2702 13030 2712 13082
rect 2712 13030 2758 13082
rect 2782 13030 2828 13082
rect 2828 13030 2838 13082
rect 2862 13030 2892 13082
rect 2892 13030 2918 13082
rect 2622 13028 2678 13030
rect 2702 13028 2758 13030
rect 2782 13028 2838 13030
rect 2862 13028 2918 13030
rect 2622 11994 2678 11996
rect 2702 11994 2758 11996
rect 2782 11994 2838 11996
rect 2862 11994 2918 11996
rect 2622 11942 2648 11994
rect 2648 11942 2678 11994
rect 2702 11942 2712 11994
rect 2712 11942 2758 11994
rect 2782 11942 2828 11994
rect 2828 11942 2838 11994
rect 2862 11942 2892 11994
rect 2892 11942 2918 11994
rect 2622 11940 2678 11942
rect 2702 11940 2758 11942
rect 2782 11940 2838 11942
rect 2862 11940 2918 11942
rect 2622 10906 2678 10908
rect 2702 10906 2758 10908
rect 2782 10906 2838 10908
rect 2862 10906 2918 10908
rect 2622 10854 2648 10906
rect 2648 10854 2678 10906
rect 2702 10854 2712 10906
rect 2712 10854 2758 10906
rect 2782 10854 2828 10906
rect 2828 10854 2838 10906
rect 2862 10854 2892 10906
rect 2892 10854 2918 10906
rect 2622 10852 2678 10854
rect 2702 10852 2758 10854
rect 2782 10852 2838 10854
rect 2862 10852 2918 10854
rect 2622 9818 2678 9820
rect 2702 9818 2758 9820
rect 2782 9818 2838 9820
rect 2862 9818 2918 9820
rect 2622 9766 2648 9818
rect 2648 9766 2678 9818
rect 2702 9766 2712 9818
rect 2712 9766 2758 9818
rect 2782 9766 2828 9818
rect 2828 9766 2838 9818
rect 2862 9766 2892 9818
rect 2892 9766 2918 9818
rect 2622 9764 2678 9766
rect 2702 9764 2758 9766
rect 2782 9764 2838 9766
rect 2862 9764 2918 9766
rect 2622 8730 2678 8732
rect 2702 8730 2758 8732
rect 2782 8730 2838 8732
rect 2862 8730 2918 8732
rect 2622 8678 2648 8730
rect 2648 8678 2678 8730
rect 2702 8678 2712 8730
rect 2712 8678 2758 8730
rect 2782 8678 2828 8730
rect 2828 8678 2838 8730
rect 2862 8678 2892 8730
rect 2892 8678 2918 8730
rect 2622 8676 2678 8678
rect 2702 8676 2758 8678
rect 2782 8676 2838 8678
rect 2862 8676 2918 8678
rect 2622 7642 2678 7644
rect 2702 7642 2758 7644
rect 2782 7642 2838 7644
rect 2862 7642 2918 7644
rect 2622 7590 2648 7642
rect 2648 7590 2678 7642
rect 2702 7590 2712 7642
rect 2712 7590 2758 7642
rect 2782 7590 2828 7642
rect 2828 7590 2838 7642
rect 2862 7590 2892 7642
rect 2892 7590 2918 7642
rect 2622 7588 2678 7590
rect 2702 7588 2758 7590
rect 2782 7588 2838 7590
rect 2862 7588 2918 7590
rect 2622 6554 2678 6556
rect 2702 6554 2758 6556
rect 2782 6554 2838 6556
rect 2862 6554 2918 6556
rect 2622 6502 2648 6554
rect 2648 6502 2678 6554
rect 2702 6502 2712 6554
rect 2712 6502 2758 6554
rect 2782 6502 2828 6554
rect 2828 6502 2838 6554
rect 2862 6502 2892 6554
rect 2892 6502 2918 6554
rect 2622 6500 2678 6502
rect 2702 6500 2758 6502
rect 2782 6500 2838 6502
rect 2862 6500 2918 6502
rect 2622 5466 2678 5468
rect 2702 5466 2758 5468
rect 2782 5466 2838 5468
rect 2862 5466 2918 5468
rect 2622 5414 2648 5466
rect 2648 5414 2678 5466
rect 2702 5414 2712 5466
rect 2712 5414 2758 5466
rect 2782 5414 2828 5466
rect 2828 5414 2838 5466
rect 2862 5414 2892 5466
rect 2892 5414 2918 5466
rect 2622 5412 2678 5414
rect 2702 5412 2758 5414
rect 2782 5412 2838 5414
rect 2862 5412 2918 5414
rect 2622 4378 2678 4380
rect 2702 4378 2758 4380
rect 2782 4378 2838 4380
rect 2862 4378 2918 4380
rect 2622 4326 2648 4378
rect 2648 4326 2678 4378
rect 2702 4326 2712 4378
rect 2712 4326 2758 4378
rect 2782 4326 2828 4378
rect 2828 4326 2838 4378
rect 2862 4326 2892 4378
rect 2892 4326 2918 4378
rect 2622 4324 2678 4326
rect 2702 4324 2758 4326
rect 2782 4324 2838 4326
rect 2862 4324 2918 4326
rect 2622 3290 2678 3292
rect 2702 3290 2758 3292
rect 2782 3290 2838 3292
rect 2862 3290 2918 3292
rect 2622 3238 2648 3290
rect 2648 3238 2678 3290
rect 2702 3238 2712 3290
rect 2712 3238 2758 3290
rect 2782 3238 2828 3290
rect 2828 3238 2838 3290
rect 2862 3238 2892 3290
rect 2892 3238 2918 3290
rect 2622 3236 2678 3238
rect 2702 3236 2758 3238
rect 2782 3236 2838 3238
rect 2862 3236 2918 3238
rect 2622 2202 2678 2204
rect 2702 2202 2758 2204
rect 2782 2202 2838 2204
rect 2862 2202 2918 2204
rect 2622 2150 2648 2202
rect 2648 2150 2678 2202
rect 2702 2150 2712 2202
rect 2712 2150 2758 2202
rect 2782 2150 2828 2202
rect 2828 2150 2838 2202
rect 2862 2150 2892 2202
rect 2892 2150 2918 2202
rect 2622 2148 2678 2150
rect 2702 2148 2758 2150
rect 2782 2148 2838 2150
rect 2862 2148 2918 2150
rect 3422 165824 3478 165880
rect 3514 150320 3570 150376
rect 4289 330234 4345 330236
rect 4369 330234 4425 330236
rect 4449 330234 4505 330236
rect 4529 330234 4585 330236
rect 4289 330182 4315 330234
rect 4315 330182 4345 330234
rect 4369 330182 4379 330234
rect 4379 330182 4425 330234
rect 4449 330182 4495 330234
rect 4495 330182 4505 330234
rect 4529 330182 4559 330234
rect 4559 330182 4585 330234
rect 4289 330180 4345 330182
rect 4369 330180 4425 330182
rect 4449 330180 4505 330182
rect 4529 330180 4585 330182
rect 4289 329146 4345 329148
rect 4369 329146 4425 329148
rect 4449 329146 4505 329148
rect 4529 329146 4585 329148
rect 4289 329094 4315 329146
rect 4315 329094 4345 329146
rect 4369 329094 4379 329146
rect 4379 329094 4425 329146
rect 4449 329094 4495 329146
rect 4495 329094 4505 329146
rect 4529 329094 4559 329146
rect 4559 329094 4585 329146
rect 4289 329092 4345 329094
rect 4369 329092 4425 329094
rect 4449 329092 4505 329094
rect 4529 329092 4585 329094
rect 4289 328058 4345 328060
rect 4369 328058 4425 328060
rect 4449 328058 4505 328060
rect 4529 328058 4585 328060
rect 4289 328006 4315 328058
rect 4315 328006 4345 328058
rect 4369 328006 4379 328058
rect 4379 328006 4425 328058
rect 4449 328006 4495 328058
rect 4495 328006 4505 328058
rect 4529 328006 4559 328058
rect 4559 328006 4585 328058
rect 4289 328004 4345 328006
rect 4369 328004 4425 328006
rect 4449 328004 4505 328006
rect 4529 328004 4585 328006
rect 4289 326970 4345 326972
rect 4369 326970 4425 326972
rect 4449 326970 4505 326972
rect 4529 326970 4585 326972
rect 4289 326918 4315 326970
rect 4315 326918 4345 326970
rect 4369 326918 4379 326970
rect 4379 326918 4425 326970
rect 4449 326918 4495 326970
rect 4495 326918 4505 326970
rect 4529 326918 4559 326970
rect 4559 326918 4585 326970
rect 4289 326916 4345 326918
rect 4369 326916 4425 326918
rect 4449 326916 4505 326918
rect 4529 326916 4585 326918
rect 4289 325882 4345 325884
rect 4369 325882 4425 325884
rect 4449 325882 4505 325884
rect 4529 325882 4585 325884
rect 4289 325830 4315 325882
rect 4315 325830 4345 325882
rect 4369 325830 4379 325882
rect 4379 325830 4425 325882
rect 4449 325830 4495 325882
rect 4495 325830 4505 325882
rect 4529 325830 4559 325882
rect 4559 325830 4585 325882
rect 4289 325828 4345 325830
rect 4369 325828 4425 325830
rect 4449 325828 4505 325830
rect 4529 325828 4585 325830
rect 4289 324794 4345 324796
rect 4369 324794 4425 324796
rect 4449 324794 4505 324796
rect 4529 324794 4585 324796
rect 4289 324742 4315 324794
rect 4315 324742 4345 324794
rect 4369 324742 4379 324794
rect 4379 324742 4425 324794
rect 4449 324742 4495 324794
rect 4495 324742 4505 324794
rect 4529 324742 4559 324794
rect 4559 324742 4585 324794
rect 4289 324740 4345 324742
rect 4369 324740 4425 324742
rect 4449 324740 4505 324742
rect 4529 324740 4585 324742
rect 4289 323706 4345 323708
rect 4369 323706 4425 323708
rect 4449 323706 4505 323708
rect 4529 323706 4585 323708
rect 4289 323654 4315 323706
rect 4315 323654 4345 323706
rect 4369 323654 4379 323706
rect 4379 323654 4425 323706
rect 4449 323654 4495 323706
rect 4495 323654 4505 323706
rect 4529 323654 4559 323706
rect 4559 323654 4585 323706
rect 4289 323652 4345 323654
rect 4369 323652 4425 323654
rect 4449 323652 4505 323654
rect 4529 323652 4585 323654
rect 4289 322618 4345 322620
rect 4369 322618 4425 322620
rect 4449 322618 4505 322620
rect 4529 322618 4585 322620
rect 4289 322566 4315 322618
rect 4315 322566 4345 322618
rect 4369 322566 4379 322618
rect 4379 322566 4425 322618
rect 4449 322566 4495 322618
rect 4495 322566 4505 322618
rect 4529 322566 4559 322618
rect 4559 322566 4585 322618
rect 4289 322564 4345 322566
rect 4369 322564 4425 322566
rect 4449 322564 4505 322566
rect 4529 322564 4585 322566
rect 4289 321530 4345 321532
rect 4369 321530 4425 321532
rect 4449 321530 4505 321532
rect 4529 321530 4585 321532
rect 4289 321478 4315 321530
rect 4315 321478 4345 321530
rect 4369 321478 4379 321530
rect 4379 321478 4425 321530
rect 4449 321478 4495 321530
rect 4495 321478 4505 321530
rect 4529 321478 4559 321530
rect 4559 321478 4585 321530
rect 4289 321476 4345 321478
rect 4369 321476 4425 321478
rect 4449 321476 4505 321478
rect 4529 321476 4585 321478
rect 4289 320442 4345 320444
rect 4369 320442 4425 320444
rect 4449 320442 4505 320444
rect 4529 320442 4585 320444
rect 4289 320390 4315 320442
rect 4315 320390 4345 320442
rect 4369 320390 4379 320442
rect 4379 320390 4425 320442
rect 4449 320390 4495 320442
rect 4495 320390 4505 320442
rect 4529 320390 4559 320442
rect 4559 320390 4585 320442
rect 4289 320388 4345 320390
rect 4369 320388 4425 320390
rect 4449 320388 4505 320390
rect 4529 320388 4585 320390
rect 4289 319354 4345 319356
rect 4369 319354 4425 319356
rect 4449 319354 4505 319356
rect 4529 319354 4585 319356
rect 4289 319302 4315 319354
rect 4315 319302 4345 319354
rect 4369 319302 4379 319354
rect 4379 319302 4425 319354
rect 4449 319302 4495 319354
rect 4495 319302 4505 319354
rect 4529 319302 4559 319354
rect 4559 319302 4585 319354
rect 4289 319300 4345 319302
rect 4369 319300 4425 319302
rect 4449 319300 4505 319302
rect 4529 319300 4585 319302
rect 4289 318266 4345 318268
rect 4369 318266 4425 318268
rect 4449 318266 4505 318268
rect 4529 318266 4585 318268
rect 4289 318214 4315 318266
rect 4315 318214 4345 318266
rect 4369 318214 4379 318266
rect 4379 318214 4425 318266
rect 4449 318214 4495 318266
rect 4495 318214 4505 318266
rect 4529 318214 4559 318266
rect 4559 318214 4585 318266
rect 4289 318212 4345 318214
rect 4369 318212 4425 318214
rect 4449 318212 4505 318214
rect 4529 318212 4585 318214
rect 4289 317178 4345 317180
rect 4369 317178 4425 317180
rect 4449 317178 4505 317180
rect 4529 317178 4585 317180
rect 4289 317126 4315 317178
rect 4315 317126 4345 317178
rect 4369 317126 4379 317178
rect 4379 317126 4425 317178
rect 4449 317126 4495 317178
rect 4495 317126 4505 317178
rect 4529 317126 4559 317178
rect 4559 317126 4585 317178
rect 4289 317124 4345 317126
rect 4369 317124 4425 317126
rect 4449 317124 4505 317126
rect 4529 317124 4585 317126
rect 4289 316090 4345 316092
rect 4369 316090 4425 316092
rect 4449 316090 4505 316092
rect 4529 316090 4585 316092
rect 4289 316038 4315 316090
rect 4315 316038 4345 316090
rect 4369 316038 4379 316090
rect 4379 316038 4425 316090
rect 4449 316038 4495 316090
rect 4495 316038 4505 316090
rect 4529 316038 4559 316090
rect 4559 316038 4585 316090
rect 4289 316036 4345 316038
rect 4369 316036 4425 316038
rect 4449 316036 4505 316038
rect 4529 316036 4585 316038
rect 4289 315002 4345 315004
rect 4369 315002 4425 315004
rect 4449 315002 4505 315004
rect 4529 315002 4585 315004
rect 4289 314950 4315 315002
rect 4315 314950 4345 315002
rect 4369 314950 4379 315002
rect 4379 314950 4425 315002
rect 4449 314950 4495 315002
rect 4495 314950 4505 315002
rect 4529 314950 4559 315002
rect 4559 314950 4585 315002
rect 4289 314948 4345 314950
rect 4369 314948 4425 314950
rect 4449 314948 4505 314950
rect 4529 314948 4585 314950
rect 4289 313914 4345 313916
rect 4369 313914 4425 313916
rect 4449 313914 4505 313916
rect 4529 313914 4585 313916
rect 4289 313862 4315 313914
rect 4315 313862 4345 313914
rect 4369 313862 4379 313914
rect 4379 313862 4425 313914
rect 4449 313862 4495 313914
rect 4495 313862 4505 313914
rect 4529 313862 4559 313914
rect 4559 313862 4585 313914
rect 4289 313860 4345 313862
rect 4369 313860 4425 313862
rect 4449 313860 4505 313862
rect 4529 313860 4585 313862
rect 4289 312826 4345 312828
rect 4369 312826 4425 312828
rect 4449 312826 4505 312828
rect 4529 312826 4585 312828
rect 4289 312774 4315 312826
rect 4315 312774 4345 312826
rect 4369 312774 4379 312826
rect 4379 312774 4425 312826
rect 4449 312774 4495 312826
rect 4495 312774 4505 312826
rect 4529 312774 4559 312826
rect 4559 312774 4585 312826
rect 4289 312772 4345 312774
rect 4369 312772 4425 312774
rect 4449 312772 4505 312774
rect 4529 312772 4585 312774
rect 4289 311738 4345 311740
rect 4369 311738 4425 311740
rect 4449 311738 4505 311740
rect 4529 311738 4585 311740
rect 4289 311686 4315 311738
rect 4315 311686 4345 311738
rect 4369 311686 4379 311738
rect 4379 311686 4425 311738
rect 4449 311686 4495 311738
rect 4495 311686 4505 311738
rect 4529 311686 4559 311738
rect 4559 311686 4585 311738
rect 4289 311684 4345 311686
rect 4369 311684 4425 311686
rect 4449 311684 4505 311686
rect 4529 311684 4585 311686
rect 4289 310650 4345 310652
rect 4369 310650 4425 310652
rect 4449 310650 4505 310652
rect 4529 310650 4585 310652
rect 4289 310598 4315 310650
rect 4315 310598 4345 310650
rect 4369 310598 4379 310650
rect 4379 310598 4425 310650
rect 4449 310598 4495 310650
rect 4495 310598 4505 310650
rect 4529 310598 4559 310650
rect 4559 310598 4585 310650
rect 4289 310596 4345 310598
rect 4369 310596 4425 310598
rect 4449 310596 4505 310598
rect 4529 310596 4585 310598
rect 4289 309562 4345 309564
rect 4369 309562 4425 309564
rect 4449 309562 4505 309564
rect 4529 309562 4585 309564
rect 4289 309510 4315 309562
rect 4315 309510 4345 309562
rect 4369 309510 4379 309562
rect 4379 309510 4425 309562
rect 4449 309510 4495 309562
rect 4495 309510 4505 309562
rect 4529 309510 4559 309562
rect 4559 309510 4585 309562
rect 4289 309508 4345 309510
rect 4369 309508 4425 309510
rect 4449 309508 4505 309510
rect 4529 309508 4585 309510
rect 4289 308474 4345 308476
rect 4369 308474 4425 308476
rect 4449 308474 4505 308476
rect 4529 308474 4585 308476
rect 4289 308422 4315 308474
rect 4315 308422 4345 308474
rect 4369 308422 4379 308474
rect 4379 308422 4425 308474
rect 4449 308422 4495 308474
rect 4495 308422 4505 308474
rect 4529 308422 4559 308474
rect 4559 308422 4585 308474
rect 4289 308420 4345 308422
rect 4369 308420 4425 308422
rect 4449 308420 4505 308422
rect 4529 308420 4585 308422
rect 4289 307386 4345 307388
rect 4369 307386 4425 307388
rect 4449 307386 4505 307388
rect 4529 307386 4585 307388
rect 4289 307334 4315 307386
rect 4315 307334 4345 307386
rect 4369 307334 4379 307386
rect 4379 307334 4425 307386
rect 4449 307334 4495 307386
rect 4495 307334 4505 307386
rect 4529 307334 4559 307386
rect 4559 307334 4585 307386
rect 4289 307332 4345 307334
rect 4369 307332 4425 307334
rect 4449 307332 4505 307334
rect 4529 307332 4585 307334
rect 4289 306298 4345 306300
rect 4369 306298 4425 306300
rect 4449 306298 4505 306300
rect 4529 306298 4585 306300
rect 4289 306246 4315 306298
rect 4315 306246 4345 306298
rect 4369 306246 4379 306298
rect 4379 306246 4425 306298
rect 4449 306246 4495 306298
rect 4495 306246 4505 306298
rect 4529 306246 4559 306298
rect 4559 306246 4585 306298
rect 4289 306244 4345 306246
rect 4369 306244 4425 306246
rect 4449 306244 4505 306246
rect 4529 306244 4585 306246
rect 4289 305210 4345 305212
rect 4369 305210 4425 305212
rect 4449 305210 4505 305212
rect 4529 305210 4585 305212
rect 4289 305158 4315 305210
rect 4315 305158 4345 305210
rect 4369 305158 4379 305210
rect 4379 305158 4425 305210
rect 4449 305158 4495 305210
rect 4495 305158 4505 305210
rect 4529 305158 4559 305210
rect 4559 305158 4585 305210
rect 4289 305156 4345 305158
rect 4369 305156 4425 305158
rect 4449 305156 4505 305158
rect 4529 305156 4585 305158
rect 4289 304122 4345 304124
rect 4369 304122 4425 304124
rect 4449 304122 4505 304124
rect 4529 304122 4585 304124
rect 4289 304070 4315 304122
rect 4315 304070 4345 304122
rect 4369 304070 4379 304122
rect 4379 304070 4425 304122
rect 4449 304070 4495 304122
rect 4495 304070 4505 304122
rect 4529 304070 4559 304122
rect 4559 304070 4585 304122
rect 4289 304068 4345 304070
rect 4369 304068 4425 304070
rect 4449 304068 4505 304070
rect 4529 304068 4585 304070
rect 4289 303034 4345 303036
rect 4369 303034 4425 303036
rect 4449 303034 4505 303036
rect 4529 303034 4585 303036
rect 4289 302982 4315 303034
rect 4315 302982 4345 303034
rect 4369 302982 4379 303034
rect 4379 302982 4425 303034
rect 4449 302982 4495 303034
rect 4495 302982 4505 303034
rect 4529 302982 4559 303034
rect 4559 302982 4585 303034
rect 4289 302980 4345 302982
rect 4369 302980 4425 302982
rect 4449 302980 4505 302982
rect 4529 302980 4585 302982
rect 4289 301946 4345 301948
rect 4369 301946 4425 301948
rect 4449 301946 4505 301948
rect 4529 301946 4585 301948
rect 4289 301894 4315 301946
rect 4315 301894 4345 301946
rect 4369 301894 4379 301946
rect 4379 301894 4425 301946
rect 4449 301894 4495 301946
rect 4495 301894 4505 301946
rect 4529 301894 4559 301946
rect 4559 301894 4585 301946
rect 4289 301892 4345 301894
rect 4369 301892 4425 301894
rect 4449 301892 4505 301894
rect 4529 301892 4585 301894
rect 4289 300858 4345 300860
rect 4369 300858 4425 300860
rect 4449 300858 4505 300860
rect 4529 300858 4585 300860
rect 4289 300806 4315 300858
rect 4315 300806 4345 300858
rect 4369 300806 4379 300858
rect 4379 300806 4425 300858
rect 4449 300806 4495 300858
rect 4495 300806 4505 300858
rect 4529 300806 4559 300858
rect 4559 300806 4585 300858
rect 4289 300804 4345 300806
rect 4369 300804 4425 300806
rect 4449 300804 4505 300806
rect 4529 300804 4585 300806
rect 4289 299770 4345 299772
rect 4369 299770 4425 299772
rect 4449 299770 4505 299772
rect 4529 299770 4585 299772
rect 4289 299718 4315 299770
rect 4315 299718 4345 299770
rect 4369 299718 4379 299770
rect 4379 299718 4425 299770
rect 4449 299718 4495 299770
rect 4495 299718 4505 299770
rect 4529 299718 4559 299770
rect 4559 299718 4585 299770
rect 4289 299716 4345 299718
rect 4369 299716 4425 299718
rect 4449 299716 4505 299718
rect 4529 299716 4585 299718
rect 4289 298682 4345 298684
rect 4369 298682 4425 298684
rect 4449 298682 4505 298684
rect 4529 298682 4585 298684
rect 4289 298630 4315 298682
rect 4315 298630 4345 298682
rect 4369 298630 4379 298682
rect 4379 298630 4425 298682
rect 4449 298630 4495 298682
rect 4495 298630 4505 298682
rect 4529 298630 4559 298682
rect 4559 298630 4585 298682
rect 4289 298628 4345 298630
rect 4369 298628 4425 298630
rect 4449 298628 4505 298630
rect 4529 298628 4585 298630
rect 4289 297594 4345 297596
rect 4369 297594 4425 297596
rect 4449 297594 4505 297596
rect 4529 297594 4585 297596
rect 4289 297542 4315 297594
rect 4315 297542 4345 297594
rect 4369 297542 4379 297594
rect 4379 297542 4425 297594
rect 4449 297542 4495 297594
rect 4495 297542 4505 297594
rect 4529 297542 4559 297594
rect 4559 297542 4585 297594
rect 4289 297540 4345 297542
rect 4369 297540 4425 297542
rect 4449 297540 4505 297542
rect 4529 297540 4585 297542
rect 4289 296506 4345 296508
rect 4369 296506 4425 296508
rect 4449 296506 4505 296508
rect 4529 296506 4585 296508
rect 4289 296454 4315 296506
rect 4315 296454 4345 296506
rect 4369 296454 4379 296506
rect 4379 296454 4425 296506
rect 4449 296454 4495 296506
rect 4495 296454 4505 296506
rect 4529 296454 4559 296506
rect 4559 296454 4585 296506
rect 4289 296452 4345 296454
rect 4369 296452 4425 296454
rect 4449 296452 4505 296454
rect 4529 296452 4585 296454
rect 4289 295418 4345 295420
rect 4369 295418 4425 295420
rect 4449 295418 4505 295420
rect 4529 295418 4585 295420
rect 4289 295366 4315 295418
rect 4315 295366 4345 295418
rect 4369 295366 4379 295418
rect 4379 295366 4425 295418
rect 4449 295366 4495 295418
rect 4495 295366 4505 295418
rect 4529 295366 4559 295418
rect 4559 295366 4585 295418
rect 4289 295364 4345 295366
rect 4369 295364 4425 295366
rect 4449 295364 4505 295366
rect 4529 295364 4585 295366
rect 4289 294330 4345 294332
rect 4369 294330 4425 294332
rect 4449 294330 4505 294332
rect 4529 294330 4585 294332
rect 4289 294278 4315 294330
rect 4315 294278 4345 294330
rect 4369 294278 4379 294330
rect 4379 294278 4425 294330
rect 4449 294278 4495 294330
rect 4495 294278 4505 294330
rect 4529 294278 4559 294330
rect 4559 294278 4585 294330
rect 4289 294276 4345 294278
rect 4369 294276 4425 294278
rect 4449 294276 4505 294278
rect 4529 294276 4585 294278
rect 4289 293242 4345 293244
rect 4369 293242 4425 293244
rect 4449 293242 4505 293244
rect 4529 293242 4585 293244
rect 4289 293190 4315 293242
rect 4315 293190 4345 293242
rect 4369 293190 4379 293242
rect 4379 293190 4425 293242
rect 4449 293190 4495 293242
rect 4495 293190 4505 293242
rect 4529 293190 4559 293242
rect 4559 293190 4585 293242
rect 4289 293188 4345 293190
rect 4369 293188 4425 293190
rect 4449 293188 4505 293190
rect 4529 293188 4585 293190
rect 4289 292154 4345 292156
rect 4369 292154 4425 292156
rect 4449 292154 4505 292156
rect 4529 292154 4585 292156
rect 4289 292102 4315 292154
rect 4315 292102 4345 292154
rect 4369 292102 4379 292154
rect 4379 292102 4425 292154
rect 4449 292102 4495 292154
rect 4495 292102 4505 292154
rect 4529 292102 4559 292154
rect 4559 292102 4585 292154
rect 4289 292100 4345 292102
rect 4369 292100 4425 292102
rect 4449 292100 4505 292102
rect 4529 292100 4585 292102
rect 4289 291066 4345 291068
rect 4369 291066 4425 291068
rect 4449 291066 4505 291068
rect 4529 291066 4585 291068
rect 4289 291014 4315 291066
rect 4315 291014 4345 291066
rect 4369 291014 4379 291066
rect 4379 291014 4425 291066
rect 4449 291014 4495 291066
rect 4495 291014 4505 291066
rect 4529 291014 4559 291066
rect 4559 291014 4585 291066
rect 4289 291012 4345 291014
rect 4369 291012 4425 291014
rect 4449 291012 4505 291014
rect 4529 291012 4585 291014
rect 4289 289978 4345 289980
rect 4369 289978 4425 289980
rect 4449 289978 4505 289980
rect 4529 289978 4585 289980
rect 4289 289926 4315 289978
rect 4315 289926 4345 289978
rect 4369 289926 4379 289978
rect 4379 289926 4425 289978
rect 4449 289926 4495 289978
rect 4495 289926 4505 289978
rect 4529 289926 4559 289978
rect 4559 289926 4585 289978
rect 4289 289924 4345 289926
rect 4369 289924 4425 289926
rect 4449 289924 4505 289926
rect 4529 289924 4585 289926
rect 4289 288890 4345 288892
rect 4369 288890 4425 288892
rect 4449 288890 4505 288892
rect 4529 288890 4585 288892
rect 4289 288838 4315 288890
rect 4315 288838 4345 288890
rect 4369 288838 4379 288890
rect 4379 288838 4425 288890
rect 4449 288838 4495 288890
rect 4495 288838 4505 288890
rect 4529 288838 4559 288890
rect 4559 288838 4585 288890
rect 4289 288836 4345 288838
rect 4369 288836 4425 288838
rect 4449 288836 4505 288838
rect 4529 288836 4585 288838
rect 4289 287802 4345 287804
rect 4369 287802 4425 287804
rect 4449 287802 4505 287804
rect 4529 287802 4585 287804
rect 4289 287750 4315 287802
rect 4315 287750 4345 287802
rect 4369 287750 4379 287802
rect 4379 287750 4425 287802
rect 4449 287750 4495 287802
rect 4495 287750 4505 287802
rect 4529 287750 4559 287802
rect 4559 287750 4585 287802
rect 4289 287748 4345 287750
rect 4369 287748 4425 287750
rect 4449 287748 4505 287750
rect 4529 287748 4585 287750
rect 4289 286714 4345 286716
rect 4369 286714 4425 286716
rect 4449 286714 4505 286716
rect 4529 286714 4585 286716
rect 4289 286662 4315 286714
rect 4315 286662 4345 286714
rect 4369 286662 4379 286714
rect 4379 286662 4425 286714
rect 4449 286662 4495 286714
rect 4495 286662 4505 286714
rect 4529 286662 4559 286714
rect 4559 286662 4585 286714
rect 4289 286660 4345 286662
rect 4369 286660 4425 286662
rect 4449 286660 4505 286662
rect 4529 286660 4585 286662
rect 4289 285626 4345 285628
rect 4369 285626 4425 285628
rect 4449 285626 4505 285628
rect 4529 285626 4585 285628
rect 4289 285574 4315 285626
rect 4315 285574 4345 285626
rect 4369 285574 4379 285626
rect 4379 285574 4425 285626
rect 4449 285574 4495 285626
rect 4495 285574 4505 285626
rect 4529 285574 4559 285626
rect 4559 285574 4585 285626
rect 4289 285572 4345 285574
rect 4369 285572 4425 285574
rect 4449 285572 4505 285574
rect 4529 285572 4585 285574
rect 4289 284538 4345 284540
rect 4369 284538 4425 284540
rect 4449 284538 4505 284540
rect 4529 284538 4585 284540
rect 4289 284486 4315 284538
rect 4315 284486 4345 284538
rect 4369 284486 4379 284538
rect 4379 284486 4425 284538
rect 4449 284486 4495 284538
rect 4495 284486 4505 284538
rect 4529 284486 4559 284538
rect 4559 284486 4585 284538
rect 4289 284484 4345 284486
rect 4369 284484 4425 284486
rect 4449 284484 4505 284486
rect 4529 284484 4585 284486
rect 4289 283450 4345 283452
rect 4369 283450 4425 283452
rect 4449 283450 4505 283452
rect 4529 283450 4585 283452
rect 4289 283398 4315 283450
rect 4315 283398 4345 283450
rect 4369 283398 4379 283450
rect 4379 283398 4425 283450
rect 4449 283398 4495 283450
rect 4495 283398 4505 283450
rect 4529 283398 4559 283450
rect 4559 283398 4585 283450
rect 4289 283396 4345 283398
rect 4369 283396 4425 283398
rect 4449 283396 4505 283398
rect 4529 283396 4585 283398
rect 4289 282362 4345 282364
rect 4369 282362 4425 282364
rect 4449 282362 4505 282364
rect 4529 282362 4585 282364
rect 4289 282310 4315 282362
rect 4315 282310 4345 282362
rect 4369 282310 4379 282362
rect 4379 282310 4425 282362
rect 4449 282310 4495 282362
rect 4495 282310 4505 282362
rect 4529 282310 4559 282362
rect 4559 282310 4585 282362
rect 4289 282308 4345 282310
rect 4369 282308 4425 282310
rect 4449 282308 4505 282310
rect 4529 282308 4585 282310
rect 4289 281274 4345 281276
rect 4369 281274 4425 281276
rect 4449 281274 4505 281276
rect 4529 281274 4585 281276
rect 4289 281222 4315 281274
rect 4315 281222 4345 281274
rect 4369 281222 4379 281274
rect 4379 281222 4425 281274
rect 4449 281222 4495 281274
rect 4495 281222 4505 281274
rect 4529 281222 4559 281274
rect 4559 281222 4585 281274
rect 4289 281220 4345 281222
rect 4369 281220 4425 281222
rect 4449 281220 4505 281222
rect 4529 281220 4585 281222
rect 4289 280186 4345 280188
rect 4369 280186 4425 280188
rect 4449 280186 4505 280188
rect 4529 280186 4585 280188
rect 4289 280134 4315 280186
rect 4315 280134 4345 280186
rect 4369 280134 4379 280186
rect 4379 280134 4425 280186
rect 4449 280134 4495 280186
rect 4495 280134 4505 280186
rect 4529 280134 4559 280186
rect 4559 280134 4585 280186
rect 4289 280132 4345 280134
rect 4369 280132 4425 280134
rect 4449 280132 4505 280134
rect 4529 280132 4585 280134
rect 4289 279098 4345 279100
rect 4369 279098 4425 279100
rect 4449 279098 4505 279100
rect 4529 279098 4585 279100
rect 4289 279046 4315 279098
rect 4315 279046 4345 279098
rect 4369 279046 4379 279098
rect 4379 279046 4425 279098
rect 4449 279046 4495 279098
rect 4495 279046 4505 279098
rect 4529 279046 4559 279098
rect 4559 279046 4585 279098
rect 4289 279044 4345 279046
rect 4369 279044 4425 279046
rect 4449 279044 4505 279046
rect 4529 279044 4585 279046
rect 4289 278010 4345 278012
rect 4369 278010 4425 278012
rect 4449 278010 4505 278012
rect 4529 278010 4585 278012
rect 4289 277958 4315 278010
rect 4315 277958 4345 278010
rect 4369 277958 4379 278010
rect 4379 277958 4425 278010
rect 4449 277958 4495 278010
rect 4495 277958 4505 278010
rect 4529 277958 4559 278010
rect 4559 277958 4585 278010
rect 4289 277956 4345 277958
rect 4369 277956 4425 277958
rect 4449 277956 4505 277958
rect 4529 277956 4585 277958
rect 4289 276922 4345 276924
rect 4369 276922 4425 276924
rect 4449 276922 4505 276924
rect 4529 276922 4585 276924
rect 4289 276870 4315 276922
rect 4315 276870 4345 276922
rect 4369 276870 4379 276922
rect 4379 276870 4425 276922
rect 4449 276870 4495 276922
rect 4495 276870 4505 276922
rect 4529 276870 4559 276922
rect 4559 276870 4585 276922
rect 4289 276868 4345 276870
rect 4369 276868 4425 276870
rect 4449 276868 4505 276870
rect 4529 276868 4585 276870
rect 4289 275834 4345 275836
rect 4369 275834 4425 275836
rect 4449 275834 4505 275836
rect 4529 275834 4585 275836
rect 4289 275782 4315 275834
rect 4315 275782 4345 275834
rect 4369 275782 4379 275834
rect 4379 275782 4425 275834
rect 4449 275782 4495 275834
rect 4495 275782 4505 275834
rect 4529 275782 4559 275834
rect 4559 275782 4585 275834
rect 4289 275780 4345 275782
rect 4369 275780 4425 275782
rect 4449 275780 4505 275782
rect 4529 275780 4585 275782
rect 4289 274746 4345 274748
rect 4369 274746 4425 274748
rect 4449 274746 4505 274748
rect 4529 274746 4585 274748
rect 4289 274694 4315 274746
rect 4315 274694 4345 274746
rect 4369 274694 4379 274746
rect 4379 274694 4425 274746
rect 4449 274694 4495 274746
rect 4495 274694 4505 274746
rect 4529 274694 4559 274746
rect 4559 274694 4585 274746
rect 4289 274692 4345 274694
rect 4369 274692 4425 274694
rect 4449 274692 4505 274694
rect 4529 274692 4585 274694
rect 4289 273658 4345 273660
rect 4369 273658 4425 273660
rect 4449 273658 4505 273660
rect 4529 273658 4585 273660
rect 4289 273606 4315 273658
rect 4315 273606 4345 273658
rect 4369 273606 4379 273658
rect 4379 273606 4425 273658
rect 4449 273606 4495 273658
rect 4495 273606 4505 273658
rect 4529 273606 4559 273658
rect 4559 273606 4585 273658
rect 4289 273604 4345 273606
rect 4369 273604 4425 273606
rect 4449 273604 4505 273606
rect 4529 273604 4585 273606
rect 4289 272570 4345 272572
rect 4369 272570 4425 272572
rect 4449 272570 4505 272572
rect 4529 272570 4585 272572
rect 4289 272518 4315 272570
rect 4315 272518 4345 272570
rect 4369 272518 4379 272570
rect 4379 272518 4425 272570
rect 4449 272518 4495 272570
rect 4495 272518 4505 272570
rect 4529 272518 4559 272570
rect 4559 272518 4585 272570
rect 4289 272516 4345 272518
rect 4369 272516 4425 272518
rect 4449 272516 4505 272518
rect 4529 272516 4585 272518
rect 4289 271482 4345 271484
rect 4369 271482 4425 271484
rect 4449 271482 4505 271484
rect 4529 271482 4585 271484
rect 4289 271430 4315 271482
rect 4315 271430 4345 271482
rect 4369 271430 4379 271482
rect 4379 271430 4425 271482
rect 4449 271430 4495 271482
rect 4495 271430 4505 271482
rect 4529 271430 4559 271482
rect 4559 271430 4585 271482
rect 4289 271428 4345 271430
rect 4369 271428 4425 271430
rect 4449 271428 4505 271430
rect 4529 271428 4585 271430
rect 4289 270394 4345 270396
rect 4369 270394 4425 270396
rect 4449 270394 4505 270396
rect 4529 270394 4585 270396
rect 4289 270342 4315 270394
rect 4315 270342 4345 270394
rect 4369 270342 4379 270394
rect 4379 270342 4425 270394
rect 4449 270342 4495 270394
rect 4495 270342 4505 270394
rect 4529 270342 4559 270394
rect 4559 270342 4585 270394
rect 4289 270340 4345 270342
rect 4369 270340 4425 270342
rect 4449 270340 4505 270342
rect 4529 270340 4585 270342
rect 4289 269306 4345 269308
rect 4369 269306 4425 269308
rect 4449 269306 4505 269308
rect 4529 269306 4585 269308
rect 4289 269254 4315 269306
rect 4315 269254 4345 269306
rect 4369 269254 4379 269306
rect 4379 269254 4425 269306
rect 4449 269254 4495 269306
rect 4495 269254 4505 269306
rect 4529 269254 4559 269306
rect 4559 269254 4585 269306
rect 4289 269252 4345 269254
rect 4369 269252 4425 269254
rect 4449 269252 4505 269254
rect 4529 269252 4585 269254
rect 4289 268218 4345 268220
rect 4369 268218 4425 268220
rect 4449 268218 4505 268220
rect 4529 268218 4585 268220
rect 4289 268166 4315 268218
rect 4315 268166 4345 268218
rect 4369 268166 4379 268218
rect 4379 268166 4425 268218
rect 4449 268166 4495 268218
rect 4495 268166 4505 268218
rect 4529 268166 4559 268218
rect 4559 268166 4585 268218
rect 4289 268164 4345 268166
rect 4369 268164 4425 268166
rect 4449 268164 4505 268166
rect 4529 268164 4585 268166
rect 4289 267130 4345 267132
rect 4369 267130 4425 267132
rect 4449 267130 4505 267132
rect 4529 267130 4585 267132
rect 4289 267078 4315 267130
rect 4315 267078 4345 267130
rect 4369 267078 4379 267130
rect 4379 267078 4425 267130
rect 4449 267078 4495 267130
rect 4495 267078 4505 267130
rect 4529 267078 4559 267130
rect 4559 267078 4585 267130
rect 4289 267076 4345 267078
rect 4369 267076 4425 267078
rect 4449 267076 4505 267078
rect 4529 267076 4585 267078
rect 4289 266042 4345 266044
rect 4369 266042 4425 266044
rect 4449 266042 4505 266044
rect 4529 266042 4585 266044
rect 4289 265990 4315 266042
rect 4315 265990 4345 266042
rect 4369 265990 4379 266042
rect 4379 265990 4425 266042
rect 4449 265990 4495 266042
rect 4495 265990 4505 266042
rect 4529 265990 4559 266042
rect 4559 265990 4585 266042
rect 4289 265988 4345 265990
rect 4369 265988 4425 265990
rect 4449 265988 4505 265990
rect 4529 265988 4585 265990
rect 4289 264954 4345 264956
rect 4369 264954 4425 264956
rect 4449 264954 4505 264956
rect 4529 264954 4585 264956
rect 4289 264902 4315 264954
rect 4315 264902 4345 264954
rect 4369 264902 4379 264954
rect 4379 264902 4425 264954
rect 4449 264902 4495 264954
rect 4495 264902 4505 264954
rect 4529 264902 4559 264954
rect 4559 264902 4585 264954
rect 4289 264900 4345 264902
rect 4369 264900 4425 264902
rect 4449 264900 4505 264902
rect 4529 264900 4585 264902
rect 4289 263866 4345 263868
rect 4369 263866 4425 263868
rect 4449 263866 4505 263868
rect 4529 263866 4585 263868
rect 4289 263814 4315 263866
rect 4315 263814 4345 263866
rect 4369 263814 4379 263866
rect 4379 263814 4425 263866
rect 4449 263814 4495 263866
rect 4495 263814 4505 263866
rect 4529 263814 4559 263866
rect 4559 263814 4585 263866
rect 4289 263812 4345 263814
rect 4369 263812 4425 263814
rect 4449 263812 4505 263814
rect 4529 263812 4585 263814
rect 4289 262778 4345 262780
rect 4369 262778 4425 262780
rect 4449 262778 4505 262780
rect 4529 262778 4585 262780
rect 4289 262726 4315 262778
rect 4315 262726 4345 262778
rect 4369 262726 4379 262778
rect 4379 262726 4425 262778
rect 4449 262726 4495 262778
rect 4495 262726 4505 262778
rect 4529 262726 4559 262778
rect 4559 262726 4585 262778
rect 4289 262724 4345 262726
rect 4369 262724 4425 262726
rect 4449 262724 4505 262726
rect 4529 262724 4585 262726
rect 4289 261690 4345 261692
rect 4369 261690 4425 261692
rect 4449 261690 4505 261692
rect 4529 261690 4585 261692
rect 4289 261638 4315 261690
rect 4315 261638 4345 261690
rect 4369 261638 4379 261690
rect 4379 261638 4425 261690
rect 4449 261638 4495 261690
rect 4495 261638 4505 261690
rect 4529 261638 4559 261690
rect 4559 261638 4585 261690
rect 4289 261636 4345 261638
rect 4369 261636 4425 261638
rect 4449 261636 4505 261638
rect 4529 261636 4585 261638
rect 4289 260602 4345 260604
rect 4369 260602 4425 260604
rect 4449 260602 4505 260604
rect 4529 260602 4585 260604
rect 4289 260550 4315 260602
rect 4315 260550 4345 260602
rect 4369 260550 4379 260602
rect 4379 260550 4425 260602
rect 4449 260550 4495 260602
rect 4495 260550 4505 260602
rect 4529 260550 4559 260602
rect 4559 260550 4585 260602
rect 4289 260548 4345 260550
rect 4369 260548 4425 260550
rect 4449 260548 4505 260550
rect 4529 260548 4585 260550
rect 4289 259514 4345 259516
rect 4369 259514 4425 259516
rect 4449 259514 4505 259516
rect 4529 259514 4585 259516
rect 4289 259462 4315 259514
rect 4315 259462 4345 259514
rect 4369 259462 4379 259514
rect 4379 259462 4425 259514
rect 4449 259462 4495 259514
rect 4495 259462 4505 259514
rect 4529 259462 4559 259514
rect 4559 259462 4585 259514
rect 4289 259460 4345 259462
rect 4369 259460 4425 259462
rect 4449 259460 4505 259462
rect 4529 259460 4585 259462
rect 4289 258426 4345 258428
rect 4369 258426 4425 258428
rect 4449 258426 4505 258428
rect 4529 258426 4585 258428
rect 4289 258374 4315 258426
rect 4315 258374 4345 258426
rect 4369 258374 4379 258426
rect 4379 258374 4425 258426
rect 4449 258374 4495 258426
rect 4495 258374 4505 258426
rect 4529 258374 4559 258426
rect 4559 258374 4585 258426
rect 4289 258372 4345 258374
rect 4369 258372 4425 258374
rect 4449 258372 4505 258374
rect 4529 258372 4585 258374
rect 4289 257338 4345 257340
rect 4369 257338 4425 257340
rect 4449 257338 4505 257340
rect 4529 257338 4585 257340
rect 4289 257286 4315 257338
rect 4315 257286 4345 257338
rect 4369 257286 4379 257338
rect 4379 257286 4425 257338
rect 4449 257286 4495 257338
rect 4495 257286 4505 257338
rect 4529 257286 4559 257338
rect 4559 257286 4585 257338
rect 4289 257284 4345 257286
rect 4369 257284 4425 257286
rect 4449 257284 4505 257286
rect 4529 257284 4585 257286
rect 4289 256250 4345 256252
rect 4369 256250 4425 256252
rect 4449 256250 4505 256252
rect 4529 256250 4585 256252
rect 4289 256198 4315 256250
rect 4315 256198 4345 256250
rect 4369 256198 4379 256250
rect 4379 256198 4425 256250
rect 4449 256198 4495 256250
rect 4495 256198 4505 256250
rect 4529 256198 4559 256250
rect 4559 256198 4585 256250
rect 4289 256196 4345 256198
rect 4369 256196 4425 256198
rect 4449 256196 4505 256198
rect 4529 256196 4585 256198
rect 4289 255162 4345 255164
rect 4369 255162 4425 255164
rect 4449 255162 4505 255164
rect 4529 255162 4585 255164
rect 4289 255110 4315 255162
rect 4315 255110 4345 255162
rect 4369 255110 4379 255162
rect 4379 255110 4425 255162
rect 4449 255110 4495 255162
rect 4495 255110 4505 255162
rect 4529 255110 4559 255162
rect 4559 255110 4585 255162
rect 4289 255108 4345 255110
rect 4369 255108 4425 255110
rect 4449 255108 4505 255110
rect 4529 255108 4585 255110
rect 4289 254074 4345 254076
rect 4369 254074 4425 254076
rect 4449 254074 4505 254076
rect 4529 254074 4585 254076
rect 4289 254022 4315 254074
rect 4315 254022 4345 254074
rect 4369 254022 4379 254074
rect 4379 254022 4425 254074
rect 4449 254022 4495 254074
rect 4495 254022 4505 254074
rect 4529 254022 4559 254074
rect 4559 254022 4585 254074
rect 4289 254020 4345 254022
rect 4369 254020 4425 254022
rect 4449 254020 4505 254022
rect 4529 254020 4585 254022
rect 4289 252986 4345 252988
rect 4369 252986 4425 252988
rect 4449 252986 4505 252988
rect 4529 252986 4585 252988
rect 4289 252934 4315 252986
rect 4315 252934 4345 252986
rect 4369 252934 4379 252986
rect 4379 252934 4425 252986
rect 4449 252934 4495 252986
rect 4495 252934 4505 252986
rect 4529 252934 4559 252986
rect 4559 252934 4585 252986
rect 4289 252932 4345 252934
rect 4369 252932 4425 252934
rect 4449 252932 4505 252934
rect 4529 252932 4585 252934
rect 4289 251898 4345 251900
rect 4369 251898 4425 251900
rect 4449 251898 4505 251900
rect 4529 251898 4585 251900
rect 4289 251846 4315 251898
rect 4315 251846 4345 251898
rect 4369 251846 4379 251898
rect 4379 251846 4425 251898
rect 4449 251846 4495 251898
rect 4495 251846 4505 251898
rect 4529 251846 4559 251898
rect 4559 251846 4585 251898
rect 4289 251844 4345 251846
rect 4369 251844 4425 251846
rect 4449 251844 4505 251846
rect 4529 251844 4585 251846
rect 4289 250810 4345 250812
rect 4369 250810 4425 250812
rect 4449 250810 4505 250812
rect 4529 250810 4585 250812
rect 4289 250758 4315 250810
rect 4315 250758 4345 250810
rect 4369 250758 4379 250810
rect 4379 250758 4425 250810
rect 4449 250758 4495 250810
rect 4495 250758 4505 250810
rect 4529 250758 4559 250810
rect 4559 250758 4585 250810
rect 4289 250756 4345 250758
rect 4369 250756 4425 250758
rect 4449 250756 4505 250758
rect 4529 250756 4585 250758
rect 4289 249722 4345 249724
rect 4369 249722 4425 249724
rect 4449 249722 4505 249724
rect 4529 249722 4585 249724
rect 4289 249670 4315 249722
rect 4315 249670 4345 249722
rect 4369 249670 4379 249722
rect 4379 249670 4425 249722
rect 4449 249670 4495 249722
rect 4495 249670 4505 249722
rect 4529 249670 4559 249722
rect 4559 249670 4585 249722
rect 4289 249668 4345 249670
rect 4369 249668 4425 249670
rect 4449 249668 4505 249670
rect 4529 249668 4585 249670
rect 4289 248634 4345 248636
rect 4369 248634 4425 248636
rect 4449 248634 4505 248636
rect 4529 248634 4585 248636
rect 4289 248582 4315 248634
rect 4315 248582 4345 248634
rect 4369 248582 4379 248634
rect 4379 248582 4425 248634
rect 4449 248582 4495 248634
rect 4495 248582 4505 248634
rect 4529 248582 4559 248634
rect 4559 248582 4585 248634
rect 4289 248580 4345 248582
rect 4369 248580 4425 248582
rect 4449 248580 4505 248582
rect 4529 248580 4585 248582
rect 4289 247546 4345 247548
rect 4369 247546 4425 247548
rect 4449 247546 4505 247548
rect 4529 247546 4585 247548
rect 4289 247494 4315 247546
rect 4315 247494 4345 247546
rect 4369 247494 4379 247546
rect 4379 247494 4425 247546
rect 4449 247494 4495 247546
rect 4495 247494 4505 247546
rect 4529 247494 4559 247546
rect 4559 247494 4585 247546
rect 4289 247492 4345 247494
rect 4369 247492 4425 247494
rect 4449 247492 4505 247494
rect 4529 247492 4585 247494
rect 4289 246458 4345 246460
rect 4369 246458 4425 246460
rect 4449 246458 4505 246460
rect 4529 246458 4585 246460
rect 4289 246406 4315 246458
rect 4315 246406 4345 246458
rect 4369 246406 4379 246458
rect 4379 246406 4425 246458
rect 4449 246406 4495 246458
rect 4495 246406 4505 246458
rect 4529 246406 4559 246458
rect 4559 246406 4585 246458
rect 4289 246404 4345 246406
rect 4369 246404 4425 246406
rect 4449 246404 4505 246406
rect 4529 246404 4585 246406
rect 4289 245370 4345 245372
rect 4369 245370 4425 245372
rect 4449 245370 4505 245372
rect 4529 245370 4585 245372
rect 4289 245318 4315 245370
rect 4315 245318 4345 245370
rect 4369 245318 4379 245370
rect 4379 245318 4425 245370
rect 4449 245318 4495 245370
rect 4495 245318 4505 245370
rect 4529 245318 4559 245370
rect 4559 245318 4585 245370
rect 4289 245316 4345 245318
rect 4369 245316 4425 245318
rect 4449 245316 4505 245318
rect 4529 245316 4585 245318
rect 4289 244282 4345 244284
rect 4369 244282 4425 244284
rect 4449 244282 4505 244284
rect 4529 244282 4585 244284
rect 4289 244230 4315 244282
rect 4315 244230 4345 244282
rect 4369 244230 4379 244282
rect 4379 244230 4425 244282
rect 4449 244230 4495 244282
rect 4495 244230 4505 244282
rect 4529 244230 4559 244282
rect 4559 244230 4585 244282
rect 4289 244228 4345 244230
rect 4369 244228 4425 244230
rect 4449 244228 4505 244230
rect 4529 244228 4585 244230
rect 4289 243194 4345 243196
rect 4369 243194 4425 243196
rect 4449 243194 4505 243196
rect 4529 243194 4585 243196
rect 4289 243142 4315 243194
rect 4315 243142 4345 243194
rect 4369 243142 4379 243194
rect 4379 243142 4425 243194
rect 4449 243142 4495 243194
rect 4495 243142 4505 243194
rect 4529 243142 4559 243194
rect 4559 243142 4585 243194
rect 4289 243140 4345 243142
rect 4369 243140 4425 243142
rect 4449 243140 4505 243142
rect 4529 243140 4585 243142
rect 4289 242106 4345 242108
rect 4369 242106 4425 242108
rect 4449 242106 4505 242108
rect 4529 242106 4585 242108
rect 4289 242054 4315 242106
rect 4315 242054 4345 242106
rect 4369 242054 4379 242106
rect 4379 242054 4425 242106
rect 4449 242054 4495 242106
rect 4495 242054 4505 242106
rect 4529 242054 4559 242106
rect 4559 242054 4585 242106
rect 4289 242052 4345 242054
rect 4369 242052 4425 242054
rect 4449 242052 4505 242054
rect 4529 242052 4585 242054
rect 4289 241018 4345 241020
rect 4369 241018 4425 241020
rect 4449 241018 4505 241020
rect 4529 241018 4585 241020
rect 4289 240966 4315 241018
rect 4315 240966 4345 241018
rect 4369 240966 4379 241018
rect 4379 240966 4425 241018
rect 4449 240966 4495 241018
rect 4495 240966 4505 241018
rect 4529 240966 4559 241018
rect 4559 240966 4585 241018
rect 4289 240964 4345 240966
rect 4369 240964 4425 240966
rect 4449 240964 4505 240966
rect 4529 240964 4585 240966
rect 4289 239930 4345 239932
rect 4369 239930 4425 239932
rect 4449 239930 4505 239932
rect 4529 239930 4585 239932
rect 4289 239878 4315 239930
rect 4315 239878 4345 239930
rect 4369 239878 4379 239930
rect 4379 239878 4425 239930
rect 4449 239878 4495 239930
rect 4495 239878 4505 239930
rect 4529 239878 4559 239930
rect 4559 239878 4585 239930
rect 4289 239876 4345 239878
rect 4369 239876 4425 239878
rect 4449 239876 4505 239878
rect 4529 239876 4585 239878
rect 4289 238842 4345 238844
rect 4369 238842 4425 238844
rect 4449 238842 4505 238844
rect 4529 238842 4585 238844
rect 4289 238790 4315 238842
rect 4315 238790 4345 238842
rect 4369 238790 4379 238842
rect 4379 238790 4425 238842
rect 4449 238790 4495 238842
rect 4495 238790 4505 238842
rect 4529 238790 4559 238842
rect 4559 238790 4585 238842
rect 4289 238788 4345 238790
rect 4369 238788 4425 238790
rect 4449 238788 4505 238790
rect 4529 238788 4585 238790
rect 4289 237754 4345 237756
rect 4369 237754 4425 237756
rect 4449 237754 4505 237756
rect 4529 237754 4585 237756
rect 4289 237702 4315 237754
rect 4315 237702 4345 237754
rect 4369 237702 4379 237754
rect 4379 237702 4425 237754
rect 4449 237702 4495 237754
rect 4495 237702 4505 237754
rect 4529 237702 4559 237754
rect 4559 237702 4585 237754
rect 4289 237700 4345 237702
rect 4369 237700 4425 237702
rect 4449 237700 4505 237702
rect 4529 237700 4585 237702
rect 4289 236666 4345 236668
rect 4369 236666 4425 236668
rect 4449 236666 4505 236668
rect 4529 236666 4585 236668
rect 4289 236614 4315 236666
rect 4315 236614 4345 236666
rect 4369 236614 4379 236666
rect 4379 236614 4425 236666
rect 4449 236614 4495 236666
rect 4495 236614 4505 236666
rect 4529 236614 4559 236666
rect 4559 236614 4585 236666
rect 4289 236612 4345 236614
rect 4369 236612 4425 236614
rect 4449 236612 4505 236614
rect 4529 236612 4585 236614
rect 4289 235578 4345 235580
rect 4369 235578 4425 235580
rect 4449 235578 4505 235580
rect 4529 235578 4585 235580
rect 4289 235526 4315 235578
rect 4315 235526 4345 235578
rect 4369 235526 4379 235578
rect 4379 235526 4425 235578
rect 4449 235526 4495 235578
rect 4495 235526 4505 235578
rect 4529 235526 4559 235578
rect 4559 235526 4585 235578
rect 4289 235524 4345 235526
rect 4369 235524 4425 235526
rect 4449 235524 4505 235526
rect 4529 235524 4585 235526
rect 4289 234490 4345 234492
rect 4369 234490 4425 234492
rect 4449 234490 4505 234492
rect 4529 234490 4585 234492
rect 4289 234438 4315 234490
rect 4315 234438 4345 234490
rect 4369 234438 4379 234490
rect 4379 234438 4425 234490
rect 4449 234438 4495 234490
rect 4495 234438 4505 234490
rect 4529 234438 4559 234490
rect 4559 234438 4585 234490
rect 4289 234436 4345 234438
rect 4369 234436 4425 234438
rect 4449 234436 4505 234438
rect 4529 234436 4585 234438
rect 4289 233402 4345 233404
rect 4369 233402 4425 233404
rect 4449 233402 4505 233404
rect 4529 233402 4585 233404
rect 4289 233350 4315 233402
rect 4315 233350 4345 233402
rect 4369 233350 4379 233402
rect 4379 233350 4425 233402
rect 4449 233350 4495 233402
rect 4495 233350 4505 233402
rect 4529 233350 4559 233402
rect 4559 233350 4585 233402
rect 4289 233348 4345 233350
rect 4369 233348 4425 233350
rect 4449 233348 4505 233350
rect 4529 233348 4585 233350
rect 4289 232314 4345 232316
rect 4369 232314 4425 232316
rect 4449 232314 4505 232316
rect 4529 232314 4585 232316
rect 4289 232262 4315 232314
rect 4315 232262 4345 232314
rect 4369 232262 4379 232314
rect 4379 232262 4425 232314
rect 4449 232262 4495 232314
rect 4495 232262 4505 232314
rect 4529 232262 4559 232314
rect 4559 232262 4585 232314
rect 4289 232260 4345 232262
rect 4369 232260 4425 232262
rect 4449 232260 4505 232262
rect 4529 232260 4585 232262
rect 4289 231226 4345 231228
rect 4369 231226 4425 231228
rect 4449 231226 4505 231228
rect 4529 231226 4585 231228
rect 4289 231174 4315 231226
rect 4315 231174 4345 231226
rect 4369 231174 4379 231226
rect 4379 231174 4425 231226
rect 4449 231174 4495 231226
rect 4495 231174 4505 231226
rect 4529 231174 4559 231226
rect 4559 231174 4585 231226
rect 4289 231172 4345 231174
rect 4369 231172 4425 231174
rect 4449 231172 4505 231174
rect 4529 231172 4585 231174
rect 4289 230138 4345 230140
rect 4369 230138 4425 230140
rect 4449 230138 4505 230140
rect 4529 230138 4585 230140
rect 4289 230086 4315 230138
rect 4315 230086 4345 230138
rect 4369 230086 4379 230138
rect 4379 230086 4425 230138
rect 4449 230086 4495 230138
rect 4495 230086 4505 230138
rect 4529 230086 4559 230138
rect 4559 230086 4585 230138
rect 4289 230084 4345 230086
rect 4369 230084 4425 230086
rect 4449 230084 4505 230086
rect 4529 230084 4585 230086
rect 4289 229050 4345 229052
rect 4369 229050 4425 229052
rect 4449 229050 4505 229052
rect 4529 229050 4585 229052
rect 4289 228998 4315 229050
rect 4315 228998 4345 229050
rect 4369 228998 4379 229050
rect 4379 228998 4425 229050
rect 4449 228998 4495 229050
rect 4495 228998 4505 229050
rect 4529 228998 4559 229050
rect 4559 228998 4585 229050
rect 4289 228996 4345 228998
rect 4369 228996 4425 228998
rect 4449 228996 4505 228998
rect 4529 228996 4585 228998
rect 4289 227962 4345 227964
rect 4369 227962 4425 227964
rect 4449 227962 4505 227964
rect 4529 227962 4585 227964
rect 4289 227910 4315 227962
rect 4315 227910 4345 227962
rect 4369 227910 4379 227962
rect 4379 227910 4425 227962
rect 4449 227910 4495 227962
rect 4495 227910 4505 227962
rect 4529 227910 4559 227962
rect 4559 227910 4585 227962
rect 4289 227908 4345 227910
rect 4369 227908 4425 227910
rect 4449 227908 4505 227910
rect 4529 227908 4585 227910
rect 4289 226874 4345 226876
rect 4369 226874 4425 226876
rect 4449 226874 4505 226876
rect 4529 226874 4585 226876
rect 4289 226822 4315 226874
rect 4315 226822 4345 226874
rect 4369 226822 4379 226874
rect 4379 226822 4425 226874
rect 4449 226822 4495 226874
rect 4495 226822 4505 226874
rect 4529 226822 4559 226874
rect 4559 226822 4585 226874
rect 4289 226820 4345 226822
rect 4369 226820 4425 226822
rect 4449 226820 4505 226822
rect 4529 226820 4585 226822
rect 4289 225786 4345 225788
rect 4369 225786 4425 225788
rect 4449 225786 4505 225788
rect 4529 225786 4585 225788
rect 4289 225734 4315 225786
rect 4315 225734 4345 225786
rect 4369 225734 4379 225786
rect 4379 225734 4425 225786
rect 4449 225734 4495 225786
rect 4495 225734 4505 225786
rect 4529 225734 4559 225786
rect 4559 225734 4585 225786
rect 4289 225732 4345 225734
rect 4369 225732 4425 225734
rect 4449 225732 4505 225734
rect 4529 225732 4585 225734
rect 4289 224698 4345 224700
rect 4369 224698 4425 224700
rect 4449 224698 4505 224700
rect 4529 224698 4585 224700
rect 4289 224646 4315 224698
rect 4315 224646 4345 224698
rect 4369 224646 4379 224698
rect 4379 224646 4425 224698
rect 4449 224646 4495 224698
rect 4495 224646 4505 224698
rect 4529 224646 4559 224698
rect 4559 224646 4585 224698
rect 4289 224644 4345 224646
rect 4369 224644 4425 224646
rect 4449 224644 4505 224646
rect 4529 224644 4585 224646
rect 4289 223610 4345 223612
rect 4369 223610 4425 223612
rect 4449 223610 4505 223612
rect 4529 223610 4585 223612
rect 4289 223558 4315 223610
rect 4315 223558 4345 223610
rect 4369 223558 4379 223610
rect 4379 223558 4425 223610
rect 4449 223558 4495 223610
rect 4495 223558 4505 223610
rect 4529 223558 4559 223610
rect 4559 223558 4585 223610
rect 4289 223556 4345 223558
rect 4369 223556 4425 223558
rect 4449 223556 4505 223558
rect 4529 223556 4585 223558
rect 4289 222522 4345 222524
rect 4369 222522 4425 222524
rect 4449 222522 4505 222524
rect 4529 222522 4585 222524
rect 4289 222470 4315 222522
rect 4315 222470 4345 222522
rect 4369 222470 4379 222522
rect 4379 222470 4425 222522
rect 4449 222470 4495 222522
rect 4495 222470 4505 222522
rect 4529 222470 4559 222522
rect 4559 222470 4585 222522
rect 4289 222468 4345 222470
rect 4369 222468 4425 222470
rect 4449 222468 4505 222470
rect 4529 222468 4585 222470
rect 4289 221434 4345 221436
rect 4369 221434 4425 221436
rect 4449 221434 4505 221436
rect 4529 221434 4585 221436
rect 4289 221382 4315 221434
rect 4315 221382 4345 221434
rect 4369 221382 4379 221434
rect 4379 221382 4425 221434
rect 4449 221382 4495 221434
rect 4495 221382 4505 221434
rect 4529 221382 4559 221434
rect 4559 221382 4585 221434
rect 4289 221380 4345 221382
rect 4369 221380 4425 221382
rect 4449 221380 4505 221382
rect 4529 221380 4585 221382
rect 4289 220346 4345 220348
rect 4369 220346 4425 220348
rect 4449 220346 4505 220348
rect 4529 220346 4585 220348
rect 4289 220294 4315 220346
rect 4315 220294 4345 220346
rect 4369 220294 4379 220346
rect 4379 220294 4425 220346
rect 4449 220294 4495 220346
rect 4495 220294 4505 220346
rect 4529 220294 4559 220346
rect 4559 220294 4585 220346
rect 4289 220292 4345 220294
rect 4369 220292 4425 220294
rect 4449 220292 4505 220294
rect 4529 220292 4585 220294
rect 4289 219258 4345 219260
rect 4369 219258 4425 219260
rect 4449 219258 4505 219260
rect 4529 219258 4585 219260
rect 4289 219206 4315 219258
rect 4315 219206 4345 219258
rect 4369 219206 4379 219258
rect 4379 219206 4425 219258
rect 4449 219206 4495 219258
rect 4495 219206 4505 219258
rect 4529 219206 4559 219258
rect 4559 219206 4585 219258
rect 4289 219204 4345 219206
rect 4369 219204 4425 219206
rect 4449 219204 4505 219206
rect 4529 219204 4585 219206
rect 4289 218170 4345 218172
rect 4369 218170 4425 218172
rect 4449 218170 4505 218172
rect 4529 218170 4585 218172
rect 4289 218118 4315 218170
rect 4315 218118 4345 218170
rect 4369 218118 4379 218170
rect 4379 218118 4425 218170
rect 4449 218118 4495 218170
rect 4495 218118 4505 218170
rect 4529 218118 4559 218170
rect 4559 218118 4585 218170
rect 4289 218116 4345 218118
rect 4369 218116 4425 218118
rect 4449 218116 4505 218118
rect 4529 218116 4585 218118
rect 4289 217082 4345 217084
rect 4369 217082 4425 217084
rect 4449 217082 4505 217084
rect 4529 217082 4585 217084
rect 4289 217030 4315 217082
rect 4315 217030 4345 217082
rect 4369 217030 4379 217082
rect 4379 217030 4425 217082
rect 4449 217030 4495 217082
rect 4495 217030 4505 217082
rect 4529 217030 4559 217082
rect 4559 217030 4585 217082
rect 4289 217028 4345 217030
rect 4369 217028 4425 217030
rect 4449 217028 4505 217030
rect 4529 217028 4585 217030
rect 4289 215994 4345 215996
rect 4369 215994 4425 215996
rect 4449 215994 4505 215996
rect 4529 215994 4585 215996
rect 4289 215942 4315 215994
rect 4315 215942 4345 215994
rect 4369 215942 4379 215994
rect 4379 215942 4425 215994
rect 4449 215942 4495 215994
rect 4495 215942 4505 215994
rect 4529 215942 4559 215994
rect 4559 215942 4585 215994
rect 4289 215940 4345 215942
rect 4369 215940 4425 215942
rect 4449 215940 4505 215942
rect 4529 215940 4585 215942
rect 4289 214906 4345 214908
rect 4369 214906 4425 214908
rect 4449 214906 4505 214908
rect 4529 214906 4585 214908
rect 4289 214854 4315 214906
rect 4315 214854 4345 214906
rect 4369 214854 4379 214906
rect 4379 214854 4425 214906
rect 4449 214854 4495 214906
rect 4495 214854 4505 214906
rect 4529 214854 4559 214906
rect 4559 214854 4585 214906
rect 4289 214852 4345 214854
rect 4369 214852 4425 214854
rect 4449 214852 4505 214854
rect 4529 214852 4585 214854
rect 4289 213818 4345 213820
rect 4369 213818 4425 213820
rect 4449 213818 4505 213820
rect 4529 213818 4585 213820
rect 4289 213766 4315 213818
rect 4315 213766 4345 213818
rect 4369 213766 4379 213818
rect 4379 213766 4425 213818
rect 4449 213766 4495 213818
rect 4495 213766 4505 213818
rect 4529 213766 4559 213818
rect 4559 213766 4585 213818
rect 4289 213764 4345 213766
rect 4369 213764 4425 213766
rect 4449 213764 4505 213766
rect 4529 213764 4585 213766
rect 4289 212730 4345 212732
rect 4369 212730 4425 212732
rect 4449 212730 4505 212732
rect 4529 212730 4585 212732
rect 4289 212678 4315 212730
rect 4315 212678 4345 212730
rect 4369 212678 4379 212730
rect 4379 212678 4425 212730
rect 4449 212678 4495 212730
rect 4495 212678 4505 212730
rect 4529 212678 4559 212730
rect 4559 212678 4585 212730
rect 4289 212676 4345 212678
rect 4369 212676 4425 212678
rect 4449 212676 4505 212678
rect 4529 212676 4585 212678
rect 4289 211642 4345 211644
rect 4369 211642 4425 211644
rect 4449 211642 4505 211644
rect 4529 211642 4585 211644
rect 4289 211590 4315 211642
rect 4315 211590 4345 211642
rect 4369 211590 4379 211642
rect 4379 211590 4425 211642
rect 4449 211590 4495 211642
rect 4495 211590 4505 211642
rect 4529 211590 4559 211642
rect 4559 211590 4585 211642
rect 4289 211588 4345 211590
rect 4369 211588 4425 211590
rect 4449 211588 4505 211590
rect 4529 211588 4585 211590
rect 4289 210554 4345 210556
rect 4369 210554 4425 210556
rect 4449 210554 4505 210556
rect 4529 210554 4585 210556
rect 4289 210502 4315 210554
rect 4315 210502 4345 210554
rect 4369 210502 4379 210554
rect 4379 210502 4425 210554
rect 4449 210502 4495 210554
rect 4495 210502 4505 210554
rect 4529 210502 4559 210554
rect 4559 210502 4585 210554
rect 4289 210500 4345 210502
rect 4369 210500 4425 210502
rect 4449 210500 4505 210502
rect 4529 210500 4585 210502
rect 4289 209466 4345 209468
rect 4369 209466 4425 209468
rect 4449 209466 4505 209468
rect 4529 209466 4585 209468
rect 4289 209414 4315 209466
rect 4315 209414 4345 209466
rect 4369 209414 4379 209466
rect 4379 209414 4425 209466
rect 4449 209414 4495 209466
rect 4495 209414 4505 209466
rect 4529 209414 4559 209466
rect 4559 209414 4585 209466
rect 4289 209412 4345 209414
rect 4369 209412 4425 209414
rect 4449 209412 4505 209414
rect 4529 209412 4585 209414
rect 4289 208378 4345 208380
rect 4369 208378 4425 208380
rect 4449 208378 4505 208380
rect 4529 208378 4585 208380
rect 4289 208326 4315 208378
rect 4315 208326 4345 208378
rect 4369 208326 4379 208378
rect 4379 208326 4425 208378
rect 4449 208326 4495 208378
rect 4495 208326 4505 208378
rect 4529 208326 4559 208378
rect 4559 208326 4585 208378
rect 4289 208324 4345 208326
rect 4369 208324 4425 208326
rect 4449 208324 4505 208326
rect 4529 208324 4585 208326
rect 4289 207290 4345 207292
rect 4369 207290 4425 207292
rect 4449 207290 4505 207292
rect 4529 207290 4585 207292
rect 4289 207238 4315 207290
rect 4315 207238 4345 207290
rect 4369 207238 4379 207290
rect 4379 207238 4425 207290
rect 4449 207238 4495 207290
rect 4495 207238 4505 207290
rect 4529 207238 4559 207290
rect 4559 207238 4585 207290
rect 4289 207236 4345 207238
rect 4369 207236 4425 207238
rect 4449 207236 4505 207238
rect 4529 207236 4585 207238
rect 4289 206202 4345 206204
rect 4369 206202 4425 206204
rect 4449 206202 4505 206204
rect 4529 206202 4585 206204
rect 4289 206150 4315 206202
rect 4315 206150 4345 206202
rect 4369 206150 4379 206202
rect 4379 206150 4425 206202
rect 4449 206150 4495 206202
rect 4495 206150 4505 206202
rect 4529 206150 4559 206202
rect 4559 206150 4585 206202
rect 4289 206148 4345 206150
rect 4369 206148 4425 206150
rect 4449 206148 4505 206150
rect 4529 206148 4585 206150
rect 4289 205114 4345 205116
rect 4369 205114 4425 205116
rect 4449 205114 4505 205116
rect 4529 205114 4585 205116
rect 4289 205062 4315 205114
rect 4315 205062 4345 205114
rect 4369 205062 4379 205114
rect 4379 205062 4425 205114
rect 4449 205062 4495 205114
rect 4495 205062 4505 205114
rect 4529 205062 4559 205114
rect 4559 205062 4585 205114
rect 4289 205060 4345 205062
rect 4369 205060 4425 205062
rect 4449 205060 4505 205062
rect 4529 205060 4585 205062
rect 4289 204026 4345 204028
rect 4369 204026 4425 204028
rect 4449 204026 4505 204028
rect 4529 204026 4585 204028
rect 4289 203974 4315 204026
rect 4315 203974 4345 204026
rect 4369 203974 4379 204026
rect 4379 203974 4425 204026
rect 4449 203974 4495 204026
rect 4495 203974 4505 204026
rect 4529 203974 4559 204026
rect 4559 203974 4585 204026
rect 4289 203972 4345 203974
rect 4369 203972 4425 203974
rect 4449 203972 4505 203974
rect 4529 203972 4585 203974
rect 4289 202938 4345 202940
rect 4369 202938 4425 202940
rect 4449 202938 4505 202940
rect 4529 202938 4585 202940
rect 4289 202886 4315 202938
rect 4315 202886 4345 202938
rect 4369 202886 4379 202938
rect 4379 202886 4425 202938
rect 4449 202886 4495 202938
rect 4495 202886 4505 202938
rect 4529 202886 4559 202938
rect 4559 202886 4585 202938
rect 4289 202884 4345 202886
rect 4369 202884 4425 202886
rect 4449 202884 4505 202886
rect 4529 202884 4585 202886
rect 4289 201850 4345 201852
rect 4369 201850 4425 201852
rect 4449 201850 4505 201852
rect 4529 201850 4585 201852
rect 4289 201798 4315 201850
rect 4315 201798 4345 201850
rect 4369 201798 4379 201850
rect 4379 201798 4425 201850
rect 4449 201798 4495 201850
rect 4495 201798 4505 201850
rect 4529 201798 4559 201850
rect 4559 201798 4585 201850
rect 4289 201796 4345 201798
rect 4369 201796 4425 201798
rect 4449 201796 4505 201798
rect 4529 201796 4585 201798
rect 4289 200762 4345 200764
rect 4369 200762 4425 200764
rect 4449 200762 4505 200764
rect 4529 200762 4585 200764
rect 4289 200710 4315 200762
rect 4315 200710 4345 200762
rect 4369 200710 4379 200762
rect 4379 200710 4425 200762
rect 4449 200710 4495 200762
rect 4495 200710 4505 200762
rect 4529 200710 4559 200762
rect 4559 200710 4585 200762
rect 4289 200708 4345 200710
rect 4369 200708 4425 200710
rect 4449 200708 4505 200710
rect 4529 200708 4585 200710
rect 4289 199674 4345 199676
rect 4369 199674 4425 199676
rect 4449 199674 4505 199676
rect 4529 199674 4585 199676
rect 4289 199622 4315 199674
rect 4315 199622 4345 199674
rect 4369 199622 4379 199674
rect 4379 199622 4425 199674
rect 4449 199622 4495 199674
rect 4495 199622 4505 199674
rect 4529 199622 4559 199674
rect 4559 199622 4585 199674
rect 4289 199620 4345 199622
rect 4369 199620 4425 199622
rect 4449 199620 4505 199622
rect 4529 199620 4585 199622
rect 4289 198586 4345 198588
rect 4369 198586 4425 198588
rect 4449 198586 4505 198588
rect 4529 198586 4585 198588
rect 4289 198534 4315 198586
rect 4315 198534 4345 198586
rect 4369 198534 4379 198586
rect 4379 198534 4425 198586
rect 4449 198534 4495 198586
rect 4495 198534 4505 198586
rect 4529 198534 4559 198586
rect 4559 198534 4585 198586
rect 4289 198532 4345 198534
rect 4369 198532 4425 198534
rect 4449 198532 4505 198534
rect 4529 198532 4585 198534
rect 4289 197498 4345 197500
rect 4369 197498 4425 197500
rect 4449 197498 4505 197500
rect 4529 197498 4585 197500
rect 4289 197446 4315 197498
rect 4315 197446 4345 197498
rect 4369 197446 4379 197498
rect 4379 197446 4425 197498
rect 4449 197446 4495 197498
rect 4495 197446 4505 197498
rect 4529 197446 4559 197498
rect 4559 197446 4585 197498
rect 4289 197444 4345 197446
rect 4369 197444 4425 197446
rect 4449 197444 4505 197446
rect 4529 197444 4585 197446
rect 4289 196410 4345 196412
rect 4369 196410 4425 196412
rect 4449 196410 4505 196412
rect 4529 196410 4585 196412
rect 4289 196358 4315 196410
rect 4315 196358 4345 196410
rect 4369 196358 4379 196410
rect 4379 196358 4425 196410
rect 4449 196358 4495 196410
rect 4495 196358 4505 196410
rect 4529 196358 4559 196410
rect 4559 196358 4585 196410
rect 4289 196356 4345 196358
rect 4369 196356 4425 196358
rect 4449 196356 4505 196358
rect 4529 196356 4585 196358
rect 4289 195322 4345 195324
rect 4369 195322 4425 195324
rect 4449 195322 4505 195324
rect 4529 195322 4585 195324
rect 4289 195270 4315 195322
rect 4315 195270 4345 195322
rect 4369 195270 4379 195322
rect 4379 195270 4425 195322
rect 4449 195270 4495 195322
rect 4495 195270 4505 195322
rect 4529 195270 4559 195322
rect 4559 195270 4585 195322
rect 4289 195268 4345 195270
rect 4369 195268 4425 195270
rect 4449 195268 4505 195270
rect 4529 195268 4585 195270
rect 4289 194234 4345 194236
rect 4369 194234 4425 194236
rect 4449 194234 4505 194236
rect 4529 194234 4585 194236
rect 4289 194182 4315 194234
rect 4315 194182 4345 194234
rect 4369 194182 4379 194234
rect 4379 194182 4425 194234
rect 4449 194182 4495 194234
rect 4495 194182 4505 194234
rect 4529 194182 4559 194234
rect 4559 194182 4585 194234
rect 4289 194180 4345 194182
rect 4369 194180 4425 194182
rect 4449 194180 4505 194182
rect 4529 194180 4585 194182
rect 4289 193146 4345 193148
rect 4369 193146 4425 193148
rect 4449 193146 4505 193148
rect 4529 193146 4585 193148
rect 4289 193094 4315 193146
rect 4315 193094 4345 193146
rect 4369 193094 4379 193146
rect 4379 193094 4425 193146
rect 4449 193094 4495 193146
rect 4495 193094 4505 193146
rect 4529 193094 4559 193146
rect 4559 193094 4585 193146
rect 4289 193092 4345 193094
rect 4369 193092 4425 193094
rect 4449 193092 4505 193094
rect 4529 193092 4585 193094
rect 4289 192058 4345 192060
rect 4369 192058 4425 192060
rect 4449 192058 4505 192060
rect 4529 192058 4585 192060
rect 4289 192006 4315 192058
rect 4315 192006 4345 192058
rect 4369 192006 4379 192058
rect 4379 192006 4425 192058
rect 4449 192006 4495 192058
rect 4495 192006 4505 192058
rect 4529 192006 4559 192058
rect 4559 192006 4585 192058
rect 4289 192004 4345 192006
rect 4369 192004 4425 192006
rect 4449 192004 4505 192006
rect 4529 192004 4585 192006
rect 4289 190970 4345 190972
rect 4369 190970 4425 190972
rect 4449 190970 4505 190972
rect 4529 190970 4585 190972
rect 4289 190918 4315 190970
rect 4315 190918 4345 190970
rect 4369 190918 4379 190970
rect 4379 190918 4425 190970
rect 4449 190918 4495 190970
rect 4495 190918 4505 190970
rect 4529 190918 4559 190970
rect 4559 190918 4585 190970
rect 4289 190916 4345 190918
rect 4369 190916 4425 190918
rect 4449 190916 4505 190918
rect 4529 190916 4585 190918
rect 4289 189882 4345 189884
rect 4369 189882 4425 189884
rect 4449 189882 4505 189884
rect 4529 189882 4585 189884
rect 4289 189830 4315 189882
rect 4315 189830 4345 189882
rect 4369 189830 4379 189882
rect 4379 189830 4425 189882
rect 4449 189830 4495 189882
rect 4495 189830 4505 189882
rect 4529 189830 4559 189882
rect 4559 189830 4585 189882
rect 4289 189828 4345 189830
rect 4369 189828 4425 189830
rect 4449 189828 4505 189830
rect 4529 189828 4585 189830
rect 4289 188794 4345 188796
rect 4369 188794 4425 188796
rect 4449 188794 4505 188796
rect 4529 188794 4585 188796
rect 4289 188742 4315 188794
rect 4315 188742 4345 188794
rect 4369 188742 4379 188794
rect 4379 188742 4425 188794
rect 4449 188742 4495 188794
rect 4495 188742 4505 188794
rect 4529 188742 4559 188794
rect 4559 188742 4585 188794
rect 4289 188740 4345 188742
rect 4369 188740 4425 188742
rect 4449 188740 4505 188742
rect 4529 188740 4585 188742
rect 4289 187706 4345 187708
rect 4369 187706 4425 187708
rect 4449 187706 4505 187708
rect 4529 187706 4585 187708
rect 4289 187654 4315 187706
rect 4315 187654 4345 187706
rect 4369 187654 4379 187706
rect 4379 187654 4425 187706
rect 4449 187654 4495 187706
rect 4495 187654 4505 187706
rect 4529 187654 4559 187706
rect 4559 187654 4585 187706
rect 4289 187652 4345 187654
rect 4369 187652 4425 187654
rect 4449 187652 4505 187654
rect 4529 187652 4585 187654
rect 4289 186618 4345 186620
rect 4369 186618 4425 186620
rect 4449 186618 4505 186620
rect 4529 186618 4585 186620
rect 4289 186566 4315 186618
rect 4315 186566 4345 186618
rect 4369 186566 4379 186618
rect 4379 186566 4425 186618
rect 4449 186566 4495 186618
rect 4495 186566 4505 186618
rect 4529 186566 4559 186618
rect 4559 186566 4585 186618
rect 4289 186564 4345 186566
rect 4369 186564 4425 186566
rect 4449 186564 4505 186566
rect 4529 186564 4585 186566
rect 4289 185530 4345 185532
rect 4369 185530 4425 185532
rect 4449 185530 4505 185532
rect 4529 185530 4585 185532
rect 4289 185478 4315 185530
rect 4315 185478 4345 185530
rect 4369 185478 4379 185530
rect 4379 185478 4425 185530
rect 4449 185478 4495 185530
rect 4495 185478 4505 185530
rect 4529 185478 4559 185530
rect 4559 185478 4585 185530
rect 4289 185476 4345 185478
rect 4369 185476 4425 185478
rect 4449 185476 4505 185478
rect 4529 185476 4585 185478
rect 4289 184442 4345 184444
rect 4369 184442 4425 184444
rect 4449 184442 4505 184444
rect 4529 184442 4585 184444
rect 4289 184390 4315 184442
rect 4315 184390 4345 184442
rect 4369 184390 4379 184442
rect 4379 184390 4425 184442
rect 4449 184390 4495 184442
rect 4495 184390 4505 184442
rect 4529 184390 4559 184442
rect 4559 184390 4585 184442
rect 4289 184388 4345 184390
rect 4369 184388 4425 184390
rect 4449 184388 4505 184390
rect 4529 184388 4585 184390
rect 4289 183354 4345 183356
rect 4369 183354 4425 183356
rect 4449 183354 4505 183356
rect 4529 183354 4585 183356
rect 4289 183302 4315 183354
rect 4315 183302 4345 183354
rect 4369 183302 4379 183354
rect 4379 183302 4425 183354
rect 4449 183302 4495 183354
rect 4495 183302 4505 183354
rect 4529 183302 4559 183354
rect 4559 183302 4585 183354
rect 4289 183300 4345 183302
rect 4369 183300 4425 183302
rect 4449 183300 4505 183302
rect 4529 183300 4585 183302
rect 4289 182266 4345 182268
rect 4369 182266 4425 182268
rect 4449 182266 4505 182268
rect 4529 182266 4585 182268
rect 4289 182214 4315 182266
rect 4315 182214 4345 182266
rect 4369 182214 4379 182266
rect 4379 182214 4425 182266
rect 4449 182214 4495 182266
rect 4495 182214 4505 182266
rect 4529 182214 4559 182266
rect 4559 182214 4585 182266
rect 4289 182212 4345 182214
rect 4369 182212 4425 182214
rect 4449 182212 4505 182214
rect 4529 182212 4585 182214
rect 4289 181178 4345 181180
rect 4369 181178 4425 181180
rect 4449 181178 4505 181180
rect 4529 181178 4585 181180
rect 4289 181126 4315 181178
rect 4315 181126 4345 181178
rect 4369 181126 4379 181178
rect 4379 181126 4425 181178
rect 4449 181126 4495 181178
rect 4495 181126 4505 181178
rect 4529 181126 4559 181178
rect 4559 181126 4585 181178
rect 4289 181124 4345 181126
rect 4369 181124 4425 181126
rect 4449 181124 4505 181126
rect 4529 181124 4585 181126
rect 4289 180090 4345 180092
rect 4369 180090 4425 180092
rect 4449 180090 4505 180092
rect 4529 180090 4585 180092
rect 4289 180038 4315 180090
rect 4315 180038 4345 180090
rect 4369 180038 4379 180090
rect 4379 180038 4425 180090
rect 4449 180038 4495 180090
rect 4495 180038 4505 180090
rect 4529 180038 4559 180090
rect 4559 180038 4585 180090
rect 4289 180036 4345 180038
rect 4369 180036 4425 180038
rect 4449 180036 4505 180038
rect 4529 180036 4585 180038
rect 4289 179002 4345 179004
rect 4369 179002 4425 179004
rect 4449 179002 4505 179004
rect 4529 179002 4585 179004
rect 4289 178950 4315 179002
rect 4315 178950 4345 179002
rect 4369 178950 4379 179002
rect 4379 178950 4425 179002
rect 4449 178950 4495 179002
rect 4495 178950 4505 179002
rect 4529 178950 4559 179002
rect 4559 178950 4585 179002
rect 4289 178948 4345 178950
rect 4369 178948 4425 178950
rect 4449 178948 4505 178950
rect 4529 178948 4585 178950
rect 4289 177914 4345 177916
rect 4369 177914 4425 177916
rect 4449 177914 4505 177916
rect 4529 177914 4585 177916
rect 4289 177862 4315 177914
rect 4315 177862 4345 177914
rect 4369 177862 4379 177914
rect 4379 177862 4425 177914
rect 4449 177862 4495 177914
rect 4495 177862 4505 177914
rect 4529 177862 4559 177914
rect 4559 177862 4585 177914
rect 4289 177860 4345 177862
rect 4369 177860 4425 177862
rect 4449 177860 4505 177862
rect 4529 177860 4585 177862
rect 4289 176826 4345 176828
rect 4369 176826 4425 176828
rect 4449 176826 4505 176828
rect 4529 176826 4585 176828
rect 4289 176774 4315 176826
rect 4315 176774 4345 176826
rect 4369 176774 4379 176826
rect 4379 176774 4425 176826
rect 4449 176774 4495 176826
rect 4495 176774 4505 176826
rect 4529 176774 4559 176826
rect 4559 176774 4585 176826
rect 4289 176772 4345 176774
rect 4369 176772 4425 176774
rect 4449 176772 4505 176774
rect 4529 176772 4585 176774
rect 4289 175738 4345 175740
rect 4369 175738 4425 175740
rect 4449 175738 4505 175740
rect 4529 175738 4585 175740
rect 4289 175686 4315 175738
rect 4315 175686 4345 175738
rect 4369 175686 4379 175738
rect 4379 175686 4425 175738
rect 4449 175686 4495 175738
rect 4495 175686 4505 175738
rect 4529 175686 4559 175738
rect 4559 175686 4585 175738
rect 4289 175684 4345 175686
rect 4369 175684 4425 175686
rect 4449 175684 4505 175686
rect 4529 175684 4585 175686
rect 4289 174650 4345 174652
rect 4369 174650 4425 174652
rect 4449 174650 4505 174652
rect 4529 174650 4585 174652
rect 4289 174598 4315 174650
rect 4315 174598 4345 174650
rect 4369 174598 4379 174650
rect 4379 174598 4425 174650
rect 4449 174598 4495 174650
rect 4495 174598 4505 174650
rect 4529 174598 4559 174650
rect 4559 174598 4585 174650
rect 4289 174596 4345 174598
rect 4369 174596 4425 174598
rect 4449 174596 4505 174598
rect 4529 174596 4585 174598
rect 4289 173562 4345 173564
rect 4369 173562 4425 173564
rect 4449 173562 4505 173564
rect 4529 173562 4585 173564
rect 4289 173510 4315 173562
rect 4315 173510 4345 173562
rect 4369 173510 4379 173562
rect 4379 173510 4425 173562
rect 4449 173510 4495 173562
rect 4495 173510 4505 173562
rect 4529 173510 4559 173562
rect 4559 173510 4585 173562
rect 4289 173508 4345 173510
rect 4369 173508 4425 173510
rect 4449 173508 4505 173510
rect 4529 173508 4585 173510
rect 4289 172474 4345 172476
rect 4369 172474 4425 172476
rect 4449 172474 4505 172476
rect 4529 172474 4585 172476
rect 4289 172422 4315 172474
rect 4315 172422 4345 172474
rect 4369 172422 4379 172474
rect 4379 172422 4425 172474
rect 4449 172422 4495 172474
rect 4495 172422 4505 172474
rect 4529 172422 4559 172474
rect 4559 172422 4585 172474
rect 4289 172420 4345 172422
rect 4369 172420 4425 172422
rect 4449 172420 4505 172422
rect 4529 172420 4585 172422
rect 4289 171386 4345 171388
rect 4369 171386 4425 171388
rect 4449 171386 4505 171388
rect 4529 171386 4585 171388
rect 4289 171334 4315 171386
rect 4315 171334 4345 171386
rect 4369 171334 4379 171386
rect 4379 171334 4425 171386
rect 4449 171334 4495 171386
rect 4495 171334 4505 171386
rect 4529 171334 4559 171386
rect 4559 171334 4585 171386
rect 4289 171332 4345 171334
rect 4369 171332 4425 171334
rect 4449 171332 4505 171334
rect 4529 171332 4585 171334
rect 4289 170298 4345 170300
rect 4369 170298 4425 170300
rect 4449 170298 4505 170300
rect 4529 170298 4585 170300
rect 4289 170246 4315 170298
rect 4315 170246 4345 170298
rect 4369 170246 4379 170298
rect 4379 170246 4425 170298
rect 4449 170246 4495 170298
rect 4495 170246 4505 170298
rect 4529 170246 4559 170298
rect 4559 170246 4585 170298
rect 4289 170244 4345 170246
rect 4369 170244 4425 170246
rect 4449 170244 4505 170246
rect 4529 170244 4585 170246
rect 4289 169210 4345 169212
rect 4369 169210 4425 169212
rect 4449 169210 4505 169212
rect 4529 169210 4585 169212
rect 4289 169158 4315 169210
rect 4315 169158 4345 169210
rect 4369 169158 4379 169210
rect 4379 169158 4425 169210
rect 4449 169158 4495 169210
rect 4495 169158 4505 169210
rect 4529 169158 4559 169210
rect 4559 169158 4585 169210
rect 4289 169156 4345 169158
rect 4369 169156 4425 169158
rect 4449 169156 4505 169158
rect 4529 169156 4585 169158
rect 4289 168122 4345 168124
rect 4369 168122 4425 168124
rect 4449 168122 4505 168124
rect 4529 168122 4585 168124
rect 4289 168070 4315 168122
rect 4315 168070 4345 168122
rect 4369 168070 4379 168122
rect 4379 168070 4425 168122
rect 4449 168070 4495 168122
rect 4495 168070 4505 168122
rect 4529 168070 4559 168122
rect 4559 168070 4585 168122
rect 4289 168068 4345 168070
rect 4369 168068 4425 168070
rect 4449 168068 4505 168070
rect 4529 168068 4585 168070
rect 4289 167034 4345 167036
rect 4369 167034 4425 167036
rect 4449 167034 4505 167036
rect 4529 167034 4585 167036
rect 4289 166982 4315 167034
rect 4315 166982 4345 167034
rect 4369 166982 4379 167034
rect 4379 166982 4425 167034
rect 4449 166982 4495 167034
rect 4495 166982 4505 167034
rect 4529 166982 4559 167034
rect 4559 166982 4585 167034
rect 4289 166980 4345 166982
rect 4369 166980 4425 166982
rect 4449 166980 4505 166982
rect 4529 166980 4585 166982
rect 4289 165946 4345 165948
rect 4369 165946 4425 165948
rect 4449 165946 4505 165948
rect 4529 165946 4585 165948
rect 4289 165894 4315 165946
rect 4315 165894 4345 165946
rect 4369 165894 4379 165946
rect 4379 165894 4425 165946
rect 4449 165894 4495 165946
rect 4495 165894 4505 165946
rect 4529 165894 4559 165946
rect 4559 165894 4585 165946
rect 4289 165892 4345 165894
rect 4369 165892 4425 165894
rect 4449 165892 4505 165894
rect 4529 165892 4585 165894
rect 4289 164858 4345 164860
rect 4369 164858 4425 164860
rect 4449 164858 4505 164860
rect 4529 164858 4585 164860
rect 4289 164806 4315 164858
rect 4315 164806 4345 164858
rect 4369 164806 4379 164858
rect 4379 164806 4425 164858
rect 4449 164806 4495 164858
rect 4495 164806 4505 164858
rect 4529 164806 4559 164858
rect 4559 164806 4585 164858
rect 4289 164804 4345 164806
rect 4369 164804 4425 164806
rect 4449 164804 4505 164806
rect 4529 164804 4585 164806
rect 4289 163770 4345 163772
rect 4369 163770 4425 163772
rect 4449 163770 4505 163772
rect 4529 163770 4585 163772
rect 4289 163718 4315 163770
rect 4315 163718 4345 163770
rect 4369 163718 4379 163770
rect 4379 163718 4425 163770
rect 4449 163718 4495 163770
rect 4495 163718 4505 163770
rect 4529 163718 4559 163770
rect 4559 163718 4585 163770
rect 4289 163716 4345 163718
rect 4369 163716 4425 163718
rect 4449 163716 4505 163718
rect 4529 163716 4585 163718
rect 4289 162682 4345 162684
rect 4369 162682 4425 162684
rect 4449 162682 4505 162684
rect 4529 162682 4585 162684
rect 4289 162630 4315 162682
rect 4315 162630 4345 162682
rect 4369 162630 4379 162682
rect 4379 162630 4425 162682
rect 4449 162630 4495 162682
rect 4495 162630 4505 162682
rect 4529 162630 4559 162682
rect 4559 162630 4585 162682
rect 4289 162628 4345 162630
rect 4369 162628 4425 162630
rect 4449 162628 4505 162630
rect 4529 162628 4585 162630
rect 4289 161594 4345 161596
rect 4369 161594 4425 161596
rect 4449 161594 4505 161596
rect 4529 161594 4585 161596
rect 4289 161542 4315 161594
rect 4315 161542 4345 161594
rect 4369 161542 4379 161594
rect 4379 161542 4425 161594
rect 4449 161542 4495 161594
rect 4495 161542 4505 161594
rect 4529 161542 4559 161594
rect 4559 161542 4585 161594
rect 4289 161540 4345 161542
rect 4369 161540 4425 161542
rect 4449 161540 4505 161542
rect 4529 161540 4585 161542
rect 4289 160506 4345 160508
rect 4369 160506 4425 160508
rect 4449 160506 4505 160508
rect 4529 160506 4585 160508
rect 4289 160454 4315 160506
rect 4315 160454 4345 160506
rect 4369 160454 4379 160506
rect 4379 160454 4425 160506
rect 4449 160454 4495 160506
rect 4495 160454 4505 160506
rect 4529 160454 4559 160506
rect 4559 160454 4585 160506
rect 4289 160452 4345 160454
rect 4369 160452 4425 160454
rect 4449 160452 4505 160454
rect 4529 160452 4585 160454
rect 4289 159418 4345 159420
rect 4369 159418 4425 159420
rect 4449 159418 4505 159420
rect 4529 159418 4585 159420
rect 4289 159366 4315 159418
rect 4315 159366 4345 159418
rect 4369 159366 4379 159418
rect 4379 159366 4425 159418
rect 4449 159366 4495 159418
rect 4495 159366 4505 159418
rect 4529 159366 4559 159418
rect 4559 159366 4585 159418
rect 4289 159364 4345 159366
rect 4369 159364 4425 159366
rect 4449 159364 4505 159366
rect 4529 159364 4585 159366
rect 4289 158330 4345 158332
rect 4369 158330 4425 158332
rect 4449 158330 4505 158332
rect 4529 158330 4585 158332
rect 4289 158278 4315 158330
rect 4315 158278 4345 158330
rect 4369 158278 4379 158330
rect 4379 158278 4425 158330
rect 4449 158278 4495 158330
rect 4495 158278 4505 158330
rect 4529 158278 4559 158330
rect 4559 158278 4585 158330
rect 4289 158276 4345 158278
rect 4369 158276 4425 158278
rect 4449 158276 4505 158278
rect 4529 158276 4585 158278
rect 4289 157242 4345 157244
rect 4369 157242 4425 157244
rect 4449 157242 4505 157244
rect 4529 157242 4585 157244
rect 4289 157190 4315 157242
rect 4315 157190 4345 157242
rect 4369 157190 4379 157242
rect 4379 157190 4425 157242
rect 4449 157190 4495 157242
rect 4495 157190 4505 157242
rect 4529 157190 4559 157242
rect 4559 157190 4585 157242
rect 4289 157188 4345 157190
rect 4369 157188 4425 157190
rect 4449 157188 4505 157190
rect 4529 157188 4585 157190
rect 4289 156154 4345 156156
rect 4369 156154 4425 156156
rect 4449 156154 4505 156156
rect 4529 156154 4585 156156
rect 4289 156102 4315 156154
rect 4315 156102 4345 156154
rect 4369 156102 4379 156154
rect 4379 156102 4425 156154
rect 4449 156102 4495 156154
rect 4495 156102 4505 156154
rect 4529 156102 4559 156154
rect 4559 156102 4585 156154
rect 4289 156100 4345 156102
rect 4369 156100 4425 156102
rect 4449 156100 4505 156102
rect 4529 156100 4585 156102
rect 4289 155066 4345 155068
rect 4369 155066 4425 155068
rect 4449 155066 4505 155068
rect 4529 155066 4585 155068
rect 4289 155014 4315 155066
rect 4315 155014 4345 155066
rect 4369 155014 4379 155066
rect 4379 155014 4425 155066
rect 4449 155014 4495 155066
rect 4495 155014 4505 155066
rect 4529 155014 4559 155066
rect 4559 155014 4585 155066
rect 4289 155012 4345 155014
rect 4369 155012 4425 155014
rect 4449 155012 4505 155014
rect 4529 155012 4585 155014
rect 4289 153978 4345 153980
rect 4369 153978 4425 153980
rect 4449 153978 4505 153980
rect 4529 153978 4585 153980
rect 4289 153926 4315 153978
rect 4315 153926 4345 153978
rect 4369 153926 4379 153978
rect 4379 153926 4425 153978
rect 4449 153926 4495 153978
rect 4495 153926 4505 153978
rect 4529 153926 4559 153978
rect 4559 153926 4585 153978
rect 4289 153924 4345 153926
rect 4369 153924 4425 153926
rect 4449 153924 4505 153926
rect 4529 153924 4585 153926
rect 4289 152890 4345 152892
rect 4369 152890 4425 152892
rect 4449 152890 4505 152892
rect 4529 152890 4585 152892
rect 4289 152838 4315 152890
rect 4315 152838 4345 152890
rect 4369 152838 4379 152890
rect 4379 152838 4425 152890
rect 4449 152838 4495 152890
rect 4495 152838 4505 152890
rect 4529 152838 4559 152890
rect 4559 152838 4585 152890
rect 4289 152836 4345 152838
rect 4369 152836 4425 152838
rect 4449 152836 4505 152838
rect 4529 152836 4585 152838
rect 4289 151802 4345 151804
rect 4369 151802 4425 151804
rect 4449 151802 4505 151804
rect 4529 151802 4585 151804
rect 4289 151750 4315 151802
rect 4315 151750 4345 151802
rect 4369 151750 4379 151802
rect 4379 151750 4425 151802
rect 4449 151750 4495 151802
rect 4495 151750 4505 151802
rect 4529 151750 4559 151802
rect 4559 151750 4585 151802
rect 4289 151748 4345 151750
rect 4369 151748 4425 151750
rect 4449 151748 4505 151750
rect 4529 151748 4585 151750
rect 4289 150714 4345 150716
rect 4369 150714 4425 150716
rect 4449 150714 4505 150716
rect 4529 150714 4585 150716
rect 4289 150662 4315 150714
rect 4315 150662 4345 150714
rect 4369 150662 4379 150714
rect 4379 150662 4425 150714
rect 4449 150662 4495 150714
rect 4495 150662 4505 150714
rect 4529 150662 4559 150714
rect 4559 150662 4585 150714
rect 4289 150660 4345 150662
rect 4369 150660 4425 150662
rect 4449 150660 4505 150662
rect 4529 150660 4585 150662
rect 4289 149626 4345 149628
rect 4369 149626 4425 149628
rect 4449 149626 4505 149628
rect 4529 149626 4585 149628
rect 4289 149574 4315 149626
rect 4315 149574 4345 149626
rect 4369 149574 4379 149626
rect 4379 149574 4425 149626
rect 4449 149574 4495 149626
rect 4495 149574 4505 149626
rect 4529 149574 4559 149626
rect 4559 149574 4585 149626
rect 4289 149572 4345 149574
rect 4369 149572 4425 149574
rect 4449 149572 4505 149574
rect 4529 149572 4585 149574
rect 4289 148538 4345 148540
rect 4369 148538 4425 148540
rect 4449 148538 4505 148540
rect 4529 148538 4585 148540
rect 4289 148486 4315 148538
rect 4315 148486 4345 148538
rect 4369 148486 4379 148538
rect 4379 148486 4425 148538
rect 4449 148486 4495 148538
rect 4495 148486 4505 148538
rect 4529 148486 4559 148538
rect 4559 148486 4585 148538
rect 4289 148484 4345 148486
rect 4369 148484 4425 148486
rect 4449 148484 4505 148486
rect 4529 148484 4585 148486
rect 4289 147450 4345 147452
rect 4369 147450 4425 147452
rect 4449 147450 4505 147452
rect 4529 147450 4585 147452
rect 4289 147398 4315 147450
rect 4315 147398 4345 147450
rect 4369 147398 4379 147450
rect 4379 147398 4425 147450
rect 4449 147398 4495 147450
rect 4495 147398 4505 147450
rect 4529 147398 4559 147450
rect 4559 147398 4585 147450
rect 4289 147396 4345 147398
rect 4369 147396 4425 147398
rect 4449 147396 4505 147398
rect 4529 147396 4585 147398
rect 4289 146362 4345 146364
rect 4369 146362 4425 146364
rect 4449 146362 4505 146364
rect 4529 146362 4585 146364
rect 4289 146310 4315 146362
rect 4315 146310 4345 146362
rect 4369 146310 4379 146362
rect 4379 146310 4425 146362
rect 4449 146310 4495 146362
rect 4495 146310 4505 146362
rect 4529 146310 4559 146362
rect 4559 146310 4585 146362
rect 4289 146308 4345 146310
rect 4369 146308 4425 146310
rect 4449 146308 4505 146310
rect 4529 146308 4585 146310
rect 4289 145274 4345 145276
rect 4369 145274 4425 145276
rect 4449 145274 4505 145276
rect 4529 145274 4585 145276
rect 4289 145222 4315 145274
rect 4315 145222 4345 145274
rect 4369 145222 4379 145274
rect 4379 145222 4425 145274
rect 4449 145222 4495 145274
rect 4495 145222 4505 145274
rect 4529 145222 4559 145274
rect 4559 145222 4585 145274
rect 4289 145220 4345 145222
rect 4369 145220 4425 145222
rect 4449 145220 4505 145222
rect 4529 145220 4585 145222
rect 4289 144186 4345 144188
rect 4369 144186 4425 144188
rect 4449 144186 4505 144188
rect 4529 144186 4585 144188
rect 4289 144134 4315 144186
rect 4315 144134 4345 144186
rect 4369 144134 4379 144186
rect 4379 144134 4425 144186
rect 4449 144134 4495 144186
rect 4495 144134 4505 144186
rect 4529 144134 4559 144186
rect 4559 144134 4585 144186
rect 4289 144132 4345 144134
rect 4369 144132 4425 144134
rect 4449 144132 4505 144134
rect 4529 144132 4585 144134
rect 4289 143098 4345 143100
rect 4369 143098 4425 143100
rect 4449 143098 4505 143100
rect 4529 143098 4585 143100
rect 4289 143046 4315 143098
rect 4315 143046 4345 143098
rect 4369 143046 4379 143098
rect 4379 143046 4425 143098
rect 4449 143046 4495 143098
rect 4495 143046 4505 143098
rect 4529 143046 4559 143098
rect 4559 143046 4585 143098
rect 4289 143044 4345 143046
rect 4369 143044 4425 143046
rect 4449 143044 4505 143046
rect 4529 143044 4585 143046
rect 4289 142010 4345 142012
rect 4369 142010 4425 142012
rect 4449 142010 4505 142012
rect 4529 142010 4585 142012
rect 4289 141958 4315 142010
rect 4315 141958 4345 142010
rect 4369 141958 4379 142010
rect 4379 141958 4425 142010
rect 4449 141958 4495 142010
rect 4495 141958 4505 142010
rect 4529 141958 4559 142010
rect 4559 141958 4585 142010
rect 4289 141956 4345 141958
rect 4369 141956 4425 141958
rect 4449 141956 4505 141958
rect 4529 141956 4585 141958
rect 4289 140922 4345 140924
rect 4369 140922 4425 140924
rect 4449 140922 4505 140924
rect 4529 140922 4585 140924
rect 4289 140870 4315 140922
rect 4315 140870 4345 140922
rect 4369 140870 4379 140922
rect 4379 140870 4425 140922
rect 4449 140870 4495 140922
rect 4495 140870 4505 140922
rect 4529 140870 4559 140922
rect 4559 140870 4585 140922
rect 4289 140868 4345 140870
rect 4369 140868 4425 140870
rect 4449 140868 4505 140870
rect 4529 140868 4585 140870
rect 4289 139834 4345 139836
rect 4369 139834 4425 139836
rect 4449 139834 4505 139836
rect 4529 139834 4585 139836
rect 4289 139782 4315 139834
rect 4315 139782 4345 139834
rect 4369 139782 4379 139834
rect 4379 139782 4425 139834
rect 4449 139782 4495 139834
rect 4495 139782 4505 139834
rect 4529 139782 4559 139834
rect 4559 139782 4585 139834
rect 4289 139780 4345 139782
rect 4369 139780 4425 139782
rect 4449 139780 4505 139782
rect 4529 139780 4585 139782
rect 4289 138746 4345 138748
rect 4369 138746 4425 138748
rect 4449 138746 4505 138748
rect 4529 138746 4585 138748
rect 4289 138694 4315 138746
rect 4315 138694 4345 138746
rect 4369 138694 4379 138746
rect 4379 138694 4425 138746
rect 4449 138694 4495 138746
rect 4495 138694 4505 138746
rect 4529 138694 4559 138746
rect 4559 138694 4585 138746
rect 4289 138692 4345 138694
rect 4369 138692 4425 138694
rect 4449 138692 4505 138694
rect 4529 138692 4585 138694
rect 4289 137658 4345 137660
rect 4369 137658 4425 137660
rect 4449 137658 4505 137660
rect 4529 137658 4585 137660
rect 4289 137606 4315 137658
rect 4315 137606 4345 137658
rect 4369 137606 4379 137658
rect 4379 137606 4425 137658
rect 4449 137606 4495 137658
rect 4495 137606 4505 137658
rect 4529 137606 4559 137658
rect 4559 137606 4585 137658
rect 4289 137604 4345 137606
rect 4369 137604 4425 137606
rect 4449 137604 4505 137606
rect 4529 137604 4585 137606
rect 4289 136570 4345 136572
rect 4369 136570 4425 136572
rect 4449 136570 4505 136572
rect 4529 136570 4585 136572
rect 4289 136518 4315 136570
rect 4315 136518 4345 136570
rect 4369 136518 4379 136570
rect 4379 136518 4425 136570
rect 4449 136518 4495 136570
rect 4495 136518 4505 136570
rect 4529 136518 4559 136570
rect 4559 136518 4585 136570
rect 4289 136516 4345 136518
rect 4369 136516 4425 136518
rect 4449 136516 4505 136518
rect 4529 136516 4585 136518
rect 4289 135482 4345 135484
rect 4369 135482 4425 135484
rect 4449 135482 4505 135484
rect 4529 135482 4585 135484
rect 4289 135430 4315 135482
rect 4315 135430 4345 135482
rect 4369 135430 4379 135482
rect 4379 135430 4425 135482
rect 4449 135430 4495 135482
rect 4495 135430 4505 135482
rect 4529 135430 4559 135482
rect 4559 135430 4585 135482
rect 4289 135428 4345 135430
rect 4369 135428 4425 135430
rect 4449 135428 4505 135430
rect 4529 135428 4585 135430
rect 4289 134394 4345 134396
rect 4369 134394 4425 134396
rect 4449 134394 4505 134396
rect 4529 134394 4585 134396
rect 4289 134342 4315 134394
rect 4315 134342 4345 134394
rect 4369 134342 4379 134394
rect 4379 134342 4425 134394
rect 4449 134342 4495 134394
rect 4495 134342 4505 134394
rect 4529 134342 4559 134394
rect 4559 134342 4585 134394
rect 4289 134340 4345 134342
rect 4369 134340 4425 134342
rect 4449 134340 4505 134342
rect 4529 134340 4585 134342
rect 4289 133306 4345 133308
rect 4369 133306 4425 133308
rect 4449 133306 4505 133308
rect 4529 133306 4585 133308
rect 4289 133254 4315 133306
rect 4315 133254 4345 133306
rect 4369 133254 4379 133306
rect 4379 133254 4425 133306
rect 4449 133254 4495 133306
rect 4495 133254 4505 133306
rect 4529 133254 4559 133306
rect 4559 133254 4585 133306
rect 4289 133252 4345 133254
rect 4369 133252 4425 133254
rect 4449 133252 4505 133254
rect 4529 133252 4585 133254
rect 4289 132218 4345 132220
rect 4369 132218 4425 132220
rect 4449 132218 4505 132220
rect 4529 132218 4585 132220
rect 4289 132166 4315 132218
rect 4315 132166 4345 132218
rect 4369 132166 4379 132218
rect 4379 132166 4425 132218
rect 4449 132166 4495 132218
rect 4495 132166 4505 132218
rect 4529 132166 4559 132218
rect 4559 132166 4585 132218
rect 4289 132164 4345 132166
rect 4369 132164 4425 132166
rect 4449 132164 4505 132166
rect 4529 132164 4585 132166
rect 4289 131130 4345 131132
rect 4369 131130 4425 131132
rect 4449 131130 4505 131132
rect 4529 131130 4585 131132
rect 4289 131078 4315 131130
rect 4315 131078 4345 131130
rect 4369 131078 4379 131130
rect 4379 131078 4425 131130
rect 4449 131078 4495 131130
rect 4495 131078 4505 131130
rect 4529 131078 4559 131130
rect 4559 131078 4585 131130
rect 4289 131076 4345 131078
rect 4369 131076 4425 131078
rect 4449 131076 4505 131078
rect 4529 131076 4585 131078
rect 4289 130042 4345 130044
rect 4369 130042 4425 130044
rect 4449 130042 4505 130044
rect 4529 130042 4585 130044
rect 4289 129990 4315 130042
rect 4315 129990 4345 130042
rect 4369 129990 4379 130042
rect 4379 129990 4425 130042
rect 4449 129990 4495 130042
rect 4495 129990 4505 130042
rect 4529 129990 4559 130042
rect 4559 129990 4585 130042
rect 4289 129988 4345 129990
rect 4369 129988 4425 129990
rect 4449 129988 4505 129990
rect 4529 129988 4585 129990
rect 4289 128954 4345 128956
rect 4369 128954 4425 128956
rect 4449 128954 4505 128956
rect 4529 128954 4585 128956
rect 4289 128902 4315 128954
rect 4315 128902 4345 128954
rect 4369 128902 4379 128954
rect 4379 128902 4425 128954
rect 4449 128902 4495 128954
rect 4495 128902 4505 128954
rect 4529 128902 4559 128954
rect 4559 128902 4585 128954
rect 4289 128900 4345 128902
rect 4369 128900 4425 128902
rect 4449 128900 4505 128902
rect 4529 128900 4585 128902
rect 4289 127866 4345 127868
rect 4369 127866 4425 127868
rect 4449 127866 4505 127868
rect 4529 127866 4585 127868
rect 4289 127814 4315 127866
rect 4315 127814 4345 127866
rect 4369 127814 4379 127866
rect 4379 127814 4425 127866
rect 4449 127814 4495 127866
rect 4495 127814 4505 127866
rect 4529 127814 4559 127866
rect 4559 127814 4585 127866
rect 4289 127812 4345 127814
rect 4369 127812 4425 127814
rect 4449 127812 4505 127814
rect 4529 127812 4585 127814
rect 4289 126778 4345 126780
rect 4369 126778 4425 126780
rect 4449 126778 4505 126780
rect 4529 126778 4585 126780
rect 4289 126726 4315 126778
rect 4315 126726 4345 126778
rect 4369 126726 4379 126778
rect 4379 126726 4425 126778
rect 4449 126726 4495 126778
rect 4495 126726 4505 126778
rect 4529 126726 4559 126778
rect 4559 126726 4585 126778
rect 4289 126724 4345 126726
rect 4369 126724 4425 126726
rect 4449 126724 4505 126726
rect 4529 126724 4585 126726
rect 4289 125690 4345 125692
rect 4369 125690 4425 125692
rect 4449 125690 4505 125692
rect 4529 125690 4585 125692
rect 4289 125638 4315 125690
rect 4315 125638 4345 125690
rect 4369 125638 4379 125690
rect 4379 125638 4425 125690
rect 4449 125638 4495 125690
rect 4495 125638 4505 125690
rect 4529 125638 4559 125690
rect 4559 125638 4585 125690
rect 4289 125636 4345 125638
rect 4369 125636 4425 125638
rect 4449 125636 4505 125638
rect 4529 125636 4585 125638
rect 4289 124602 4345 124604
rect 4369 124602 4425 124604
rect 4449 124602 4505 124604
rect 4529 124602 4585 124604
rect 4289 124550 4315 124602
rect 4315 124550 4345 124602
rect 4369 124550 4379 124602
rect 4379 124550 4425 124602
rect 4449 124550 4495 124602
rect 4495 124550 4505 124602
rect 4529 124550 4559 124602
rect 4559 124550 4585 124602
rect 4289 124548 4345 124550
rect 4369 124548 4425 124550
rect 4449 124548 4505 124550
rect 4529 124548 4585 124550
rect 4289 123514 4345 123516
rect 4369 123514 4425 123516
rect 4449 123514 4505 123516
rect 4529 123514 4585 123516
rect 4289 123462 4315 123514
rect 4315 123462 4345 123514
rect 4369 123462 4379 123514
rect 4379 123462 4425 123514
rect 4449 123462 4495 123514
rect 4495 123462 4505 123514
rect 4529 123462 4559 123514
rect 4559 123462 4585 123514
rect 4289 123460 4345 123462
rect 4369 123460 4425 123462
rect 4449 123460 4505 123462
rect 4529 123460 4585 123462
rect 4289 122426 4345 122428
rect 4369 122426 4425 122428
rect 4449 122426 4505 122428
rect 4529 122426 4585 122428
rect 4289 122374 4315 122426
rect 4315 122374 4345 122426
rect 4369 122374 4379 122426
rect 4379 122374 4425 122426
rect 4449 122374 4495 122426
rect 4495 122374 4505 122426
rect 4529 122374 4559 122426
rect 4559 122374 4585 122426
rect 4289 122372 4345 122374
rect 4369 122372 4425 122374
rect 4449 122372 4505 122374
rect 4529 122372 4585 122374
rect 4289 121338 4345 121340
rect 4369 121338 4425 121340
rect 4449 121338 4505 121340
rect 4529 121338 4585 121340
rect 4289 121286 4315 121338
rect 4315 121286 4345 121338
rect 4369 121286 4379 121338
rect 4379 121286 4425 121338
rect 4449 121286 4495 121338
rect 4495 121286 4505 121338
rect 4529 121286 4559 121338
rect 4559 121286 4585 121338
rect 4289 121284 4345 121286
rect 4369 121284 4425 121286
rect 4449 121284 4505 121286
rect 4529 121284 4585 121286
rect 4289 120250 4345 120252
rect 4369 120250 4425 120252
rect 4449 120250 4505 120252
rect 4529 120250 4585 120252
rect 4289 120198 4315 120250
rect 4315 120198 4345 120250
rect 4369 120198 4379 120250
rect 4379 120198 4425 120250
rect 4449 120198 4495 120250
rect 4495 120198 4505 120250
rect 4529 120198 4559 120250
rect 4559 120198 4585 120250
rect 4289 120196 4345 120198
rect 4369 120196 4425 120198
rect 4449 120196 4505 120198
rect 4529 120196 4585 120198
rect 4289 119162 4345 119164
rect 4369 119162 4425 119164
rect 4449 119162 4505 119164
rect 4529 119162 4585 119164
rect 4289 119110 4315 119162
rect 4315 119110 4345 119162
rect 4369 119110 4379 119162
rect 4379 119110 4425 119162
rect 4449 119110 4495 119162
rect 4495 119110 4505 119162
rect 4529 119110 4559 119162
rect 4559 119110 4585 119162
rect 4289 119108 4345 119110
rect 4369 119108 4425 119110
rect 4449 119108 4505 119110
rect 4529 119108 4585 119110
rect 4289 118074 4345 118076
rect 4369 118074 4425 118076
rect 4449 118074 4505 118076
rect 4529 118074 4585 118076
rect 4289 118022 4315 118074
rect 4315 118022 4345 118074
rect 4369 118022 4379 118074
rect 4379 118022 4425 118074
rect 4449 118022 4495 118074
rect 4495 118022 4505 118074
rect 4529 118022 4559 118074
rect 4559 118022 4585 118074
rect 4289 118020 4345 118022
rect 4369 118020 4425 118022
rect 4449 118020 4505 118022
rect 4529 118020 4585 118022
rect 4289 116986 4345 116988
rect 4369 116986 4425 116988
rect 4449 116986 4505 116988
rect 4529 116986 4585 116988
rect 4289 116934 4315 116986
rect 4315 116934 4345 116986
rect 4369 116934 4379 116986
rect 4379 116934 4425 116986
rect 4449 116934 4495 116986
rect 4495 116934 4505 116986
rect 4529 116934 4559 116986
rect 4559 116934 4585 116986
rect 4289 116932 4345 116934
rect 4369 116932 4425 116934
rect 4449 116932 4505 116934
rect 4529 116932 4585 116934
rect 4289 115898 4345 115900
rect 4369 115898 4425 115900
rect 4449 115898 4505 115900
rect 4529 115898 4585 115900
rect 4289 115846 4315 115898
rect 4315 115846 4345 115898
rect 4369 115846 4379 115898
rect 4379 115846 4425 115898
rect 4449 115846 4495 115898
rect 4495 115846 4505 115898
rect 4529 115846 4559 115898
rect 4559 115846 4585 115898
rect 4289 115844 4345 115846
rect 4369 115844 4425 115846
rect 4449 115844 4505 115846
rect 4529 115844 4585 115846
rect 4289 114810 4345 114812
rect 4369 114810 4425 114812
rect 4449 114810 4505 114812
rect 4529 114810 4585 114812
rect 4289 114758 4315 114810
rect 4315 114758 4345 114810
rect 4369 114758 4379 114810
rect 4379 114758 4425 114810
rect 4449 114758 4495 114810
rect 4495 114758 4505 114810
rect 4529 114758 4559 114810
rect 4559 114758 4585 114810
rect 4289 114756 4345 114758
rect 4369 114756 4425 114758
rect 4449 114756 4505 114758
rect 4529 114756 4585 114758
rect 4289 113722 4345 113724
rect 4369 113722 4425 113724
rect 4449 113722 4505 113724
rect 4529 113722 4585 113724
rect 4289 113670 4315 113722
rect 4315 113670 4345 113722
rect 4369 113670 4379 113722
rect 4379 113670 4425 113722
rect 4449 113670 4495 113722
rect 4495 113670 4505 113722
rect 4529 113670 4559 113722
rect 4559 113670 4585 113722
rect 4289 113668 4345 113670
rect 4369 113668 4425 113670
rect 4449 113668 4505 113670
rect 4529 113668 4585 113670
rect 4289 112634 4345 112636
rect 4369 112634 4425 112636
rect 4449 112634 4505 112636
rect 4529 112634 4585 112636
rect 4289 112582 4315 112634
rect 4315 112582 4345 112634
rect 4369 112582 4379 112634
rect 4379 112582 4425 112634
rect 4449 112582 4495 112634
rect 4495 112582 4505 112634
rect 4529 112582 4559 112634
rect 4559 112582 4585 112634
rect 4289 112580 4345 112582
rect 4369 112580 4425 112582
rect 4449 112580 4505 112582
rect 4529 112580 4585 112582
rect 4289 111546 4345 111548
rect 4369 111546 4425 111548
rect 4449 111546 4505 111548
rect 4529 111546 4585 111548
rect 4289 111494 4315 111546
rect 4315 111494 4345 111546
rect 4369 111494 4379 111546
rect 4379 111494 4425 111546
rect 4449 111494 4495 111546
rect 4495 111494 4505 111546
rect 4529 111494 4559 111546
rect 4559 111494 4585 111546
rect 4289 111492 4345 111494
rect 4369 111492 4425 111494
rect 4449 111492 4505 111494
rect 4529 111492 4585 111494
rect 4289 110458 4345 110460
rect 4369 110458 4425 110460
rect 4449 110458 4505 110460
rect 4529 110458 4585 110460
rect 4289 110406 4315 110458
rect 4315 110406 4345 110458
rect 4369 110406 4379 110458
rect 4379 110406 4425 110458
rect 4449 110406 4495 110458
rect 4495 110406 4505 110458
rect 4529 110406 4559 110458
rect 4559 110406 4585 110458
rect 4289 110404 4345 110406
rect 4369 110404 4425 110406
rect 4449 110404 4505 110406
rect 4529 110404 4585 110406
rect 4289 109370 4345 109372
rect 4369 109370 4425 109372
rect 4449 109370 4505 109372
rect 4529 109370 4585 109372
rect 4289 109318 4315 109370
rect 4315 109318 4345 109370
rect 4369 109318 4379 109370
rect 4379 109318 4425 109370
rect 4449 109318 4495 109370
rect 4495 109318 4505 109370
rect 4529 109318 4559 109370
rect 4559 109318 4585 109370
rect 4289 109316 4345 109318
rect 4369 109316 4425 109318
rect 4449 109316 4505 109318
rect 4529 109316 4585 109318
rect 4289 108282 4345 108284
rect 4369 108282 4425 108284
rect 4449 108282 4505 108284
rect 4529 108282 4585 108284
rect 4289 108230 4315 108282
rect 4315 108230 4345 108282
rect 4369 108230 4379 108282
rect 4379 108230 4425 108282
rect 4449 108230 4495 108282
rect 4495 108230 4505 108282
rect 4529 108230 4559 108282
rect 4559 108230 4585 108282
rect 4289 108228 4345 108230
rect 4369 108228 4425 108230
rect 4449 108228 4505 108230
rect 4529 108228 4585 108230
rect 4289 107194 4345 107196
rect 4369 107194 4425 107196
rect 4449 107194 4505 107196
rect 4529 107194 4585 107196
rect 4289 107142 4315 107194
rect 4315 107142 4345 107194
rect 4369 107142 4379 107194
rect 4379 107142 4425 107194
rect 4449 107142 4495 107194
rect 4495 107142 4505 107194
rect 4529 107142 4559 107194
rect 4559 107142 4585 107194
rect 4289 107140 4345 107142
rect 4369 107140 4425 107142
rect 4449 107140 4505 107142
rect 4529 107140 4585 107142
rect 4289 106106 4345 106108
rect 4369 106106 4425 106108
rect 4449 106106 4505 106108
rect 4529 106106 4585 106108
rect 4289 106054 4315 106106
rect 4315 106054 4345 106106
rect 4369 106054 4379 106106
rect 4379 106054 4425 106106
rect 4449 106054 4495 106106
rect 4495 106054 4505 106106
rect 4529 106054 4559 106106
rect 4559 106054 4585 106106
rect 4289 106052 4345 106054
rect 4369 106052 4425 106054
rect 4449 106052 4505 106054
rect 4529 106052 4585 106054
rect 4289 105018 4345 105020
rect 4369 105018 4425 105020
rect 4449 105018 4505 105020
rect 4529 105018 4585 105020
rect 4289 104966 4315 105018
rect 4315 104966 4345 105018
rect 4369 104966 4379 105018
rect 4379 104966 4425 105018
rect 4449 104966 4495 105018
rect 4495 104966 4505 105018
rect 4529 104966 4559 105018
rect 4559 104966 4585 105018
rect 4289 104964 4345 104966
rect 4369 104964 4425 104966
rect 4449 104964 4505 104966
rect 4529 104964 4585 104966
rect 4289 103930 4345 103932
rect 4369 103930 4425 103932
rect 4449 103930 4505 103932
rect 4529 103930 4585 103932
rect 4289 103878 4315 103930
rect 4315 103878 4345 103930
rect 4369 103878 4379 103930
rect 4379 103878 4425 103930
rect 4449 103878 4495 103930
rect 4495 103878 4505 103930
rect 4529 103878 4559 103930
rect 4559 103878 4585 103930
rect 4289 103876 4345 103878
rect 4369 103876 4425 103878
rect 4449 103876 4505 103878
rect 4529 103876 4585 103878
rect 4289 102842 4345 102844
rect 4369 102842 4425 102844
rect 4449 102842 4505 102844
rect 4529 102842 4585 102844
rect 4289 102790 4315 102842
rect 4315 102790 4345 102842
rect 4369 102790 4379 102842
rect 4379 102790 4425 102842
rect 4449 102790 4495 102842
rect 4495 102790 4505 102842
rect 4529 102790 4559 102842
rect 4559 102790 4585 102842
rect 4289 102788 4345 102790
rect 4369 102788 4425 102790
rect 4449 102788 4505 102790
rect 4529 102788 4585 102790
rect 4289 101754 4345 101756
rect 4369 101754 4425 101756
rect 4449 101754 4505 101756
rect 4529 101754 4585 101756
rect 4289 101702 4315 101754
rect 4315 101702 4345 101754
rect 4369 101702 4379 101754
rect 4379 101702 4425 101754
rect 4449 101702 4495 101754
rect 4495 101702 4505 101754
rect 4529 101702 4559 101754
rect 4559 101702 4585 101754
rect 4289 101700 4345 101702
rect 4369 101700 4425 101702
rect 4449 101700 4505 101702
rect 4529 101700 4585 101702
rect 4289 100666 4345 100668
rect 4369 100666 4425 100668
rect 4449 100666 4505 100668
rect 4529 100666 4585 100668
rect 4289 100614 4315 100666
rect 4315 100614 4345 100666
rect 4369 100614 4379 100666
rect 4379 100614 4425 100666
rect 4449 100614 4495 100666
rect 4495 100614 4505 100666
rect 4529 100614 4559 100666
rect 4559 100614 4585 100666
rect 4289 100612 4345 100614
rect 4369 100612 4425 100614
rect 4449 100612 4505 100614
rect 4529 100612 4585 100614
rect 4289 99578 4345 99580
rect 4369 99578 4425 99580
rect 4449 99578 4505 99580
rect 4529 99578 4585 99580
rect 4289 99526 4315 99578
rect 4315 99526 4345 99578
rect 4369 99526 4379 99578
rect 4379 99526 4425 99578
rect 4449 99526 4495 99578
rect 4495 99526 4505 99578
rect 4529 99526 4559 99578
rect 4559 99526 4585 99578
rect 4289 99524 4345 99526
rect 4369 99524 4425 99526
rect 4449 99524 4505 99526
rect 4529 99524 4585 99526
rect 4289 98490 4345 98492
rect 4369 98490 4425 98492
rect 4449 98490 4505 98492
rect 4529 98490 4585 98492
rect 4289 98438 4315 98490
rect 4315 98438 4345 98490
rect 4369 98438 4379 98490
rect 4379 98438 4425 98490
rect 4449 98438 4495 98490
rect 4495 98438 4505 98490
rect 4529 98438 4559 98490
rect 4559 98438 4585 98490
rect 4289 98436 4345 98438
rect 4369 98436 4425 98438
rect 4449 98436 4505 98438
rect 4529 98436 4585 98438
rect 4289 97402 4345 97404
rect 4369 97402 4425 97404
rect 4449 97402 4505 97404
rect 4529 97402 4585 97404
rect 4289 97350 4315 97402
rect 4315 97350 4345 97402
rect 4369 97350 4379 97402
rect 4379 97350 4425 97402
rect 4449 97350 4495 97402
rect 4495 97350 4505 97402
rect 4529 97350 4559 97402
rect 4559 97350 4585 97402
rect 4289 97348 4345 97350
rect 4369 97348 4425 97350
rect 4449 97348 4505 97350
rect 4529 97348 4585 97350
rect 4289 96314 4345 96316
rect 4369 96314 4425 96316
rect 4449 96314 4505 96316
rect 4529 96314 4585 96316
rect 4289 96262 4315 96314
rect 4315 96262 4345 96314
rect 4369 96262 4379 96314
rect 4379 96262 4425 96314
rect 4449 96262 4495 96314
rect 4495 96262 4505 96314
rect 4529 96262 4559 96314
rect 4559 96262 4585 96314
rect 4289 96260 4345 96262
rect 4369 96260 4425 96262
rect 4449 96260 4505 96262
rect 4529 96260 4585 96262
rect 4289 95226 4345 95228
rect 4369 95226 4425 95228
rect 4449 95226 4505 95228
rect 4529 95226 4585 95228
rect 4289 95174 4315 95226
rect 4315 95174 4345 95226
rect 4369 95174 4379 95226
rect 4379 95174 4425 95226
rect 4449 95174 4495 95226
rect 4495 95174 4505 95226
rect 4529 95174 4559 95226
rect 4559 95174 4585 95226
rect 4289 95172 4345 95174
rect 4369 95172 4425 95174
rect 4449 95172 4505 95174
rect 4529 95172 4585 95174
rect 4289 94138 4345 94140
rect 4369 94138 4425 94140
rect 4449 94138 4505 94140
rect 4529 94138 4585 94140
rect 4289 94086 4315 94138
rect 4315 94086 4345 94138
rect 4369 94086 4379 94138
rect 4379 94086 4425 94138
rect 4449 94086 4495 94138
rect 4495 94086 4505 94138
rect 4529 94086 4559 94138
rect 4559 94086 4585 94138
rect 4289 94084 4345 94086
rect 4369 94084 4425 94086
rect 4449 94084 4505 94086
rect 4529 94084 4585 94086
rect 4289 93050 4345 93052
rect 4369 93050 4425 93052
rect 4449 93050 4505 93052
rect 4529 93050 4585 93052
rect 4289 92998 4315 93050
rect 4315 92998 4345 93050
rect 4369 92998 4379 93050
rect 4379 92998 4425 93050
rect 4449 92998 4495 93050
rect 4495 92998 4505 93050
rect 4529 92998 4559 93050
rect 4559 92998 4585 93050
rect 4289 92996 4345 92998
rect 4369 92996 4425 92998
rect 4449 92996 4505 92998
rect 4529 92996 4585 92998
rect 4289 91962 4345 91964
rect 4369 91962 4425 91964
rect 4449 91962 4505 91964
rect 4529 91962 4585 91964
rect 4289 91910 4315 91962
rect 4315 91910 4345 91962
rect 4369 91910 4379 91962
rect 4379 91910 4425 91962
rect 4449 91910 4495 91962
rect 4495 91910 4505 91962
rect 4529 91910 4559 91962
rect 4559 91910 4585 91962
rect 4289 91908 4345 91910
rect 4369 91908 4425 91910
rect 4449 91908 4505 91910
rect 4529 91908 4585 91910
rect 4289 90874 4345 90876
rect 4369 90874 4425 90876
rect 4449 90874 4505 90876
rect 4529 90874 4585 90876
rect 4289 90822 4315 90874
rect 4315 90822 4345 90874
rect 4369 90822 4379 90874
rect 4379 90822 4425 90874
rect 4449 90822 4495 90874
rect 4495 90822 4505 90874
rect 4529 90822 4559 90874
rect 4559 90822 4585 90874
rect 4289 90820 4345 90822
rect 4369 90820 4425 90822
rect 4449 90820 4505 90822
rect 4529 90820 4585 90822
rect 4289 89786 4345 89788
rect 4369 89786 4425 89788
rect 4449 89786 4505 89788
rect 4529 89786 4585 89788
rect 4289 89734 4315 89786
rect 4315 89734 4345 89786
rect 4369 89734 4379 89786
rect 4379 89734 4425 89786
rect 4449 89734 4495 89786
rect 4495 89734 4505 89786
rect 4529 89734 4559 89786
rect 4559 89734 4585 89786
rect 4289 89732 4345 89734
rect 4369 89732 4425 89734
rect 4449 89732 4505 89734
rect 4529 89732 4585 89734
rect 4289 88698 4345 88700
rect 4369 88698 4425 88700
rect 4449 88698 4505 88700
rect 4529 88698 4585 88700
rect 4289 88646 4315 88698
rect 4315 88646 4345 88698
rect 4369 88646 4379 88698
rect 4379 88646 4425 88698
rect 4449 88646 4495 88698
rect 4495 88646 4505 88698
rect 4529 88646 4559 88698
rect 4559 88646 4585 88698
rect 4289 88644 4345 88646
rect 4369 88644 4425 88646
rect 4449 88644 4505 88646
rect 4529 88644 4585 88646
rect 4289 87610 4345 87612
rect 4369 87610 4425 87612
rect 4449 87610 4505 87612
rect 4529 87610 4585 87612
rect 4289 87558 4315 87610
rect 4315 87558 4345 87610
rect 4369 87558 4379 87610
rect 4379 87558 4425 87610
rect 4449 87558 4495 87610
rect 4495 87558 4505 87610
rect 4529 87558 4559 87610
rect 4559 87558 4585 87610
rect 4289 87556 4345 87558
rect 4369 87556 4425 87558
rect 4449 87556 4505 87558
rect 4529 87556 4585 87558
rect 4289 86522 4345 86524
rect 4369 86522 4425 86524
rect 4449 86522 4505 86524
rect 4529 86522 4585 86524
rect 4289 86470 4315 86522
rect 4315 86470 4345 86522
rect 4369 86470 4379 86522
rect 4379 86470 4425 86522
rect 4449 86470 4495 86522
rect 4495 86470 4505 86522
rect 4529 86470 4559 86522
rect 4559 86470 4585 86522
rect 4289 86468 4345 86470
rect 4369 86468 4425 86470
rect 4449 86468 4505 86470
rect 4529 86468 4585 86470
rect 4289 85434 4345 85436
rect 4369 85434 4425 85436
rect 4449 85434 4505 85436
rect 4529 85434 4585 85436
rect 4289 85382 4315 85434
rect 4315 85382 4345 85434
rect 4369 85382 4379 85434
rect 4379 85382 4425 85434
rect 4449 85382 4495 85434
rect 4495 85382 4505 85434
rect 4529 85382 4559 85434
rect 4559 85382 4585 85434
rect 4289 85380 4345 85382
rect 4369 85380 4425 85382
rect 4449 85380 4505 85382
rect 4529 85380 4585 85382
rect 4289 84346 4345 84348
rect 4369 84346 4425 84348
rect 4449 84346 4505 84348
rect 4529 84346 4585 84348
rect 4289 84294 4315 84346
rect 4315 84294 4345 84346
rect 4369 84294 4379 84346
rect 4379 84294 4425 84346
rect 4449 84294 4495 84346
rect 4495 84294 4505 84346
rect 4529 84294 4559 84346
rect 4559 84294 4585 84346
rect 4289 84292 4345 84294
rect 4369 84292 4425 84294
rect 4449 84292 4505 84294
rect 4529 84292 4585 84294
rect 4289 83258 4345 83260
rect 4369 83258 4425 83260
rect 4449 83258 4505 83260
rect 4529 83258 4585 83260
rect 4289 83206 4315 83258
rect 4315 83206 4345 83258
rect 4369 83206 4379 83258
rect 4379 83206 4425 83258
rect 4449 83206 4495 83258
rect 4495 83206 4505 83258
rect 4529 83206 4559 83258
rect 4559 83206 4585 83258
rect 4289 83204 4345 83206
rect 4369 83204 4425 83206
rect 4449 83204 4505 83206
rect 4529 83204 4585 83206
rect 4289 82170 4345 82172
rect 4369 82170 4425 82172
rect 4449 82170 4505 82172
rect 4529 82170 4585 82172
rect 4289 82118 4315 82170
rect 4315 82118 4345 82170
rect 4369 82118 4379 82170
rect 4379 82118 4425 82170
rect 4449 82118 4495 82170
rect 4495 82118 4505 82170
rect 4529 82118 4559 82170
rect 4559 82118 4585 82170
rect 4289 82116 4345 82118
rect 4369 82116 4425 82118
rect 4449 82116 4505 82118
rect 4529 82116 4585 82118
rect 4289 81082 4345 81084
rect 4369 81082 4425 81084
rect 4449 81082 4505 81084
rect 4529 81082 4585 81084
rect 4289 81030 4315 81082
rect 4315 81030 4345 81082
rect 4369 81030 4379 81082
rect 4379 81030 4425 81082
rect 4449 81030 4495 81082
rect 4495 81030 4505 81082
rect 4529 81030 4559 81082
rect 4559 81030 4585 81082
rect 4289 81028 4345 81030
rect 4369 81028 4425 81030
rect 4449 81028 4505 81030
rect 4529 81028 4585 81030
rect 4289 79994 4345 79996
rect 4369 79994 4425 79996
rect 4449 79994 4505 79996
rect 4529 79994 4585 79996
rect 4289 79942 4315 79994
rect 4315 79942 4345 79994
rect 4369 79942 4379 79994
rect 4379 79942 4425 79994
rect 4449 79942 4495 79994
rect 4495 79942 4505 79994
rect 4529 79942 4559 79994
rect 4559 79942 4585 79994
rect 4289 79940 4345 79942
rect 4369 79940 4425 79942
rect 4449 79940 4505 79942
rect 4529 79940 4585 79942
rect 4289 78906 4345 78908
rect 4369 78906 4425 78908
rect 4449 78906 4505 78908
rect 4529 78906 4585 78908
rect 4289 78854 4315 78906
rect 4315 78854 4345 78906
rect 4369 78854 4379 78906
rect 4379 78854 4425 78906
rect 4449 78854 4495 78906
rect 4495 78854 4505 78906
rect 4529 78854 4559 78906
rect 4559 78854 4585 78906
rect 4289 78852 4345 78854
rect 4369 78852 4425 78854
rect 4449 78852 4505 78854
rect 4529 78852 4585 78854
rect 4289 77818 4345 77820
rect 4369 77818 4425 77820
rect 4449 77818 4505 77820
rect 4529 77818 4585 77820
rect 4289 77766 4315 77818
rect 4315 77766 4345 77818
rect 4369 77766 4379 77818
rect 4379 77766 4425 77818
rect 4449 77766 4495 77818
rect 4495 77766 4505 77818
rect 4529 77766 4559 77818
rect 4559 77766 4585 77818
rect 4289 77764 4345 77766
rect 4369 77764 4425 77766
rect 4449 77764 4505 77766
rect 4529 77764 4585 77766
rect 4289 76730 4345 76732
rect 4369 76730 4425 76732
rect 4449 76730 4505 76732
rect 4529 76730 4585 76732
rect 4289 76678 4315 76730
rect 4315 76678 4345 76730
rect 4369 76678 4379 76730
rect 4379 76678 4425 76730
rect 4449 76678 4495 76730
rect 4495 76678 4505 76730
rect 4529 76678 4559 76730
rect 4559 76678 4585 76730
rect 4289 76676 4345 76678
rect 4369 76676 4425 76678
rect 4449 76676 4505 76678
rect 4529 76676 4585 76678
rect 4289 75642 4345 75644
rect 4369 75642 4425 75644
rect 4449 75642 4505 75644
rect 4529 75642 4585 75644
rect 4289 75590 4315 75642
rect 4315 75590 4345 75642
rect 4369 75590 4379 75642
rect 4379 75590 4425 75642
rect 4449 75590 4495 75642
rect 4495 75590 4505 75642
rect 4529 75590 4559 75642
rect 4559 75590 4585 75642
rect 4289 75588 4345 75590
rect 4369 75588 4425 75590
rect 4449 75588 4505 75590
rect 4529 75588 4585 75590
rect 4289 74554 4345 74556
rect 4369 74554 4425 74556
rect 4449 74554 4505 74556
rect 4529 74554 4585 74556
rect 4289 74502 4315 74554
rect 4315 74502 4345 74554
rect 4369 74502 4379 74554
rect 4379 74502 4425 74554
rect 4449 74502 4495 74554
rect 4495 74502 4505 74554
rect 4529 74502 4559 74554
rect 4559 74502 4585 74554
rect 4289 74500 4345 74502
rect 4369 74500 4425 74502
rect 4449 74500 4505 74502
rect 4529 74500 4585 74502
rect 4289 73466 4345 73468
rect 4369 73466 4425 73468
rect 4449 73466 4505 73468
rect 4529 73466 4585 73468
rect 4289 73414 4315 73466
rect 4315 73414 4345 73466
rect 4369 73414 4379 73466
rect 4379 73414 4425 73466
rect 4449 73414 4495 73466
rect 4495 73414 4505 73466
rect 4529 73414 4559 73466
rect 4559 73414 4585 73466
rect 4289 73412 4345 73414
rect 4369 73412 4425 73414
rect 4449 73412 4505 73414
rect 4529 73412 4585 73414
rect 4289 72378 4345 72380
rect 4369 72378 4425 72380
rect 4449 72378 4505 72380
rect 4529 72378 4585 72380
rect 4289 72326 4315 72378
rect 4315 72326 4345 72378
rect 4369 72326 4379 72378
rect 4379 72326 4425 72378
rect 4449 72326 4495 72378
rect 4495 72326 4505 72378
rect 4529 72326 4559 72378
rect 4559 72326 4585 72378
rect 4289 72324 4345 72326
rect 4369 72324 4425 72326
rect 4449 72324 4505 72326
rect 4529 72324 4585 72326
rect 4289 71290 4345 71292
rect 4369 71290 4425 71292
rect 4449 71290 4505 71292
rect 4529 71290 4585 71292
rect 4289 71238 4315 71290
rect 4315 71238 4345 71290
rect 4369 71238 4379 71290
rect 4379 71238 4425 71290
rect 4449 71238 4495 71290
rect 4495 71238 4505 71290
rect 4529 71238 4559 71290
rect 4559 71238 4585 71290
rect 4289 71236 4345 71238
rect 4369 71236 4425 71238
rect 4449 71236 4505 71238
rect 4529 71236 4585 71238
rect 4289 70202 4345 70204
rect 4369 70202 4425 70204
rect 4449 70202 4505 70204
rect 4529 70202 4585 70204
rect 4289 70150 4315 70202
rect 4315 70150 4345 70202
rect 4369 70150 4379 70202
rect 4379 70150 4425 70202
rect 4449 70150 4495 70202
rect 4495 70150 4505 70202
rect 4529 70150 4559 70202
rect 4559 70150 4585 70202
rect 4289 70148 4345 70150
rect 4369 70148 4425 70150
rect 4449 70148 4505 70150
rect 4529 70148 4585 70150
rect 4289 69114 4345 69116
rect 4369 69114 4425 69116
rect 4449 69114 4505 69116
rect 4529 69114 4585 69116
rect 4289 69062 4315 69114
rect 4315 69062 4345 69114
rect 4369 69062 4379 69114
rect 4379 69062 4425 69114
rect 4449 69062 4495 69114
rect 4495 69062 4505 69114
rect 4529 69062 4559 69114
rect 4559 69062 4585 69114
rect 4289 69060 4345 69062
rect 4369 69060 4425 69062
rect 4449 69060 4505 69062
rect 4529 69060 4585 69062
rect 4289 68026 4345 68028
rect 4369 68026 4425 68028
rect 4449 68026 4505 68028
rect 4529 68026 4585 68028
rect 4289 67974 4315 68026
rect 4315 67974 4345 68026
rect 4369 67974 4379 68026
rect 4379 67974 4425 68026
rect 4449 67974 4495 68026
rect 4495 67974 4505 68026
rect 4529 67974 4559 68026
rect 4559 67974 4585 68026
rect 4289 67972 4345 67974
rect 4369 67972 4425 67974
rect 4449 67972 4505 67974
rect 4529 67972 4585 67974
rect 4289 66938 4345 66940
rect 4369 66938 4425 66940
rect 4449 66938 4505 66940
rect 4529 66938 4585 66940
rect 4289 66886 4315 66938
rect 4315 66886 4345 66938
rect 4369 66886 4379 66938
rect 4379 66886 4425 66938
rect 4449 66886 4495 66938
rect 4495 66886 4505 66938
rect 4529 66886 4559 66938
rect 4559 66886 4585 66938
rect 4289 66884 4345 66886
rect 4369 66884 4425 66886
rect 4449 66884 4505 66886
rect 4529 66884 4585 66886
rect 4289 65850 4345 65852
rect 4369 65850 4425 65852
rect 4449 65850 4505 65852
rect 4529 65850 4585 65852
rect 4289 65798 4315 65850
rect 4315 65798 4345 65850
rect 4369 65798 4379 65850
rect 4379 65798 4425 65850
rect 4449 65798 4495 65850
rect 4495 65798 4505 65850
rect 4529 65798 4559 65850
rect 4559 65798 4585 65850
rect 4289 65796 4345 65798
rect 4369 65796 4425 65798
rect 4449 65796 4505 65798
rect 4529 65796 4585 65798
rect 4289 64762 4345 64764
rect 4369 64762 4425 64764
rect 4449 64762 4505 64764
rect 4529 64762 4585 64764
rect 4289 64710 4315 64762
rect 4315 64710 4345 64762
rect 4369 64710 4379 64762
rect 4379 64710 4425 64762
rect 4449 64710 4495 64762
rect 4495 64710 4505 64762
rect 4529 64710 4559 64762
rect 4559 64710 4585 64762
rect 4289 64708 4345 64710
rect 4369 64708 4425 64710
rect 4449 64708 4505 64710
rect 4529 64708 4585 64710
rect 4289 63674 4345 63676
rect 4369 63674 4425 63676
rect 4449 63674 4505 63676
rect 4529 63674 4585 63676
rect 4289 63622 4315 63674
rect 4315 63622 4345 63674
rect 4369 63622 4379 63674
rect 4379 63622 4425 63674
rect 4449 63622 4495 63674
rect 4495 63622 4505 63674
rect 4529 63622 4559 63674
rect 4559 63622 4585 63674
rect 4289 63620 4345 63622
rect 4369 63620 4425 63622
rect 4449 63620 4505 63622
rect 4529 63620 4585 63622
rect 4289 62586 4345 62588
rect 4369 62586 4425 62588
rect 4449 62586 4505 62588
rect 4529 62586 4585 62588
rect 4289 62534 4315 62586
rect 4315 62534 4345 62586
rect 4369 62534 4379 62586
rect 4379 62534 4425 62586
rect 4449 62534 4495 62586
rect 4495 62534 4505 62586
rect 4529 62534 4559 62586
rect 4559 62534 4585 62586
rect 4289 62532 4345 62534
rect 4369 62532 4425 62534
rect 4449 62532 4505 62534
rect 4529 62532 4585 62534
rect 4289 61498 4345 61500
rect 4369 61498 4425 61500
rect 4449 61498 4505 61500
rect 4529 61498 4585 61500
rect 4289 61446 4315 61498
rect 4315 61446 4345 61498
rect 4369 61446 4379 61498
rect 4379 61446 4425 61498
rect 4449 61446 4495 61498
rect 4495 61446 4505 61498
rect 4529 61446 4559 61498
rect 4559 61446 4585 61498
rect 4289 61444 4345 61446
rect 4369 61444 4425 61446
rect 4449 61444 4505 61446
rect 4529 61444 4585 61446
rect 4289 60410 4345 60412
rect 4369 60410 4425 60412
rect 4449 60410 4505 60412
rect 4529 60410 4585 60412
rect 4289 60358 4315 60410
rect 4315 60358 4345 60410
rect 4369 60358 4379 60410
rect 4379 60358 4425 60410
rect 4449 60358 4495 60410
rect 4495 60358 4505 60410
rect 4529 60358 4559 60410
rect 4559 60358 4585 60410
rect 4289 60356 4345 60358
rect 4369 60356 4425 60358
rect 4449 60356 4505 60358
rect 4529 60356 4585 60358
rect 4289 59322 4345 59324
rect 4369 59322 4425 59324
rect 4449 59322 4505 59324
rect 4529 59322 4585 59324
rect 4289 59270 4315 59322
rect 4315 59270 4345 59322
rect 4369 59270 4379 59322
rect 4379 59270 4425 59322
rect 4449 59270 4495 59322
rect 4495 59270 4505 59322
rect 4529 59270 4559 59322
rect 4559 59270 4585 59322
rect 4289 59268 4345 59270
rect 4369 59268 4425 59270
rect 4449 59268 4505 59270
rect 4529 59268 4585 59270
rect 4289 58234 4345 58236
rect 4369 58234 4425 58236
rect 4449 58234 4505 58236
rect 4529 58234 4585 58236
rect 4289 58182 4315 58234
rect 4315 58182 4345 58234
rect 4369 58182 4379 58234
rect 4379 58182 4425 58234
rect 4449 58182 4495 58234
rect 4495 58182 4505 58234
rect 4529 58182 4559 58234
rect 4559 58182 4585 58234
rect 4289 58180 4345 58182
rect 4369 58180 4425 58182
rect 4449 58180 4505 58182
rect 4529 58180 4585 58182
rect 4289 57146 4345 57148
rect 4369 57146 4425 57148
rect 4449 57146 4505 57148
rect 4529 57146 4585 57148
rect 4289 57094 4315 57146
rect 4315 57094 4345 57146
rect 4369 57094 4379 57146
rect 4379 57094 4425 57146
rect 4449 57094 4495 57146
rect 4495 57094 4505 57146
rect 4529 57094 4559 57146
rect 4559 57094 4585 57146
rect 4289 57092 4345 57094
rect 4369 57092 4425 57094
rect 4449 57092 4505 57094
rect 4529 57092 4585 57094
rect 4289 56058 4345 56060
rect 4369 56058 4425 56060
rect 4449 56058 4505 56060
rect 4529 56058 4585 56060
rect 4289 56006 4315 56058
rect 4315 56006 4345 56058
rect 4369 56006 4379 56058
rect 4379 56006 4425 56058
rect 4449 56006 4495 56058
rect 4495 56006 4505 56058
rect 4529 56006 4559 56058
rect 4559 56006 4585 56058
rect 4289 56004 4345 56006
rect 4369 56004 4425 56006
rect 4449 56004 4505 56006
rect 4529 56004 4585 56006
rect 4289 54970 4345 54972
rect 4369 54970 4425 54972
rect 4449 54970 4505 54972
rect 4529 54970 4585 54972
rect 4289 54918 4315 54970
rect 4315 54918 4345 54970
rect 4369 54918 4379 54970
rect 4379 54918 4425 54970
rect 4449 54918 4495 54970
rect 4495 54918 4505 54970
rect 4529 54918 4559 54970
rect 4559 54918 4585 54970
rect 4289 54916 4345 54918
rect 4369 54916 4425 54918
rect 4449 54916 4505 54918
rect 4529 54916 4585 54918
rect 4289 53882 4345 53884
rect 4369 53882 4425 53884
rect 4449 53882 4505 53884
rect 4529 53882 4585 53884
rect 4289 53830 4315 53882
rect 4315 53830 4345 53882
rect 4369 53830 4379 53882
rect 4379 53830 4425 53882
rect 4449 53830 4495 53882
rect 4495 53830 4505 53882
rect 4529 53830 4559 53882
rect 4559 53830 4585 53882
rect 4289 53828 4345 53830
rect 4369 53828 4425 53830
rect 4449 53828 4505 53830
rect 4529 53828 4585 53830
rect 4289 52794 4345 52796
rect 4369 52794 4425 52796
rect 4449 52794 4505 52796
rect 4529 52794 4585 52796
rect 4289 52742 4315 52794
rect 4315 52742 4345 52794
rect 4369 52742 4379 52794
rect 4379 52742 4425 52794
rect 4449 52742 4495 52794
rect 4495 52742 4505 52794
rect 4529 52742 4559 52794
rect 4559 52742 4585 52794
rect 4289 52740 4345 52742
rect 4369 52740 4425 52742
rect 4449 52740 4505 52742
rect 4529 52740 4585 52742
rect 4289 51706 4345 51708
rect 4369 51706 4425 51708
rect 4449 51706 4505 51708
rect 4529 51706 4585 51708
rect 4289 51654 4315 51706
rect 4315 51654 4345 51706
rect 4369 51654 4379 51706
rect 4379 51654 4425 51706
rect 4449 51654 4495 51706
rect 4495 51654 4505 51706
rect 4529 51654 4559 51706
rect 4559 51654 4585 51706
rect 4289 51652 4345 51654
rect 4369 51652 4425 51654
rect 4449 51652 4505 51654
rect 4529 51652 4585 51654
rect 4289 50618 4345 50620
rect 4369 50618 4425 50620
rect 4449 50618 4505 50620
rect 4529 50618 4585 50620
rect 4289 50566 4315 50618
rect 4315 50566 4345 50618
rect 4369 50566 4379 50618
rect 4379 50566 4425 50618
rect 4449 50566 4495 50618
rect 4495 50566 4505 50618
rect 4529 50566 4559 50618
rect 4559 50566 4585 50618
rect 4289 50564 4345 50566
rect 4369 50564 4425 50566
rect 4449 50564 4505 50566
rect 4529 50564 4585 50566
rect 4289 49530 4345 49532
rect 4369 49530 4425 49532
rect 4449 49530 4505 49532
rect 4529 49530 4585 49532
rect 4289 49478 4315 49530
rect 4315 49478 4345 49530
rect 4369 49478 4379 49530
rect 4379 49478 4425 49530
rect 4449 49478 4495 49530
rect 4495 49478 4505 49530
rect 4529 49478 4559 49530
rect 4559 49478 4585 49530
rect 4289 49476 4345 49478
rect 4369 49476 4425 49478
rect 4449 49476 4505 49478
rect 4529 49476 4585 49478
rect 4289 48442 4345 48444
rect 4369 48442 4425 48444
rect 4449 48442 4505 48444
rect 4529 48442 4585 48444
rect 4289 48390 4315 48442
rect 4315 48390 4345 48442
rect 4369 48390 4379 48442
rect 4379 48390 4425 48442
rect 4449 48390 4495 48442
rect 4495 48390 4505 48442
rect 4529 48390 4559 48442
rect 4559 48390 4585 48442
rect 4289 48388 4345 48390
rect 4369 48388 4425 48390
rect 4449 48388 4505 48390
rect 4529 48388 4585 48390
rect 4289 47354 4345 47356
rect 4369 47354 4425 47356
rect 4449 47354 4505 47356
rect 4529 47354 4585 47356
rect 4289 47302 4315 47354
rect 4315 47302 4345 47354
rect 4369 47302 4379 47354
rect 4379 47302 4425 47354
rect 4449 47302 4495 47354
rect 4495 47302 4505 47354
rect 4529 47302 4559 47354
rect 4559 47302 4585 47354
rect 4289 47300 4345 47302
rect 4369 47300 4425 47302
rect 4449 47300 4505 47302
rect 4529 47300 4585 47302
rect 4289 46266 4345 46268
rect 4369 46266 4425 46268
rect 4449 46266 4505 46268
rect 4529 46266 4585 46268
rect 4289 46214 4315 46266
rect 4315 46214 4345 46266
rect 4369 46214 4379 46266
rect 4379 46214 4425 46266
rect 4449 46214 4495 46266
rect 4495 46214 4505 46266
rect 4529 46214 4559 46266
rect 4559 46214 4585 46266
rect 4289 46212 4345 46214
rect 4369 46212 4425 46214
rect 4449 46212 4505 46214
rect 4529 46212 4585 46214
rect 4289 45178 4345 45180
rect 4369 45178 4425 45180
rect 4449 45178 4505 45180
rect 4529 45178 4585 45180
rect 4289 45126 4315 45178
rect 4315 45126 4345 45178
rect 4369 45126 4379 45178
rect 4379 45126 4425 45178
rect 4449 45126 4495 45178
rect 4495 45126 4505 45178
rect 4529 45126 4559 45178
rect 4559 45126 4585 45178
rect 4289 45124 4345 45126
rect 4369 45124 4425 45126
rect 4449 45124 4505 45126
rect 4529 45124 4585 45126
rect 4289 44090 4345 44092
rect 4369 44090 4425 44092
rect 4449 44090 4505 44092
rect 4529 44090 4585 44092
rect 4289 44038 4315 44090
rect 4315 44038 4345 44090
rect 4369 44038 4379 44090
rect 4379 44038 4425 44090
rect 4449 44038 4495 44090
rect 4495 44038 4505 44090
rect 4529 44038 4559 44090
rect 4559 44038 4585 44090
rect 4289 44036 4345 44038
rect 4369 44036 4425 44038
rect 4449 44036 4505 44038
rect 4529 44036 4585 44038
rect 4289 43002 4345 43004
rect 4369 43002 4425 43004
rect 4449 43002 4505 43004
rect 4529 43002 4585 43004
rect 4289 42950 4315 43002
rect 4315 42950 4345 43002
rect 4369 42950 4379 43002
rect 4379 42950 4425 43002
rect 4449 42950 4495 43002
rect 4495 42950 4505 43002
rect 4529 42950 4559 43002
rect 4559 42950 4585 43002
rect 4289 42948 4345 42950
rect 4369 42948 4425 42950
rect 4449 42948 4505 42950
rect 4529 42948 4585 42950
rect 4289 41914 4345 41916
rect 4369 41914 4425 41916
rect 4449 41914 4505 41916
rect 4529 41914 4585 41916
rect 4289 41862 4315 41914
rect 4315 41862 4345 41914
rect 4369 41862 4379 41914
rect 4379 41862 4425 41914
rect 4449 41862 4495 41914
rect 4495 41862 4505 41914
rect 4529 41862 4559 41914
rect 4559 41862 4585 41914
rect 4289 41860 4345 41862
rect 4369 41860 4425 41862
rect 4449 41860 4505 41862
rect 4529 41860 4585 41862
rect 4289 40826 4345 40828
rect 4369 40826 4425 40828
rect 4449 40826 4505 40828
rect 4529 40826 4585 40828
rect 4289 40774 4315 40826
rect 4315 40774 4345 40826
rect 4369 40774 4379 40826
rect 4379 40774 4425 40826
rect 4449 40774 4495 40826
rect 4495 40774 4505 40826
rect 4529 40774 4559 40826
rect 4559 40774 4585 40826
rect 4289 40772 4345 40774
rect 4369 40772 4425 40774
rect 4449 40772 4505 40774
rect 4529 40772 4585 40774
rect 4289 39738 4345 39740
rect 4369 39738 4425 39740
rect 4449 39738 4505 39740
rect 4529 39738 4585 39740
rect 4289 39686 4315 39738
rect 4315 39686 4345 39738
rect 4369 39686 4379 39738
rect 4379 39686 4425 39738
rect 4449 39686 4495 39738
rect 4495 39686 4505 39738
rect 4529 39686 4559 39738
rect 4559 39686 4585 39738
rect 4289 39684 4345 39686
rect 4369 39684 4425 39686
rect 4449 39684 4505 39686
rect 4529 39684 4585 39686
rect 4289 38650 4345 38652
rect 4369 38650 4425 38652
rect 4449 38650 4505 38652
rect 4529 38650 4585 38652
rect 4289 38598 4315 38650
rect 4315 38598 4345 38650
rect 4369 38598 4379 38650
rect 4379 38598 4425 38650
rect 4449 38598 4495 38650
rect 4495 38598 4505 38650
rect 4529 38598 4559 38650
rect 4559 38598 4585 38650
rect 4289 38596 4345 38598
rect 4369 38596 4425 38598
rect 4449 38596 4505 38598
rect 4529 38596 4585 38598
rect 4289 37562 4345 37564
rect 4369 37562 4425 37564
rect 4449 37562 4505 37564
rect 4529 37562 4585 37564
rect 4289 37510 4315 37562
rect 4315 37510 4345 37562
rect 4369 37510 4379 37562
rect 4379 37510 4425 37562
rect 4449 37510 4495 37562
rect 4495 37510 4505 37562
rect 4529 37510 4559 37562
rect 4559 37510 4585 37562
rect 4289 37508 4345 37510
rect 4369 37508 4425 37510
rect 4449 37508 4505 37510
rect 4529 37508 4585 37510
rect 4289 36474 4345 36476
rect 4369 36474 4425 36476
rect 4449 36474 4505 36476
rect 4529 36474 4585 36476
rect 4289 36422 4315 36474
rect 4315 36422 4345 36474
rect 4369 36422 4379 36474
rect 4379 36422 4425 36474
rect 4449 36422 4495 36474
rect 4495 36422 4505 36474
rect 4529 36422 4559 36474
rect 4559 36422 4585 36474
rect 4289 36420 4345 36422
rect 4369 36420 4425 36422
rect 4449 36420 4505 36422
rect 4529 36420 4585 36422
rect 4289 35386 4345 35388
rect 4369 35386 4425 35388
rect 4449 35386 4505 35388
rect 4529 35386 4585 35388
rect 4289 35334 4315 35386
rect 4315 35334 4345 35386
rect 4369 35334 4379 35386
rect 4379 35334 4425 35386
rect 4449 35334 4495 35386
rect 4495 35334 4505 35386
rect 4529 35334 4559 35386
rect 4559 35334 4585 35386
rect 4289 35332 4345 35334
rect 4369 35332 4425 35334
rect 4449 35332 4505 35334
rect 4529 35332 4585 35334
rect 4289 34298 4345 34300
rect 4369 34298 4425 34300
rect 4449 34298 4505 34300
rect 4529 34298 4585 34300
rect 4289 34246 4315 34298
rect 4315 34246 4345 34298
rect 4369 34246 4379 34298
rect 4379 34246 4425 34298
rect 4449 34246 4495 34298
rect 4495 34246 4505 34298
rect 4529 34246 4559 34298
rect 4559 34246 4585 34298
rect 4289 34244 4345 34246
rect 4369 34244 4425 34246
rect 4449 34244 4505 34246
rect 4529 34244 4585 34246
rect 4289 33210 4345 33212
rect 4369 33210 4425 33212
rect 4449 33210 4505 33212
rect 4529 33210 4585 33212
rect 4289 33158 4315 33210
rect 4315 33158 4345 33210
rect 4369 33158 4379 33210
rect 4379 33158 4425 33210
rect 4449 33158 4495 33210
rect 4495 33158 4505 33210
rect 4529 33158 4559 33210
rect 4559 33158 4585 33210
rect 4289 33156 4345 33158
rect 4369 33156 4425 33158
rect 4449 33156 4505 33158
rect 4529 33156 4585 33158
rect 4289 32122 4345 32124
rect 4369 32122 4425 32124
rect 4449 32122 4505 32124
rect 4529 32122 4585 32124
rect 4289 32070 4315 32122
rect 4315 32070 4345 32122
rect 4369 32070 4379 32122
rect 4379 32070 4425 32122
rect 4449 32070 4495 32122
rect 4495 32070 4505 32122
rect 4529 32070 4559 32122
rect 4559 32070 4585 32122
rect 4289 32068 4345 32070
rect 4369 32068 4425 32070
rect 4449 32068 4505 32070
rect 4529 32068 4585 32070
rect 4289 31034 4345 31036
rect 4369 31034 4425 31036
rect 4449 31034 4505 31036
rect 4529 31034 4585 31036
rect 4289 30982 4315 31034
rect 4315 30982 4345 31034
rect 4369 30982 4379 31034
rect 4379 30982 4425 31034
rect 4449 30982 4495 31034
rect 4495 30982 4505 31034
rect 4529 30982 4559 31034
rect 4559 30982 4585 31034
rect 4289 30980 4345 30982
rect 4369 30980 4425 30982
rect 4449 30980 4505 30982
rect 4529 30980 4585 30982
rect 4289 29946 4345 29948
rect 4369 29946 4425 29948
rect 4449 29946 4505 29948
rect 4529 29946 4585 29948
rect 4289 29894 4315 29946
rect 4315 29894 4345 29946
rect 4369 29894 4379 29946
rect 4379 29894 4425 29946
rect 4449 29894 4495 29946
rect 4495 29894 4505 29946
rect 4529 29894 4559 29946
rect 4559 29894 4585 29946
rect 4289 29892 4345 29894
rect 4369 29892 4425 29894
rect 4449 29892 4505 29894
rect 4529 29892 4585 29894
rect 4289 28858 4345 28860
rect 4369 28858 4425 28860
rect 4449 28858 4505 28860
rect 4529 28858 4585 28860
rect 4289 28806 4315 28858
rect 4315 28806 4345 28858
rect 4369 28806 4379 28858
rect 4379 28806 4425 28858
rect 4449 28806 4495 28858
rect 4495 28806 4505 28858
rect 4529 28806 4559 28858
rect 4559 28806 4585 28858
rect 4289 28804 4345 28806
rect 4369 28804 4425 28806
rect 4449 28804 4505 28806
rect 4529 28804 4585 28806
rect 4289 27770 4345 27772
rect 4369 27770 4425 27772
rect 4449 27770 4505 27772
rect 4529 27770 4585 27772
rect 4289 27718 4315 27770
rect 4315 27718 4345 27770
rect 4369 27718 4379 27770
rect 4379 27718 4425 27770
rect 4449 27718 4495 27770
rect 4495 27718 4505 27770
rect 4529 27718 4559 27770
rect 4559 27718 4585 27770
rect 4289 27716 4345 27718
rect 4369 27716 4425 27718
rect 4449 27716 4505 27718
rect 4529 27716 4585 27718
rect 4289 26682 4345 26684
rect 4369 26682 4425 26684
rect 4449 26682 4505 26684
rect 4529 26682 4585 26684
rect 4289 26630 4315 26682
rect 4315 26630 4345 26682
rect 4369 26630 4379 26682
rect 4379 26630 4425 26682
rect 4449 26630 4495 26682
rect 4495 26630 4505 26682
rect 4529 26630 4559 26682
rect 4559 26630 4585 26682
rect 4289 26628 4345 26630
rect 4369 26628 4425 26630
rect 4449 26628 4505 26630
rect 4529 26628 4585 26630
rect 4289 25594 4345 25596
rect 4369 25594 4425 25596
rect 4449 25594 4505 25596
rect 4529 25594 4585 25596
rect 4289 25542 4315 25594
rect 4315 25542 4345 25594
rect 4369 25542 4379 25594
rect 4379 25542 4425 25594
rect 4449 25542 4495 25594
rect 4495 25542 4505 25594
rect 4529 25542 4559 25594
rect 4559 25542 4585 25594
rect 4289 25540 4345 25542
rect 4369 25540 4425 25542
rect 4449 25540 4505 25542
rect 4529 25540 4585 25542
rect 4289 24506 4345 24508
rect 4369 24506 4425 24508
rect 4449 24506 4505 24508
rect 4529 24506 4585 24508
rect 4289 24454 4315 24506
rect 4315 24454 4345 24506
rect 4369 24454 4379 24506
rect 4379 24454 4425 24506
rect 4449 24454 4495 24506
rect 4495 24454 4505 24506
rect 4529 24454 4559 24506
rect 4559 24454 4585 24506
rect 4289 24452 4345 24454
rect 4369 24452 4425 24454
rect 4449 24452 4505 24454
rect 4529 24452 4585 24454
rect 3790 24248 3846 24304
rect 4289 23418 4345 23420
rect 4369 23418 4425 23420
rect 4449 23418 4505 23420
rect 4529 23418 4585 23420
rect 4289 23366 4315 23418
rect 4315 23366 4345 23418
rect 4369 23366 4379 23418
rect 4379 23366 4425 23418
rect 4449 23366 4495 23418
rect 4495 23366 4505 23418
rect 4529 23366 4559 23418
rect 4559 23366 4585 23418
rect 4289 23364 4345 23366
rect 4369 23364 4425 23366
rect 4449 23364 4505 23366
rect 4529 23364 4585 23366
rect 4289 22330 4345 22332
rect 4369 22330 4425 22332
rect 4449 22330 4505 22332
rect 4529 22330 4585 22332
rect 4289 22278 4315 22330
rect 4315 22278 4345 22330
rect 4369 22278 4379 22330
rect 4379 22278 4425 22330
rect 4449 22278 4495 22330
rect 4495 22278 4505 22330
rect 4529 22278 4559 22330
rect 4559 22278 4585 22330
rect 4289 22276 4345 22278
rect 4369 22276 4425 22278
rect 4449 22276 4505 22278
rect 4529 22276 4585 22278
rect 4289 21242 4345 21244
rect 4369 21242 4425 21244
rect 4449 21242 4505 21244
rect 4529 21242 4585 21244
rect 4289 21190 4315 21242
rect 4315 21190 4345 21242
rect 4369 21190 4379 21242
rect 4379 21190 4425 21242
rect 4449 21190 4495 21242
rect 4495 21190 4505 21242
rect 4529 21190 4559 21242
rect 4559 21190 4585 21242
rect 4289 21188 4345 21190
rect 4369 21188 4425 21190
rect 4449 21188 4505 21190
rect 4529 21188 4585 21190
rect 4289 20154 4345 20156
rect 4369 20154 4425 20156
rect 4449 20154 4505 20156
rect 4529 20154 4585 20156
rect 4289 20102 4315 20154
rect 4315 20102 4345 20154
rect 4369 20102 4379 20154
rect 4379 20102 4425 20154
rect 4449 20102 4495 20154
rect 4495 20102 4505 20154
rect 4529 20102 4559 20154
rect 4559 20102 4585 20154
rect 4289 20100 4345 20102
rect 4369 20100 4425 20102
rect 4449 20100 4505 20102
rect 4529 20100 4585 20102
rect 4289 19066 4345 19068
rect 4369 19066 4425 19068
rect 4449 19066 4505 19068
rect 4529 19066 4585 19068
rect 4289 19014 4315 19066
rect 4315 19014 4345 19066
rect 4369 19014 4379 19066
rect 4379 19014 4425 19066
rect 4449 19014 4495 19066
rect 4495 19014 4505 19066
rect 4529 19014 4559 19066
rect 4559 19014 4585 19066
rect 4289 19012 4345 19014
rect 4369 19012 4425 19014
rect 4449 19012 4505 19014
rect 4529 19012 4585 19014
rect 4289 17978 4345 17980
rect 4369 17978 4425 17980
rect 4449 17978 4505 17980
rect 4529 17978 4585 17980
rect 4289 17926 4315 17978
rect 4315 17926 4345 17978
rect 4369 17926 4379 17978
rect 4379 17926 4425 17978
rect 4449 17926 4495 17978
rect 4495 17926 4505 17978
rect 4529 17926 4559 17978
rect 4559 17926 4585 17978
rect 4289 17924 4345 17926
rect 4369 17924 4425 17926
rect 4449 17924 4505 17926
rect 4529 17924 4585 17926
rect 5956 330778 6012 330780
rect 6036 330778 6092 330780
rect 6116 330778 6172 330780
rect 6196 330778 6252 330780
rect 5956 330726 5982 330778
rect 5982 330726 6012 330778
rect 6036 330726 6046 330778
rect 6046 330726 6092 330778
rect 6116 330726 6162 330778
rect 6162 330726 6172 330778
rect 6196 330726 6226 330778
rect 6226 330726 6252 330778
rect 5956 330724 6012 330726
rect 6036 330724 6092 330726
rect 6116 330724 6172 330726
rect 6196 330724 6252 330726
rect 5956 329690 6012 329692
rect 6036 329690 6092 329692
rect 6116 329690 6172 329692
rect 6196 329690 6252 329692
rect 5956 329638 5982 329690
rect 5982 329638 6012 329690
rect 6036 329638 6046 329690
rect 6046 329638 6092 329690
rect 6116 329638 6162 329690
rect 6162 329638 6172 329690
rect 6196 329638 6226 329690
rect 6226 329638 6252 329690
rect 5956 329636 6012 329638
rect 6036 329636 6092 329638
rect 6116 329636 6172 329638
rect 6196 329636 6252 329638
rect 5956 328602 6012 328604
rect 6036 328602 6092 328604
rect 6116 328602 6172 328604
rect 6196 328602 6252 328604
rect 5956 328550 5982 328602
rect 5982 328550 6012 328602
rect 6036 328550 6046 328602
rect 6046 328550 6092 328602
rect 6116 328550 6162 328602
rect 6162 328550 6172 328602
rect 6196 328550 6226 328602
rect 6226 328550 6252 328602
rect 5956 328548 6012 328550
rect 6036 328548 6092 328550
rect 6116 328548 6172 328550
rect 6196 328548 6252 328550
rect 5956 327514 6012 327516
rect 6036 327514 6092 327516
rect 6116 327514 6172 327516
rect 6196 327514 6252 327516
rect 5956 327462 5982 327514
rect 5982 327462 6012 327514
rect 6036 327462 6046 327514
rect 6046 327462 6092 327514
rect 6116 327462 6162 327514
rect 6162 327462 6172 327514
rect 6196 327462 6226 327514
rect 6226 327462 6252 327514
rect 5956 327460 6012 327462
rect 6036 327460 6092 327462
rect 6116 327460 6172 327462
rect 6196 327460 6252 327462
rect 5956 326426 6012 326428
rect 6036 326426 6092 326428
rect 6116 326426 6172 326428
rect 6196 326426 6252 326428
rect 5956 326374 5982 326426
rect 5982 326374 6012 326426
rect 6036 326374 6046 326426
rect 6046 326374 6092 326426
rect 6116 326374 6162 326426
rect 6162 326374 6172 326426
rect 6196 326374 6226 326426
rect 6226 326374 6252 326426
rect 5956 326372 6012 326374
rect 6036 326372 6092 326374
rect 6116 326372 6172 326374
rect 6196 326372 6252 326374
rect 5956 325338 6012 325340
rect 6036 325338 6092 325340
rect 6116 325338 6172 325340
rect 6196 325338 6252 325340
rect 5956 325286 5982 325338
rect 5982 325286 6012 325338
rect 6036 325286 6046 325338
rect 6046 325286 6092 325338
rect 6116 325286 6162 325338
rect 6162 325286 6172 325338
rect 6196 325286 6226 325338
rect 6226 325286 6252 325338
rect 5956 325284 6012 325286
rect 6036 325284 6092 325286
rect 6116 325284 6172 325286
rect 6196 325284 6252 325286
rect 5956 324250 6012 324252
rect 6036 324250 6092 324252
rect 6116 324250 6172 324252
rect 6196 324250 6252 324252
rect 5956 324198 5982 324250
rect 5982 324198 6012 324250
rect 6036 324198 6046 324250
rect 6046 324198 6092 324250
rect 6116 324198 6162 324250
rect 6162 324198 6172 324250
rect 6196 324198 6226 324250
rect 6226 324198 6252 324250
rect 5956 324196 6012 324198
rect 6036 324196 6092 324198
rect 6116 324196 6172 324198
rect 6196 324196 6252 324198
rect 5956 323162 6012 323164
rect 6036 323162 6092 323164
rect 6116 323162 6172 323164
rect 6196 323162 6252 323164
rect 5956 323110 5982 323162
rect 5982 323110 6012 323162
rect 6036 323110 6046 323162
rect 6046 323110 6092 323162
rect 6116 323110 6162 323162
rect 6162 323110 6172 323162
rect 6196 323110 6226 323162
rect 6226 323110 6252 323162
rect 5956 323108 6012 323110
rect 6036 323108 6092 323110
rect 6116 323108 6172 323110
rect 6196 323108 6252 323110
rect 5956 322074 6012 322076
rect 6036 322074 6092 322076
rect 6116 322074 6172 322076
rect 6196 322074 6252 322076
rect 5956 322022 5982 322074
rect 5982 322022 6012 322074
rect 6036 322022 6046 322074
rect 6046 322022 6092 322074
rect 6116 322022 6162 322074
rect 6162 322022 6172 322074
rect 6196 322022 6226 322074
rect 6226 322022 6252 322074
rect 5956 322020 6012 322022
rect 6036 322020 6092 322022
rect 6116 322020 6172 322022
rect 6196 322020 6252 322022
rect 5956 320986 6012 320988
rect 6036 320986 6092 320988
rect 6116 320986 6172 320988
rect 6196 320986 6252 320988
rect 5956 320934 5982 320986
rect 5982 320934 6012 320986
rect 6036 320934 6046 320986
rect 6046 320934 6092 320986
rect 6116 320934 6162 320986
rect 6162 320934 6172 320986
rect 6196 320934 6226 320986
rect 6226 320934 6252 320986
rect 5956 320932 6012 320934
rect 6036 320932 6092 320934
rect 6116 320932 6172 320934
rect 6196 320932 6252 320934
rect 5956 319898 6012 319900
rect 6036 319898 6092 319900
rect 6116 319898 6172 319900
rect 6196 319898 6252 319900
rect 5956 319846 5982 319898
rect 5982 319846 6012 319898
rect 6036 319846 6046 319898
rect 6046 319846 6092 319898
rect 6116 319846 6162 319898
rect 6162 319846 6172 319898
rect 6196 319846 6226 319898
rect 6226 319846 6252 319898
rect 5956 319844 6012 319846
rect 6036 319844 6092 319846
rect 6116 319844 6172 319846
rect 6196 319844 6252 319846
rect 5956 318810 6012 318812
rect 6036 318810 6092 318812
rect 6116 318810 6172 318812
rect 6196 318810 6252 318812
rect 5956 318758 5982 318810
rect 5982 318758 6012 318810
rect 6036 318758 6046 318810
rect 6046 318758 6092 318810
rect 6116 318758 6162 318810
rect 6162 318758 6172 318810
rect 6196 318758 6226 318810
rect 6226 318758 6252 318810
rect 5956 318756 6012 318758
rect 6036 318756 6092 318758
rect 6116 318756 6172 318758
rect 6196 318756 6252 318758
rect 5956 317722 6012 317724
rect 6036 317722 6092 317724
rect 6116 317722 6172 317724
rect 6196 317722 6252 317724
rect 5956 317670 5982 317722
rect 5982 317670 6012 317722
rect 6036 317670 6046 317722
rect 6046 317670 6092 317722
rect 6116 317670 6162 317722
rect 6162 317670 6172 317722
rect 6196 317670 6226 317722
rect 6226 317670 6252 317722
rect 5956 317668 6012 317670
rect 6036 317668 6092 317670
rect 6116 317668 6172 317670
rect 6196 317668 6252 317670
rect 5956 316634 6012 316636
rect 6036 316634 6092 316636
rect 6116 316634 6172 316636
rect 6196 316634 6252 316636
rect 5956 316582 5982 316634
rect 5982 316582 6012 316634
rect 6036 316582 6046 316634
rect 6046 316582 6092 316634
rect 6116 316582 6162 316634
rect 6162 316582 6172 316634
rect 6196 316582 6226 316634
rect 6226 316582 6252 316634
rect 5956 316580 6012 316582
rect 6036 316580 6092 316582
rect 6116 316580 6172 316582
rect 6196 316580 6252 316582
rect 5956 315546 6012 315548
rect 6036 315546 6092 315548
rect 6116 315546 6172 315548
rect 6196 315546 6252 315548
rect 5956 315494 5982 315546
rect 5982 315494 6012 315546
rect 6036 315494 6046 315546
rect 6046 315494 6092 315546
rect 6116 315494 6162 315546
rect 6162 315494 6172 315546
rect 6196 315494 6226 315546
rect 6226 315494 6252 315546
rect 5956 315492 6012 315494
rect 6036 315492 6092 315494
rect 6116 315492 6172 315494
rect 6196 315492 6252 315494
rect 5956 314458 6012 314460
rect 6036 314458 6092 314460
rect 6116 314458 6172 314460
rect 6196 314458 6252 314460
rect 5956 314406 5982 314458
rect 5982 314406 6012 314458
rect 6036 314406 6046 314458
rect 6046 314406 6092 314458
rect 6116 314406 6162 314458
rect 6162 314406 6172 314458
rect 6196 314406 6226 314458
rect 6226 314406 6252 314458
rect 5956 314404 6012 314406
rect 6036 314404 6092 314406
rect 6116 314404 6172 314406
rect 6196 314404 6252 314406
rect 5956 313370 6012 313372
rect 6036 313370 6092 313372
rect 6116 313370 6172 313372
rect 6196 313370 6252 313372
rect 5956 313318 5982 313370
rect 5982 313318 6012 313370
rect 6036 313318 6046 313370
rect 6046 313318 6092 313370
rect 6116 313318 6162 313370
rect 6162 313318 6172 313370
rect 6196 313318 6226 313370
rect 6226 313318 6252 313370
rect 5956 313316 6012 313318
rect 6036 313316 6092 313318
rect 6116 313316 6172 313318
rect 6196 313316 6252 313318
rect 5956 312282 6012 312284
rect 6036 312282 6092 312284
rect 6116 312282 6172 312284
rect 6196 312282 6252 312284
rect 5956 312230 5982 312282
rect 5982 312230 6012 312282
rect 6036 312230 6046 312282
rect 6046 312230 6092 312282
rect 6116 312230 6162 312282
rect 6162 312230 6172 312282
rect 6196 312230 6226 312282
rect 6226 312230 6252 312282
rect 5956 312228 6012 312230
rect 6036 312228 6092 312230
rect 6116 312228 6172 312230
rect 6196 312228 6252 312230
rect 5956 311194 6012 311196
rect 6036 311194 6092 311196
rect 6116 311194 6172 311196
rect 6196 311194 6252 311196
rect 5956 311142 5982 311194
rect 5982 311142 6012 311194
rect 6036 311142 6046 311194
rect 6046 311142 6092 311194
rect 6116 311142 6162 311194
rect 6162 311142 6172 311194
rect 6196 311142 6226 311194
rect 6226 311142 6252 311194
rect 5956 311140 6012 311142
rect 6036 311140 6092 311142
rect 6116 311140 6172 311142
rect 6196 311140 6252 311142
rect 5956 310106 6012 310108
rect 6036 310106 6092 310108
rect 6116 310106 6172 310108
rect 6196 310106 6252 310108
rect 5956 310054 5982 310106
rect 5982 310054 6012 310106
rect 6036 310054 6046 310106
rect 6046 310054 6092 310106
rect 6116 310054 6162 310106
rect 6162 310054 6172 310106
rect 6196 310054 6226 310106
rect 6226 310054 6252 310106
rect 5956 310052 6012 310054
rect 6036 310052 6092 310054
rect 6116 310052 6172 310054
rect 6196 310052 6252 310054
rect 5956 309018 6012 309020
rect 6036 309018 6092 309020
rect 6116 309018 6172 309020
rect 6196 309018 6252 309020
rect 5956 308966 5982 309018
rect 5982 308966 6012 309018
rect 6036 308966 6046 309018
rect 6046 308966 6092 309018
rect 6116 308966 6162 309018
rect 6162 308966 6172 309018
rect 6196 308966 6226 309018
rect 6226 308966 6252 309018
rect 5956 308964 6012 308966
rect 6036 308964 6092 308966
rect 6116 308964 6172 308966
rect 6196 308964 6252 308966
rect 5956 307930 6012 307932
rect 6036 307930 6092 307932
rect 6116 307930 6172 307932
rect 6196 307930 6252 307932
rect 5956 307878 5982 307930
rect 5982 307878 6012 307930
rect 6036 307878 6046 307930
rect 6046 307878 6092 307930
rect 6116 307878 6162 307930
rect 6162 307878 6172 307930
rect 6196 307878 6226 307930
rect 6226 307878 6252 307930
rect 5956 307876 6012 307878
rect 6036 307876 6092 307878
rect 6116 307876 6172 307878
rect 6196 307876 6252 307878
rect 5956 306842 6012 306844
rect 6036 306842 6092 306844
rect 6116 306842 6172 306844
rect 6196 306842 6252 306844
rect 5956 306790 5982 306842
rect 5982 306790 6012 306842
rect 6036 306790 6046 306842
rect 6046 306790 6092 306842
rect 6116 306790 6162 306842
rect 6162 306790 6172 306842
rect 6196 306790 6226 306842
rect 6226 306790 6252 306842
rect 5956 306788 6012 306790
rect 6036 306788 6092 306790
rect 6116 306788 6172 306790
rect 6196 306788 6252 306790
rect 5956 305754 6012 305756
rect 6036 305754 6092 305756
rect 6116 305754 6172 305756
rect 6196 305754 6252 305756
rect 5956 305702 5982 305754
rect 5982 305702 6012 305754
rect 6036 305702 6046 305754
rect 6046 305702 6092 305754
rect 6116 305702 6162 305754
rect 6162 305702 6172 305754
rect 6196 305702 6226 305754
rect 6226 305702 6252 305754
rect 5956 305700 6012 305702
rect 6036 305700 6092 305702
rect 6116 305700 6172 305702
rect 6196 305700 6252 305702
rect 5956 304666 6012 304668
rect 6036 304666 6092 304668
rect 6116 304666 6172 304668
rect 6196 304666 6252 304668
rect 5956 304614 5982 304666
rect 5982 304614 6012 304666
rect 6036 304614 6046 304666
rect 6046 304614 6092 304666
rect 6116 304614 6162 304666
rect 6162 304614 6172 304666
rect 6196 304614 6226 304666
rect 6226 304614 6252 304666
rect 5956 304612 6012 304614
rect 6036 304612 6092 304614
rect 6116 304612 6172 304614
rect 6196 304612 6252 304614
rect 5956 303578 6012 303580
rect 6036 303578 6092 303580
rect 6116 303578 6172 303580
rect 6196 303578 6252 303580
rect 5956 303526 5982 303578
rect 5982 303526 6012 303578
rect 6036 303526 6046 303578
rect 6046 303526 6092 303578
rect 6116 303526 6162 303578
rect 6162 303526 6172 303578
rect 6196 303526 6226 303578
rect 6226 303526 6252 303578
rect 5956 303524 6012 303526
rect 6036 303524 6092 303526
rect 6116 303524 6172 303526
rect 6196 303524 6252 303526
rect 5956 302490 6012 302492
rect 6036 302490 6092 302492
rect 6116 302490 6172 302492
rect 6196 302490 6252 302492
rect 5956 302438 5982 302490
rect 5982 302438 6012 302490
rect 6036 302438 6046 302490
rect 6046 302438 6092 302490
rect 6116 302438 6162 302490
rect 6162 302438 6172 302490
rect 6196 302438 6226 302490
rect 6226 302438 6252 302490
rect 5956 302436 6012 302438
rect 6036 302436 6092 302438
rect 6116 302436 6172 302438
rect 6196 302436 6252 302438
rect 5956 301402 6012 301404
rect 6036 301402 6092 301404
rect 6116 301402 6172 301404
rect 6196 301402 6252 301404
rect 5956 301350 5982 301402
rect 5982 301350 6012 301402
rect 6036 301350 6046 301402
rect 6046 301350 6092 301402
rect 6116 301350 6162 301402
rect 6162 301350 6172 301402
rect 6196 301350 6226 301402
rect 6226 301350 6252 301402
rect 5956 301348 6012 301350
rect 6036 301348 6092 301350
rect 6116 301348 6172 301350
rect 6196 301348 6252 301350
rect 5956 300314 6012 300316
rect 6036 300314 6092 300316
rect 6116 300314 6172 300316
rect 6196 300314 6252 300316
rect 5956 300262 5982 300314
rect 5982 300262 6012 300314
rect 6036 300262 6046 300314
rect 6046 300262 6092 300314
rect 6116 300262 6162 300314
rect 6162 300262 6172 300314
rect 6196 300262 6226 300314
rect 6226 300262 6252 300314
rect 5956 300260 6012 300262
rect 6036 300260 6092 300262
rect 6116 300260 6172 300262
rect 6196 300260 6252 300262
rect 5956 299226 6012 299228
rect 6036 299226 6092 299228
rect 6116 299226 6172 299228
rect 6196 299226 6252 299228
rect 5956 299174 5982 299226
rect 5982 299174 6012 299226
rect 6036 299174 6046 299226
rect 6046 299174 6092 299226
rect 6116 299174 6162 299226
rect 6162 299174 6172 299226
rect 6196 299174 6226 299226
rect 6226 299174 6252 299226
rect 5956 299172 6012 299174
rect 6036 299172 6092 299174
rect 6116 299172 6172 299174
rect 6196 299172 6252 299174
rect 5956 298138 6012 298140
rect 6036 298138 6092 298140
rect 6116 298138 6172 298140
rect 6196 298138 6252 298140
rect 5956 298086 5982 298138
rect 5982 298086 6012 298138
rect 6036 298086 6046 298138
rect 6046 298086 6092 298138
rect 6116 298086 6162 298138
rect 6162 298086 6172 298138
rect 6196 298086 6226 298138
rect 6226 298086 6252 298138
rect 5956 298084 6012 298086
rect 6036 298084 6092 298086
rect 6116 298084 6172 298086
rect 6196 298084 6252 298086
rect 5956 297050 6012 297052
rect 6036 297050 6092 297052
rect 6116 297050 6172 297052
rect 6196 297050 6252 297052
rect 5956 296998 5982 297050
rect 5982 296998 6012 297050
rect 6036 296998 6046 297050
rect 6046 296998 6092 297050
rect 6116 296998 6162 297050
rect 6162 296998 6172 297050
rect 6196 296998 6226 297050
rect 6226 296998 6252 297050
rect 5956 296996 6012 296998
rect 6036 296996 6092 296998
rect 6116 296996 6172 296998
rect 6196 296996 6252 296998
rect 5956 295962 6012 295964
rect 6036 295962 6092 295964
rect 6116 295962 6172 295964
rect 6196 295962 6252 295964
rect 5956 295910 5982 295962
rect 5982 295910 6012 295962
rect 6036 295910 6046 295962
rect 6046 295910 6092 295962
rect 6116 295910 6162 295962
rect 6162 295910 6172 295962
rect 6196 295910 6226 295962
rect 6226 295910 6252 295962
rect 5956 295908 6012 295910
rect 6036 295908 6092 295910
rect 6116 295908 6172 295910
rect 6196 295908 6252 295910
rect 5956 294874 6012 294876
rect 6036 294874 6092 294876
rect 6116 294874 6172 294876
rect 6196 294874 6252 294876
rect 5956 294822 5982 294874
rect 5982 294822 6012 294874
rect 6036 294822 6046 294874
rect 6046 294822 6092 294874
rect 6116 294822 6162 294874
rect 6162 294822 6172 294874
rect 6196 294822 6226 294874
rect 6226 294822 6252 294874
rect 5956 294820 6012 294822
rect 6036 294820 6092 294822
rect 6116 294820 6172 294822
rect 6196 294820 6252 294822
rect 5956 293786 6012 293788
rect 6036 293786 6092 293788
rect 6116 293786 6172 293788
rect 6196 293786 6252 293788
rect 5956 293734 5982 293786
rect 5982 293734 6012 293786
rect 6036 293734 6046 293786
rect 6046 293734 6092 293786
rect 6116 293734 6162 293786
rect 6162 293734 6172 293786
rect 6196 293734 6226 293786
rect 6226 293734 6252 293786
rect 5956 293732 6012 293734
rect 6036 293732 6092 293734
rect 6116 293732 6172 293734
rect 6196 293732 6252 293734
rect 5956 292698 6012 292700
rect 6036 292698 6092 292700
rect 6116 292698 6172 292700
rect 6196 292698 6252 292700
rect 5956 292646 5982 292698
rect 5982 292646 6012 292698
rect 6036 292646 6046 292698
rect 6046 292646 6092 292698
rect 6116 292646 6162 292698
rect 6162 292646 6172 292698
rect 6196 292646 6226 292698
rect 6226 292646 6252 292698
rect 5956 292644 6012 292646
rect 6036 292644 6092 292646
rect 6116 292644 6172 292646
rect 6196 292644 6252 292646
rect 5956 291610 6012 291612
rect 6036 291610 6092 291612
rect 6116 291610 6172 291612
rect 6196 291610 6252 291612
rect 5956 291558 5982 291610
rect 5982 291558 6012 291610
rect 6036 291558 6046 291610
rect 6046 291558 6092 291610
rect 6116 291558 6162 291610
rect 6162 291558 6172 291610
rect 6196 291558 6226 291610
rect 6226 291558 6252 291610
rect 5956 291556 6012 291558
rect 6036 291556 6092 291558
rect 6116 291556 6172 291558
rect 6196 291556 6252 291558
rect 5956 290522 6012 290524
rect 6036 290522 6092 290524
rect 6116 290522 6172 290524
rect 6196 290522 6252 290524
rect 5956 290470 5982 290522
rect 5982 290470 6012 290522
rect 6036 290470 6046 290522
rect 6046 290470 6092 290522
rect 6116 290470 6162 290522
rect 6162 290470 6172 290522
rect 6196 290470 6226 290522
rect 6226 290470 6252 290522
rect 5956 290468 6012 290470
rect 6036 290468 6092 290470
rect 6116 290468 6172 290470
rect 6196 290468 6252 290470
rect 5956 289434 6012 289436
rect 6036 289434 6092 289436
rect 6116 289434 6172 289436
rect 6196 289434 6252 289436
rect 5956 289382 5982 289434
rect 5982 289382 6012 289434
rect 6036 289382 6046 289434
rect 6046 289382 6092 289434
rect 6116 289382 6162 289434
rect 6162 289382 6172 289434
rect 6196 289382 6226 289434
rect 6226 289382 6252 289434
rect 5956 289380 6012 289382
rect 6036 289380 6092 289382
rect 6116 289380 6172 289382
rect 6196 289380 6252 289382
rect 5956 288346 6012 288348
rect 6036 288346 6092 288348
rect 6116 288346 6172 288348
rect 6196 288346 6252 288348
rect 5956 288294 5982 288346
rect 5982 288294 6012 288346
rect 6036 288294 6046 288346
rect 6046 288294 6092 288346
rect 6116 288294 6162 288346
rect 6162 288294 6172 288346
rect 6196 288294 6226 288346
rect 6226 288294 6252 288346
rect 5956 288292 6012 288294
rect 6036 288292 6092 288294
rect 6116 288292 6172 288294
rect 6196 288292 6252 288294
rect 5956 287258 6012 287260
rect 6036 287258 6092 287260
rect 6116 287258 6172 287260
rect 6196 287258 6252 287260
rect 5956 287206 5982 287258
rect 5982 287206 6012 287258
rect 6036 287206 6046 287258
rect 6046 287206 6092 287258
rect 6116 287206 6162 287258
rect 6162 287206 6172 287258
rect 6196 287206 6226 287258
rect 6226 287206 6252 287258
rect 5956 287204 6012 287206
rect 6036 287204 6092 287206
rect 6116 287204 6172 287206
rect 6196 287204 6252 287206
rect 5956 286170 6012 286172
rect 6036 286170 6092 286172
rect 6116 286170 6172 286172
rect 6196 286170 6252 286172
rect 5956 286118 5982 286170
rect 5982 286118 6012 286170
rect 6036 286118 6046 286170
rect 6046 286118 6092 286170
rect 6116 286118 6162 286170
rect 6162 286118 6172 286170
rect 6196 286118 6226 286170
rect 6226 286118 6252 286170
rect 5956 286116 6012 286118
rect 6036 286116 6092 286118
rect 6116 286116 6172 286118
rect 6196 286116 6252 286118
rect 5956 285082 6012 285084
rect 6036 285082 6092 285084
rect 6116 285082 6172 285084
rect 6196 285082 6252 285084
rect 5956 285030 5982 285082
rect 5982 285030 6012 285082
rect 6036 285030 6046 285082
rect 6046 285030 6092 285082
rect 6116 285030 6162 285082
rect 6162 285030 6172 285082
rect 6196 285030 6226 285082
rect 6226 285030 6252 285082
rect 5956 285028 6012 285030
rect 6036 285028 6092 285030
rect 6116 285028 6172 285030
rect 6196 285028 6252 285030
rect 5956 283994 6012 283996
rect 6036 283994 6092 283996
rect 6116 283994 6172 283996
rect 6196 283994 6252 283996
rect 5956 283942 5982 283994
rect 5982 283942 6012 283994
rect 6036 283942 6046 283994
rect 6046 283942 6092 283994
rect 6116 283942 6162 283994
rect 6162 283942 6172 283994
rect 6196 283942 6226 283994
rect 6226 283942 6252 283994
rect 5956 283940 6012 283942
rect 6036 283940 6092 283942
rect 6116 283940 6172 283942
rect 6196 283940 6252 283942
rect 5956 282906 6012 282908
rect 6036 282906 6092 282908
rect 6116 282906 6172 282908
rect 6196 282906 6252 282908
rect 5956 282854 5982 282906
rect 5982 282854 6012 282906
rect 6036 282854 6046 282906
rect 6046 282854 6092 282906
rect 6116 282854 6162 282906
rect 6162 282854 6172 282906
rect 6196 282854 6226 282906
rect 6226 282854 6252 282906
rect 5956 282852 6012 282854
rect 6036 282852 6092 282854
rect 6116 282852 6172 282854
rect 6196 282852 6252 282854
rect 6274 282512 6330 282568
rect 5956 281818 6012 281820
rect 6036 281818 6092 281820
rect 6116 281818 6172 281820
rect 6196 281818 6252 281820
rect 5956 281766 5982 281818
rect 5982 281766 6012 281818
rect 6036 281766 6046 281818
rect 6046 281766 6092 281818
rect 6116 281766 6162 281818
rect 6162 281766 6172 281818
rect 6196 281766 6226 281818
rect 6226 281766 6252 281818
rect 5956 281764 6012 281766
rect 6036 281764 6092 281766
rect 6116 281764 6172 281766
rect 6196 281764 6252 281766
rect 5956 280730 6012 280732
rect 6036 280730 6092 280732
rect 6116 280730 6172 280732
rect 6196 280730 6252 280732
rect 5956 280678 5982 280730
rect 5982 280678 6012 280730
rect 6036 280678 6046 280730
rect 6046 280678 6092 280730
rect 6116 280678 6162 280730
rect 6162 280678 6172 280730
rect 6196 280678 6226 280730
rect 6226 280678 6252 280730
rect 5956 280676 6012 280678
rect 6036 280676 6092 280678
rect 6116 280676 6172 280678
rect 6196 280676 6252 280678
rect 5956 279642 6012 279644
rect 6036 279642 6092 279644
rect 6116 279642 6172 279644
rect 6196 279642 6252 279644
rect 5956 279590 5982 279642
rect 5982 279590 6012 279642
rect 6036 279590 6046 279642
rect 6046 279590 6092 279642
rect 6116 279590 6162 279642
rect 6162 279590 6172 279642
rect 6196 279590 6226 279642
rect 6226 279590 6252 279642
rect 5956 279588 6012 279590
rect 6036 279588 6092 279590
rect 6116 279588 6172 279590
rect 6196 279588 6252 279590
rect 5956 278554 6012 278556
rect 6036 278554 6092 278556
rect 6116 278554 6172 278556
rect 6196 278554 6252 278556
rect 5956 278502 5982 278554
rect 5982 278502 6012 278554
rect 6036 278502 6046 278554
rect 6046 278502 6092 278554
rect 6116 278502 6162 278554
rect 6162 278502 6172 278554
rect 6196 278502 6226 278554
rect 6226 278502 6252 278554
rect 5956 278500 6012 278502
rect 6036 278500 6092 278502
rect 6116 278500 6172 278502
rect 6196 278500 6252 278502
rect 5956 277466 6012 277468
rect 6036 277466 6092 277468
rect 6116 277466 6172 277468
rect 6196 277466 6252 277468
rect 5956 277414 5982 277466
rect 5982 277414 6012 277466
rect 6036 277414 6046 277466
rect 6046 277414 6092 277466
rect 6116 277414 6162 277466
rect 6162 277414 6172 277466
rect 6196 277414 6226 277466
rect 6226 277414 6252 277466
rect 5956 277412 6012 277414
rect 6036 277412 6092 277414
rect 6116 277412 6172 277414
rect 6196 277412 6252 277414
rect 5956 276378 6012 276380
rect 6036 276378 6092 276380
rect 6116 276378 6172 276380
rect 6196 276378 6252 276380
rect 5956 276326 5982 276378
rect 5982 276326 6012 276378
rect 6036 276326 6046 276378
rect 6046 276326 6092 276378
rect 6116 276326 6162 276378
rect 6162 276326 6172 276378
rect 6196 276326 6226 276378
rect 6226 276326 6252 276378
rect 5956 276324 6012 276326
rect 6036 276324 6092 276326
rect 6116 276324 6172 276326
rect 6196 276324 6252 276326
rect 5956 275290 6012 275292
rect 6036 275290 6092 275292
rect 6116 275290 6172 275292
rect 6196 275290 6252 275292
rect 5956 275238 5982 275290
rect 5982 275238 6012 275290
rect 6036 275238 6046 275290
rect 6046 275238 6092 275290
rect 6116 275238 6162 275290
rect 6162 275238 6172 275290
rect 6196 275238 6226 275290
rect 6226 275238 6252 275290
rect 5956 275236 6012 275238
rect 6036 275236 6092 275238
rect 6116 275236 6172 275238
rect 6196 275236 6252 275238
rect 5956 274202 6012 274204
rect 6036 274202 6092 274204
rect 6116 274202 6172 274204
rect 6196 274202 6252 274204
rect 5956 274150 5982 274202
rect 5982 274150 6012 274202
rect 6036 274150 6046 274202
rect 6046 274150 6092 274202
rect 6116 274150 6162 274202
rect 6162 274150 6172 274202
rect 6196 274150 6226 274202
rect 6226 274150 6252 274202
rect 5956 274148 6012 274150
rect 6036 274148 6092 274150
rect 6116 274148 6172 274150
rect 6196 274148 6252 274150
rect 5956 273114 6012 273116
rect 6036 273114 6092 273116
rect 6116 273114 6172 273116
rect 6196 273114 6252 273116
rect 5956 273062 5982 273114
rect 5982 273062 6012 273114
rect 6036 273062 6046 273114
rect 6046 273062 6092 273114
rect 6116 273062 6162 273114
rect 6162 273062 6172 273114
rect 6196 273062 6226 273114
rect 6226 273062 6252 273114
rect 5956 273060 6012 273062
rect 6036 273060 6092 273062
rect 6116 273060 6172 273062
rect 6196 273060 6252 273062
rect 5956 272026 6012 272028
rect 6036 272026 6092 272028
rect 6116 272026 6172 272028
rect 6196 272026 6252 272028
rect 5956 271974 5982 272026
rect 5982 271974 6012 272026
rect 6036 271974 6046 272026
rect 6046 271974 6092 272026
rect 6116 271974 6162 272026
rect 6162 271974 6172 272026
rect 6196 271974 6226 272026
rect 6226 271974 6252 272026
rect 5956 271972 6012 271974
rect 6036 271972 6092 271974
rect 6116 271972 6172 271974
rect 6196 271972 6252 271974
rect 5956 270938 6012 270940
rect 6036 270938 6092 270940
rect 6116 270938 6172 270940
rect 6196 270938 6252 270940
rect 5956 270886 5982 270938
rect 5982 270886 6012 270938
rect 6036 270886 6046 270938
rect 6046 270886 6092 270938
rect 6116 270886 6162 270938
rect 6162 270886 6172 270938
rect 6196 270886 6226 270938
rect 6226 270886 6252 270938
rect 5956 270884 6012 270886
rect 6036 270884 6092 270886
rect 6116 270884 6172 270886
rect 6196 270884 6252 270886
rect 5956 269850 6012 269852
rect 6036 269850 6092 269852
rect 6116 269850 6172 269852
rect 6196 269850 6252 269852
rect 5956 269798 5982 269850
rect 5982 269798 6012 269850
rect 6036 269798 6046 269850
rect 6046 269798 6092 269850
rect 6116 269798 6162 269850
rect 6162 269798 6172 269850
rect 6196 269798 6226 269850
rect 6226 269798 6252 269850
rect 5956 269796 6012 269798
rect 6036 269796 6092 269798
rect 6116 269796 6172 269798
rect 6196 269796 6252 269798
rect 5956 268762 6012 268764
rect 6036 268762 6092 268764
rect 6116 268762 6172 268764
rect 6196 268762 6252 268764
rect 5956 268710 5982 268762
rect 5982 268710 6012 268762
rect 6036 268710 6046 268762
rect 6046 268710 6092 268762
rect 6116 268710 6162 268762
rect 6162 268710 6172 268762
rect 6196 268710 6226 268762
rect 6226 268710 6252 268762
rect 5956 268708 6012 268710
rect 6036 268708 6092 268710
rect 6116 268708 6172 268710
rect 6196 268708 6252 268710
rect 5956 267674 6012 267676
rect 6036 267674 6092 267676
rect 6116 267674 6172 267676
rect 6196 267674 6252 267676
rect 5956 267622 5982 267674
rect 5982 267622 6012 267674
rect 6036 267622 6046 267674
rect 6046 267622 6092 267674
rect 6116 267622 6162 267674
rect 6162 267622 6172 267674
rect 6196 267622 6226 267674
rect 6226 267622 6252 267674
rect 5956 267620 6012 267622
rect 6036 267620 6092 267622
rect 6116 267620 6172 267622
rect 6196 267620 6252 267622
rect 5956 266586 6012 266588
rect 6036 266586 6092 266588
rect 6116 266586 6172 266588
rect 6196 266586 6252 266588
rect 5956 266534 5982 266586
rect 5982 266534 6012 266586
rect 6036 266534 6046 266586
rect 6046 266534 6092 266586
rect 6116 266534 6162 266586
rect 6162 266534 6172 266586
rect 6196 266534 6226 266586
rect 6226 266534 6252 266586
rect 5956 266532 6012 266534
rect 6036 266532 6092 266534
rect 6116 266532 6172 266534
rect 6196 266532 6252 266534
rect 5956 265498 6012 265500
rect 6036 265498 6092 265500
rect 6116 265498 6172 265500
rect 6196 265498 6252 265500
rect 5956 265446 5982 265498
rect 5982 265446 6012 265498
rect 6036 265446 6046 265498
rect 6046 265446 6092 265498
rect 6116 265446 6162 265498
rect 6162 265446 6172 265498
rect 6196 265446 6226 265498
rect 6226 265446 6252 265498
rect 5956 265444 6012 265446
rect 6036 265444 6092 265446
rect 6116 265444 6172 265446
rect 6196 265444 6252 265446
rect 5956 264410 6012 264412
rect 6036 264410 6092 264412
rect 6116 264410 6172 264412
rect 6196 264410 6252 264412
rect 5956 264358 5982 264410
rect 5982 264358 6012 264410
rect 6036 264358 6046 264410
rect 6046 264358 6092 264410
rect 6116 264358 6162 264410
rect 6162 264358 6172 264410
rect 6196 264358 6226 264410
rect 6226 264358 6252 264410
rect 5956 264356 6012 264358
rect 6036 264356 6092 264358
rect 6116 264356 6172 264358
rect 6196 264356 6252 264358
rect 5956 263322 6012 263324
rect 6036 263322 6092 263324
rect 6116 263322 6172 263324
rect 6196 263322 6252 263324
rect 5956 263270 5982 263322
rect 5982 263270 6012 263322
rect 6036 263270 6046 263322
rect 6046 263270 6092 263322
rect 6116 263270 6162 263322
rect 6162 263270 6172 263322
rect 6196 263270 6226 263322
rect 6226 263270 6252 263322
rect 5956 263268 6012 263270
rect 6036 263268 6092 263270
rect 6116 263268 6172 263270
rect 6196 263268 6252 263270
rect 5956 262234 6012 262236
rect 6036 262234 6092 262236
rect 6116 262234 6172 262236
rect 6196 262234 6252 262236
rect 5956 262182 5982 262234
rect 5982 262182 6012 262234
rect 6036 262182 6046 262234
rect 6046 262182 6092 262234
rect 6116 262182 6162 262234
rect 6162 262182 6172 262234
rect 6196 262182 6226 262234
rect 6226 262182 6252 262234
rect 5956 262180 6012 262182
rect 6036 262180 6092 262182
rect 6116 262180 6172 262182
rect 6196 262180 6252 262182
rect 5956 261146 6012 261148
rect 6036 261146 6092 261148
rect 6116 261146 6172 261148
rect 6196 261146 6252 261148
rect 5956 261094 5982 261146
rect 5982 261094 6012 261146
rect 6036 261094 6046 261146
rect 6046 261094 6092 261146
rect 6116 261094 6162 261146
rect 6162 261094 6172 261146
rect 6196 261094 6226 261146
rect 6226 261094 6252 261146
rect 5956 261092 6012 261094
rect 6036 261092 6092 261094
rect 6116 261092 6172 261094
rect 6196 261092 6252 261094
rect 5956 260058 6012 260060
rect 6036 260058 6092 260060
rect 6116 260058 6172 260060
rect 6196 260058 6252 260060
rect 5956 260006 5982 260058
rect 5982 260006 6012 260058
rect 6036 260006 6046 260058
rect 6046 260006 6092 260058
rect 6116 260006 6162 260058
rect 6162 260006 6172 260058
rect 6196 260006 6226 260058
rect 6226 260006 6252 260058
rect 5956 260004 6012 260006
rect 6036 260004 6092 260006
rect 6116 260004 6172 260006
rect 6196 260004 6252 260006
rect 5956 258970 6012 258972
rect 6036 258970 6092 258972
rect 6116 258970 6172 258972
rect 6196 258970 6252 258972
rect 5956 258918 5982 258970
rect 5982 258918 6012 258970
rect 6036 258918 6046 258970
rect 6046 258918 6092 258970
rect 6116 258918 6162 258970
rect 6162 258918 6172 258970
rect 6196 258918 6226 258970
rect 6226 258918 6252 258970
rect 5956 258916 6012 258918
rect 6036 258916 6092 258918
rect 6116 258916 6172 258918
rect 6196 258916 6252 258918
rect 5956 257882 6012 257884
rect 6036 257882 6092 257884
rect 6116 257882 6172 257884
rect 6196 257882 6252 257884
rect 5956 257830 5982 257882
rect 5982 257830 6012 257882
rect 6036 257830 6046 257882
rect 6046 257830 6092 257882
rect 6116 257830 6162 257882
rect 6162 257830 6172 257882
rect 6196 257830 6226 257882
rect 6226 257830 6252 257882
rect 5956 257828 6012 257830
rect 6036 257828 6092 257830
rect 6116 257828 6172 257830
rect 6196 257828 6252 257830
rect 5956 256794 6012 256796
rect 6036 256794 6092 256796
rect 6116 256794 6172 256796
rect 6196 256794 6252 256796
rect 5956 256742 5982 256794
rect 5982 256742 6012 256794
rect 6036 256742 6046 256794
rect 6046 256742 6092 256794
rect 6116 256742 6162 256794
rect 6162 256742 6172 256794
rect 6196 256742 6226 256794
rect 6226 256742 6252 256794
rect 5956 256740 6012 256742
rect 6036 256740 6092 256742
rect 6116 256740 6172 256742
rect 6196 256740 6252 256742
rect 5956 255706 6012 255708
rect 6036 255706 6092 255708
rect 6116 255706 6172 255708
rect 6196 255706 6252 255708
rect 5956 255654 5982 255706
rect 5982 255654 6012 255706
rect 6036 255654 6046 255706
rect 6046 255654 6092 255706
rect 6116 255654 6162 255706
rect 6162 255654 6172 255706
rect 6196 255654 6226 255706
rect 6226 255654 6252 255706
rect 5956 255652 6012 255654
rect 6036 255652 6092 255654
rect 6116 255652 6172 255654
rect 6196 255652 6252 255654
rect 5956 254618 6012 254620
rect 6036 254618 6092 254620
rect 6116 254618 6172 254620
rect 6196 254618 6252 254620
rect 5956 254566 5982 254618
rect 5982 254566 6012 254618
rect 6036 254566 6046 254618
rect 6046 254566 6092 254618
rect 6116 254566 6162 254618
rect 6162 254566 6172 254618
rect 6196 254566 6226 254618
rect 6226 254566 6252 254618
rect 5956 254564 6012 254566
rect 6036 254564 6092 254566
rect 6116 254564 6172 254566
rect 6196 254564 6252 254566
rect 5956 253530 6012 253532
rect 6036 253530 6092 253532
rect 6116 253530 6172 253532
rect 6196 253530 6252 253532
rect 5956 253478 5982 253530
rect 5982 253478 6012 253530
rect 6036 253478 6046 253530
rect 6046 253478 6092 253530
rect 6116 253478 6162 253530
rect 6162 253478 6172 253530
rect 6196 253478 6226 253530
rect 6226 253478 6252 253530
rect 5956 253476 6012 253478
rect 6036 253476 6092 253478
rect 6116 253476 6172 253478
rect 6196 253476 6252 253478
rect 5956 252442 6012 252444
rect 6036 252442 6092 252444
rect 6116 252442 6172 252444
rect 6196 252442 6252 252444
rect 5956 252390 5982 252442
rect 5982 252390 6012 252442
rect 6036 252390 6046 252442
rect 6046 252390 6092 252442
rect 6116 252390 6162 252442
rect 6162 252390 6172 252442
rect 6196 252390 6226 252442
rect 6226 252390 6252 252442
rect 5956 252388 6012 252390
rect 6036 252388 6092 252390
rect 6116 252388 6172 252390
rect 6196 252388 6252 252390
rect 5956 251354 6012 251356
rect 6036 251354 6092 251356
rect 6116 251354 6172 251356
rect 6196 251354 6252 251356
rect 5956 251302 5982 251354
rect 5982 251302 6012 251354
rect 6036 251302 6046 251354
rect 6046 251302 6092 251354
rect 6116 251302 6162 251354
rect 6162 251302 6172 251354
rect 6196 251302 6226 251354
rect 6226 251302 6252 251354
rect 5956 251300 6012 251302
rect 6036 251300 6092 251302
rect 6116 251300 6172 251302
rect 6196 251300 6252 251302
rect 5956 250266 6012 250268
rect 6036 250266 6092 250268
rect 6116 250266 6172 250268
rect 6196 250266 6252 250268
rect 5956 250214 5982 250266
rect 5982 250214 6012 250266
rect 6036 250214 6046 250266
rect 6046 250214 6092 250266
rect 6116 250214 6162 250266
rect 6162 250214 6172 250266
rect 6196 250214 6226 250266
rect 6226 250214 6252 250266
rect 5956 250212 6012 250214
rect 6036 250212 6092 250214
rect 6116 250212 6172 250214
rect 6196 250212 6252 250214
rect 5956 249178 6012 249180
rect 6036 249178 6092 249180
rect 6116 249178 6172 249180
rect 6196 249178 6252 249180
rect 5956 249126 5982 249178
rect 5982 249126 6012 249178
rect 6036 249126 6046 249178
rect 6046 249126 6092 249178
rect 6116 249126 6162 249178
rect 6162 249126 6172 249178
rect 6196 249126 6226 249178
rect 6226 249126 6252 249178
rect 5956 249124 6012 249126
rect 6036 249124 6092 249126
rect 6116 249124 6172 249126
rect 6196 249124 6252 249126
rect 5956 248090 6012 248092
rect 6036 248090 6092 248092
rect 6116 248090 6172 248092
rect 6196 248090 6252 248092
rect 5956 248038 5982 248090
rect 5982 248038 6012 248090
rect 6036 248038 6046 248090
rect 6046 248038 6092 248090
rect 6116 248038 6162 248090
rect 6162 248038 6172 248090
rect 6196 248038 6226 248090
rect 6226 248038 6252 248090
rect 5956 248036 6012 248038
rect 6036 248036 6092 248038
rect 6116 248036 6172 248038
rect 6196 248036 6252 248038
rect 5956 247002 6012 247004
rect 6036 247002 6092 247004
rect 6116 247002 6172 247004
rect 6196 247002 6252 247004
rect 5956 246950 5982 247002
rect 5982 246950 6012 247002
rect 6036 246950 6046 247002
rect 6046 246950 6092 247002
rect 6116 246950 6162 247002
rect 6162 246950 6172 247002
rect 6196 246950 6226 247002
rect 6226 246950 6252 247002
rect 5956 246948 6012 246950
rect 6036 246948 6092 246950
rect 6116 246948 6172 246950
rect 6196 246948 6252 246950
rect 5956 245914 6012 245916
rect 6036 245914 6092 245916
rect 6116 245914 6172 245916
rect 6196 245914 6252 245916
rect 5956 245862 5982 245914
rect 5982 245862 6012 245914
rect 6036 245862 6046 245914
rect 6046 245862 6092 245914
rect 6116 245862 6162 245914
rect 6162 245862 6172 245914
rect 6196 245862 6226 245914
rect 6226 245862 6252 245914
rect 5956 245860 6012 245862
rect 6036 245860 6092 245862
rect 6116 245860 6172 245862
rect 6196 245860 6252 245862
rect 5956 244826 6012 244828
rect 6036 244826 6092 244828
rect 6116 244826 6172 244828
rect 6196 244826 6252 244828
rect 5956 244774 5982 244826
rect 5982 244774 6012 244826
rect 6036 244774 6046 244826
rect 6046 244774 6092 244826
rect 6116 244774 6162 244826
rect 6162 244774 6172 244826
rect 6196 244774 6226 244826
rect 6226 244774 6252 244826
rect 5956 244772 6012 244774
rect 6036 244772 6092 244774
rect 6116 244772 6172 244774
rect 6196 244772 6252 244774
rect 5956 243738 6012 243740
rect 6036 243738 6092 243740
rect 6116 243738 6172 243740
rect 6196 243738 6252 243740
rect 5956 243686 5982 243738
rect 5982 243686 6012 243738
rect 6036 243686 6046 243738
rect 6046 243686 6092 243738
rect 6116 243686 6162 243738
rect 6162 243686 6172 243738
rect 6196 243686 6226 243738
rect 6226 243686 6252 243738
rect 5956 243684 6012 243686
rect 6036 243684 6092 243686
rect 6116 243684 6172 243686
rect 6196 243684 6252 243686
rect 5956 242650 6012 242652
rect 6036 242650 6092 242652
rect 6116 242650 6172 242652
rect 6196 242650 6252 242652
rect 5956 242598 5982 242650
rect 5982 242598 6012 242650
rect 6036 242598 6046 242650
rect 6046 242598 6092 242650
rect 6116 242598 6162 242650
rect 6162 242598 6172 242650
rect 6196 242598 6226 242650
rect 6226 242598 6252 242650
rect 5956 242596 6012 242598
rect 6036 242596 6092 242598
rect 6116 242596 6172 242598
rect 6196 242596 6252 242598
rect 5956 241562 6012 241564
rect 6036 241562 6092 241564
rect 6116 241562 6172 241564
rect 6196 241562 6252 241564
rect 5956 241510 5982 241562
rect 5982 241510 6012 241562
rect 6036 241510 6046 241562
rect 6046 241510 6092 241562
rect 6116 241510 6162 241562
rect 6162 241510 6172 241562
rect 6196 241510 6226 241562
rect 6226 241510 6252 241562
rect 5956 241508 6012 241510
rect 6036 241508 6092 241510
rect 6116 241508 6172 241510
rect 6196 241508 6252 241510
rect 5956 240474 6012 240476
rect 6036 240474 6092 240476
rect 6116 240474 6172 240476
rect 6196 240474 6252 240476
rect 5956 240422 5982 240474
rect 5982 240422 6012 240474
rect 6036 240422 6046 240474
rect 6046 240422 6092 240474
rect 6116 240422 6162 240474
rect 6162 240422 6172 240474
rect 6196 240422 6226 240474
rect 6226 240422 6252 240474
rect 5956 240420 6012 240422
rect 6036 240420 6092 240422
rect 6116 240420 6172 240422
rect 6196 240420 6252 240422
rect 5956 239386 6012 239388
rect 6036 239386 6092 239388
rect 6116 239386 6172 239388
rect 6196 239386 6252 239388
rect 5956 239334 5982 239386
rect 5982 239334 6012 239386
rect 6036 239334 6046 239386
rect 6046 239334 6092 239386
rect 6116 239334 6162 239386
rect 6162 239334 6172 239386
rect 6196 239334 6226 239386
rect 6226 239334 6252 239386
rect 5956 239332 6012 239334
rect 6036 239332 6092 239334
rect 6116 239332 6172 239334
rect 6196 239332 6252 239334
rect 5956 238298 6012 238300
rect 6036 238298 6092 238300
rect 6116 238298 6172 238300
rect 6196 238298 6252 238300
rect 5956 238246 5982 238298
rect 5982 238246 6012 238298
rect 6036 238246 6046 238298
rect 6046 238246 6092 238298
rect 6116 238246 6162 238298
rect 6162 238246 6172 238298
rect 6196 238246 6226 238298
rect 6226 238246 6252 238298
rect 5956 238244 6012 238246
rect 6036 238244 6092 238246
rect 6116 238244 6172 238246
rect 6196 238244 6252 238246
rect 5956 237210 6012 237212
rect 6036 237210 6092 237212
rect 6116 237210 6172 237212
rect 6196 237210 6252 237212
rect 5956 237158 5982 237210
rect 5982 237158 6012 237210
rect 6036 237158 6046 237210
rect 6046 237158 6092 237210
rect 6116 237158 6162 237210
rect 6162 237158 6172 237210
rect 6196 237158 6226 237210
rect 6226 237158 6252 237210
rect 5956 237156 6012 237158
rect 6036 237156 6092 237158
rect 6116 237156 6172 237158
rect 6196 237156 6252 237158
rect 5956 236122 6012 236124
rect 6036 236122 6092 236124
rect 6116 236122 6172 236124
rect 6196 236122 6252 236124
rect 5956 236070 5982 236122
rect 5982 236070 6012 236122
rect 6036 236070 6046 236122
rect 6046 236070 6092 236122
rect 6116 236070 6162 236122
rect 6162 236070 6172 236122
rect 6196 236070 6226 236122
rect 6226 236070 6252 236122
rect 5956 236068 6012 236070
rect 6036 236068 6092 236070
rect 6116 236068 6172 236070
rect 6196 236068 6252 236070
rect 5956 235034 6012 235036
rect 6036 235034 6092 235036
rect 6116 235034 6172 235036
rect 6196 235034 6252 235036
rect 5956 234982 5982 235034
rect 5982 234982 6012 235034
rect 6036 234982 6046 235034
rect 6046 234982 6092 235034
rect 6116 234982 6162 235034
rect 6162 234982 6172 235034
rect 6196 234982 6226 235034
rect 6226 234982 6252 235034
rect 5956 234980 6012 234982
rect 6036 234980 6092 234982
rect 6116 234980 6172 234982
rect 6196 234980 6252 234982
rect 5956 233946 6012 233948
rect 6036 233946 6092 233948
rect 6116 233946 6172 233948
rect 6196 233946 6252 233948
rect 5956 233894 5982 233946
rect 5982 233894 6012 233946
rect 6036 233894 6046 233946
rect 6046 233894 6092 233946
rect 6116 233894 6162 233946
rect 6162 233894 6172 233946
rect 6196 233894 6226 233946
rect 6226 233894 6252 233946
rect 5956 233892 6012 233894
rect 6036 233892 6092 233894
rect 6116 233892 6172 233894
rect 6196 233892 6252 233894
rect 5956 232858 6012 232860
rect 6036 232858 6092 232860
rect 6116 232858 6172 232860
rect 6196 232858 6252 232860
rect 5956 232806 5982 232858
rect 5982 232806 6012 232858
rect 6036 232806 6046 232858
rect 6046 232806 6092 232858
rect 6116 232806 6162 232858
rect 6162 232806 6172 232858
rect 6196 232806 6226 232858
rect 6226 232806 6252 232858
rect 5956 232804 6012 232806
rect 6036 232804 6092 232806
rect 6116 232804 6172 232806
rect 6196 232804 6252 232806
rect 5956 231770 6012 231772
rect 6036 231770 6092 231772
rect 6116 231770 6172 231772
rect 6196 231770 6252 231772
rect 5956 231718 5982 231770
rect 5982 231718 6012 231770
rect 6036 231718 6046 231770
rect 6046 231718 6092 231770
rect 6116 231718 6162 231770
rect 6162 231718 6172 231770
rect 6196 231718 6226 231770
rect 6226 231718 6252 231770
rect 5956 231716 6012 231718
rect 6036 231716 6092 231718
rect 6116 231716 6172 231718
rect 6196 231716 6252 231718
rect 5956 230682 6012 230684
rect 6036 230682 6092 230684
rect 6116 230682 6172 230684
rect 6196 230682 6252 230684
rect 5956 230630 5982 230682
rect 5982 230630 6012 230682
rect 6036 230630 6046 230682
rect 6046 230630 6092 230682
rect 6116 230630 6162 230682
rect 6162 230630 6172 230682
rect 6196 230630 6226 230682
rect 6226 230630 6252 230682
rect 5956 230628 6012 230630
rect 6036 230628 6092 230630
rect 6116 230628 6172 230630
rect 6196 230628 6252 230630
rect 5956 229594 6012 229596
rect 6036 229594 6092 229596
rect 6116 229594 6172 229596
rect 6196 229594 6252 229596
rect 5956 229542 5982 229594
rect 5982 229542 6012 229594
rect 6036 229542 6046 229594
rect 6046 229542 6092 229594
rect 6116 229542 6162 229594
rect 6162 229542 6172 229594
rect 6196 229542 6226 229594
rect 6226 229542 6252 229594
rect 5956 229540 6012 229542
rect 6036 229540 6092 229542
rect 6116 229540 6172 229542
rect 6196 229540 6252 229542
rect 5956 228506 6012 228508
rect 6036 228506 6092 228508
rect 6116 228506 6172 228508
rect 6196 228506 6252 228508
rect 5956 228454 5982 228506
rect 5982 228454 6012 228506
rect 6036 228454 6046 228506
rect 6046 228454 6092 228506
rect 6116 228454 6162 228506
rect 6162 228454 6172 228506
rect 6196 228454 6226 228506
rect 6226 228454 6252 228506
rect 5956 228452 6012 228454
rect 6036 228452 6092 228454
rect 6116 228452 6172 228454
rect 6196 228452 6252 228454
rect 5956 227418 6012 227420
rect 6036 227418 6092 227420
rect 6116 227418 6172 227420
rect 6196 227418 6252 227420
rect 5956 227366 5982 227418
rect 5982 227366 6012 227418
rect 6036 227366 6046 227418
rect 6046 227366 6092 227418
rect 6116 227366 6162 227418
rect 6162 227366 6172 227418
rect 6196 227366 6226 227418
rect 6226 227366 6252 227418
rect 5956 227364 6012 227366
rect 6036 227364 6092 227366
rect 6116 227364 6172 227366
rect 6196 227364 6252 227366
rect 5956 226330 6012 226332
rect 6036 226330 6092 226332
rect 6116 226330 6172 226332
rect 6196 226330 6252 226332
rect 5956 226278 5982 226330
rect 5982 226278 6012 226330
rect 6036 226278 6046 226330
rect 6046 226278 6092 226330
rect 6116 226278 6162 226330
rect 6162 226278 6172 226330
rect 6196 226278 6226 226330
rect 6226 226278 6252 226330
rect 5956 226276 6012 226278
rect 6036 226276 6092 226278
rect 6116 226276 6172 226278
rect 6196 226276 6252 226278
rect 6366 249192 6422 249248
rect 7622 330234 7678 330236
rect 7702 330234 7758 330236
rect 7782 330234 7838 330236
rect 7862 330234 7918 330236
rect 7622 330182 7648 330234
rect 7648 330182 7678 330234
rect 7702 330182 7712 330234
rect 7712 330182 7758 330234
rect 7782 330182 7828 330234
rect 7828 330182 7838 330234
rect 7862 330182 7892 330234
rect 7892 330182 7918 330234
rect 7622 330180 7678 330182
rect 7702 330180 7758 330182
rect 7782 330180 7838 330182
rect 7862 330180 7918 330182
rect 7622 329146 7678 329148
rect 7702 329146 7758 329148
rect 7782 329146 7838 329148
rect 7862 329146 7918 329148
rect 7622 329094 7648 329146
rect 7648 329094 7678 329146
rect 7702 329094 7712 329146
rect 7712 329094 7758 329146
rect 7782 329094 7828 329146
rect 7828 329094 7838 329146
rect 7862 329094 7892 329146
rect 7892 329094 7918 329146
rect 7622 329092 7678 329094
rect 7702 329092 7758 329094
rect 7782 329092 7838 329094
rect 7862 329092 7918 329094
rect 7622 328058 7678 328060
rect 7702 328058 7758 328060
rect 7782 328058 7838 328060
rect 7862 328058 7918 328060
rect 7622 328006 7648 328058
rect 7648 328006 7678 328058
rect 7702 328006 7712 328058
rect 7712 328006 7758 328058
rect 7782 328006 7828 328058
rect 7828 328006 7838 328058
rect 7862 328006 7892 328058
rect 7892 328006 7918 328058
rect 7622 328004 7678 328006
rect 7702 328004 7758 328006
rect 7782 328004 7838 328006
rect 7862 328004 7918 328006
rect 7622 326970 7678 326972
rect 7702 326970 7758 326972
rect 7782 326970 7838 326972
rect 7862 326970 7918 326972
rect 7622 326918 7648 326970
rect 7648 326918 7678 326970
rect 7702 326918 7712 326970
rect 7712 326918 7758 326970
rect 7782 326918 7828 326970
rect 7828 326918 7838 326970
rect 7862 326918 7892 326970
rect 7892 326918 7918 326970
rect 7622 326916 7678 326918
rect 7702 326916 7758 326918
rect 7782 326916 7838 326918
rect 7862 326916 7918 326918
rect 7622 325882 7678 325884
rect 7702 325882 7758 325884
rect 7782 325882 7838 325884
rect 7862 325882 7918 325884
rect 7622 325830 7648 325882
rect 7648 325830 7678 325882
rect 7702 325830 7712 325882
rect 7712 325830 7758 325882
rect 7782 325830 7828 325882
rect 7828 325830 7838 325882
rect 7862 325830 7892 325882
rect 7892 325830 7918 325882
rect 7622 325828 7678 325830
rect 7702 325828 7758 325830
rect 7782 325828 7838 325830
rect 7862 325828 7918 325830
rect 7622 324794 7678 324796
rect 7702 324794 7758 324796
rect 7782 324794 7838 324796
rect 7862 324794 7918 324796
rect 7622 324742 7648 324794
rect 7648 324742 7678 324794
rect 7702 324742 7712 324794
rect 7712 324742 7758 324794
rect 7782 324742 7828 324794
rect 7828 324742 7838 324794
rect 7862 324742 7892 324794
rect 7892 324742 7918 324794
rect 7622 324740 7678 324742
rect 7702 324740 7758 324742
rect 7782 324740 7838 324742
rect 7862 324740 7918 324742
rect 7622 323706 7678 323708
rect 7702 323706 7758 323708
rect 7782 323706 7838 323708
rect 7862 323706 7918 323708
rect 7622 323654 7648 323706
rect 7648 323654 7678 323706
rect 7702 323654 7712 323706
rect 7712 323654 7758 323706
rect 7782 323654 7828 323706
rect 7828 323654 7838 323706
rect 7862 323654 7892 323706
rect 7892 323654 7918 323706
rect 7622 323652 7678 323654
rect 7702 323652 7758 323654
rect 7782 323652 7838 323654
rect 7862 323652 7918 323654
rect 7622 322618 7678 322620
rect 7702 322618 7758 322620
rect 7782 322618 7838 322620
rect 7862 322618 7918 322620
rect 7622 322566 7648 322618
rect 7648 322566 7678 322618
rect 7702 322566 7712 322618
rect 7712 322566 7758 322618
rect 7782 322566 7828 322618
rect 7828 322566 7838 322618
rect 7862 322566 7892 322618
rect 7892 322566 7918 322618
rect 7622 322564 7678 322566
rect 7702 322564 7758 322566
rect 7782 322564 7838 322566
rect 7862 322564 7918 322566
rect 7622 321530 7678 321532
rect 7702 321530 7758 321532
rect 7782 321530 7838 321532
rect 7862 321530 7918 321532
rect 7622 321478 7648 321530
rect 7648 321478 7678 321530
rect 7702 321478 7712 321530
rect 7712 321478 7758 321530
rect 7782 321478 7828 321530
rect 7828 321478 7838 321530
rect 7862 321478 7892 321530
rect 7892 321478 7918 321530
rect 7622 321476 7678 321478
rect 7702 321476 7758 321478
rect 7782 321476 7838 321478
rect 7862 321476 7918 321478
rect 7622 320442 7678 320444
rect 7702 320442 7758 320444
rect 7782 320442 7838 320444
rect 7862 320442 7918 320444
rect 7622 320390 7648 320442
rect 7648 320390 7678 320442
rect 7702 320390 7712 320442
rect 7712 320390 7758 320442
rect 7782 320390 7828 320442
rect 7828 320390 7838 320442
rect 7862 320390 7892 320442
rect 7892 320390 7918 320442
rect 7622 320388 7678 320390
rect 7702 320388 7758 320390
rect 7782 320388 7838 320390
rect 7862 320388 7918 320390
rect 7622 319354 7678 319356
rect 7702 319354 7758 319356
rect 7782 319354 7838 319356
rect 7862 319354 7918 319356
rect 7622 319302 7648 319354
rect 7648 319302 7678 319354
rect 7702 319302 7712 319354
rect 7712 319302 7758 319354
rect 7782 319302 7828 319354
rect 7828 319302 7838 319354
rect 7862 319302 7892 319354
rect 7892 319302 7918 319354
rect 7622 319300 7678 319302
rect 7702 319300 7758 319302
rect 7782 319300 7838 319302
rect 7862 319300 7918 319302
rect 7622 318266 7678 318268
rect 7702 318266 7758 318268
rect 7782 318266 7838 318268
rect 7862 318266 7918 318268
rect 7622 318214 7648 318266
rect 7648 318214 7678 318266
rect 7702 318214 7712 318266
rect 7712 318214 7758 318266
rect 7782 318214 7828 318266
rect 7828 318214 7838 318266
rect 7862 318214 7892 318266
rect 7892 318214 7918 318266
rect 7622 318212 7678 318214
rect 7702 318212 7758 318214
rect 7782 318212 7838 318214
rect 7862 318212 7918 318214
rect 7622 317178 7678 317180
rect 7702 317178 7758 317180
rect 7782 317178 7838 317180
rect 7862 317178 7918 317180
rect 7622 317126 7648 317178
rect 7648 317126 7678 317178
rect 7702 317126 7712 317178
rect 7712 317126 7758 317178
rect 7782 317126 7828 317178
rect 7828 317126 7838 317178
rect 7862 317126 7892 317178
rect 7892 317126 7918 317178
rect 7622 317124 7678 317126
rect 7702 317124 7758 317126
rect 7782 317124 7838 317126
rect 7862 317124 7918 317126
rect 7622 316090 7678 316092
rect 7702 316090 7758 316092
rect 7782 316090 7838 316092
rect 7862 316090 7918 316092
rect 7622 316038 7648 316090
rect 7648 316038 7678 316090
rect 7702 316038 7712 316090
rect 7712 316038 7758 316090
rect 7782 316038 7828 316090
rect 7828 316038 7838 316090
rect 7862 316038 7892 316090
rect 7892 316038 7918 316090
rect 7622 316036 7678 316038
rect 7702 316036 7758 316038
rect 7782 316036 7838 316038
rect 7862 316036 7918 316038
rect 7286 315832 7342 315888
rect 5956 225242 6012 225244
rect 6036 225242 6092 225244
rect 6116 225242 6172 225244
rect 6196 225242 6252 225244
rect 5956 225190 5982 225242
rect 5982 225190 6012 225242
rect 6036 225190 6046 225242
rect 6046 225190 6092 225242
rect 6116 225190 6162 225242
rect 6162 225190 6172 225242
rect 6196 225190 6226 225242
rect 6226 225190 6252 225242
rect 5956 225188 6012 225190
rect 6036 225188 6092 225190
rect 6116 225188 6172 225190
rect 6196 225188 6252 225190
rect 5956 224154 6012 224156
rect 6036 224154 6092 224156
rect 6116 224154 6172 224156
rect 6196 224154 6252 224156
rect 5956 224102 5982 224154
rect 5982 224102 6012 224154
rect 6036 224102 6046 224154
rect 6046 224102 6092 224154
rect 6116 224102 6162 224154
rect 6162 224102 6172 224154
rect 6196 224102 6226 224154
rect 6226 224102 6252 224154
rect 5956 224100 6012 224102
rect 6036 224100 6092 224102
rect 6116 224100 6172 224102
rect 6196 224100 6252 224102
rect 5956 223066 6012 223068
rect 6036 223066 6092 223068
rect 6116 223066 6172 223068
rect 6196 223066 6252 223068
rect 5956 223014 5982 223066
rect 5982 223014 6012 223066
rect 6036 223014 6046 223066
rect 6046 223014 6092 223066
rect 6116 223014 6162 223066
rect 6162 223014 6172 223066
rect 6196 223014 6226 223066
rect 6226 223014 6252 223066
rect 5956 223012 6012 223014
rect 6036 223012 6092 223014
rect 6116 223012 6172 223014
rect 6196 223012 6252 223014
rect 5956 221978 6012 221980
rect 6036 221978 6092 221980
rect 6116 221978 6172 221980
rect 6196 221978 6252 221980
rect 5956 221926 5982 221978
rect 5982 221926 6012 221978
rect 6036 221926 6046 221978
rect 6046 221926 6092 221978
rect 6116 221926 6162 221978
rect 6162 221926 6172 221978
rect 6196 221926 6226 221978
rect 6226 221926 6252 221978
rect 5956 221924 6012 221926
rect 6036 221924 6092 221926
rect 6116 221924 6172 221926
rect 6196 221924 6252 221926
rect 5956 220890 6012 220892
rect 6036 220890 6092 220892
rect 6116 220890 6172 220892
rect 6196 220890 6252 220892
rect 5956 220838 5982 220890
rect 5982 220838 6012 220890
rect 6036 220838 6046 220890
rect 6046 220838 6092 220890
rect 6116 220838 6162 220890
rect 6162 220838 6172 220890
rect 6196 220838 6226 220890
rect 6226 220838 6252 220890
rect 5956 220836 6012 220838
rect 6036 220836 6092 220838
rect 6116 220836 6172 220838
rect 6196 220836 6252 220838
rect 5956 219802 6012 219804
rect 6036 219802 6092 219804
rect 6116 219802 6172 219804
rect 6196 219802 6252 219804
rect 5956 219750 5982 219802
rect 5982 219750 6012 219802
rect 6036 219750 6046 219802
rect 6046 219750 6092 219802
rect 6116 219750 6162 219802
rect 6162 219750 6172 219802
rect 6196 219750 6226 219802
rect 6226 219750 6252 219802
rect 5956 219748 6012 219750
rect 6036 219748 6092 219750
rect 6116 219748 6172 219750
rect 6196 219748 6252 219750
rect 5956 218714 6012 218716
rect 6036 218714 6092 218716
rect 6116 218714 6172 218716
rect 6196 218714 6252 218716
rect 5956 218662 5982 218714
rect 5982 218662 6012 218714
rect 6036 218662 6046 218714
rect 6046 218662 6092 218714
rect 6116 218662 6162 218714
rect 6162 218662 6172 218714
rect 6196 218662 6226 218714
rect 6226 218662 6252 218714
rect 5956 218660 6012 218662
rect 6036 218660 6092 218662
rect 6116 218660 6172 218662
rect 6196 218660 6252 218662
rect 5956 217626 6012 217628
rect 6036 217626 6092 217628
rect 6116 217626 6172 217628
rect 6196 217626 6252 217628
rect 5956 217574 5982 217626
rect 5982 217574 6012 217626
rect 6036 217574 6046 217626
rect 6046 217574 6092 217626
rect 6116 217574 6162 217626
rect 6162 217574 6172 217626
rect 6196 217574 6226 217626
rect 6226 217574 6252 217626
rect 5956 217572 6012 217574
rect 6036 217572 6092 217574
rect 6116 217572 6172 217574
rect 6196 217572 6252 217574
rect 5956 216538 6012 216540
rect 6036 216538 6092 216540
rect 6116 216538 6172 216540
rect 6196 216538 6252 216540
rect 5956 216486 5982 216538
rect 5982 216486 6012 216538
rect 6036 216486 6046 216538
rect 6046 216486 6092 216538
rect 6116 216486 6162 216538
rect 6162 216486 6172 216538
rect 6196 216486 6226 216538
rect 6226 216486 6252 216538
rect 5956 216484 6012 216486
rect 6036 216484 6092 216486
rect 6116 216484 6172 216486
rect 6196 216484 6252 216486
rect 5956 215450 6012 215452
rect 6036 215450 6092 215452
rect 6116 215450 6172 215452
rect 6196 215450 6252 215452
rect 5956 215398 5982 215450
rect 5982 215398 6012 215450
rect 6036 215398 6046 215450
rect 6046 215398 6092 215450
rect 6116 215398 6162 215450
rect 6162 215398 6172 215450
rect 6196 215398 6226 215450
rect 6226 215398 6252 215450
rect 5956 215396 6012 215398
rect 6036 215396 6092 215398
rect 6116 215396 6172 215398
rect 6196 215396 6252 215398
rect 5956 214362 6012 214364
rect 6036 214362 6092 214364
rect 6116 214362 6172 214364
rect 6196 214362 6252 214364
rect 5956 214310 5982 214362
rect 5982 214310 6012 214362
rect 6036 214310 6046 214362
rect 6046 214310 6092 214362
rect 6116 214310 6162 214362
rect 6162 214310 6172 214362
rect 6196 214310 6226 214362
rect 6226 214310 6252 214362
rect 5956 214308 6012 214310
rect 6036 214308 6092 214310
rect 6116 214308 6172 214310
rect 6196 214308 6252 214310
rect 5956 213274 6012 213276
rect 6036 213274 6092 213276
rect 6116 213274 6172 213276
rect 6196 213274 6252 213276
rect 5956 213222 5982 213274
rect 5982 213222 6012 213274
rect 6036 213222 6046 213274
rect 6046 213222 6092 213274
rect 6116 213222 6162 213274
rect 6162 213222 6172 213274
rect 6196 213222 6226 213274
rect 6226 213222 6252 213274
rect 5956 213220 6012 213222
rect 6036 213220 6092 213222
rect 6116 213220 6172 213222
rect 6196 213220 6252 213222
rect 5956 212186 6012 212188
rect 6036 212186 6092 212188
rect 6116 212186 6172 212188
rect 6196 212186 6252 212188
rect 5956 212134 5982 212186
rect 5982 212134 6012 212186
rect 6036 212134 6046 212186
rect 6046 212134 6092 212186
rect 6116 212134 6162 212186
rect 6162 212134 6172 212186
rect 6196 212134 6226 212186
rect 6226 212134 6252 212186
rect 5956 212132 6012 212134
rect 6036 212132 6092 212134
rect 6116 212132 6172 212134
rect 6196 212132 6252 212134
rect 5956 211098 6012 211100
rect 6036 211098 6092 211100
rect 6116 211098 6172 211100
rect 6196 211098 6252 211100
rect 5956 211046 5982 211098
rect 5982 211046 6012 211098
rect 6036 211046 6046 211098
rect 6046 211046 6092 211098
rect 6116 211046 6162 211098
rect 6162 211046 6172 211098
rect 6196 211046 6226 211098
rect 6226 211046 6252 211098
rect 5956 211044 6012 211046
rect 6036 211044 6092 211046
rect 6116 211044 6172 211046
rect 6196 211044 6252 211046
rect 5956 210010 6012 210012
rect 6036 210010 6092 210012
rect 6116 210010 6172 210012
rect 6196 210010 6252 210012
rect 5956 209958 5982 210010
rect 5982 209958 6012 210010
rect 6036 209958 6046 210010
rect 6046 209958 6092 210010
rect 6116 209958 6162 210010
rect 6162 209958 6172 210010
rect 6196 209958 6226 210010
rect 6226 209958 6252 210010
rect 5956 209956 6012 209958
rect 6036 209956 6092 209958
rect 6116 209956 6172 209958
rect 6196 209956 6252 209958
rect 5956 208922 6012 208924
rect 6036 208922 6092 208924
rect 6116 208922 6172 208924
rect 6196 208922 6252 208924
rect 5956 208870 5982 208922
rect 5982 208870 6012 208922
rect 6036 208870 6046 208922
rect 6046 208870 6092 208922
rect 6116 208870 6162 208922
rect 6162 208870 6172 208922
rect 6196 208870 6226 208922
rect 6226 208870 6252 208922
rect 5956 208868 6012 208870
rect 6036 208868 6092 208870
rect 6116 208868 6172 208870
rect 6196 208868 6252 208870
rect 5956 207834 6012 207836
rect 6036 207834 6092 207836
rect 6116 207834 6172 207836
rect 6196 207834 6252 207836
rect 5956 207782 5982 207834
rect 5982 207782 6012 207834
rect 6036 207782 6046 207834
rect 6046 207782 6092 207834
rect 6116 207782 6162 207834
rect 6162 207782 6172 207834
rect 6196 207782 6226 207834
rect 6226 207782 6252 207834
rect 5956 207780 6012 207782
rect 6036 207780 6092 207782
rect 6116 207780 6172 207782
rect 6196 207780 6252 207782
rect 5956 206746 6012 206748
rect 6036 206746 6092 206748
rect 6116 206746 6172 206748
rect 6196 206746 6252 206748
rect 5956 206694 5982 206746
rect 5982 206694 6012 206746
rect 6036 206694 6046 206746
rect 6046 206694 6092 206746
rect 6116 206694 6162 206746
rect 6162 206694 6172 206746
rect 6196 206694 6226 206746
rect 6226 206694 6252 206746
rect 5956 206692 6012 206694
rect 6036 206692 6092 206694
rect 6116 206692 6172 206694
rect 6196 206692 6252 206694
rect 5956 205658 6012 205660
rect 6036 205658 6092 205660
rect 6116 205658 6172 205660
rect 6196 205658 6252 205660
rect 5956 205606 5982 205658
rect 5982 205606 6012 205658
rect 6036 205606 6046 205658
rect 6046 205606 6092 205658
rect 6116 205606 6162 205658
rect 6162 205606 6172 205658
rect 6196 205606 6226 205658
rect 6226 205606 6252 205658
rect 5956 205604 6012 205606
rect 6036 205604 6092 205606
rect 6116 205604 6172 205606
rect 6196 205604 6252 205606
rect 5956 204570 6012 204572
rect 6036 204570 6092 204572
rect 6116 204570 6172 204572
rect 6196 204570 6252 204572
rect 5956 204518 5982 204570
rect 5982 204518 6012 204570
rect 6036 204518 6046 204570
rect 6046 204518 6092 204570
rect 6116 204518 6162 204570
rect 6162 204518 6172 204570
rect 6196 204518 6226 204570
rect 6226 204518 6252 204570
rect 5956 204516 6012 204518
rect 6036 204516 6092 204518
rect 6116 204516 6172 204518
rect 6196 204516 6252 204518
rect 5956 203482 6012 203484
rect 6036 203482 6092 203484
rect 6116 203482 6172 203484
rect 6196 203482 6252 203484
rect 5956 203430 5982 203482
rect 5982 203430 6012 203482
rect 6036 203430 6046 203482
rect 6046 203430 6092 203482
rect 6116 203430 6162 203482
rect 6162 203430 6172 203482
rect 6196 203430 6226 203482
rect 6226 203430 6252 203482
rect 5956 203428 6012 203430
rect 6036 203428 6092 203430
rect 6116 203428 6172 203430
rect 6196 203428 6252 203430
rect 5956 202394 6012 202396
rect 6036 202394 6092 202396
rect 6116 202394 6172 202396
rect 6196 202394 6252 202396
rect 5956 202342 5982 202394
rect 5982 202342 6012 202394
rect 6036 202342 6046 202394
rect 6046 202342 6092 202394
rect 6116 202342 6162 202394
rect 6162 202342 6172 202394
rect 6196 202342 6226 202394
rect 6226 202342 6252 202394
rect 5956 202340 6012 202342
rect 6036 202340 6092 202342
rect 6116 202340 6172 202342
rect 6196 202340 6252 202342
rect 5956 201306 6012 201308
rect 6036 201306 6092 201308
rect 6116 201306 6172 201308
rect 6196 201306 6252 201308
rect 5956 201254 5982 201306
rect 5982 201254 6012 201306
rect 6036 201254 6046 201306
rect 6046 201254 6092 201306
rect 6116 201254 6162 201306
rect 6162 201254 6172 201306
rect 6196 201254 6226 201306
rect 6226 201254 6252 201306
rect 5956 201252 6012 201254
rect 6036 201252 6092 201254
rect 6116 201252 6172 201254
rect 6196 201252 6252 201254
rect 5956 200218 6012 200220
rect 6036 200218 6092 200220
rect 6116 200218 6172 200220
rect 6196 200218 6252 200220
rect 5956 200166 5982 200218
rect 5982 200166 6012 200218
rect 6036 200166 6046 200218
rect 6046 200166 6092 200218
rect 6116 200166 6162 200218
rect 6162 200166 6172 200218
rect 6196 200166 6226 200218
rect 6226 200166 6252 200218
rect 5956 200164 6012 200166
rect 6036 200164 6092 200166
rect 6116 200164 6172 200166
rect 6196 200164 6252 200166
rect 5956 199130 6012 199132
rect 6036 199130 6092 199132
rect 6116 199130 6172 199132
rect 6196 199130 6252 199132
rect 5956 199078 5982 199130
rect 5982 199078 6012 199130
rect 6036 199078 6046 199130
rect 6046 199078 6092 199130
rect 6116 199078 6162 199130
rect 6162 199078 6172 199130
rect 6196 199078 6226 199130
rect 6226 199078 6252 199130
rect 5956 199076 6012 199078
rect 6036 199076 6092 199078
rect 6116 199076 6172 199078
rect 6196 199076 6252 199078
rect 5956 198042 6012 198044
rect 6036 198042 6092 198044
rect 6116 198042 6172 198044
rect 6196 198042 6252 198044
rect 5956 197990 5982 198042
rect 5982 197990 6012 198042
rect 6036 197990 6046 198042
rect 6046 197990 6092 198042
rect 6116 197990 6162 198042
rect 6162 197990 6172 198042
rect 6196 197990 6226 198042
rect 6226 197990 6252 198042
rect 5956 197988 6012 197990
rect 6036 197988 6092 197990
rect 6116 197988 6172 197990
rect 6196 197988 6252 197990
rect 5956 196954 6012 196956
rect 6036 196954 6092 196956
rect 6116 196954 6172 196956
rect 6196 196954 6252 196956
rect 5956 196902 5982 196954
rect 5982 196902 6012 196954
rect 6036 196902 6046 196954
rect 6046 196902 6092 196954
rect 6116 196902 6162 196954
rect 6162 196902 6172 196954
rect 6196 196902 6226 196954
rect 6226 196902 6252 196954
rect 5956 196900 6012 196902
rect 6036 196900 6092 196902
rect 6116 196900 6172 196902
rect 6196 196900 6252 196902
rect 5956 195866 6012 195868
rect 6036 195866 6092 195868
rect 6116 195866 6172 195868
rect 6196 195866 6252 195868
rect 5956 195814 5982 195866
rect 5982 195814 6012 195866
rect 6036 195814 6046 195866
rect 6046 195814 6092 195866
rect 6116 195814 6162 195866
rect 6162 195814 6172 195866
rect 6196 195814 6226 195866
rect 6226 195814 6252 195866
rect 5956 195812 6012 195814
rect 6036 195812 6092 195814
rect 6116 195812 6172 195814
rect 6196 195812 6252 195814
rect 5956 194778 6012 194780
rect 6036 194778 6092 194780
rect 6116 194778 6172 194780
rect 6196 194778 6252 194780
rect 5956 194726 5982 194778
rect 5982 194726 6012 194778
rect 6036 194726 6046 194778
rect 6046 194726 6092 194778
rect 6116 194726 6162 194778
rect 6162 194726 6172 194778
rect 6196 194726 6226 194778
rect 6226 194726 6252 194778
rect 5956 194724 6012 194726
rect 6036 194724 6092 194726
rect 6116 194724 6172 194726
rect 6196 194724 6252 194726
rect 5956 193690 6012 193692
rect 6036 193690 6092 193692
rect 6116 193690 6172 193692
rect 6196 193690 6252 193692
rect 5956 193638 5982 193690
rect 5982 193638 6012 193690
rect 6036 193638 6046 193690
rect 6046 193638 6092 193690
rect 6116 193638 6162 193690
rect 6162 193638 6172 193690
rect 6196 193638 6226 193690
rect 6226 193638 6252 193690
rect 5956 193636 6012 193638
rect 6036 193636 6092 193638
rect 6116 193636 6172 193638
rect 6196 193636 6252 193638
rect 5956 192602 6012 192604
rect 6036 192602 6092 192604
rect 6116 192602 6172 192604
rect 6196 192602 6252 192604
rect 5956 192550 5982 192602
rect 5982 192550 6012 192602
rect 6036 192550 6046 192602
rect 6046 192550 6092 192602
rect 6116 192550 6162 192602
rect 6162 192550 6172 192602
rect 6196 192550 6226 192602
rect 6226 192550 6252 192602
rect 5956 192548 6012 192550
rect 6036 192548 6092 192550
rect 6116 192548 6172 192550
rect 6196 192548 6252 192550
rect 5956 191514 6012 191516
rect 6036 191514 6092 191516
rect 6116 191514 6172 191516
rect 6196 191514 6252 191516
rect 5956 191462 5982 191514
rect 5982 191462 6012 191514
rect 6036 191462 6046 191514
rect 6046 191462 6092 191514
rect 6116 191462 6162 191514
rect 6162 191462 6172 191514
rect 6196 191462 6226 191514
rect 6226 191462 6252 191514
rect 5956 191460 6012 191462
rect 6036 191460 6092 191462
rect 6116 191460 6172 191462
rect 6196 191460 6252 191462
rect 5956 190426 6012 190428
rect 6036 190426 6092 190428
rect 6116 190426 6172 190428
rect 6196 190426 6252 190428
rect 5956 190374 5982 190426
rect 5982 190374 6012 190426
rect 6036 190374 6046 190426
rect 6046 190374 6092 190426
rect 6116 190374 6162 190426
rect 6162 190374 6172 190426
rect 6196 190374 6226 190426
rect 6226 190374 6252 190426
rect 5956 190372 6012 190374
rect 6036 190372 6092 190374
rect 6116 190372 6172 190374
rect 6196 190372 6252 190374
rect 5956 189338 6012 189340
rect 6036 189338 6092 189340
rect 6116 189338 6172 189340
rect 6196 189338 6252 189340
rect 5956 189286 5982 189338
rect 5982 189286 6012 189338
rect 6036 189286 6046 189338
rect 6046 189286 6092 189338
rect 6116 189286 6162 189338
rect 6162 189286 6172 189338
rect 6196 189286 6226 189338
rect 6226 189286 6252 189338
rect 5956 189284 6012 189286
rect 6036 189284 6092 189286
rect 6116 189284 6172 189286
rect 6196 189284 6252 189286
rect 5956 188250 6012 188252
rect 6036 188250 6092 188252
rect 6116 188250 6172 188252
rect 6196 188250 6252 188252
rect 5956 188198 5982 188250
rect 5982 188198 6012 188250
rect 6036 188198 6046 188250
rect 6046 188198 6092 188250
rect 6116 188198 6162 188250
rect 6162 188198 6172 188250
rect 6196 188198 6226 188250
rect 6226 188198 6252 188250
rect 5956 188196 6012 188198
rect 6036 188196 6092 188198
rect 6116 188196 6172 188198
rect 6196 188196 6252 188198
rect 5956 187162 6012 187164
rect 6036 187162 6092 187164
rect 6116 187162 6172 187164
rect 6196 187162 6252 187164
rect 5956 187110 5982 187162
rect 5982 187110 6012 187162
rect 6036 187110 6046 187162
rect 6046 187110 6092 187162
rect 6116 187110 6162 187162
rect 6162 187110 6172 187162
rect 6196 187110 6226 187162
rect 6226 187110 6252 187162
rect 5956 187108 6012 187110
rect 6036 187108 6092 187110
rect 6116 187108 6172 187110
rect 6196 187108 6252 187110
rect 5956 186074 6012 186076
rect 6036 186074 6092 186076
rect 6116 186074 6172 186076
rect 6196 186074 6252 186076
rect 5956 186022 5982 186074
rect 5982 186022 6012 186074
rect 6036 186022 6046 186074
rect 6046 186022 6092 186074
rect 6116 186022 6162 186074
rect 6162 186022 6172 186074
rect 6196 186022 6226 186074
rect 6226 186022 6252 186074
rect 5956 186020 6012 186022
rect 6036 186020 6092 186022
rect 6116 186020 6172 186022
rect 6196 186020 6252 186022
rect 5956 184986 6012 184988
rect 6036 184986 6092 184988
rect 6116 184986 6172 184988
rect 6196 184986 6252 184988
rect 5956 184934 5982 184986
rect 5982 184934 6012 184986
rect 6036 184934 6046 184986
rect 6046 184934 6092 184986
rect 6116 184934 6162 184986
rect 6162 184934 6172 184986
rect 6196 184934 6226 184986
rect 6226 184934 6252 184986
rect 5956 184932 6012 184934
rect 6036 184932 6092 184934
rect 6116 184932 6172 184934
rect 6196 184932 6252 184934
rect 5956 183898 6012 183900
rect 6036 183898 6092 183900
rect 6116 183898 6172 183900
rect 6196 183898 6252 183900
rect 5956 183846 5982 183898
rect 5982 183846 6012 183898
rect 6036 183846 6046 183898
rect 6046 183846 6092 183898
rect 6116 183846 6162 183898
rect 6162 183846 6172 183898
rect 6196 183846 6226 183898
rect 6226 183846 6252 183898
rect 5956 183844 6012 183846
rect 6036 183844 6092 183846
rect 6116 183844 6172 183846
rect 6196 183844 6252 183846
rect 5956 182810 6012 182812
rect 6036 182810 6092 182812
rect 6116 182810 6172 182812
rect 6196 182810 6252 182812
rect 5956 182758 5982 182810
rect 5982 182758 6012 182810
rect 6036 182758 6046 182810
rect 6046 182758 6092 182810
rect 6116 182758 6162 182810
rect 6162 182758 6172 182810
rect 6196 182758 6226 182810
rect 6226 182758 6252 182810
rect 5956 182756 6012 182758
rect 6036 182756 6092 182758
rect 6116 182756 6172 182758
rect 6196 182756 6252 182758
rect 5956 181722 6012 181724
rect 6036 181722 6092 181724
rect 6116 181722 6172 181724
rect 6196 181722 6252 181724
rect 5956 181670 5982 181722
rect 5982 181670 6012 181722
rect 6036 181670 6046 181722
rect 6046 181670 6092 181722
rect 6116 181670 6162 181722
rect 6162 181670 6172 181722
rect 6196 181670 6226 181722
rect 6226 181670 6252 181722
rect 5956 181668 6012 181670
rect 6036 181668 6092 181670
rect 6116 181668 6172 181670
rect 6196 181668 6252 181670
rect 5956 180634 6012 180636
rect 6036 180634 6092 180636
rect 6116 180634 6172 180636
rect 6196 180634 6252 180636
rect 5956 180582 5982 180634
rect 5982 180582 6012 180634
rect 6036 180582 6046 180634
rect 6046 180582 6092 180634
rect 6116 180582 6162 180634
rect 6162 180582 6172 180634
rect 6196 180582 6226 180634
rect 6226 180582 6252 180634
rect 5956 180580 6012 180582
rect 6036 180580 6092 180582
rect 6116 180580 6172 180582
rect 6196 180580 6252 180582
rect 5956 179546 6012 179548
rect 6036 179546 6092 179548
rect 6116 179546 6172 179548
rect 6196 179546 6252 179548
rect 5956 179494 5982 179546
rect 5982 179494 6012 179546
rect 6036 179494 6046 179546
rect 6046 179494 6092 179546
rect 6116 179494 6162 179546
rect 6162 179494 6172 179546
rect 6196 179494 6226 179546
rect 6226 179494 6252 179546
rect 5956 179492 6012 179494
rect 6036 179492 6092 179494
rect 6116 179492 6172 179494
rect 6196 179492 6252 179494
rect 5956 178458 6012 178460
rect 6036 178458 6092 178460
rect 6116 178458 6172 178460
rect 6196 178458 6252 178460
rect 5956 178406 5982 178458
rect 5982 178406 6012 178458
rect 6036 178406 6046 178458
rect 6046 178406 6092 178458
rect 6116 178406 6162 178458
rect 6162 178406 6172 178458
rect 6196 178406 6226 178458
rect 6226 178406 6252 178458
rect 5956 178404 6012 178406
rect 6036 178404 6092 178406
rect 6116 178404 6172 178406
rect 6196 178404 6252 178406
rect 5956 177370 6012 177372
rect 6036 177370 6092 177372
rect 6116 177370 6172 177372
rect 6196 177370 6252 177372
rect 5956 177318 5982 177370
rect 5982 177318 6012 177370
rect 6036 177318 6046 177370
rect 6046 177318 6092 177370
rect 6116 177318 6162 177370
rect 6162 177318 6172 177370
rect 6196 177318 6226 177370
rect 6226 177318 6252 177370
rect 5956 177316 6012 177318
rect 6036 177316 6092 177318
rect 6116 177316 6172 177318
rect 6196 177316 6252 177318
rect 5956 176282 6012 176284
rect 6036 176282 6092 176284
rect 6116 176282 6172 176284
rect 6196 176282 6252 176284
rect 5956 176230 5982 176282
rect 5982 176230 6012 176282
rect 6036 176230 6046 176282
rect 6046 176230 6092 176282
rect 6116 176230 6162 176282
rect 6162 176230 6172 176282
rect 6196 176230 6226 176282
rect 6226 176230 6252 176282
rect 5956 176228 6012 176230
rect 6036 176228 6092 176230
rect 6116 176228 6172 176230
rect 6196 176228 6252 176230
rect 5956 175194 6012 175196
rect 6036 175194 6092 175196
rect 6116 175194 6172 175196
rect 6196 175194 6252 175196
rect 5956 175142 5982 175194
rect 5982 175142 6012 175194
rect 6036 175142 6046 175194
rect 6046 175142 6092 175194
rect 6116 175142 6162 175194
rect 6162 175142 6172 175194
rect 6196 175142 6226 175194
rect 6226 175142 6252 175194
rect 5956 175140 6012 175142
rect 6036 175140 6092 175142
rect 6116 175140 6172 175142
rect 6196 175140 6252 175142
rect 5956 174106 6012 174108
rect 6036 174106 6092 174108
rect 6116 174106 6172 174108
rect 6196 174106 6252 174108
rect 5956 174054 5982 174106
rect 5982 174054 6012 174106
rect 6036 174054 6046 174106
rect 6046 174054 6092 174106
rect 6116 174054 6162 174106
rect 6162 174054 6172 174106
rect 6196 174054 6226 174106
rect 6226 174054 6252 174106
rect 5956 174052 6012 174054
rect 6036 174052 6092 174054
rect 6116 174052 6172 174054
rect 6196 174052 6252 174054
rect 5956 173018 6012 173020
rect 6036 173018 6092 173020
rect 6116 173018 6172 173020
rect 6196 173018 6252 173020
rect 5956 172966 5982 173018
rect 5982 172966 6012 173018
rect 6036 172966 6046 173018
rect 6046 172966 6092 173018
rect 6116 172966 6162 173018
rect 6162 172966 6172 173018
rect 6196 172966 6226 173018
rect 6226 172966 6252 173018
rect 5956 172964 6012 172966
rect 6036 172964 6092 172966
rect 6116 172964 6172 172966
rect 6196 172964 6252 172966
rect 7010 216144 7066 216200
rect 6642 182552 6698 182608
rect 5956 171930 6012 171932
rect 6036 171930 6092 171932
rect 6116 171930 6172 171932
rect 6196 171930 6252 171932
rect 5956 171878 5982 171930
rect 5982 171878 6012 171930
rect 6036 171878 6046 171930
rect 6046 171878 6092 171930
rect 6116 171878 6162 171930
rect 6162 171878 6172 171930
rect 6196 171878 6226 171930
rect 6226 171878 6252 171930
rect 5956 171876 6012 171878
rect 6036 171876 6092 171878
rect 6116 171876 6172 171878
rect 6196 171876 6252 171878
rect 5956 170842 6012 170844
rect 6036 170842 6092 170844
rect 6116 170842 6172 170844
rect 6196 170842 6252 170844
rect 5956 170790 5982 170842
rect 5982 170790 6012 170842
rect 6036 170790 6046 170842
rect 6046 170790 6092 170842
rect 6116 170790 6162 170842
rect 6162 170790 6172 170842
rect 6196 170790 6226 170842
rect 6226 170790 6252 170842
rect 5956 170788 6012 170790
rect 6036 170788 6092 170790
rect 6116 170788 6172 170790
rect 6196 170788 6252 170790
rect 5956 169754 6012 169756
rect 6036 169754 6092 169756
rect 6116 169754 6172 169756
rect 6196 169754 6252 169756
rect 5956 169702 5982 169754
rect 5982 169702 6012 169754
rect 6036 169702 6046 169754
rect 6046 169702 6092 169754
rect 6116 169702 6162 169754
rect 6162 169702 6172 169754
rect 6196 169702 6226 169754
rect 6226 169702 6252 169754
rect 5956 169700 6012 169702
rect 6036 169700 6092 169702
rect 6116 169700 6172 169702
rect 6196 169700 6252 169702
rect 5956 168666 6012 168668
rect 6036 168666 6092 168668
rect 6116 168666 6172 168668
rect 6196 168666 6252 168668
rect 5956 168614 5982 168666
rect 5982 168614 6012 168666
rect 6036 168614 6046 168666
rect 6046 168614 6092 168666
rect 6116 168614 6162 168666
rect 6162 168614 6172 168666
rect 6196 168614 6226 168666
rect 6226 168614 6252 168666
rect 5956 168612 6012 168614
rect 6036 168612 6092 168614
rect 6116 168612 6172 168614
rect 6196 168612 6252 168614
rect 5956 167578 6012 167580
rect 6036 167578 6092 167580
rect 6116 167578 6172 167580
rect 6196 167578 6252 167580
rect 5956 167526 5982 167578
rect 5982 167526 6012 167578
rect 6036 167526 6046 167578
rect 6046 167526 6092 167578
rect 6116 167526 6162 167578
rect 6162 167526 6172 167578
rect 6196 167526 6226 167578
rect 6226 167526 6252 167578
rect 5956 167524 6012 167526
rect 6036 167524 6092 167526
rect 6116 167524 6172 167526
rect 6196 167524 6252 167526
rect 5956 166490 6012 166492
rect 6036 166490 6092 166492
rect 6116 166490 6172 166492
rect 6196 166490 6252 166492
rect 5956 166438 5982 166490
rect 5982 166438 6012 166490
rect 6036 166438 6046 166490
rect 6046 166438 6092 166490
rect 6116 166438 6162 166490
rect 6162 166438 6172 166490
rect 6196 166438 6226 166490
rect 6226 166438 6252 166490
rect 5956 166436 6012 166438
rect 6036 166436 6092 166438
rect 6116 166436 6172 166438
rect 6196 166436 6252 166438
rect 5956 165402 6012 165404
rect 6036 165402 6092 165404
rect 6116 165402 6172 165404
rect 6196 165402 6252 165404
rect 5956 165350 5982 165402
rect 5982 165350 6012 165402
rect 6036 165350 6046 165402
rect 6046 165350 6092 165402
rect 6116 165350 6162 165402
rect 6162 165350 6172 165402
rect 6196 165350 6226 165402
rect 6226 165350 6252 165402
rect 5956 165348 6012 165350
rect 6036 165348 6092 165350
rect 6116 165348 6172 165350
rect 6196 165348 6252 165350
rect 5956 164314 6012 164316
rect 6036 164314 6092 164316
rect 6116 164314 6172 164316
rect 6196 164314 6252 164316
rect 5956 164262 5982 164314
rect 5982 164262 6012 164314
rect 6036 164262 6046 164314
rect 6046 164262 6092 164314
rect 6116 164262 6162 164314
rect 6162 164262 6172 164314
rect 6196 164262 6226 164314
rect 6226 164262 6252 164314
rect 5956 164260 6012 164262
rect 6036 164260 6092 164262
rect 6116 164260 6172 164262
rect 6196 164260 6252 164262
rect 5956 163226 6012 163228
rect 6036 163226 6092 163228
rect 6116 163226 6172 163228
rect 6196 163226 6252 163228
rect 5956 163174 5982 163226
rect 5982 163174 6012 163226
rect 6036 163174 6046 163226
rect 6046 163174 6092 163226
rect 6116 163174 6162 163226
rect 6162 163174 6172 163226
rect 6196 163174 6226 163226
rect 6226 163174 6252 163226
rect 5956 163172 6012 163174
rect 6036 163172 6092 163174
rect 6116 163172 6172 163174
rect 6196 163172 6252 163174
rect 5956 162138 6012 162140
rect 6036 162138 6092 162140
rect 6116 162138 6172 162140
rect 6196 162138 6252 162140
rect 5956 162086 5982 162138
rect 5982 162086 6012 162138
rect 6036 162086 6046 162138
rect 6046 162086 6092 162138
rect 6116 162086 6162 162138
rect 6162 162086 6172 162138
rect 6196 162086 6226 162138
rect 6226 162086 6252 162138
rect 5956 162084 6012 162086
rect 6036 162084 6092 162086
rect 6116 162084 6172 162086
rect 6196 162084 6252 162086
rect 5956 161050 6012 161052
rect 6036 161050 6092 161052
rect 6116 161050 6172 161052
rect 6196 161050 6252 161052
rect 5956 160998 5982 161050
rect 5982 160998 6012 161050
rect 6036 160998 6046 161050
rect 6046 160998 6092 161050
rect 6116 160998 6162 161050
rect 6162 160998 6172 161050
rect 6196 160998 6226 161050
rect 6226 160998 6252 161050
rect 5956 160996 6012 160998
rect 6036 160996 6092 160998
rect 6116 160996 6172 160998
rect 6196 160996 6252 160998
rect 5956 159962 6012 159964
rect 6036 159962 6092 159964
rect 6116 159962 6172 159964
rect 6196 159962 6252 159964
rect 5956 159910 5982 159962
rect 5982 159910 6012 159962
rect 6036 159910 6046 159962
rect 6046 159910 6092 159962
rect 6116 159910 6162 159962
rect 6162 159910 6172 159962
rect 6196 159910 6226 159962
rect 6226 159910 6252 159962
rect 5956 159908 6012 159910
rect 6036 159908 6092 159910
rect 6116 159908 6172 159910
rect 6196 159908 6252 159910
rect 5956 158874 6012 158876
rect 6036 158874 6092 158876
rect 6116 158874 6172 158876
rect 6196 158874 6252 158876
rect 5956 158822 5982 158874
rect 5982 158822 6012 158874
rect 6036 158822 6046 158874
rect 6046 158822 6092 158874
rect 6116 158822 6162 158874
rect 6162 158822 6172 158874
rect 6196 158822 6226 158874
rect 6226 158822 6252 158874
rect 5956 158820 6012 158822
rect 6036 158820 6092 158822
rect 6116 158820 6172 158822
rect 6196 158820 6252 158822
rect 5956 157786 6012 157788
rect 6036 157786 6092 157788
rect 6116 157786 6172 157788
rect 6196 157786 6252 157788
rect 5956 157734 5982 157786
rect 5982 157734 6012 157786
rect 6036 157734 6046 157786
rect 6046 157734 6092 157786
rect 6116 157734 6162 157786
rect 6162 157734 6172 157786
rect 6196 157734 6226 157786
rect 6226 157734 6252 157786
rect 5956 157732 6012 157734
rect 6036 157732 6092 157734
rect 6116 157732 6172 157734
rect 6196 157732 6252 157734
rect 5956 156698 6012 156700
rect 6036 156698 6092 156700
rect 6116 156698 6172 156700
rect 6196 156698 6252 156700
rect 5956 156646 5982 156698
rect 5982 156646 6012 156698
rect 6036 156646 6046 156698
rect 6046 156646 6092 156698
rect 6116 156646 6162 156698
rect 6162 156646 6172 156698
rect 6196 156646 6226 156698
rect 6226 156646 6252 156698
rect 5956 156644 6012 156646
rect 6036 156644 6092 156646
rect 6116 156644 6172 156646
rect 6196 156644 6252 156646
rect 5956 155610 6012 155612
rect 6036 155610 6092 155612
rect 6116 155610 6172 155612
rect 6196 155610 6252 155612
rect 5956 155558 5982 155610
rect 5982 155558 6012 155610
rect 6036 155558 6046 155610
rect 6046 155558 6092 155610
rect 6116 155558 6162 155610
rect 6162 155558 6172 155610
rect 6196 155558 6226 155610
rect 6226 155558 6252 155610
rect 5956 155556 6012 155558
rect 6036 155556 6092 155558
rect 6116 155556 6172 155558
rect 6196 155556 6252 155558
rect 5956 154522 6012 154524
rect 6036 154522 6092 154524
rect 6116 154522 6172 154524
rect 6196 154522 6252 154524
rect 5956 154470 5982 154522
rect 5982 154470 6012 154522
rect 6036 154470 6046 154522
rect 6046 154470 6092 154522
rect 6116 154470 6162 154522
rect 6162 154470 6172 154522
rect 6196 154470 6226 154522
rect 6226 154470 6252 154522
rect 5956 154468 6012 154470
rect 6036 154468 6092 154470
rect 6116 154468 6172 154470
rect 6196 154468 6252 154470
rect 5956 153434 6012 153436
rect 6036 153434 6092 153436
rect 6116 153434 6172 153436
rect 6196 153434 6252 153436
rect 5956 153382 5982 153434
rect 5982 153382 6012 153434
rect 6036 153382 6046 153434
rect 6046 153382 6092 153434
rect 6116 153382 6162 153434
rect 6162 153382 6172 153434
rect 6196 153382 6226 153434
rect 6226 153382 6252 153434
rect 5956 153380 6012 153382
rect 6036 153380 6092 153382
rect 6116 153380 6172 153382
rect 6196 153380 6252 153382
rect 5956 152346 6012 152348
rect 6036 152346 6092 152348
rect 6116 152346 6172 152348
rect 6196 152346 6252 152348
rect 5956 152294 5982 152346
rect 5982 152294 6012 152346
rect 6036 152294 6046 152346
rect 6046 152294 6092 152346
rect 6116 152294 6162 152346
rect 6162 152294 6172 152346
rect 6196 152294 6226 152346
rect 6226 152294 6252 152346
rect 5956 152292 6012 152294
rect 6036 152292 6092 152294
rect 6116 152292 6172 152294
rect 6196 152292 6252 152294
rect 5956 151258 6012 151260
rect 6036 151258 6092 151260
rect 6116 151258 6172 151260
rect 6196 151258 6252 151260
rect 5956 151206 5982 151258
rect 5982 151206 6012 151258
rect 6036 151206 6046 151258
rect 6046 151206 6092 151258
rect 6116 151206 6162 151258
rect 6162 151206 6172 151258
rect 6196 151206 6226 151258
rect 6226 151206 6252 151258
rect 5956 151204 6012 151206
rect 6036 151204 6092 151206
rect 6116 151204 6172 151206
rect 6196 151204 6252 151206
rect 5956 150170 6012 150172
rect 6036 150170 6092 150172
rect 6116 150170 6172 150172
rect 6196 150170 6252 150172
rect 5956 150118 5982 150170
rect 5982 150118 6012 150170
rect 6036 150118 6046 150170
rect 6046 150118 6092 150170
rect 6116 150118 6162 150170
rect 6162 150118 6172 150170
rect 6196 150118 6226 150170
rect 6226 150118 6252 150170
rect 5956 150116 6012 150118
rect 6036 150116 6092 150118
rect 6116 150116 6172 150118
rect 6196 150116 6252 150118
rect 5956 149082 6012 149084
rect 6036 149082 6092 149084
rect 6116 149082 6172 149084
rect 6196 149082 6252 149084
rect 5956 149030 5982 149082
rect 5982 149030 6012 149082
rect 6036 149030 6046 149082
rect 6046 149030 6092 149082
rect 6116 149030 6162 149082
rect 6162 149030 6172 149082
rect 6196 149030 6226 149082
rect 6226 149030 6252 149082
rect 5956 149028 6012 149030
rect 6036 149028 6092 149030
rect 6116 149028 6172 149030
rect 6196 149028 6252 149030
rect 5956 147994 6012 147996
rect 6036 147994 6092 147996
rect 6116 147994 6172 147996
rect 6196 147994 6252 147996
rect 5956 147942 5982 147994
rect 5982 147942 6012 147994
rect 6036 147942 6046 147994
rect 6046 147942 6092 147994
rect 6116 147942 6162 147994
rect 6162 147942 6172 147994
rect 6196 147942 6226 147994
rect 6226 147942 6252 147994
rect 5956 147940 6012 147942
rect 6036 147940 6092 147942
rect 6116 147940 6172 147942
rect 6196 147940 6252 147942
rect 5956 146906 6012 146908
rect 6036 146906 6092 146908
rect 6116 146906 6172 146908
rect 6196 146906 6252 146908
rect 5956 146854 5982 146906
rect 5982 146854 6012 146906
rect 6036 146854 6046 146906
rect 6046 146854 6092 146906
rect 6116 146854 6162 146906
rect 6162 146854 6172 146906
rect 6196 146854 6226 146906
rect 6226 146854 6252 146906
rect 5956 146852 6012 146854
rect 6036 146852 6092 146854
rect 6116 146852 6172 146854
rect 6196 146852 6252 146854
rect 5956 145818 6012 145820
rect 6036 145818 6092 145820
rect 6116 145818 6172 145820
rect 6196 145818 6252 145820
rect 5956 145766 5982 145818
rect 5982 145766 6012 145818
rect 6036 145766 6046 145818
rect 6046 145766 6092 145818
rect 6116 145766 6162 145818
rect 6162 145766 6172 145818
rect 6196 145766 6226 145818
rect 6226 145766 6252 145818
rect 5956 145764 6012 145766
rect 6036 145764 6092 145766
rect 6116 145764 6172 145766
rect 6196 145764 6252 145766
rect 5956 144730 6012 144732
rect 6036 144730 6092 144732
rect 6116 144730 6172 144732
rect 6196 144730 6252 144732
rect 5956 144678 5982 144730
rect 5982 144678 6012 144730
rect 6036 144678 6046 144730
rect 6046 144678 6092 144730
rect 6116 144678 6162 144730
rect 6162 144678 6172 144730
rect 6196 144678 6226 144730
rect 6226 144678 6252 144730
rect 5956 144676 6012 144678
rect 6036 144676 6092 144678
rect 6116 144676 6172 144678
rect 6196 144676 6252 144678
rect 5956 143642 6012 143644
rect 6036 143642 6092 143644
rect 6116 143642 6172 143644
rect 6196 143642 6252 143644
rect 5956 143590 5982 143642
rect 5982 143590 6012 143642
rect 6036 143590 6046 143642
rect 6046 143590 6092 143642
rect 6116 143590 6162 143642
rect 6162 143590 6172 143642
rect 6196 143590 6226 143642
rect 6226 143590 6252 143642
rect 5956 143588 6012 143590
rect 6036 143588 6092 143590
rect 6116 143588 6172 143590
rect 6196 143588 6252 143590
rect 5956 142554 6012 142556
rect 6036 142554 6092 142556
rect 6116 142554 6172 142556
rect 6196 142554 6252 142556
rect 5956 142502 5982 142554
rect 5982 142502 6012 142554
rect 6036 142502 6046 142554
rect 6046 142502 6092 142554
rect 6116 142502 6162 142554
rect 6162 142502 6172 142554
rect 6196 142502 6226 142554
rect 6226 142502 6252 142554
rect 5956 142500 6012 142502
rect 6036 142500 6092 142502
rect 6116 142500 6172 142502
rect 6196 142500 6252 142502
rect 5956 141466 6012 141468
rect 6036 141466 6092 141468
rect 6116 141466 6172 141468
rect 6196 141466 6252 141468
rect 5956 141414 5982 141466
rect 5982 141414 6012 141466
rect 6036 141414 6046 141466
rect 6046 141414 6092 141466
rect 6116 141414 6162 141466
rect 6162 141414 6172 141466
rect 6196 141414 6226 141466
rect 6226 141414 6252 141466
rect 5956 141412 6012 141414
rect 6036 141412 6092 141414
rect 6116 141412 6172 141414
rect 6196 141412 6252 141414
rect 5956 140378 6012 140380
rect 6036 140378 6092 140380
rect 6116 140378 6172 140380
rect 6196 140378 6252 140380
rect 5956 140326 5982 140378
rect 5982 140326 6012 140378
rect 6036 140326 6046 140378
rect 6046 140326 6092 140378
rect 6116 140326 6162 140378
rect 6162 140326 6172 140378
rect 6196 140326 6226 140378
rect 6226 140326 6252 140378
rect 5956 140324 6012 140326
rect 6036 140324 6092 140326
rect 6116 140324 6172 140326
rect 6196 140324 6252 140326
rect 5956 139290 6012 139292
rect 6036 139290 6092 139292
rect 6116 139290 6172 139292
rect 6196 139290 6252 139292
rect 5956 139238 5982 139290
rect 5982 139238 6012 139290
rect 6036 139238 6046 139290
rect 6046 139238 6092 139290
rect 6116 139238 6162 139290
rect 6162 139238 6172 139290
rect 6196 139238 6226 139290
rect 6226 139238 6252 139290
rect 5956 139236 6012 139238
rect 6036 139236 6092 139238
rect 6116 139236 6172 139238
rect 6196 139236 6252 139238
rect 5956 138202 6012 138204
rect 6036 138202 6092 138204
rect 6116 138202 6172 138204
rect 6196 138202 6252 138204
rect 5956 138150 5982 138202
rect 5982 138150 6012 138202
rect 6036 138150 6046 138202
rect 6046 138150 6092 138202
rect 6116 138150 6162 138202
rect 6162 138150 6172 138202
rect 6196 138150 6226 138202
rect 6226 138150 6252 138202
rect 5956 138148 6012 138150
rect 6036 138148 6092 138150
rect 6116 138148 6172 138150
rect 6196 138148 6252 138150
rect 5956 137114 6012 137116
rect 6036 137114 6092 137116
rect 6116 137114 6172 137116
rect 6196 137114 6252 137116
rect 5956 137062 5982 137114
rect 5982 137062 6012 137114
rect 6036 137062 6046 137114
rect 6046 137062 6092 137114
rect 6116 137062 6162 137114
rect 6162 137062 6172 137114
rect 6196 137062 6226 137114
rect 6226 137062 6252 137114
rect 5956 137060 6012 137062
rect 6036 137060 6092 137062
rect 6116 137060 6172 137062
rect 6196 137060 6252 137062
rect 5956 136026 6012 136028
rect 6036 136026 6092 136028
rect 6116 136026 6172 136028
rect 6196 136026 6252 136028
rect 5956 135974 5982 136026
rect 5982 135974 6012 136026
rect 6036 135974 6046 136026
rect 6046 135974 6092 136026
rect 6116 135974 6162 136026
rect 6162 135974 6172 136026
rect 6196 135974 6226 136026
rect 6226 135974 6252 136026
rect 5956 135972 6012 135974
rect 6036 135972 6092 135974
rect 6116 135972 6172 135974
rect 6196 135972 6252 135974
rect 5956 134938 6012 134940
rect 6036 134938 6092 134940
rect 6116 134938 6172 134940
rect 6196 134938 6252 134940
rect 5956 134886 5982 134938
rect 5982 134886 6012 134938
rect 6036 134886 6046 134938
rect 6046 134886 6092 134938
rect 6116 134886 6162 134938
rect 6162 134886 6172 134938
rect 6196 134886 6226 134938
rect 6226 134886 6252 134938
rect 5956 134884 6012 134886
rect 6036 134884 6092 134886
rect 6116 134884 6172 134886
rect 6196 134884 6252 134886
rect 5956 133850 6012 133852
rect 6036 133850 6092 133852
rect 6116 133850 6172 133852
rect 6196 133850 6252 133852
rect 5956 133798 5982 133850
rect 5982 133798 6012 133850
rect 6036 133798 6046 133850
rect 6046 133798 6092 133850
rect 6116 133798 6162 133850
rect 6162 133798 6172 133850
rect 6196 133798 6226 133850
rect 6226 133798 6252 133850
rect 5956 133796 6012 133798
rect 6036 133796 6092 133798
rect 6116 133796 6172 133798
rect 6196 133796 6252 133798
rect 5956 132762 6012 132764
rect 6036 132762 6092 132764
rect 6116 132762 6172 132764
rect 6196 132762 6252 132764
rect 5956 132710 5982 132762
rect 5982 132710 6012 132762
rect 6036 132710 6046 132762
rect 6046 132710 6092 132762
rect 6116 132710 6162 132762
rect 6162 132710 6172 132762
rect 6196 132710 6226 132762
rect 6226 132710 6252 132762
rect 5956 132708 6012 132710
rect 6036 132708 6092 132710
rect 6116 132708 6172 132710
rect 6196 132708 6252 132710
rect 5956 131674 6012 131676
rect 6036 131674 6092 131676
rect 6116 131674 6172 131676
rect 6196 131674 6252 131676
rect 5956 131622 5982 131674
rect 5982 131622 6012 131674
rect 6036 131622 6046 131674
rect 6046 131622 6092 131674
rect 6116 131622 6162 131674
rect 6162 131622 6172 131674
rect 6196 131622 6226 131674
rect 6226 131622 6252 131674
rect 5956 131620 6012 131622
rect 6036 131620 6092 131622
rect 6116 131620 6172 131622
rect 6196 131620 6252 131622
rect 5956 130586 6012 130588
rect 6036 130586 6092 130588
rect 6116 130586 6172 130588
rect 6196 130586 6252 130588
rect 5956 130534 5982 130586
rect 5982 130534 6012 130586
rect 6036 130534 6046 130586
rect 6046 130534 6092 130586
rect 6116 130534 6162 130586
rect 6162 130534 6172 130586
rect 6196 130534 6226 130586
rect 6226 130534 6252 130586
rect 5956 130532 6012 130534
rect 6036 130532 6092 130534
rect 6116 130532 6172 130534
rect 6196 130532 6252 130534
rect 5956 129498 6012 129500
rect 6036 129498 6092 129500
rect 6116 129498 6172 129500
rect 6196 129498 6252 129500
rect 5956 129446 5982 129498
rect 5982 129446 6012 129498
rect 6036 129446 6046 129498
rect 6046 129446 6092 129498
rect 6116 129446 6162 129498
rect 6162 129446 6172 129498
rect 6196 129446 6226 129498
rect 6226 129446 6252 129498
rect 5956 129444 6012 129446
rect 6036 129444 6092 129446
rect 6116 129444 6172 129446
rect 6196 129444 6252 129446
rect 5956 128410 6012 128412
rect 6036 128410 6092 128412
rect 6116 128410 6172 128412
rect 6196 128410 6252 128412
rect 5956 128358 5982 128410
rect 5982 128358 6012 128410
rect 6036 128358 6046 128410
rect 6046 128358 6092 128410
rect 6116 128358 6162 128410
rect 6162 128358 6172 128410
rect 6196 128358 6226 128410
rect 6226 128358 6252 128410
rect 5956 128356 6012 128358
rect 6036 128356 6092 128358
rect 6116 128356 6172 128358
rect 6196 128356 6252 128358
rect 5956 127322 6012 127324
rect 6036 127322 6092 127324
rect 6116 127322 6172 127324
rect 6196 127322 6252 127324
rect 5956 127270 5982 127322
rect 5982 127270 6012 127322
rect 6036 127270 6046 127322
rect 6046 127270 6092 127322
rect 6116 127270 6162 127322
rect 6162 127270 6172 127322
rect 6196 127270 6226 127322
rect 6226 127270 6252 127322
rect 5956 127268 6012 127270
rect 6036 127268 6092 127270
rect 6116 127268 6172 127270
rect 6196 127268 6252 127270
rect 5956 126234 6012 126236
rect 6036 126234 6092 126236
rect 6116 126234 6172 126236
rect 6196 126234 6252 126236
rect 5956 126182 5982 126234
rect 5982 126182 6012 126234
rect 6036 126182 6046 126234
rect 6046 126182 6092 126234
rect 6116 126182 6162 126234
rect 6162 126182 6172 126234
rect 6196 126182 6226 126234
rect 6226 126182 6252 126234
rect 5956 126180 6012 126182
rect 6036 126180 6092 126182
rect 6116 126180 6172 126182
rect 6196 126180 6252 126182
rect 5956 125146 6012 125148
rect 6036 125146 6092 125148
rect 6116 125146 6172 125148
rect 6196 125146 6252 125148
rect 5956 125094 5982 125146
rect 5982 125094 6012 125146
rect 6036 125094 6046 125146
rect 6046 125094 6092 125146
rect 6116 125094 6162 125146
rect 6162 125094 6172 125146
rect 6196 125094 6226 125146
rect 6226 125094 6252 125146
rect 5956 125092 6012 125094
rect 6036 125092 6092 125094
rect 6116 125092 6172 125094
rect 6196 125092 6252 125094
rect 5956 124058 6012 124060
rect 6036 124058 6092 124060
rect 6116 124058 6172 124060
rect 6196 124058 6252 124060
rect 5956 124006 5982 124058
rect 5982 124006 6012 124058
rect 6036 124006 6046 124058
rect 6046 124006 6092 124058
rect 6116 124006 6162 124058
rect 6162 124006 6172 124058
rect 6196 124006 6226 124058
rect 6226 124006 6252 124058
rect 5956 124004 6012 124006
rect 6036 124004 6092 124006
rect 6116 124004 6172 124006
rect 6196 124004 6252 124006
rect 5956 122970 6012 122972
rect 6036 122970 6092 122972
rect 6116 122970 6172 122972
rect 6196 122970 6252 122972
rect 5956 122918 5982 122970
rect 5982 122918 6012 122970
rect 6036 122918 6046 122970
rect 6046 122918 6092 122970
rect 6116 122918 6162 122970
rect 6162 122918 6172 122970
rect 6196 122918 6226 122970
rect 6226 122918 6252 122970
rect 5956 122916 6012 122918
rect 6036 122916 6092 122918
rect 6116 122916 6172 122918
rect 6196 122916 6252 122918
rect 5956 121882 6012 121884
rect 6036 121882 6092 121884
rect 6116 121882 6172 121884
rect 6196 121882 6252 121884
rect 5956 121830 5982 121882
rect 5982 121830 6012 121882
rect 6036 121830 6046 121882
rect 6046 121830 6092 121882
rect 6116 121830 6162 121882
rect 6162 121830 6172 121882
rect 6196 121830 6226 121882
rect 6226 121830 6252 121882
rect 5956 121828 6012 121830
rect 6036 121828 6092 121830
rect 6116 121828 6172 121830
rect 6196 121828 6252 121830
rect 5956 120794 6012 120796
rect 6036 120794 6092 120796
rect 6116 120794 6172 120796
rect 6196 120794 6252 120796
rect 5956 120742 5982 120794
rect 5982 120742 6012 120794
rect 6036 120742 6046 120794
rect 6046 120742 6092 120794
rect 6116 120742 6162 120794
rect 6162 120742 6172 120794
rect 6196 120742 6226 120794
rect 6226 120742 6252 120794
rect 5956 120740 6012 120742
rect 6036 120740 6092 120742
rect 6116 120740 6172 120742
rect 6196 120740 6252 120742
rect 5956 119706 6012 119708
rect 6036 119706 6092 119708
rect 6116 119706 6172 119708
rect 6196 119706 6252 119708
rect 5956 119654 5982 119706
rect 5982 119654 6012 119706
rect 6036 119654 6046 119706
rect 6046 119654 6092 119706
rect 6116 119654 6162 119706
rect 6162 119654 6172 119706
rect 6196 119654 6226 119706
rect 6226 119654 6252 119706
rect 5956 119652 6012 119654
rect 6036 119652 6092 119654
rect 6116 119652 6172 119654
rect 6196 119652 6252 119654
rect 5956 118618 6012 118620
rect 6036 118618 6092 118620
rect 6116 118618 6172 118620
rect 6196 118618 6252 118620
rect 5956 118566 5982 118618
rect 5982 118566 6012 118618
rect 6036 118566 6046 118618
rect 6046 118566 6092 118618
rect 6116 118566 6162 118618
rect 6162 118566 6172 118618
rect 6196 118566 6226 118618
rect 6226 118566 6252 118618
rect 5956 118564 6012 118566
rect 6036 118564 6092 118566
rect 6116 118564 6172 118566
rect 6196 118564 6252 118566
rect 5956 117530 6012 117532
rect 6036 117530 6092 117532
rect 6116 117530 6172 117532
rect 6196 117530 6252 117532
rect 5956 117478 5982 117530
rect 5982 117478 6012 117530
rect 6036 117478 6046 117530
rect 6046 117478 6092 117530
rect 6116 117478 6162 117530
rect 6162 117478 6172 117530
rect 6196 117478 6226 117530
rect 6226 117478 6252 117530
rect 5956 117476 6012 117478
rect 6036 117476 6092 117478
rect 6116 117476 6172 117478
rect 6196 117476 6252 117478
rect 7622 315002 7678 315004
rect 7702 315002 7758 315004
rect 7782 315002 7838 315004
rect 7862 315002 7918 315004
rect 7622 314950 7648 315002
rect 7648 314950 7678 315002
rect 7702 314950 7712 315002
rect 7712 314950 7758 315002
rect 7782 314950 7828 315002
rect 7828 314950 7838 315002
rect 7862 314950 7892 315002
rect 7892 314950 7918 315002
rect 7622 314948 7678 314950
rect 7702 314948 7758 314950
rect 7782 314948 7838 314950
rect 7862 314948 7918 314950
rect 7622 313914 7678 313916
rect 7702 313914 7758 313916
rect 7782 313914 7838 313916
rect 7862 313914 7918 313916
rect 7622 313862 7648 313914
rect 7648 313862 7678 313914
rect 7702 313862 7712 313914
rect 7712 313862 7758 313914
rect 7782 313862 7828 313914
rect 7828 313862 7838 313914
rect 7862 313862 7892 313914
rect 7892 313862 7918 313914
rect 7622 313860 7678 313862
rect 7702 313860 7758 313862
rect 7782 313860 7838 313862
rect 7862 313860 7918 313862
rect 7622 312826 7678 312828
rect 7702 312826 7758 312828
rect 7782 312826 7838 312828
rect 7862 312826 7918 312828
rect 7622 312774 7648 312826
rect 7648 312774 7678 312826
rect 7702 312774 7712 312826
rect 7712 312774 7758 312826
rect 7782 312774 7828 312826
rect 7828 312774 7838 312826
rect 7862 312774 7892 312826
rect 7892 312774 7918 312826
rect 7622 312772 7678 312774
rect 7702 312772 7758 312774
rect 7782 312772 7838 312774
rect 7862 312772 7918 312774
rect 7622 311738 7678 311740
rect 7702 311738 7758 311740
rect 7782 311738 7838 311740
rect 7862 311738 7918 311740
rect 7622 311686 7648 311738
rect 7648 311686 7678 311738
rect 7702 311686 7712 311738
rect 7712 311686 7758 311738
rect 7782 311686 7828 311738
rect 7828 311686 7838 311738
rect 7862 311686 7892 311738
rect 7892 311686 7918 311738
rect 7622 311684 7678 311686
rect 7702 311684 7758 311686
rect 7782 311684 7838 311686
rect 7862 311684 7918 311686
rect 7622 310650 7678 310652
rect 7702 310650 7758 310652
rect 7782 310650 7838 310652
rect 7862 310650 7918 310652
rect 7622 310598 7648 310650
rect 7648 310598 7678 310650
rect 7702 310598 7712 310650
rect 7712 310598 7758 310650
rect 7782 310598 7828 310650
rect 7828 310598 7838 310650
rect 7862 310598 7892 310650
rect 7892 310598 7918 310650
rect 7622 310596 7678 310598
rect 7702 310596 7758 310598
rect 7782 310596 7838 310598
rect 7862 310596 7918 310598
rect 7622 309562 7678 309564
rect 7702 309562 7758 309564
rect 7782 309562 7838 309564
rect 7862 309562 7918 309564
rect 7622 309510 7648 309562
rect 7648 309510 7678 309562
rect 7702 309510 7712 309562
rect 7712 309510 7758 309562
rect 7782 309510 7828 309562
rect 7828 309510 7838 309562
rect 7862 309510 7892 309562
rect 7892 309510 7918 309562
rect 7622 309508 7678 309510
rect 7702 309508 7758 309510
rect 7782 309508 7838 309510
rect 7862 309508 7918 309510
rect 7622 308474 7678 308476
rect 7702 308474 7758 308476
rect 7782 308474 7838 308476
rect 7862 308474 7918 308476
rect 7622 308422 7648 308474
rect 7648 308422 7678 308474
rect 7702 308422 7712 308474
rect 7712 308422 7758 308474
rect 7782 308422 7828 308474
rect 7828 308422 7838 308474
rect 7862 308422 7892 308474
rect 7892 308422 7918 308474
rect 7622 308420 7678 308422
rect 7702 308420 7758 308422
rect 7782 308420 7838 308422
rect 7862 308420 7918 308422
rect 7622 307386 7678 307388
rect 7702 307386 7758 307388
rect 7782 307386 7838 307388
rect 7862 307386 7918 307388
rect 7622 307334 7648 307386
rect 7648 307334 7678 307386
rect 7702 307334 7712 307386
rect 7712 307334 7758 307386
rect 7782 307334 7828 307386
rect 7828 307334 7838 307386
rect 7862 307334 7892 307386
rect 7892 307334 7918 307386
rect 7622 307332 7678 307334
rect 7702 307332 7758 307334
rect 7782 307332 7838 307334
rect 7862 307332 7918 307334
rect 7622 306298 7678 306300
rect 7702 306298 7758 306300
rect 7782 306298 7838 306300
rect 7862 306298 7918 306300
rect 7622 306246 7648 306298
rect 7648 306246 7678 306298
rect 7702 306246 7712 306298
rect 7712 306246 7758 306298
rect 7782 306246 7828 306298
rect 7828 306246 7838 306298
rect 7862 306246 7892 306298
rect 7892 306246 7918 306298
rect 7622 306244 7678 306246
rect 7702 306244 7758 306246
rect 7782 306244 7838 306246
rect 7862 306244 7918 306246
rect 7622 305210 7678 305212
rect 7702 305210 7758 305212
rect 7782 305210 7838 305212
rect 7862 305210 7918 305212
rect 7622 305158 7648 305210
rect 7648 305158 7678 305210
rect 7702 305158 7712 305210
rect 7712 305158 7758 305210
rect 7782 305158 7828 305210
rect 7828 305158 7838 305210
rect 7862 305158 7892 305210
rect 7892 305158 7918 305210
rect 7622 305156 7678 305158
rect 7702 305156 7758 305158
rect 7782 305156 7838 305158
rect 7862 305156 7918 305158
rect 7622 304122 7678 304124
rect 7702 304122 7758 304124
rect 7782 304122 7838 304124
rect 7862 304122 7918 304124
rect 7622 304070 7648 304122
rect 7648 304070 7678 304122
rect 7702 304070 7712 304122
rect 7712 304070 7758 304122
rect 7782 304070 7828 304122
rect 7828 304070 7838 304122
rect 7862 304070 7892 304122
rect 7892 304070 7918 304122
rect 7622 304068 7678 304070
rect 7702 304068 7758 304070
rect 7782 304068 7838 304070
rect 7862 304068 7918 304070
rect 7622 303034 7678 303036
rect 7702 303034 7758 303036
rect 7782 303034 7838 303036
rect 7862 303034 7918 303036
rect 7622 302982 7648 303034
rect 7648 302982 7678 303034
rect 7702 302982 7712 303034
rect 7712 302982 7758 303034
rect 7782 302982 7828 303034
rect 7828 302982 7838 303034
rect 7862 302982 7892 303034
rect 7892 302982 7918 303034
rect 7622 302980 7678 302982
rect 7702 302980 7758 302982
rect 7782 302980 7838 302982
rect 7862 302980 7918 302982
rect 7622 301946 7678 301948
rect 7702 301946 7758 301948
rect 7782 301946 7838 301948
rect 7862 301946 7918 301948
rect 7622 301894 7648 301946
rect 7648 301894 7678 301946
rect 7702 301894 7712 301946
rect 7712 301894 7758 301946
rect 7782 301894 7828 301946
rect 7828 301894 7838 301946
rect 7862 301894 7892 301946
rect 7892 301894 7918 301946
rect 7622 301892 7678 301894
rect 7702 301892 7758 301894
rect 7782 301892 7838 301894
rect 7862 301892 7918 301894
rect 7622 300858 7678 300860
rect 7702 300858 7758 300860
rect 7782 300858 7838 300860
rect 7862 300858 7918 300860
rect 7622 300806 7648 300858
rect 7648 300806 7678 300858
rect 7702 300806 7712 300858
rect 7712 300806 7758 300858
rect 7782 300806 7828 300858
rect 7828 300806 7838 300858
rect 7862 300806 7892 300858
rect 7892 300806 7918 300858
rect 7622 300804 7678 300806
rect 7702 300804 7758 300806
rect 7782 300804 7838 300806
rect 7862 300804 7918 300806
rect 7622 299770 7678 299772
rect 7702 299770 7758 299772
rect 7782 299770 7838 299772
rect 7862 299770 7918 299772
rect 7622 299718 7648 299770
rect 7648 299718 7678 299770
rect 7702 299718 7712 299770
rect 7712 299718 7758 299770
rect 7782 299718 7828 299770
rect 7828 299718 7838 299770
rect 7862 299718 7892 299770
rect 7892 299718 7918 299770
rect 7622 299716 7678 299718
rect 7702 299716 7758 299718
rect 7782 299716 7838 299718
rect 7862 299716 7918 299718
rect 7622 298682 7678 298684
rect 7702 298682 7758 298684
rect 7782 298682 7838 298684
rect 7862 298682 7918 298684
rect 7622 298630 7648 298682
rect 7648 298630 7678 298682
rect 7702 298630 7712 298682
rect 7712 298630 7758 298682
rect 7782 298630 7828 298682
rect 7828 298630 7838 298682
rect 7862 298630 7892 298682
rect 7892 298630 7918 298682
rect 7622 298628 7678 298630
rect 7702 298628 7758 298630
rect 7782 298628 7838 298630
rect 7862 298628 7918 298630
rect 7622 297594 7678 297596
rect 7702 297594 7758 297596
rect 7782 297594 7838 297596
rect 7862 297594 7918 297596
rect 7622 297542 7648 297594
rect 7648 297542 7678 297594
rect 7702 297542 7712 297594
rect 7712 297542 7758 297594
rect 7782 297542 7828 297594
rect 7828 297542 7838 297594
rect 7862 297542 7892 297594
rect 7892 297542 7918 297594
rect 7622 297540 7678 297542
rect 7702 297540 7758 297542
rect 7782 297540 7838 297542
rect 7862 297540 7918 297542
rect 7622 296506 7678 296508
rect 7702 296506 7758 296508
rect 7782 296506 7838 296508
rect 7862 296506 7918 296508
rect 7622 296454 7648 296506
rect 7648 296454 7678 296506
rect 7702 296454 7712 296506
rect 7712 296454 7758 296506
rect 7782 296454 7828 296506
rect 7828 296454 7838 296506
rect 7862 296454 7892 296506
rect 7892 296454 7918 296506
rect 7622 296452 7678 296454
rect 7702 296452 7758 296454
rect 7782 296452 7838 296454
rect 7862 296452 7918 296454
rect 7622 295418 7678 295420
rect 7702 295418 7758 295420
rect 7782 295418 7838 295420
rect 7862 295418 7918 295420
rect 7622 295366 7648 295418
rect 7648 295366 7678 295418
rect 7702 295366 7712 295418
rect 7712 295366 7758 295418
rect 7782 295366 7828 295418
rect 7828 295366 7838 295418
rect 7862 295366 7892 295418
rect 7892 295366 7918 295418
rect 7622 295364 7678 295366
rect 7702 295364 7758 295366
rect 7782 295364 7838 295366
rect 7862 295364 7918 295366
rect 7622 294330 7678 294332
rect 7702 294330 7758 294332
rect 7782 294330 7838 294332
rect 7862 294330 7918 294332
rect 7622 294278 7648 294330
rect 7648 294278 7678 294330
rect 7702 294278 7712 294330
rect 7712 294278 7758 294330
rect 7782 294278 7828 294330
rect 7828 294278 7838 294330
rect 7862 294278 7892 294330
rect 7892 294278 7918 294330
rect 7622 294276 7678 294278
rect 7702 294276 7758 294278
rect 7782 294276 7838 294278
rect 7862 294276 7918 294278
rect 7622 293242 7678 293244
rect 7702 293242 7758 293244
rect 7782 293242 7838 293244
rect 7862 293242 7918 293244
rect 7622 293190 7648 293242
rect 7648 293190 7678 293242
rect 7702 293190 7712 293242
rect 7712 293190 7758 293242
rect 7782 293190 7828 293242
rect 7828 293190 7838 293242
rect 7862 293190 7892 293242
rect 7892 293190 7918 293242
rect 7622 293188 7678 293190
rect 7702 293188 7758 293190
rect 7782 293188 7838 293190
rect 7862 293188 7918 293190
rect 7622 292154 7678 292156
rect 7702 292154 7758 292156
rect 7782 292154 7838 292156
rect 7862 292154 7918 292156
rect 7622 292102 7648 292154
rect 7648 292102 7678 292154
rect 7702 292102 7712 292154
rect 7712 292102 7758 292154
rect 7782 292102 7828 292154
rect 7828 292102 7838 292154
rect 7862 292102 7892 292154
rect 7892 292102 7918 292154
rect 7622 292100 7678 292102
rect 7702 292100 7758 292102
rect 7782 292100 7838 292102
rect 7862 292100 7918 292102
rect 7622 291066 7678 291068
rect 7702 291066 7758 291068
rect 7782 291066 7838 291068
rect 7862 291066 7918 291068
rect 7622 291014 7648 291066
rect 7648 291014 7678 291066
rect 7702 291014 7712 291066
rect 7712 291014 7758 291066
rect 7782 291014 7828 291066
rect 7828 291014 7838 291066
rect 7862 291014 7892 291066
rect 7892 291014 7918 291066
rect 7622 291012 7678 291014
rect 7702 291012 7758 291014
rect 7782 291012 7838 291014
rect 7862 291012 7918 291014
rect 7622 289978 7678 289980
rect 7702 289978 7758 289980
rect 7782 289978 7838 289980
rect 7862 289978 7918 289980
rect 7622 289926 7648 289978
rect 7648 289926 7678 289978
rect 7702 289926 7712 289978
rect 7712 289926 7758 289978
rect 7782 289926 7828 289978
rect 7828 289926 7838 289978
rect 7862 289926 7892 289978
rect 7892 289926 7918 289978
rect 7622 289924 7678 289926
rect 7702 289924 7758 289926
rect 7782 289924 7838 289926
rect 7862 289924 7918 289926
rect 7622 288890 7678 288892
rect 7702 288890 7758 288892
rect 7782 288890 7838 288892
rect 7862 288890 7918 288892
rect 7622 288838 7648 288890
rect 7648 288838 7678 288890
rect 7702 288838 7712 288890
rect 7712 288838 7758 288890
rect 7782 288838 7828 288890
rect 7828 288838 7838 288890
rect 7862 288838 7892 288890
rect 7892 288838 7918 288890
rect 7622 288836 7678 288838
rect 7702 288836 7758 288838
rect 7782 288836 7838 288838
rect 7862 288836 7918 288838
rect 7622 287802 7678 287804
rect 7702 287802 7758 287804
rect 7782 287802 7838 287804
rect 7862 287802 7918 287804
rect 7622 287750 7648 287802
rect 7648 287750 7678 287802
rect 7702 287750 7712 287802
rect 7712 287750 7758 287802
rect 7782 287750 7828 287802
rect 7828 287750 7838 287802
rect 7862 287750 7892 287802
rect 7892 287750 7918 287802
rect 7622 287748 7678 287750
rect 7702 287748 7758 287750
rect 7782 287748 7838 287750
rect 7862 287748 7918 287750
rect 7622 286714 7678 286716
rect 7702 286714 7758 286716
rect 7782 286714 7838 286716
rect 7862 286714 7918 286716
rect 7622 286662 7648 286714
rect 7648 286662 7678 286714
rect 7702 286662 7712 286714
rect 7712 286662 7758 286714
rect 7782 286662 7828 286714
rect 7828 286662 7838 286714
rect 7862 286662 7892 286714
rect 7892 286662 7918 286714
rect 7622 286660 7678 286662
rect 7702 286660 7758 286662
rect 7782 286660 7838 286662
rect 7862 286660 7918 286662
rect 7622 285626 7678 285628
rect 7702 285626 7758 285628
rect 7782 285626 7838 285628
rect 7862 285626 7918 285628
rect 7622 285574 7648 285626
rect 7648 285574 7678 285626
rect 7702 285574 7712 285626
rect 7712 285574 7758 285626
rect 7782 285574 7828 285626
rect 7828 285574 7838 285626
rect 7862 285574 7892 285626
rect 7892 285574 7918 285626
rect 7622 285572 7678 285574
rect 7702 285572 7758 285574
rect 7782 285572 7838 285574
rect 7862 285572 7918 285574
rect 7622 284538 7678 284540
rect 7702 284538 7758 284540
rect 7782 284538 7838 284540
rect 7862 284538 7918 284540
rect 7622 284486 7648 284538
rect 7648 284486 7678 284538
rect 7702 284486 7712 284538
rect 7712 284486 7758 284538
rect 7782 284486 7828 284538
rect 7828 284486 7838 284538
rect 7862 284486 7892 284538
rect 7892 284486 7918 284538
rect 7622 284484 7678 284486
rect 7702 284484 7758 284486
rect 7782 284484 7838 284486
rect 7862 284484 7918 284486
rect 7622 283450 7678 283452
rect 7702 283450 7758 283452
rect 7782 283450 7838 283452
rect 7862 283450 7918 283452
rect 7622 283398 7648 283450
rect 7648 283398 7678 283450
rect 7702 283398 7712 283450
rect 7712 283398 7758 283450
rect 7782 283398 7828 283450
rect 7828 283398 7838 283450
rect 7862 283398 7892 283450
rect 7892 283398 7918 283450
rect 7622 283396 7678 283398
rect 7702 283396 7758 283398
rect 7782 283396 7838 283398
rect 7862 283396 7918 283398
rect 7622 282362 7678 282364
rect 7702 282362 7758 282364
rect 7782 282362 7838 282364
rect 7862 282362 7918 282364
rect 7622 282310 7648 282362
rect 7648 282310 7678 282362
rect 7702 282310 7712 282362
rect 7712 282310 7758 282362
rect 7782 282310 7828 282362
rect 7828 282310 7838 282362
rect 7862 282310 7892 282362
rect 7892 282310 7918 282362
rect 7622 282308 7678 282310
rect 7702 282308 7758 282310
rect 7782 282308 7838 282310
rect 7862 282308 7918 282310
rect 7622 281274 7678 281276
rect 7702 281274 7758 281276
rect 7782 281274 7838 281276
rect 7862 281274 7918 281276
rect 7622 281222 7648 281274
rect 7648 281222 7678 281274
rect 7702 281222 7712 281274
rect 7712 281222 7758 281274
rect 7782 281222 7828 281274
rect 7828 281222 7838 281274
rect 7862 281222 7892 281274
rect 7892 281222 7918 281274
rect 7622 281220 7678 281222
rect 7702 281220 7758 281222
rect 7782 281220 7838 281222
rect 7862 281220 7918 281222
rect 7622 280186 7678 280188
rect 7702 280186 7758 280188
rect 7782 280186 7838 280188
rect 7862 280186 7918 280188
rect 7622 280134 7648 280186
rect 7648 280134 7678 280186
rect 7702 280134 7712 280186
rect 7712 280134 7758 280186
rect 7782 280134 7828 280186
rect 7828 280134 7838 280186
rect 7862 280134 7892 280186
rect 7892 280134 7918 280186
rect 7622 280132 7678 280134
rect 7702 280132 7758 280134
rect 7782 280132 7838 280134
rect 7862 280132 7918 280134
rect 7622 279098 7678 279100
rect 7702 279098 7758 279100
rect 7782 279098 7838 279100
rect 7862 279098 7918 279100
rect 7622 279046 7648 279098
rect 7648 279046 7678 279098
rect 7702 279046 7712 279098
rect 7712 279046 7758 279098
rect 7782 279046 7828 279098
rect 7828 279046 7838 279098
rect 7862 279046 7892 279098
rect 7892 279046 7918 279098
rect 7622 279044 7678 279046
rect 7702 279044 7758 279046
rect 7782 279044 7838 279046
rect 7862 279044 7918 279046
rect 7622 278010 7678 278012
rect 7702 278010 7758 278012
rect 7782 278010 7838 278012
rect 7862 278010 7918 278012
rect 7622 277958 7648 278010
rect 7648 277958 7678 278010
rect 7702 277958 7712 278010
rect 7712 277958 7758 278010
rect 7782 277958 7828 278010
rect 7828 277958 7838 278010
rect 7862 277958 7892 278010
rect 7892 277958 7918 278010
rect 7622 277956 7678 277958
rect 7702 277956 7758 277958
rect 7782 277956 7838 277958
rect 7862 277956 7918 277958
rect 7622 276922 7678 276924
rect 7702 276922 7758 276924
rect 7782 276922 7838 276924
rect 7862 276922 7918 276924
rect 7622 276870 7648 276922
rect 7648 276870 7678 276922
rect 7702 276870 7712 276922
rect 7712 276870 7758 276922
rect 7782 276870 7828 276922
rect 7828 276870 7838 276922
rect 7862 276870 7892 276922
rect 7892 276870 7918 276922
rect 7622 276868 7678 276870
rect 7702 276868 7758 276870
rect 7782 276868 7838 276870
rect 7862 276868 7918 276870
rect 7622 275834 7678 275836
rect 7702 275834 7758 275836
rect 7782 275834 7838 275836
rect 7862 275834 7918 275836
rect 7622 275782 7648 275834
rect 7648 275782 7678 275834
rect 7702 275782 7712 275834
rect 7712 275782 7758 275834
rect 7782 275782 7828 275834
rect 7828 275782 7838 275834
rect 7862 275782 7892 275834
rect 7892 275782 7918 275834
rect 7622 275780 7678 275782
rect 7702 275780 7758 275782
rect 7782 275780 7838 275782
rect 7862 275780 7918 275782
rect 7622 274746 7678 274748
rect 7702 274746 7758 274748
rect 7782 274746 7838 274748
rect 7862 274746 7918 274748
rect 7622 274694 7648 274746
rect 7648 274694 7678 274746
rect 7702 274694 7712 274746
rect 7712 274694 7758 274746
rect 7782 274694 7828 274746
rect 7828 274694 7838 274746
rect 7862 274694 7892 274746
rect 7892 274694 7918 274746
rect 7622 274692 7678 274694
rect 7702 274692 7758 274694
rect 7782 274692 7838 274694
rect 7862 274692 7918 274694
rect 7622 273658 7678 273660
rect 7702 273658 7758 273660
rect 7782 273658 7838 273660
rect 7862 273658 7918 273660
rect 7622 273606 7648 273658
rect 7648 273606 7678 273658
rect 7702 273606 7712 273658
rect 7712 273606 7758 273658
rect 7782 273606 7828 273658
rect 7828 273606 7838 273658
rect 7862 273606 7892 273658
rect 7892 273606 7918 273658
rect 7622 273604 7678 273606
rect 7702 273604 7758 273606
rect 7782 273604 7838 273606
rect 7862 273604 7918 273606
rect 7622 272570 7678 272572
rect 7702 272570 7758 272572
rect 7782 272570 7838 272572
rect 7862 272570 7918 272572
rect 7622 272518 7648 272570
rect 7648 272518 7678 272570
rect 7702 272518 7712 272570
rect 7712 272518 7758 272570
rect 7782 272518 7828 272570
rect 7828 272518 7838 272570
rect 7862 272518 7892 272570
rect 7892 272518 7918 272570
rect 7622 272516 7678 272518
rect 7702 272516 7758 272518
rect 7782 272516 7838 272518
rect 7862 272516 7918 272518
rect 7622 271482 7678 271484
rect 7702 271482 7758 271484
rect 7782 271482 7838 271484
rect 7862 271482 7918 271484
rect 7622 271430 7648 271482
rect 7648 271430 7678 271482
rect 7702 271430 7712 271482
rect 7712 271430 7758 271482
rect 7782 271430 7828 271482
rect 7828 271430 7838 271482
rect 7862 271430 7892 271482
rect 7892 271430 7918 271482
rect 7622 271428 7678 271430
rect 7702 271428 7758 271430
rect 7782 271428 7838 271430
rect 7862 271428 7918 271430
rect 7622 270394 7678 270396
rect 7702 270394 7758 270396
rect 7782 270394 7838 270396
rect 7862 270394 7918 270396
rect 7622 270342 7648 270394
rect 7648 270342 7678 270394
rect 7702 270342 7712 270394
rect 7712 270342 7758 270394
rect 7782 270342 7828 270394
rect 7828 270342 7838 270394
rect 7862 270342 7892 270394
rect 7892 270342 7918 270394
rect 7622 270340 7678 270342
rect 7702 270340 7758 270342
rect 7782 270340 7838 270342
rect 7862 270340 7918 270342
rect 7622 269306 7678 269308
rect 7702 269306 7758 269308
rect 7782 269306 7838 269308
rect 7862 269306 7918 269308
rect 7622 269254 7648 269306
rect 7648 269254 7678 269306
rect 7702 269254 7712 269306
rect 7712 269254 7758 269306
rect 7782 269254 7828 269306
rect 7828 269254 7838 269306
rect 7862 269254 7892 269306
rect 7892 269254 7918 269306
rect 7622 269252 7678 269254
rect 7702 269252 7758 269254
rect 7782 269252 7838 269254
rect 7862 269252 7918 269254
rect 7622 268218 7678 268220
rect 7702 268218 7758 268220
rect 7782 268218 7838 268220
rect 7862 268218 7918 268220
rect 7622 268166 7648 268218
rect 7648 268166 7678 268218
rect 7702 268166 7712 268218
rect 7712 268166 7758 268218
rect 7782 268166 7828 268218
rect 7828 268166 7838 268218
rect 7862 268166 7892 268218
rect 7892 268166 7918 268218
rect 7622 268164 7678 268166
rect 7702 268164 7758 268166
rect 7782 268164 7838 268166
rect 7862 268164 7918 268166
rect 7622 267130 7678 267132
rect 7702 267130 7758 267132
rect 7782 267130 7838 267132
rect 7862 267130 7918 267132
rect 7622 267078 7648 267130
rect 7648 267078 7678 267130
rect 7702 267078 7712 267130
rect 7712 267078 7758 267130
rect 7782 267078 7828 267130
rect 7828 267078 7838 267130
rect 7862 267078 7892 267130
rect 7892 267078 7918 267130
rect 7622 267076 7678 267078
rect 7702 267076 7758 267078
rect 7782 267076 7838 267078
rect 7862 267076 7918 267078
rect 7622 266042 7678 266044
rect 7702 266042 7758 266044
rect 7782 266042 7838 266044
rect 7862 266042 7918 266044
rect 7622 265990 7648 266042
rect 7648 265990 7678 266042
rect 7702 265990 7712 266042
rect 7712 265990 7758 266042
rect 7782 265990 7828 266042
rect 7828 265990 7838 266042
rect 7862 265990 7892 266042
rect 7892 265990 7918 266042
rect 7622 265988 7678 265990
rect 7702 265988 7758 265990
rect 7782 265988 7838 265990
rect 7862 265988 7918 265990
rect 7622 264954 7678 264956
rect 7702 264954 7758 264956
rect 7782 264954 7838 264956
rect 7862 264954 7918 264956
rect 7622 264902 7648 264954
rect 7648 264902 7678 264954
rect 7702 264902 7712 264954
rect 7712 264902 7758 264954
rect 7782 264902 7828 264954
rect 7828 264902 7838 264954
rect 7862 264902 7892 264954
rect 7892 264902 7918 264954
rect 7622 264900 7678 264902
rect 7702 264900 7758 264902
rect 7782 264900 7838 264902
rect 7862 264900 7918 264902
rect 7622 263866 7678 263868
rect 7702 263866 7758 263868
rect 7782 263866 7838 263868
rect 7862 263866 7918 263868
rect 7622 263814 7648 263866
rect 7648 263814 7678 263866
rect 7702 263814 7712 263866
rect 7712 263814 7758 263866
rect 7782 263814 7828 263866
rect 7828 263814 7838 263866
rect 7862 263814 7892 263866
rect 7892 263814 7918 263866
rect 7622 263812 7678 263814
rect 7702 263812 7758 263814
rect 7782 263812 7838 263814
rect 7862 263812 7918 263814
rect 7622 262778 7678 262780
rect 7702 262778 7758 262780
rect 7782 262778 7838 262780
rect 7862 262778 7918 262780
rect 7622 262726 7648 262778
rect 7648 262726 7678 262778
rect 7702 262726 7712 262778
rect 7712 262726 7758 262778
rect 7782 262726 7828 262778
rect 7828 262726 7838 262778
rect 7862 262726 7892 262778
rect 7892 262726 7918 262778
rect 7622 262724 7678 262726
rect 7702 262724 7758 262726
rect 7782 262724 7838 262726
rect 7862 262724 7918 262726
rect 7622 261690 7678 261692
rect 7702 261690 7758 261692
rect 7782 261690 7838 261692
rect 7862 261690 7918 261692
rect 7622 261638 7648 261690
rect 7648 261638 7678 261690
rect 7702 261638 7712 261690
rect 7712 261638 7758 261690
rect 7782 261638 7828 261690
rect 7828 261638 7838 261690
rect 7862 261638 7892 261690
rect 7892 261638 7918 261690
rect 7622 261636 7678 261638
rect 7702 261636 7758 261638
rect 7782 261636 7838 261638
rect 7862 261636 7918 261638
rect 7622 260602 7678 260604
rect 7702 260602 7758 260604
rect 7782 260602 7838 260604
rect 7862 260602 7918 260604
rect 7622 260550 7648 260602
rect 7648 260550 7678 260602
rect 7702 260550 7712 260602
rect 7712 260550 7758 260602
rect 7782 260550 7828 260602
rect 7828 260550 7838 260602
rect 7862 260550 7892 260602
rect 7892 260550 7918 260602
rect 7622 260548 7678 260550
rect 7702 260548 7758 260550
rect 7782 260548 7838 260550
rect 7862 260548 7918 260550
rect 7622 259514 7678 259516
rect 7702 259514 7758 259516
rect 7782 259514 7838 259516
rect 7862 259514 7918 259516
rect 7622 259462 7648 259514
rect 7648 259462 7678 259514
rect 7702 259462 7712 259514
rect 7712 259462 7758 259514
rect 7782 259462 7828 259514
rect 7828 259462 7838 259514
rect 7862 259462 7892 259514
rect 7892 259462 7918 259514
rect 7622 259460 7678 259462
rect 7702 259460 7758 259462
rect 7782 259460 7838 259462
rect 7862 259460 7918 259462
rect 7622 258426 7678 258428
rect 7702 258426 7758 258428
rect 7782 258426 7838 258428
rect 7862 258426 7918 258428
rect 7622 258374 7648 258426
rect 7648 258374 7678 258426
rect 7702 258374 7712 258426
rect 7712 258374 7758 258426
rect 7782 258374 7828 258426
rect 7828 258374 7838 258426
rect 7862 258374 7892 258426
rect 7892 258374 7918 258426
rect 7622 258372 7678 258374
rect 7702 258372 7758 258374
rect 7782 258372 7838 258374
rect 7862 258372 7918 258374
rect 7622 257338 7678 257340
rect 7702 257338 7758 257340
rect 7782 257338 7838 257340
rect 7862 257338 7918 257340
rect 7622 257286 7648 257338
rect 7648 257286 7678 257338
rect 7702 257286 7712 257338
rect 7712 257286 7758 257338
rect 7782 257286 7828 257338
rect 7828 257286 7838 257338
rect 7862 257286 7892 257338
rect 7892 257286 7918 257338
rect 7622 257284 7678 257286
rect 7702 257284 7758 257286
rect 7782 257284 7838 257286
rect 7862 257284 7918 257286
rect 7622 256250 7678 256252
rect 7702 256250 7758 256252
rect 7782 256250 7838 256252
rect 7862 256250 7918 256252
rect 7622 256198 7648 256250
rect 7648 256198 7678 256250
rect 7702 256198 7712 256250
rect 7712 256198 7758 256250
rect 7782 256198 7828 256250
rect 7828 256198 7838 256250
rect 7862 256198 7892 256250
rect 7892 256198 7918 256250
rect 7622 256196 7678 256198
rect 7702 256196 7758 256198
rect 7782 256196 7838 256198
rect 7862 256196 7918 256198
rect 7622 255162 7678 255164
rect 7702 255162 7758 255164
rect 7782 255162 7838 255164
rect 7862 255162 7918 255164
rect 7622 255110 7648 255162
rect 7648 255110 7678 255162
rect 7702 255110 7712 255162
rect 7712 255110 7758 255162
rect 7782 255110 7828 255162
rect 7828 255110 7838 255162
rect 7862 255110 7892 255162
rect 7892 255110 7918 255162
rect 7622 255108 7678 255110
rect 7702 255108 7758 255110
rect 7782 255108 7838 255110
rect 7862 255108 7918 255110
rect 7622 254074 7678 254076
rect 7702 254074 7758 254076
rect 7782 254074 7838 254076
rect 7862 254074 7918 254076
rect 7622 254022 7648 254074
rect 7648 254022 7678 254074
rect 7702 254022 7712 254074
rect 7712 254022 7758 254074
rect 7782 254022 7828 254074
rect 7828 254022 7838 254074
rect 7862 254022 7892 254074
rect 7892 254022 7918 254074
rect 7622 254020 7678 254022
rect 7702 254020 7758 254022
rect 7782 254020 7838 254022
rect 7862 254020 7918 254022
rect 7622 252986 7678 252988
rect 7702 252986 7758 252988
rect 7782 252986 7838 252988
rect 7862 252986 7918 252988
rect 7622 252934 7648 252986
rect 7648 252934 7678 252986
rect 7702 252934 7712 252986
rect 7712 252934 7758 252986
rect 7782 252934 7828 252986
rect 7828 252934 7838 252986
rect 7862 252934 7892 252986
rect 7892 252934 7918 252986
rect 7622 252932 7678 252934
rect 7702 252932 7758 252934
rect 7782 252932 7838 252934
rect 7862 252932 7918 252934
rect 7622 251898 7678 251900
rect 7702 251898 7758 251900
rect 7782 251898 7838 251900
rect 7862 251898 7918 251900
rect 7622 251846 7648 251898
rect 7648 251846 7678 251898
rect 7702 251846 7712 251898
rect 7712 251846 7758 251898
rect 7782 251846 7828 251898
rect 7828 251846 7838 251898
rect 7862 251846 7892 251898
rect 7892 251846 7918 251898
rect 7622 251844 7678 251846
rect 7702 251844 7758 251846
rect 7782 251844 7838 251846
rect 7862 251844 7918 251846
rect 7622 250810 7678 250812
rect 7702 250810 7758 250812
rect 7782 250810 7838 250812
rect 7862 250810 7918 250812
rect 7622 250758 7648 250810
rect 7648 250758 7678 250810
rect 7702 250758 7712 250810
rect 7712 250758 7758 250810
rect 7782 250758 7828 250810
rect 7828 250758 7838 250810
rect 7862 250758 7892 250810
rect 7892 250758 7918 250810
rect 7622 250756 7678 250758
rect 7702 250756 7758 250758
rect 7782 250756 7838 250758
rect 7862 250756 7918 250758
rect 7622 249722 7678 249724
rect 7702 249722 7758 249724
rect 7782 249722 7838 249724
rect 7862 249722 7918 249724
rect 7622 249670 7648 249722
rect 7648 249670 7678 249722
rect 7702 249670 7712 249722
rect 7712 249670 7758 249722
rect 7782 249670 7828 249722
rect 7828 249670 7838 249722
rect 7862 249670 7892 249722
rect 7892 249670 7918 249722
rect 7622 249668 7678 249670
rect 7702 249668 7758 249670
rect 7782 249668 7838 249670
rect 7862 249668 7918 249670
rect 7622 248634 7678 248636
rect 7702 248634 7758 248636
rect 7782 248634 7838 248636
rect 7862 248634 7918 248636
rect 7622 248582 7648 248634
rect 7648 248582 7678 248634
rect 7702 248582 7712 248634
rect 7712 248582 7758 248634
rect 7782 248582 7828 248634
rect 7828 248582 7838 248634
rect 7862 248582 7892 248634
rect 7892 248582 7918 248634
rect 7622 248580 7678 248582
rect 7702 248580 7758 248582
rect 7782 248580 7838 248582
rect 7862 248580 7918 248582
rect 7622 247546 7678 247548
rect 7702 247546 7758 247548
rect 7782 247546 7838 247548
rect 7862 247546 7918 247548
rect 7622 247494 7648 247546
rect 7648 247494 7678 247546
rect 7702 247494 7712 247546
rect 7712 247494 7758 247546
rect 7782 247494 7828 247546
rect 7828 247494 7838 247546
rect 7862 247494 7892 247546
rect 7892 247494 7918 247546
rect 7622 247492 7678 247494
rect 7702 247492 7758 247494
rect 7782 247492 7838 247494
rect 7862 247492 7918 247494
rect 7622 246458 7678 246460
rect 7702 246458 7758 246460
rect 7782 246458 7838 246460
rect 7862 246458 7918 246460
rect 7622 246406 7648 246458
rect 7648 246406 7678 246458
rect 7702 246406 7712 246458
rect 7712 246406 7758 246458
rect 7782 246406 7828 246458
rect 7828 246406 7838 246458
rect 7862 246406 7892 246458
rect 7892 246406 7918 246458
rect 7622 246404 7678 246406
rect 7702 246404 7758 246406
rect 7782 246404 7838 246406
rect 7862 246404 7918 246406
rect 7622 245370 7678 245372
rect 7702 245370 7758 245372
rect 7782 245370 7838 245372
rect 7862 245370 7918 245372
rect 7622 245318 7648 245370
rect 7648 245318 7678 245370
rect 7702 245318 7712 245370
rect 7712 245318 7758 245370
rect 7782 245318 7828 245370
rect 7828 245318 7838 245370
rect 7862 245318 7892 245370
rect 7892 245318 7918 245370
rect 7622 245316 7678 245318
rect 7702 245316 7758 245318
rect 7782 245316 7838 245318
rect 7862 245316 7918 245318
rect 7622 244282 7678 244284
rect 7702 244282 7758 244284
rect 7782 244282 7838 244284
rect 7862 244282 7918 244284
rect 7622 244230 7648 244282
rect 7648 244230 7678 244282
rect 7702 244230 7712 244282
rect 7712 244230 7758 244282
rect 7782 244230 7828 244282
rect 7828 244230 7838 244282
rect 7862 244230 7892 244282
rect 7892 244230 7918 244282
rect 7622 244228 7678 244230
rect 7702 244228 7758 244230
rect 7782 244228 7838 244230
rect 7862 244228 7918 244230
rect 7622 243194 7678 243196
rect 7702 243194 7758 243196
rect 7782 243194 7838 243196
rect 7862 243194 7918 243196
rect 7622 243142 7648 243194
rect 7648 243142 7678 243194
rect 7702 243142 7712 243194
rect 7712 243142 7758 243194
rect 7782 243142 7828 243194
rect 7828 243142 7838 243194
rect 7862 243142 7892 243194
rect 7892 243142 7918 243194
rect 7622 243140 7678 243142
rect 7702 243140 7758 243142
rect 7782 243140 7838 243142
rect 7862 243140 7918 243142
rect 7622 242106 7678 242108
rect 7702 242106 7758 242108
rect 7782 242106 7838 242108
rect 7862 242106 7918 242108
rect 7622 242054 7648 242106
rect 7648 242054 7678 242106
rect 7702 242054 7712 242106
rect 7712 242054 7758 242106
rect 7782 242054 7828 242106
rect 7828 242054 7838 242106
rect 7862 242054 7892 242106
rect 7892 242054 7918 242106
rect 7622 242052 7678 242054
rect 7702 242052 7758 242054
rect 7782 242052 7838 242054
rect 7862 242052 7918 242054
rect 7622 241018 7678 241020
rect 7702 241018 7758 241020
rect 7782 241018 7838 241020
rect 7862 241018 7918 241020
rect 7622 240966 7648 241018
rect 7648 240966 7678 241018
rect 7702 240966 7712 241018
rect 7712 240966 7758 241018
rect 7782 240966 7828 241018
rect 7828 240966 7838 241018
rect 7862 240966 7892 241018
rect 7892 240966 7918 241018
rect 7622 240964 7678 240966
rect 7702 240964 7758 240966
rect 7782 240964 7838 240966
rect 7862 240964 7918 240966
rect 7622 239930 7678 239932
rect 7702 239930 7758 239932
rect 7782 239930 7838 239932
rect 7862 239930 7918 239932
rect 7622 239878 7648 239930
rect 7648 239878 7678 239930
rect 7702 239878 7712 239930
rect 7712 239878 7758 239930
rect 7782 239878 7828 239930
rect 7828 239878 7838 239930
rect 7862 239878 7892 239930
rect 7892 239878 7918 239930
rect 7622 239876 7678 239878
rect 7702 239876 7758 239878
rect 7782 239876 7838 239878
rect 7862 239876 7918 239878
rect 7622 238842 7678 238844
rect 7702 238842 7758 238844
rect 7782 238842 7838 238844
rect 7862 238842 7918 238844
rect 7622 238790 7648 238842
rect 7648 238790 7678 238842
rect 7702 238790 7712 238842
rect 7712 238790 7758 238842
rect 7782 238790 7828 238842
rect 7828 238790 7838 238842
rect 7862 238790 7892 238842
rect 7892 238790 7918 238842
rect 7622 238788 7678 238790
rect 7702 238788 7758 238790
rect 7782 238788 7838 238790
rect 7862 238788 7918 238790
rect 7622 237754 7678 237756
rect 7702 237754 7758 237756
rect 7782 237754 7838 237756
rect 7862 237754 7918 237756
rect 7622 237702 7648 237754
rect 7648 237702 7678 237754
rect 7702 237702 7712 237754
rect 7712 237702 7758 237754
rect 7782 237702 7828 237754
rect 7828 237702 7838 237754
rect 7862 237702 7892 237754
rect 7892 237702 7918 237754
rect 7622 237700 7678 237702
rect 7702 237700 7758 237702
rect 7782 237700 7838 237702
rect 7862 237700 7918 237702
rect 7622 236666 7678 236668
rect 7702 236666 7758 236668
rect 7782 236666 7838 236668
rect 7862 236666 7918 236668
rect 7622 236614 7648 236666
rect 7648 236614 7678 236666
rect 7702 236614 7712 236666
rect 7712 236614 7758 236666
rect 7782 236614 7828 236666
rect 7828 236614 7838 236666
rect 7862 236614 7892 236666
rect 7892 236614 7918 236666
rect 7622 236612 7678 236614
rect 7702 236612 7758 236614
rect 7782 236612 7838 236614
rect 7862 236612 7918 236614
rect 7622 235578 7678 235580
rect 7702 235578 7758 235580
rect 7782 235578 7838 235580
rect 7862 235578 7918 235580
rect 7622 235526 7648 235578
rect 7648 235526 7678 235578
rect 7702 235526 7712 235578
rect 7712 235526 7758 235578
rect 7782 235526 7828 235578
rect 7828 235526 7838 235578
rect 7862 235526 7892 235578
rect 7892 235526 7918 235578
rect 7622 235524 7678 235526
rect 7702 235524 7758 235526
rect 7782 235524 7838 235526
rect 7862 235524 7918 235526
rect 7622 234490 7678 234492
rect 7702 234490 7758 234492
rect 7782 234490 7838 234492
rect 7862 234490 7918 234492
rect 7622 234438 7648 234490
rect 7648 234438 7678 234490
rect 7702 234438 7712 234490
rect 7712 234438 7758 234490
rect 7782 234438 7828 234490
rect 7828 234438 7838 234490
rect 7862 234438 7892 234490
rect 7892 234438 7918 234490
rect 7622 234436 7678 234438
rect 7702 234436 7758 234438
rect 7782 234436 7838 234438
rect 7862 234436 7918 234438
rect 7622 233402 7678 233404
rect 7702 233402 7758 233404
rect 7782 233402 7838 233404
rect 7862 233402 7918 233404
rect 7622 233350 7648 233402
rect 7648 233350 7678 233402
rect 7702 233350 7712 233402
rect 7712 233350 7758 233402
rect 7782 233350 7828 233402
rect 7828 233350 7838 233402
rect 7862 233350 7892 233402
rect 7892 233350 7918 233402
rect 7622 233348 7678 233350
rect 7702 233348 7758 233350
rect 7782 233348 7838 233350
rect 7862 233348 7918 233350
rect 7622 232314 7678 232316
rect 7702 232314 7758 232316
rect 7782 232314 7838 232316
rect 7862 232314 7918 232316
rect 7622 232262 7648 232314
rect 7648 232262 7678 232314
rect 7702 232262 7712 232314
rect 7712 232262 7758 232314
rect 7782 232262 7828 232314
rect 7828 232262 7838 232314
rect 7862 232262 7892 232314
rect 7892 232262 7918 232314
rect 7622 232260 7678 232262
rect 7702 232260 7758 232262
rect 7782 232260 7838 232262
rect 7862 232260 7918 232262
rect 7622 231226 7678 231228
rect 7702 231226 7758 231228
rect 7782 231226 7838 231228
rect 7862 231226 7918 231228
rect 7622 231174 7648 231226
rect 7648 231174 7678 231226
rect 7702 231174 7712 231226
rect 7712 231174 7758 231226
rect 7782 231174 7828 231226
rect 7828 231174 7838 231226
rect 7862 231174 7892 231226
rect 7892 231174 7918 231226
rect 7622 231172 7678 231174
rect 7702 231172 7758 231174
rect 7782 231172 7838 231174
rect 7862 231172 7918 231174
rect 7622 230138 7678 230140
rect 7702 230138 7758 230140
rect 7782 230138 7838 230140
rect 7862 230138 7918 230140
rect 7622 230086 7648 230138
rect 7648 230086 7678 230138
rect 7702 230086 7712 230138
rect 7712 230086 7758 230138
rect 7782 230086 7828 230138
rect 7828 230086 7838 230138
rect 7862 230086 7892 230138
rect 7892 230086 7918 230138
rect 7622 230084 7678 230086
rect 7702 230084 7758 230086
rect 7782 230084 7838 230086
rect 7862 230084 7918 230086
rect 7622 229050 7678 229052
rect 7702 229050 7758 229052
rect 7782 229050 7838 229052
rect 7862 229050 7918 229052
rect 7622 228998 7648 229050
rect 7648 228998 7678 229050
rect 7702 228998 7712 229050
rect 7712 228998 7758 229050
rect 7782 228998 7828 229050
rect 7828 228998 7838 229050
rect 7862 228998 7892 229050
rect 7892 228998 7918 229050
rect 7622 228996 7678 228998
rect 7702 228996 7758 228998
rect 7782 228996 7838 228998
rect 7862 228996 7918 228998
rect 7622 227962 7678 227964
rect 7702 227962 7758 227964
rect 7782 227962 7838 227964
rect 7862 227962 7918 227964
rect 7622 227910 7648 227962
rect 7648 227910 7678 227962
rect 7702 227910 7712 227962
rect 7712 227910 7758 227962
rect 7782 227910 7828 227962
rect 7828 227910 7838 227962
rect 7862 227910 7892 227962
rect 7892 227910 7918 227962
rect 7622 227908 7678 227910
rect 7702 227908 7758 227910
rect 7782 227908 7838 227910
rect 7862 227908 7918 227910
rect 7622 226874 7678 226876
rect 7702 226874 7758 226876
rect 7782 226874 7838 226876
rect 7862 226874 7918 226876
rect 7622 226822 7648 226874
rect 7648 226822 7678 226874
rect 7702 226822 7712 226874
rect 7712 226822 7758 226874
rect 7782 226822 7828 226874
rect 7828 226822 7838 226874
rect 7862 226822 7892 226874
rect 7892 226822 7918 226874
rect 7622 226820 7678 226822
rect 7702 226820 7758 226822
rect 7782 226820 7838 226822
rect 7862 226820 7918 226822
rect 7622 225786 7678 225788
rect 7702 225786 7758 225788
rect 7782 225786 7838 225788
rect 7862 225786 7918 225788
rect 7622 225734 7648 225786
rect 7648 225734 7678 225786
rect 7702 225734 7712 225786
rect 7712 225734 7758 225786
rect 7782 225734 7828 225786
rect 7828 225734 7838 225786
rect 7862 225734 7892 225786
rect 7892 225734 7918 225786
rect 7622 225732 7678 225734
rect 7702 225732 7758 225734
rect 7782 225732 7838 225734
rect 7862 225732 7918 225734
rect 7622 224698 7678 224700
rect 7702 224698 7758 224700
rect 7782 224698 7838 224700
rect 7862 224698 7918 224700
rect 7622 224646 7648 224698
rect 7648 224646 7678 224698
rect 7702 224646 7712 224698
rect 7712 224646 7758 224698
rect 7782 224646 7828 224698
rect 7828 224646 7838 224698
rect 7862 224646 7892 224698
rect 7892 224646 7918 224698
rect 7622 224644 7678 224646
rect 7702 224644 7758 224646
rect 7782 224644 7838 224646
rect 7862 224644 7918 224646
rect 7622 223610 7678 223612
rect 7702 223610 7758 223612
rect 7782 223610 7838 223612
rect 7862 223610 7918 223612
rect 7622 223558 7648 223610
rect 7648 223558 7678 223610
rect 7702 223558 7712 223610
rect 7712 223558 7758 223610
rect 7782 223558 7828 223610
rect 7828 223558 7838 223610
rect 7862 223558 7892 223610
rect 7892 223558 7918 223610
rect 7622 223556 7678 223558
rect 7702 223556 7758 223558
rect 7782 223556 7838 223558
rect 7862 223556 7918 223558
rect 7622 222522 7678 222524
rect 7702 222522 7758 222524
rect 7782 222522 7838 222524
rect 7862 222522 7918 222524
rect 7622 222470 7648 222522
rect 7648 222470 7678 222522
rect 7702 222470 7712 222522
rect 7712 222470 7758 222522
rect 7782 222470 7828 222522
rect 7828 222470 7838 222522
rect 7862 222470 7892 222522
rect 7892 222470 7918 222522
rect 7622 222468 7678 222470
rect 7702 222468 7758 222470
rect 7782 222468 7838 222470
rect 7862 222468 7918 222470
rect 7622 221434 7678 221436
rect 7702 221434 7758 221436
rect 7782 221434 7838 221436
rect 7862 221434 7918 221436
rect 7622 221382 7648 221434
rect 7648 221382 7678 221434
rect 7702 221382 7712 221434
rect 7712 221382 7758 221434
rect 7782 221382 7828 221434
rect 7828 221382 7838 221434
rect 7862 221382 7892 221434
rect 7892 221382 7918 221434
rect 7622 221380 7678 221382
rect 7702 221380 7758 221382
rect 7782 221380 7838 221382
rect 7862 221380 7918 221382
rect 7622 220346 7678 220348
rect 7702 220346 7758 220348
rect 7782 220346 7838 220348
rect 7862 220346 7918 220348
rect 7622 220294 7648 220346
rect 7648 220294 7678 220346
rect 7702 220294 7712 220346
rect 7712 220294 7758 220346
rect 7782 220294 7828 220346
rect 7828 220294 7838 220346
rect 7862 220294 7892 220346
rect 7892 220294 7918 220346
rect 7622 220292 7678 220294
rect 7702 220292 7758 220294
rect 7782 220292 7838 220294
rect 7862 220292 7918 220294
rect 7622 219258 7678 219260
rect 7702 219258 7758 219260
rect 7782 219258 7838 219260
rect 7862 219258 7918 219260
rect 7622 219206 7648 219258
rect 7648 219206 7678 219258
rect 7702 219206 7712 219258
rect 7712 219206 7758 219258
rect 7782 219206 7828 219258
rect 7828 219206 7838 219258
rect 7862 219206 7892 219258
rect 7892 219206 7918 219258
rect 7622 219204 7678 219206
rect 7702 219204 7758 219206
rect 7782 219204 7838 219206
rect 7862 219204 7918 219206
rect 7622 218170 7678 218172
rect 7702 218170 7758 218172
rect 7782 218170 7838 218172
rect 7862 218170 7918 218172
rect 7622 218118 7648 218170
rect 7648 218118 7678 218170
rect 7702 218118 7712 218170
rect 7712 218118 7758 218170
rect 7782 218118 7828 218170
rect 7828 218118 7838 218170
rect 7862 218118 7892 218170
rect 7892 218118 7918 218170
rect 7622 218116 7678 218118
rect 7702 218116 7758 218118
rect 7782 218116 7838 218118
rect 7862 218116 7918 218118
rect 7622 217082 7678 217084
rect 7702 217082 7758 217084
rect 7782 217082 7838 217084
rect 7862 217082 7918 217084
rect 7622 217030 7648 217082
rect 7648 217030 7678 217082
rect 7702 217030 7712 217082
rect 7712 217030 7758 217082
rect 7782 217030 7828 217082
rect 7828 217030 7838 217082
rect 7862 217030 7892 217082
rect 7892 217030 7918 217082
rect 7622 217028 7678 217030
rect 7702 217028 7758 217030
rect 7782 217028 7838 217030
rect 7862 217028 7918 217030
rect 7622 215994 7678 215996
rect 7702 215994 7758 215996
rect 7782 215994 7838 215996
rect 7862 215994 7918 215996
rect 7622 215942 7648 215994
rect 7648 215942 7678 215994
rect 7702 215942 7712 215994
rect 7712 215942 7758 215994
rect 7782 215942 7828 215994
rect 7828 215942 7838 215994
rect 7862 215942 7892 215994
rect 7892 215942 7918 215994
rect 7622 215940 7678 215942
rect 7702 215940 7758 215942
rect 7782 215940 7838 215942
rect 7862 215940 7918 215942
rect 7622 214906 7678 214908
rect 7702 214906 7758 214908
rect 7782 214906 7838 214908
rect 7862 214906 7918 214908
rect 7622 214854 7648 214906
rect 7648 214854 7678 214906
rect 7702 214854 7712 214906
rect 7712 214854 7758 214906
rect 7782 214854 7828 214906
rect 7828 214854 7838 214906
rect 7862 214854 7892 214906
rect 7892 214854 7918 214906
rect 7622 214852 7678 214854
rect 7702 214852 7758 214854
rect 7782 214852 7838 214854
rect 7862 214852 7918 214854
rect 7622 213818 7678 213820
rect 7702 213818 7758 213820
rect 7782 213818 7838 213820
rect 7862 213818 7918 213820
rect 7622 213766 7648 213818
rect 7648 213766 7678 213818
rect 7702 213766 7712 213818
rect 7712 213766 7758 213818
rect 7782 213766 7828 213818
rect 7828 213766 7838 213818
rect 7862 213766 7892 213818
rect 7892 213766 7918 213818
rect 7622 213764 7678 213766
rect 7702 213764 7758 213766
rect 7782 213764 7838 213766
rect 7862 213764 7918 213766
rect 7622 212730 7678 212732
rect 7702 212730 7758 212732
rect 7782 212730 7838 212732
rect 7862 212730 7918 212732
rect 7622 212678 7648 212730
rect 7648 212678 7678 212730
rect 7702 212678 7712 212730
rect 7712 212678 7758 212730
rect 7782 212678 7828 212730
rect 7828 212678 7838 212730
rect 7862 212678 7892 212730
rect 7892 212678 7918 212730
rect 7622 212676 7678 212678
rect 7702 212676 7758 212678
rect 7782 212676 7838 212678
rect 7862 212676 7918 212678
rect 7622 211642 7678 211644
rect 7702 211642 7758 211644
rect 7782 211642 7838 211644
rect 7862 211642 7918 211644
rect 7622 211590 7648 211642
rect 7648 211590 7678 211642
rect 7702 211590 7712 211642
rect 7712 211590 7758 211642
rect 7782 211590 7828 211642
rect 7828 211590 7838 211642
rect 7862 211590 7892 211642
rect 7892 211590 7918 211642
rect 7622 211588 7678 211590
rect 7702 211588 7758 211590
rect 7782 211588 7838 211590
rect 7862 211588 7918 211590
rect 7622 210554 7678 210556
rect 7702 210554 7758 210556
rect 7782 210554 7838 210556
rect 7862 210554 7918 210556
rect 7622 210502 7648 210554
rect 7648 210502 7678 210554
rect 7702 210502 7712 210554
rect 7712 210502 7758 210554
rect 7782 210502 7828 210554
rect 7828 210502 7838 210554
rect 7862 210502 7892 210554
rect 7892 210502 7918 210554
rect 7622 210500 7678 210502
rect 7702 210500 7758 210502
rect 7782 210500 7838 210502
rect 7862 210500 7918 210502
rect 7622 209466 7678 209468
rect 7702 209466 7758 209468
rect 7782 209466 7838 209468
rect 7862 209466 7918 209468
rect 7622 209414 7648 209466
rect 7648 209414 7678 209466
rect 7702 209414 7712 209466
rect 7712 209414 7758 209466
rect 7782 209414 7828 209466
rect 7828 209414 7838 209466
rect 7862 209414 7892 209466
rect 7892 209414 7918 209466
rect 7622 209412 7678 209414
rect 7702 209412 7758 209414
rect 7782 209412 7838 209414
rect 7862 209412 7918 209414
rect 7622 208378 7678 208380
rect 7702 208378 7758 208380
rect 7782 208378 7838 208380
rect 7862 208378 7918 208380
rect 7622 208326 7648 208378
rect 7648 208326 7678 208378
rect 7702 208326 7712 208378
rect 7712 208326 7758 208378
rect 7782 208326 7828 208378
rect 7828 208326 7838 208378
rect 7862 208326 7892 208378
rect 7892 208326 7918 208378
rect 7622 208324 7678 208326
rect 7702 208324 7758 208326
rect 7782 208324 7838 208326
rect 7862 208324 7918 208326
rect 7622 207290 7678 207292
rect 7702 207290 7758 207292
rect 7782 207290 7838 207292
rect 7862 207290 7918 207292
rect 7622 207238 7648 207290
rect 7648 207238 7678 207290
rect 7702 207238 7712 207290
rect 7712 207238 7758 207290
rect 7782 207238 7828 207290
rect 7828 207238 7838 207290
rect 7862 207238 7892 207290
rect 7892 207238 7918 207290
rect 7622 207236 7678 207238
rect 7702 207236 7758 207238
rect 7782 207236 7838 207238
rect 7862 207236 7918 207238
rect 7622 206202 7678 206204
rect 7702 206202 7758 206204
rect 7782 206202 7838 206204
rect 7862 206202 7918 206204
rect 7622 206150 7648 206202
rect 7648 206150 7678 206202
rect 7702 206150 7712 206202
rect 7712 206150 7758 206202
rect 7782 206150 7828 206202
rect 7828 206150 7838 206202
rect 7862 206150 7892 206202
rect 7892 206150 7918 206202
rect 7622 206148 7678 206150
rect 7702 206148 7758 206150
rect 7782 206148 7838 206150
rect 7862 206148 7918 206150
rect 7622 205114 7678 205116
rect 7702 205114 7758 205116
rect 7782 205114 7838 205116
rect 7862 205114 7918 205116
rect 7622 205062 7648 205114
rect 7648 205062 7678 205114
rect 7702 205062 7712 205114
rect 7712 205062 7758 205114
rect 7782 205062 7828 205114
rect 7828 205062 7838 205114
rect 7862 205062 7892 205114
rect 7892 205062 7918 205114
rect 7622 205060 7678 205062
rect 7702 205060 7758 205062
rect 7782 205060 7838 205062
rect 7862 205060 7918 205062
rect 7622 204026 7678 204028
rect 7702 204026 7758 204028
rect 7782 204026 7838 204028
rect 7862 204026 7918 204028
rect 7622 203974 7648 204026
rect 7648 203974 7678 204026
rect 7702 203974 7712 204026
rect 7712 203974 7758 204026
rect 7782 203974 7828 204026
rect 7828 203974 7838 204026
rect 7862 203974 7892 204026
rect 7892 203974 7918 204026
rect 7622 203972 7678 203974
rect 7702 203972 7758 203974
rect 7782 203972 7838 203974
rect 7862 203972 7918 203974
rect 7622 202938 7678 202940
rect 7702 202938 7758 202940
rect 7782 202938 7838 202940
rect 7862 202938 7918 202940
rect 7622 202886 7648 202938
rect 7648 202886 7678 202938
rect 7702 202886 7712 202938
rect 7712 202886 7758 202938
rect 7782 202886 7828 202938
rect 7828 202886 7838 202938
rect 7862 202886 7892 202938
rect 7892 202886 7918 202938
rect 7622 202884 7678 202886
rect 7702 202884 7758 202886
rect 7782 202884 7838 202886
rect 7862 202884 7918 202886
rect 7622 201850 7678 201852
rect 7702 201850 7758 201852
rect 7782 201850 7838 201852
rect 7862 201850 7918 201852
rect 7622 201798 7648 201850
rect 7648 201798 7678 201850
rect 7702 201798 7712 201850
rect 7712 201798 7758 201850
rect 7782 201798 7828 201850
rect 7828 201798 7838 201850
rect 7862 201798 7892 201850
rect 7892 201798 7918 201850
rect 7622 201796 7678 201798
rect 7702 201796 7758 201798
rect 7782 201796 7838 201798
rect 7862 201796 7918 201798
rect 7622 200762 7678 200764
rect 7702 200762 7758 200764
rect 7782 200762 7838 200764
rect 7862 200762 7918 200764
rect 7622 200710 7648 200762
rect 7648 200710 7678 200762
rect 7702 200710 7712 200762
rect 7712 200710 7758 200762
rect 7782 200710 7828 200762
rect 7828 200710 7838 200762
rect 7862 200710 7892 200762
rect 7892 200710 7918 200762
rect 7622 200708 7678 200710
rect 7702 200708 7758 200710
rect 7782 200708 7838 200710
rect 7862 200708 7918 200710
rect 7622 199674 7678 199676
rect 7702 199674 7758 199676
rect 7782 199674 7838 199676
rect 7862 199674 7918 199676
rect 7622 199622 7648 199674
rect 7648 199622 7678 199674
rect 7702 199622 7712 199674
rect 7712 199622 7758 199674
rect 7782 199622 7828 199674
rect 7828 199622 7838 199674
rect 7862 199622 7892 199674
rect 7892 199622 7918 199674
rect 7622 199620 7678 199622
rect 7702 199620 7758 199622
rect 7782 199620 7838 199622
rect 7862 199620 7918 199622
rect 7622 198586 7678 198588
rect 7702 198586 7758 198588
rect 7782 198586 7838 198588
rect 7862 198586 7918 198588
rect 7622 198534 7648 198586
rect 7648 198534 7678 198586
rect 7702 198534 7712 198586
rect 7712 198534 7758 198586
rect 7782 198534 7828 198586
rect 7828 198534 7838 198586
rect 7862 198534 7892 198586
rect 7892 198534 7918 198586
rect 7622 198532 7678 198534
rect 7702 198532 7758 198534
rect 7782 198532 7838 198534
rect 7862 198532 7918 198534
rect 7622 197498 7678 197500
rect 7702 197498 7758 197500
rect 7782 197498 7838 197500
rect 7862 197498 7918 197500
rect 7622 197446 7648 197498
rect 7648 197446 7678 197498
rect 7702 197446 7712 197498
rect 7712 197446 7758 197498
rect 7782 197446 7828 197498
rect 7828 197446 7838 197498
rect 7862 197446 7892 197498
rect 7892 197446 7918 197498
rect 7622 197444 7678 197446
rect 7702 197444 7758 197446
rect 7782 197444 7838 197446
rect 7862 197444 7918 197446
rect 7622 196410 7678 196412
rect 7702 196410 7758 196412
rect 7782 196410 7838 196412
rect 7862 196410 7918 196412
rect 7622 196358 7648 196410
rect 7648 196358 7678 196410
rect 7702 196358 7712 196410
rect 7712 196358 7758 196410
rect 7782 196358 7828 196410
rect 7828 196358 7838 196410
rect 7862 196358 7892 196410
rect 7892 196358 7918 196410
rect 7622 196356 7678 196358
rect 7702 196356 7758 196358
rect 7782 196356 7838 196358
rect 7862 196356 7918 196358
rect 7622 195322 7678 195324
rect 7702 195322 7758 195324
rect 7782 195322 7838 195324
rect 7862 195322 7918 195324
rect 7622 195270 7648 195322
rect 7648 195270 7678 195322
rect 7702 195270 7712 195322
rect 7712 195270 7758 195322
rect 7782 195270 7828 195322
rect 7828 195270 7838 195322
rect 7862 195270 7892 195322
rect 7892 195270 7918 195322
rect 7622 195268 7678 195270
rect 7702 195268 7758 195270
rect 7782 195268 7838 195270
rect 7862 195268 7918 195270
rect 7622 194234 7678 194236
rect 7702 194234 7758 194236
rect 7782 194234 7838 194236
rect 7862 194234 7918 194236
rect 7622 194182 7648 194234
rect 7648 194182 7678 194234
rect 7702 194182 7712 194234
rect 7712 194182 7758 194234
rect 7782 194182 7828 194234
rect 7828 194182 7838 194234
rect 7862 194182 7892 194234
rect 7892 194182 7918 194234
rect 7622 194180 7678 194182
rect 7702 194180 7758 194182
rect 7782 194180 7838 194182
rect 7862 194180 7918 194182
rect 7622 193146 7678 193148
rect 7702 193146 7758 193148
rect 7782 193146 7838 193148
rect 7862 193146 7918 193148
rect 7622 193094 7648 193146
rect 7648 193094 7678 193146
rect 7702 193094 7712 193146
rect 7712 193094 7758 193146
rect 7782 193094 7828 193146
rect 7828 193094 7838 193146
rect 7862 193094 7892 193146
rect 7892 193094 7918 193146
rect 7622 193092 7678 193094
rect 7702 193092 7758 193094
rect 7782 193092 7838 193094
rect 7862 193092 7918 193094
rect 7622 192058 7678 192060
rect 7702 192058 7758 192060
rect 7782 192058 7838 192060
rect 7862 192058 7918 192060
rect 7622 192006 7648 192058
rect 7648 192006 7678 192058
rect 7702 192006 7712 192058
rect 7712 192006 7758 192058
rect 7782 192006 7828 192058
rect 7828 192006 7838 192058
rect 7862 192006 7892 192058
rect 7892 192006 7918 192058
rect 7622 192004 7678 192006
rect 7702 192004 7758 192006
rect 7782 192004 7838 192006
rect 7862 192004 7918 192006
rect 7622 190970 7678 190972
rect 7702 190970 7758 190972
rect 7782 190970 7838 190972
rect 7862 190970 7918 190972
rect 7622 190918 7648 190970
rect 7648 190918 7678 190970
rect 7702 190918 7712 190970
rect 7712 190918 7758 190970
rect 7782 190918 7828 190970
rect 7828 190918 7838 190970
rect 7862 190918 7892 190970
rect 7892 190918 7918 190970
rect 7622 190916 7678 190918
rect 7702 190916 7758 190918
rect 7782 190916 7838 190918
rect 7862 190916 7918 190918
rect 7622 189882 7678 189884
rect 7702 189882 7758 189884
rect 7782 189882 7838 189884
rect 7862 189882 7918 189884
rect 7622 189830 7648 189882
rect 7648 189830 7678 189882
rect 7702 189830 7712 189882
rect 7712 189830 7758 189882
rect 7782 189830 7828 189882
rect 7828 189830 7838 189882
rect 7862 189830 7892 189882
rect 7892 189830 7918 189882
rect 7622 189828 7678 189830
rect 7702 189828 7758 189830
rect 7782 189828 7838 189830
rect 7862 189828 7918 189830
rect 7622 188794 7678 188796
rect 7702 188794 7758 188796
rect 7782 188794 7838 188796
rect 7862 188794 7918 188796
rect 7622 188742 7648 188794
rect 7648 188742 7678 188794
rect 7702 188742 7712 188794
rect 7712 188742 7758 188794
rect 7782 188742 7828 188794
rect 7828 188742 7838 188794
rect 7862 188742 7892 188794
rect 7892 188742 7918 188794
rect 7622 188740 7678 188742
rect 7702 188740 7758 188742
rect 7782 188740 7838 188742
rect 7862 188740 7918 188742
rect 7622 187706 7678 187708
rect 7702 187706 7758 187708
rect 7782 187706 7838 187708
rect 7862 187706 7918 187708
rect 7622 187654 7648 187706
rect 7648 187654 7678 187706
rect 7702 187654 7712 187706
rect 7712 187654 7758 187706
rect 7782 187654 7828 187706
rect 7828 187654 7838 187706
rect 7862 187654 7892 187706
rect 7892 187654 7918 187706
rect 7622 187652 7678 187654
rect 7702 187652 7758 187654
rect 7782 187652 7838 187654
rect 7862 187652 7918 187654
rect 7622 186618 7678 186620
rect 7702 186618 7758 186620
rect 7782 186618 7838 186620
rect 7862 186618 7918 186620
rect 7622 186566 7648 186618
rect 7648 186566 7678 186618
rect 7702 186566 7712 186618
rect 7712 186566 7758 186618
rect 7782 186566 7828 186618
rect 7828 186566 7838 186618
rect 7862 186566 7892 186618
rect 7892 186566 7918 186618
rect 7622 186564 7678 186566
rect 7702 186564 7758 186566
rect 7782 186564 7838 186566
rect 7862 186564 7918 186566
rect 7622 185530 7678 185532
rect 7702 185530 7758 185532
rect 7782 185530 7838 185532
rect 7862 185530 7918 185532
rect 7622 185478 7648 185530
rect 7648 185478 7678 185530
rect 7702 185478 7712 185530
rect 7712 185478 7758 185530
rect 7782 185478 7828 185530
rect 7828 185478 7838 185530
rect 7862 185478 7892 185530
rect 7892 185478 7918 185530
rect 7622 185476 7678 185478
rect 7702 185476 7758 185478
rect 7782 185476 7838 185478
rect 7862 185476 7918 185478
rect 7622 184442 7678 184444
rect 7702 184442 7758 184444
rect 7782 184442 7838 184444
rect 7862 184442 7918 184444
rect 7622 184390 7648 184442
rect 7648 184390 7678 184442
rect 7702 184390 7712 184442
rect 7712 184390 7758 184442
rect 7782 184390 7828 184442
rect 7828 184390 7838 184442
rect 7862 184390 7892 184442
rect 7892 184390 7918 184442
rect 7622 184388 7678 184390
rect 7702 184388 7758 184390
rect 7782 184388 7838 184390
rect 7862 184388 7918 184390
rect 7622 183354 7678 183356
rect 7702 183354 7758 183356
rect 7782 183354 7838 183356
rect 7862 183354 7918 183356
rect 7622 183302 7648 183354
rect 7648 183302 7678 183354
rect 7702 183302 7712 183354
rect 7712 183302 7758 183354
rect 7782 183302 7828 183354
rect 7828 183302 7838 183354
rect 7862 183302 7892 183354
rect 7892 183302 7918 183354
rect 7622 183300 7678 183302
rect 7702 183300 7758 183302
rect 7782 183300 7838 183302
rect 7862 183300 7918 183302
rect 7622 182266 7678 182268
rect 7702 182266 7758 182268
rect 7782 182266 7838 182268
rect 7862 182266 7918 182268
rect 7622 182214 7648 182266
rect 7648 182214 7678 182266
rect 7702 182214 7712 182266
rect 7712 182214 7758 182266
rect 7782 182214 7828 182266
rect 7828 182214 7838 182266
rect 7862 182214 7892 182266
rect 7892 182214 7918 182266
rect 7622 182212 7678 182214
rect 7702 182212 7758 182214
rect 7782 182212 7838 182214
rect 7862 182212 7918 182214
rect 7622 181178 7678 181180
rect 7702 181178 7758 181180
rect 7782 181178 7838 181180
rect 7862 181178 7918 181180
rect 7622 181126 7648 181178
rect 7648 181126 7678 181178
rect 7702 181126 7712 181178
rect 7712 181126 7758 181178
rect 7782 181126 7828 181178
rect 7828 181126 7838 181178
rect 7862 181126 7892 181178
rect 7892 181126 7918 181178
rect 7622 181124 7678 181126
rect 7702 181124 7758 181126
rect 7782 181124 7838 181126
rect 7862 181124 7918 181126
rect 7622 180090 7678 180092
rect 7702 180090 7758 180092
rect 7782 180090 7838 180092
rect 7862 180090 7918 180092
rect 7622 180038 7648 180090
rect 7648 180038 7678 180090
rect 7702 180038 7712 180090
rect 7712 180038 7758 180090
rect 7782 180038 7828 180090
rect 7828 180038 7838 180090
rect 7862 180038 7892 180090
rect 7892 180038 7918 180090
rect 7622 180036 7678 180038
rect 7702 180036 7758 180038
rect 7782 180036 7838 180038
rect 7862 180036 7918 180038
rect 7622 179002 7678 179004
rect 7702 179002 7758 179004
rect 7782 179002 7838 179004
rect 7862 179002 7918 179004
rect 7622 178950 7648 179002
rect 7648 178950 7678 179002
rect 7702 178950 7712 179002
rect 7712 178950 7758 179002
rect 7782 178950 7828 179002
rect 7828 178950 7838 179002
rect 7862 178950 7892 179002
rect 7892 178950 7918 179002
rect 7622 178948 7678 178950
rect 7702 178948 7758 178950
rect 7782 178948 7838 178950
rect 7862 178948 7918 178950
rect 7622 177914 7678 177916
rect 7702 177914 7758 177916
rect 7782 177914 7838 177916
rect 7862 177914 7918 177916
rect 7622 177862 7648 177914
rect 7648 177862 7678 177914
rect 7702 177862 7712 177914
rect 7712 177862 7758 177914
rect 7782 177862 7828 177914
rect 7828 177862 7838 177914
rect 7862 177862 7892 177914
rect 7892 177862 7918 177914
rect 7622 177860 7678 177862
rect 7702 177860 7758 177862
rect 7782 177860 7838 177862
rect 7862 177860 7918 177862
rect 7622 176826 7678 176828
rect 7702 176826 7758 176828
rect 7782 176826 7838 176828
rect 7862 176826 7918 176828
rect 7622 176774 7648 176826
rect 7648 176774 7678 176826
rect 7702 176774 7712 176826
rect 7712 176774 7758 176826
rect 7782 176774 7828 176826
rect 7828 176774 7838 176826
rect 7862 176774 7892 176826
rect 7892 176774 7918 176826
rect 7622 176772 7678 176774
rect 7702 176772 7758 176774
rect 7782 176772 7838 176774
rect 7862 176772 7918 176774
rect 7622 175738 7678 175740
rect 7702 175738 7758 175740
rect 7782 175738 7838 175740
rect 7862 175738 7918 175740
rect 7622 175686 7648 175738
rect 7648 175686 7678 175738
rect 7702 175686 7712 175738
rect 7712 175686 7758 175738
rect 7782 175686 7828 175738
rect 7828 175686 7838 175738
rect 7862 175686 7892 175738
rect 7892 175686 7918 175738
rect 7622 175684 7678 175686
rect 7702 175684 7758 175686
rect 7782 175684 7838 175686
rect 7862 175684 7918 175686
rect 7622 174650 7678 174652
rect 7702 174650 7758 174652
rect 7782 174650 7838 174652
rect 7862 174650 7918 174652
rect 7622 174598 7648 174650
rect 7648 174598 7678 174650
rect 7702 174598 7712 174650
rect 7712 174598 7758 174650
rect 7782 174598 7828 174650
rect 7828 174598 7838 174650
rect 7862 174598 7892 174650
rect 7892 174598 7918 174650
rect 7622 174596 7678 174598
rect 7702 174596 7758 174598
rect 7782 174596 7838 174598
rect 7862 174596 7918 174598
rect 7622 173562 7678 173564
rect 7702 173562 7758 173564
rect 7782 173562 7838 173564
rect 7862 173562 7918 173564
rect 7622 173510 7648 173562
rect 7648 173510 7678 173562
rect 7702 173510 7712 173562
rect 7712 173510 7758 173562
rect 7782 173510 7828 173562
rect 7828 173510 7838 173562
rect 7862 173510 7892 173562
rect 7892 173510 7918 173562
rect 7622 173508 7678 173510
rect 7702 173508 7758 173510
rect 7782 173508 7838 173510
rect 7862 173508 7918 173510
rect 7622 172474 7678 172476
rect 7702 172474 7758 172476
rect 7782 172474 7838 172476
rect 7862 172474 7918 172476
rect 7622 172422 7648 172474
rect 7648 172422 7678 172474
rect 7702 172422 7712 172474
rect 7712 172422 7758 172474
rect 7782 172422 7828 172474
rect 7828 172422 7838 172474
rect 7862 172422 7892 172474
rect 7892 172422 7918 172474
rect 7622 172420 7678 172422
rect 7702 172420 7758 172422
rect 7782 172420 7838 172422
rect 7862 172420 7918 172422
rect 6734 116728 6790 116784
rect 5956 116442 6012 116444
rect 6036 116442 6092 116444
rect 6116 116442 6172 116444
rect 6196 116442 6252 116444
rect 5956 116390 5982 116442
rect 5982 116390 6012 116442
rect 6036 116390 6046 116442
rect 6046 116390 6092 116442
rect 6116 116390 6162 116442
rect 6162 116390 6172 116442
rect 6196 116390 6226 116442
rect 6226 116390 6252 116442
rect 5956 116388 6012 116390
rect 6036 116388 6092 116390
rect 6116 116388 6172 116390
rect 6196 116388 6252 116390
rect 5956 115354 6012 115356
rect 6036 115354 6092 115356
rect 6116 115354 6172 115356
rect 6196 115354 6252 115356
rect 5956 115302 5982 115354
rect 5982 115302 6012 115354
rect 6036 115302 6046 115354
rect 6046 115302 6092 115354
rect 6116 115302 6162 115354
rect 6162 115302 6172 115354
rect 6196 115302 6226 115354
rect 6226 115302 6252 115354
rect 5956 115300 6012 115302
rect 6036 115300 6092 115302
rect 6116 115300 6172 115302
rect 6196 115300 6252 115302
rect 5956 114266 6012 114268
rect 6036 114266 6092 114268
rect 6116 114266 6172 114268
rect 6196 114266 6252 114268
rect 5956 114214 5982 114266
rect 5982 114214 6012 114266
rect 6036 114214 6046 114266
rect 6046 114214 6092 114266
rect 6116 114214 6162 114266
rect 6162 114214 6172 114266
rect 6196 114214 6226 114266
rect 6226 114214 6252 114266
rect 5956 114212 6012 114214
rect 6036 114212 6092 114214
rect 6116 114212 6172 114214
rect 6196 114212 6252 114214
rect 5956 113178 6012 113180
rect 6036 113178 6092 113180
rect 6116 113178 6172 113180
rect 6196 113178 6252 113180
rect 5956 113126 5982 113178
rect 5982 113126 6012 113178
rect 6036 113126 6046 113178
rect 6046 113126 6092 113178
rect 6116 113126 6162 113178
rect 6162 113126 6172 113178
rect 6196 113126 6226 113178
rect 6226 113126 6252 113178
rect 5956 113124 6012 113126
rect 6036 113124 6092 113126
rect 6116 113124 6172 113126
rect 6196 113124 6252 113126
rect 5956 112090 6012 112092
rect 6036 112090 6092 112092
rect 6116 112090 6172 112092
rect 6196 112090 6252 112092
rect 5956 112038 5982 112090
rect 5982 112038 6012 112090
rect 6036 112038 6046 112090
rect 6046 112038 6092 112090
rect 6116 112038 6162 112090
rect 6162 112038 6172 112090
rect 6196 112038 6226 112090
rect 6226 112038 6252 112090
rect 5956 112036 6012 112038
rect 6036 112036 6092 112038
rect 6116 112036 6172 112038
rect 6196 112036 6252 112038
rect 5956 111002 6012 111004
rect 6036 111002 6092 111004
rect 6116 111002 6172 111004
rect 6196 111002 6252 111004
rect 5956 110950 5982 111002
rect 5982 110950 6012 111002
rect 6036 110950 6046 111002
rect 6046 110950 6092 111002
rect 6116 110950 6162 111002
rect 6162 110950 6172 111002
rect 6196 110950 6226 111002
rect 6226 110950 6252 111002
rect 5956 110948 6012 110950
rect 6036 110948 6092 110950
rect 6116 110948 6172 110950
rect 6196 110948 6252 110950
rect 5956 109914 6012 109916
rect 6036 109914 6092 109916
rect 6116 109914 6172 109916
rect 6196 109914 6252 109916
rect 5956 109862 5982 109914
rect 5982 109862 6012 109914
rect 6036 109862 6046 109914
rect 6046 109862 6092 109914
rect 6116 109862 6162 109914
rect 6162 109862 6172 109914
rect 6196 109862 6226 109914
rect 6226 109862 6252 109914
rect 5956 109860 6012 109862
rect 6036 109860 6092 109862
rect 6116 109860 6172 109862
rect 6196 109860 6252 109862
rect 5956 108826 6012 108828
rect 6036 108826 6092 108828
rect 6116 108826 6172 108828
rect 6196 108826 6252 108828
rect 5956 108774 5982 108826
rect 5982 108774 6012 108826
rect 6036 108774 6046 108826
rect 6046 108774 6092 108826
rect 6116 108774 6162 108826
rect 6162 108774 6172 108826
rect 6196 108774 6226 108826
rect 6226 108774 6252 108826
rect 5956 108772 6012 108774
rect 6036 108772 6092 108774
rect 6116 108772 6172 108774
rect 6196 108772 6252 108774
rect 5956 107738 6012 107740
rect 6036 107738 6092 107740
rect 6116 107738 6172 107740
rect 6196 107738 6252 107740
rect 5956 107686 5982 107738
rect 5982 107686 6012 107738
rect 6036 107686 6046 107738
rect 6046 107686 6092 107738
rect 6116 107686 6162 107738
rect 6162 107686 6172 107738
rect 6196 107686 6226 107738
rect 6226 107686 6252 107738
rect 5956 107684 6012 107686
rect 6036 107684 6092 107686
rect 6116 107684 6172 107686
rect 6196 107684 6252 107686
rect 5956 106650 6012 106652
rect 6036 106650 6092 106652
rect 6116 106650 6172 106652
rect 6196 106650 6252 106652
rect 5956 106598 5982 106650
rect 5982 106598 6012 106650
rect 6036 106598 6046 106650
rect 6046 106598 6092 106650
rect 6116 106598 6162 106650
rect 6162 106598 6172 106650
rect 6196 106598 6226 106650
rect 6226 106598 6252 106650
rect 5956 106596 6012 106598
rect 6036 106596 6092 106598
rect 6116 106596 6172 106598
rect 6196 106596 6252 106598
rect 5956 105562 6012 105564
rect 6036 105562 6092 105564
rect 6116 105562 6172 105564
rect 6196 105562 6252 105564
rect 5956 105510 5982 105562
rect 5982 105510 6012 105562
rect 6036 105510 6046 105562
rect 6046 105510 6092 105562
rect 6116 105510 6162 105562
rect 6162 105510 6172 105562
rect 6196 105510 6226 105562
rect 6226 105510 6252 105562
rect 5956 105508 6012 105510
rect 6036 105508 6092 105510
rect 6116 105508 6172 105510
rect 6196 105508 6252 105510
rect 5956 104474 6012 104476
rect 6036 104474 6092 104476
rect 6116 104474 6172 104476
rect 6196 104474 6252 104476
rect 5956 104422 5982 104474
rect 5982 104422 6012 104474
rect 6036 104422 6046 104474
rect 6046 104422 6092 104474
rect 6116 104422 6162 104474
rect 6162 104422 6172 104474
rect 6196 104422 6226 104474
rect 6226 104422 6252 104474
rect 5956 104420 6012 104422
rect 6036 104420 6092 104422
rect 6116 104420 6172 104422
rect 6196 104420 6252 104422
rect 5956 103386 6012 103388
rect 6036 103386 6092 103388
rect 6116 103386 6172 103388
rect 6196 103386 6252 103388
rect 5956 103334 5982 103386
rect 5982 103334 6012 103386
rect 6036 103334 6046 103386
rect 6046 103334 6092 103386
rect 6116 103334 6162 103386
rect 6162 103334 6172 103386
rect 6196 103334 6226 103386
rect 6226 103334 6252 103386
rect 5956 103332 6012 103334
rect 6036 103332 6092 103334
rect 6116 103332 6172 103334
rect 6196 103332 6252 103334
rect 5956 102298 6012 102300
rect 6036 102298 6092 102300
rect 6116 102298 6172 102300
rect 6196 102298 6252 102300
rect 5956 102246 5982 102298
rect 5982 102246 6012 102298
rect 6036 102246 6046 102298
rect 6046 102246 6092 102298
rect 6116 102246 6162 102298
rect 6162 102246 6172 102298
rect 6196 102246 6226 102298
rect 6226 102246 6252 102298
rect 5956 102244 6012 102246
rect 6036 102244 6092 102246
rect 6116 102244 6172 102246
rect 6196 102244 6252 102246
rect 5956 101210 6012 101212
rect 6036 101210 6092 101212
rect 6116 101210 6172 101212
rect 6196 101210 6252 101212
rect 5956 101158 5982 101210
rect 5982 101158 6012 101210
rect 6036 101158 6046 101210
rect 6046 101158 6092 101210
rect 6116 101158 6162 101210
rect 6162 101158 6172 101210
rect 6196 101158 6226 101210
rect 6226 101158 6252 101210
rect 5956 101156 6012 101158
rect 6036 101156 6092 101158
rect 6116 101156 6172 101158
rect 6196 101156 6252 101158
rect 5956 100122 6012 100124
rect 6036 100122 6092 100124
rect 6116 100122 6172 100124
rect 6196 100122 6252 100124
rect 5956 100070 5982 100122
rect 5982 100070 6012 100122
rect 6036 100070 6046 100122
rect 6046 100070 6092 100122
rect 6116 100070 6162 100122
rect 6162 100070 6172 100122
rect 6196 100070 6226 100122
rect 6226 100070 6252 100122
rect 5956 100068 6012 100070
rect 6036 100068 6092 100070
rect 6116 100068 6172 100070
rect 6196 100068 6252 100070
rect 5956 99034 6012 99036
rect 6036 99034 6092 99036
rect 6116 99034 6172 99036
rect 6196 99034 6252 99036
rect 5956 98982 5982 99034
rect 5982 98982 6012 99034
rect 6036 98982 6046 99034
rect 6046 98982 6092 99034
rect 6116 98982 6162 99034
rect 6162 98982 6172 99034
rect 6196 98982 6226 99034
rect 6226 98982 6252 99034
rect 5956 98980 6012 98982
rect 6036 98980 6092 98982
rect 6116 98980 6172 98982
rect 6196 98980 6252 98982
rect 5956 97946 6012 97948
rect 6036 97946 6092 97948
rect 6116 97946 6172 97948
rect 6196 97946 6252 97948
rect 5956 97894 5982 97946
rect 5982 97894 6012 97946
rect 6036 97894 6046 97946
rect 6046 97894 6092 97946
rect 6116 97894 6162 97946
rect 6162 97894 6172 97946
rect 6196 97894 6226 97946
rect 6226 97894 6252 97946
rect 5956 97892 6012 97894
rect 6036 97892 6092 97894
rect 6116 97892 6172 97894
rect 6196 97892 6252 97894
rect 5956 96858 6012 96860
rect 6036 96858 6092 96860
rect 6116 96858 6172 96860
rect 6196 96858 6252 96860
rect 5956 96806 5982 96858
rect 5982 96806 6012 96858
rect 6036 96806 6046 96858
rect 6046 96806 6092 96858
rect 6116 96806 6162 96858
rect 6162 96806 6172 96858
rect 6196 96806 6226 96858
rect 6226 96806 6252 96858
rect 5956 96804 6012 96806
rect 6036 96804 6092 96806
rect 6116 96804 6172 96806
rect 6196 96804 6252 96806
rect 5956 95770 6012 95772
rect 6036 95770 6092 95772
rect 6116 95770 6172 95772
rect 6196 95770 6252 95772
rect 5956 95718 5982 95770
rect 5982 95718 6012 95770
rect 6036 95718 6046 95770
rect 6046 95718 6092 95770
rect 6116 95718 6162 95770
rect 6162 95718 6172 95770
rect 6196 95718 6226 95770
rect 6226 95718 6252 95770
rect 5956 95716 6012 95718
rect 6036 95716 6092 95718
rect 6116 95716 6172 95718
rect 6196 95716 6252 95718
rect 5956 94682 6012 94684
rect 6036 94682 6092 94684
rect 6116 94682 6172 94684
rect 6196 94682 6252 94684
rect 5956 94630 5982 94682
rect 5982 94630 6012 94682
rect 6036 94630 6046 94682
rect 6046 94630 6092 94682
rect 6116 94630 6162 94682
rect 6162 94630 6172 94682
rect 6196 94630 6226 94682
rect 6226 94630 6252 94682
rect 5956 94628 6012 94630
rect 6036 94628 6092 94630
rect 6116 94628 6172 94630
rect 6196 94628 6252 94630
rect 5956 93594 6012 93596
rect 6036 93594 6092 93596
rect 6116 93594 6172 93596
rect 6196 93594 6252 93596
rect 5956 93542 5982 93594
rect 5982 93542 6012 93594
rect 6036 93542 6046 93594
rect 6046 93542 6092 93594
rect 6116 93542 6162 93594
rect 6162 93542 6172 93594
rect 6196 93542 6226 93594
rect 6226 93542 6252 93594
rect 5956 93540 6012 93542
rect 6036 93540 6092 93542
rect 6116 93540 6172 93542
rect 6196 93540 6252 93542
rect 5956 92506 6012 92508
rect 6036 92506 6092 92508
rect 6116 92506 6172 92508
rect 6196 92506 6252 92508
rect 5956 92454 5982 92506
rect 5982 92454 6012 92506
rect 6036 92454 6046 92506
rect 6046 92454 6092 92506
rect 6116 92454 6162 92506
rect 6162 92454 6172 92506
rect 6196 92454 6226 92506
rect 6226 92454 6252 92506
rect 5956 92452 6012 92454
rect 6036 92452 6092 92454
rect 6116 92452 6172 92454
rect 6196 92452 6252 92454
rect 5956 91418 6012 91420
rect 6036 91418 6092 91420
rect 6116 91418 6172 91420
rect 6196 91418 6252 91420
rect 5956 91366 5982 91418
rect 5982 91366 6012 91418
rect 6036 91366 6046 91418
rect 6046 91366 6092 91418
rect 6116 91366 6162 91418
rect 6162 91366 6172 91418
rect 6196 91366 6226 91418
rect 6226 91366 6252 91418
rect 5956 91364 6012 91366
rect 6036 91364 6092 91366
rect 6116 91364 6172 91366
rect 6196 91364 6252 91366
rect 5956 90330 6012 90332
rect 6036 90330 6092 90332
rect 6116 90330 6172 90332
rect 6196 90330 6252 90332
rect 5956 90278 5982 90330
rect 5982 90278 6012 90330
rect 6036 90278 6046 90330
rect 6046 90278 6092 90330
rect 6116 90278 6162 90330
rect 6162 90278 6172 90330
rect 6196 90278 6226 90330
rect 6226 90278 6252 90330
rect 5956 90276 6012 90278
rect 6036 90276 6092 90278
rect 6116 90276 6172 90278
rect 6196 90276 6252 90278
rect 5956 89242 6012 89244
rect 6036 89242 6092 89244
rect 6116 89242 6172 89244
rect 6196 89242 6252 89244
rect 5956 89190 5982 89242
rect 5982 89190 6012 89242
rect 6036 89190 6046 89242
rect 6046 89190 6092 89242
rect 6116 89190 6162 89242
rect 6162 89190 6172 89242
rect 6196 89190 6226 89242
rect 6226 89190 6252 89242
rect 5956 89188 6012 89190
rect 6036 89188 6092 89190
rect 6116 89188 6172 89190
rect 6196 89188 6252 89190
rect 5956 88154 6012 88156
rect 6036 88154 6092 88156
rect 6116 88154 6172 88156
rect 6196 88154 6252 88156
rect 5956 88102 5982 88154
rect 5982 88102 6012 88154
rect 6036 88102 6046 88154
rect 6046 88102 6092 88154
rect 6116 88102 6162 88154
rect 6162 88102 6172 88154
rect 6196 88102 6226 88154
rect 6226 88102 6252 88154
rect 5956 88100 6012 88102
rect 6036 88100 6092 88102
rect 6116 88100 6172 88102
rect 6196 88100 6252 88102
rect 5956 87066 6012 87068
rect 6036 87066 6092 87068
rect 6116 87066 6172 87068
rect 6196 87066 6252 87068
rect 5956 87014 5982 87066
rect 5982 87014 6012 87066
rect 6036 87014 6046 87066
rect 6046 87014 6092 87066
rect 6116 87014 6162 87066
rect 6162 87014 6172 87066
rect 6196 87014 6226 87066
rect 6226 87014 6252 87066
rect 5956 87012 6012 87014
rect 6036 87012 6092 87014
rect 6116 87012 6172 87014
rect 6196 87012 6252 87014
rect 5956 85978 6012 85980
rect 6036 85978 6092 85980
rect 6116 85978 6172 85980
rect 6196 85978 6252 85980
rect 5956 85926 5982 85978
rect 5982 85926 6012 85978
rect 6036 85926 6046 85978
rect 6046 85926 6092 85978
rect 6116 85926 6162 85978
rect 6162 85926 6172 85978
rect 6196 85926 6226 85978
rect 6226 85926 6252 85978
rect 5956 85924 6012 85926
rect 6036 85924 6092 85926
rect 6116 85924 6172 85926
rect 6196 85924 6252 85926
rect 5956 84890 6012 84892
rect 6036 84890 6092 84892
rect 6116 84890 6172 84892
rect 6196 84890 6252 84892
rect 5956 84838 5982 84890
rect 5982 84838 6012 84890
rect 6036 84838 6046 84890
rect 6046 84838 6092 84890
rect 6116 84838 6162 84890
rect 6162 84838 6172 84890
rect 6196 84838 6226 84890
rect 6226 84838 6252 84890
rect 5956 84836 6012 84838
rect 6036 84836 6092 84838
rect 6116 84836 6172 84838
rect 6196 84836 6252 84838
rect 5956 83802 6012 83804
rect 6036 83802 6092 83804
rect 6116 83802 6172 83804
rect 6196 83802 6252 83804
rect 5956 83750 5982 83802
rect 5982 83750 6012 83802
rect 6036 83750 6046 83802
rect 6046 83750 6092 83802
rect 6116 83750 6162 83802
rect 6162 83750 6172 83802
rect 6196 83750 6226 83802
rect 6226 83750 6252 83802
rect 5956 83748 6012 83750
rect 6036 83748 6092 83750
rect 6116 83748 6172 83750
rect 6196 83748 6252 83750
rect 5956 82714 6012 82716
rect 6036 82714 6092 82716
rect 6116 82714 6172 82716
rect 6196 82714 6252 82716
rect 5956 82662 5982 82714
rect 5982 82662 6012 82714
rect 6036 82662 6046 82714
rect 6046 82662 6092 82714
rect 6116 82662 6162 82714
rect 6162 82662 6172 82714
rect 6196 82662 6226 82714
rect 6226 82662 6252 82714
rect 5956 82660 6012 82662
rect 6036 82660 6092 82662
rect 6116 82660 6172 82662
rect 6196 82660 6252 82662
rect 5956 81626 6012 81628
rect 6036 81626 6092 81628
rect 6116 81626 6172 81628
rect 6196 81626 6252 81628
rect 5956 81574 5982 81626
rect 5982 81574 6012 81626
rect 6036 81574 6046 81626
rect 6046 81574 6092 81626
rect 6116 81574 6162 81626
rect 6162 81574 6172 81626
rect 6196 81574 6226 81626
rect 6226 81574 6252 81626
rect 5956 81572 6012 81574
rect 6036 81572 6092 81574
rect 6116 81572 6172 81574
rect 6196 81572 6252 81574
rect 5956 80538 6012 80540
rect 6036 80538 6092 80540
rect 6116 80538 6172 80540
rect 6196 80538 6252 80540
rect 5956 80486 5982 80538
rect 5982 80486 6012 80538
rect 6036 80486 6046 80538
rect 6046 80486 6092 80538
rect 6116 80486 6162 80538
rect 6162 80486 6172 80538
rect 6196 80486 6226 80538
rect 6226 80486 6252 80538
rect 5956 80484 6012 80486
rect 6036 80484 6092 80486
rect 6116 80484 6172 80486
rect 6196 80484 6252 80486
rect 5956 79450 6012 79452
rect 6036 79450 6092 79452
rect 6116 79450 6172 79452
rect 6196 79450 6252 79452
rect 5956 79398 5982 79450
rect 5982 79398 6012 79450
rect 6036 79398 6046 79450
rect 6046 79398 6092 79450
rect 6116 79398 6162 79450
rect 6162 79398 6172 79450
rect 6196 79398 6226 79450
rect 6226 79398 6252 79450
rect 5956 79396 6012 79398
rect 6036 79396 6092 79398
rect 6116 79396 6172 79398
rect 6196 79396 6252 79398
rect 5956 78362 6012 78364
rect 6036 78362 6092 78364
rect 6116 78362 6172 78364
rect 6196 78362 6252 78364
rect 5956 78310 5982 78362
rect 5982 78310 6012 78362
rect 6036 78310 6046 78362
rect 6046 78310 6092 78362
rect 6116 78310 6162 78362
rect 6162 78310 6172 78362
rect 6196 78310 6226 78362
rect 6226 78310 6252 78362
rect 5956 78308 6012 78310
rect 6036 78308 6092 78310
rect 6116 78308 6172 78310
rect 6196 78308 6252 78310
rect 5956 77274 6012 77276
rect 6036 77274 6092 77276
rect 6116 77274 6172 77276
rect 6196 77274 6252 77276
rect 5956 77222 5982 77274
rect 5982 77222 6012 77274
rect 6036 77222 6046 77274
rect 6046 77222 6092 77274
rect 6116 77222 6162 77274
rect 6162 77222 6172 77274
rect 6196 77222 6226 77274
rect 6226 77222 6252 77274
rect 5956 77220 6012 77222
rect 6036 77220 6092 77222
rect 6116 77220 6172 77222
rect 6196 77220 6252 77222
rect 5956 76186 6012 76188
rect 6036 76186 6092 76188
rect 6116 76186 6172 76188
rect 6196 76186 6252 76188
rect 5956 76134 5982 76186
rect 5982 76134 6012 76186
rect 6036 76134 6046 76186
rect 6046 76134 6092 76186
rect 6116 76134 6162 76186
rect 6162 76134 6172 76186
rect 6196 76134 6226 76186
rect 6226 76134 6252 76186
rect 5956 76132 6012 76134
rect 6036 76132 6092 76134
rect 6116 76132 6172 76134
rect 6196 76132 6252 76134
rect 5956 75098 6012 75100
rect 6036 75098 6092 75100
rect 6116 75098 6172 75100
rect 6196 75098 6252 75100
rect 5956 75046 5982 75098
rect 5982 75046 6012 75098
rect 6036 75046 6046 75098
rect 6046 75046 6092 75098
rect 6116 75046 6162 75098
rect 6162 75046 6172 75098
rect 6196 75046 6226 75098
rect 6226 75046 6252 75098
rect 5956 75044 6012 75046
rect 6036 75044 6092 75046
rect 6116 75044 6172 75046
rect 6196 75044 6252 75046
rect 5956 74010 6012 74012
rect 6036 74010 6092 74012
rect 6116 74010 6172 74012
rect 6196 74010 6252 74012
rect 5956 73958 5982 74010
rect 5982 73958 6012 74010
rect 6036 73958 6046 74010
rect 6046 73958 6092 74010
rect 6116 73958 6162 74010
rect 6162 73958 6172 74010
rect 6196 73958 6226 74010
rect 6226 73958 6252 74010
rect 5956 73956 6012 73958
rect 6036 73956 6092 73958
rect 6116 73956 6172 73958
rect 6196 73956 6252 73958
rect 5956 72922 6012 72924
rect 6036 72922 6092 72924
rect 6116 72922 6172 72924
rect 6196 72922 6252 72924
rect 5956 72870 5982 72922
rect 5982 72870 6012 72922
rect 6036 72870 6046 72922
rect 6046 72870 6092 72922
rect 6116 72870 6162 72922
rect 6162 72870 6172 72922
rect 6196 72870 6226 72922
rect 6226 72870 6252 72922
rect 5956 72868 6012 72870
rect 6036 72868 6092 72870
rect 6116 72868 6172 72870
rect 6196 72868 6252 72870
rect 5956 71834 6012 71836
rect 6036 71834 6092 71836
rect 6116 71834 6172 71836
rect 6196 71834 6252 71836
rect 5956 71782 5982 71834
rect 5982 71782 6012 71834
rect 6036 71782 6046 71834
rect 6046 71782 6092 71834
rect 6116 71782 6162 71834
rect 6162 71782 6172 71834
rect 6196 71782 6226 71834
rect 6226 71782 6252 71834
rect 5956 71780 6012 71782
rect 6036 71780 6092 71782
rect 6116 71780 6172 71782
rect 6196 71780 6252 71782
rect 5956 70746 6012 70748
rect 6036 70746 6092 70748
rect 6116 70746 6172 70748
rect 6196 70746 6252 70748
rect 5956 70694 5982 70746
rect 5982 70694 6012 70746
rect 6036 70694 6046 70746
rect 6046 70694 6092 70746
rect 6116 70694 6162 70746
rect 6162 70694 6172 70746
rect 6196 70694 6226 70746
rect 6226 70694 6252 70746
rect 5956 70692 6012 70694
rect 6036 70692 6092 70694
rect 6116 70692 6172 70694
rect 6196 70692 6252 70694
rect 5956 69658 6012 69660
rect 6036 69658 6092 69660
rect 6116 69658 6172 69660
rect 6196 69658 6252 69660
rect 5956 69606 5982 69658
rect 5982 69606 6012 69658
rect 6036 69606 6046 69658
rect 6046 69606 6092 69658
rect 6116 69606 6162 69658
rect 6162 69606 6172 69658
rect 6196 69606 6226 69658
rect 6226 69606 6252 69658
rect 5956 69604 6012 69606
rect 6036 69604 6092 69606
rect 6116 69604 6172 69606
rect 6196 69604 6252 69606
rect 5956 68570 6012 68572
rect 6036 68570 6092 68572
rect 6116 68570 6172 68572
rect 6196 68570 6252 68572
rect 5956 68518 5982 68570
rect 5982 68518 6012 68570
rect 6036 68518 6046 68570
rect 6046 68518 6092 68570
rect 6116 68518 6162 68570
rect 6162 68518 6172 68570
rect 6196 68518 6226 68570
rect 6226 68518 6252 68570
rect 5956 68516 6012 68518
rect 6036 68516 6092 68518
rect 6116 68516 6172 68518
rect 6196 68516 6252 68518
rect 5956 67482 6012 67484
rect 6036 67482 6092 67484
rect 6116 67482 6172 67484
rect 6196 67482 6252 67484
rect 5956 67430 5982 67482
rect 5982 67430 6012 67482
rect 6036 67430 6046 67482
rect 6046 67430 6092 67482
rect 6116 67430 6162 67482
rect 6162 67430 6172 67482
rect 6196 67430 6226 67482
rect 6226 67430 6252 67482
rect 5956 67428 6012 67430
rect 6036 67428 6092 67430
rect 6116 67428 6172 67430
rect 6196 67428 6252 67430
rect 5956 66394 6012 66396
rect 6036 66394 6092 66396
rect 6116 66394 6172 66396
rect 6196 66394 6252 66396
rect 5956 66342 5982 66394
rect 5982 66342 6012 66394
rect 6036 66342 6046 66394
rect 6046 66342 6092 66394
rect 6116 66342 6162 66394
rect 6162 66342 6172 66394
rect 6196 66342 6226 66394
rect 6226 66342 6252 66394
rect 5956 66340 6012 66342
rect 6036 66340 6092 66342
rect 6116 66340 6172 66342
rect 6196 66340 6252 66342
rect 5956 65306 6012 65308
rect 6036 65306 6092 65308
rect 6116 65306 6172 65308
rect 6196 65306 6252 65308
rect 5956 65254 5982 65306
rect 5982 65254 6012 65306
rect 6036 65254 6046 65306
rect 6046 65254 6092 65306
rect 6116 65254 6162 65306
rect 6162 65254 6172 65306
rect 6196 65254 6226 65306
rect 6226 65254 6252 65306
rect 5956 65252 6012 65254
rect 6036 65252 6092 65254
rect 6116 65252 6172 65254
rect 6196 65252 6252 65254
rect 5956 64218 6012 64220
rect 6036 64218 6092 64220
rect 6116 64218 6172 64220
rect 6196 64218 6252 64220
rect 5956 64166 5982 64218
rect 5982 64166 6012 64218
rect 6036 64166 6046 64218
rect 6046 64166 6092 64218
rect 6116 64166 6162 64218
rect 6162 64166 6172 64218
rect 6196 64166 6226 64218
rect 6226 64166 6252 64218
rect 5956 64164 6012 64166
rect 6036 64164 6092 64166
rect 6116 64164 6172 64166
rect 6196 64164 6252 64166
rect 5956 63130 6012 63132
rect 6036 63130 6092 63132
rect 6116 63130 6172 63132
rect 6196 63130 6252 63132
rect 5956 63078 5982 63130
rect 5982 63078 6012 63130
rect 6036 63078 6046 63130
rect 6046 63078 6092 63130
rect 6116 63078 6162 63130
rect 6162 63078 6172 63130
rect 6196 63078 6226 63130
rect 6226 63078 6252 63130
rect 5956 63076 6012 63078
rect 6036 63076 6092 63078
rect 6116 63076 6172 63078
rect 6196 63076 6252 63078
rect 5956 62042 6012 62044
rect 6036 62042 6092 62044
rect 6116 62042 6172 62044
rect 6196 62042 6252 62044
rect 5956 61990 5982 62042
rect 5982 61990 6012 62042
rect 6036 61990 6046 62042
rect 6046 61990 6092 62042
rect 6116 61990 6162 62042
rect 6162 61990 6172 62042
rect 6196 61990 6226 62042
rect 6226 61990 6252 62042
rect 5956 61988 6012 61990
rect 6036 61988 6092 61990
rect 6116 61988 6172 61990
rect 6196 61988 6252 61990
rect 5956 60954 6012 60956
rect 6036 60954 6092 60956
rect 6116 60954 6172 60956
rect 6196 60954 6252 60956
rect 5956 60902 5982 60954
rect 5982 60902 6012 60954
rect 6036 60902 6046 60954
rect 6046 60902 6092 60954
rect 6116 60902 6162 60954
rect 6162 60902 6172 60954
rect 6196 60902 6226 60954
rect 6226 60902 6252 60954
rect 5956 60900 6012 60902
rect 6036 60900 6092 60902
rect 6116 60900 6172 60902
rect 6196 60900 6252 60902
rect 5956 59866 6012 59868
rect 6036 59866 6092 59868
rect 6116 59866 6172 59868
rect 6196 59866 6252 59868
rect 5956 59814 5982 59866
rect 5982 59814 6012 59866
rect 6036 59814 6046 59866
rect 6046 59814 6092 59866
rect 6116 59814 6162 59866
rect 6162 59814 6172 59866
rect 6196 59814 6226 59866
rect 6226 59814 6252 59866
rect 5956 59812 6012 59814
rect 6036 59812 6092 59814
rect 6116 59812 6172 59814
rect 6196 59812 6252 59814
rect 5956 58778 6012 58780
rect 6036 58778 6092 58780
rect 6116 58778 6172 58780
rect 6196 58778 6252 58780
rect 5956 58726 5982 58778
rect 5982 58726 6012 58778
rect 6036 58726 6046 58778
rect 6046 58726 6092 58778
rect 6116 58726 6162 58778
rect 6162 58726 6172 58778
rect 6196 58726 6226 58778
rect 6226 58726 6252 58778
rect 5956 58724 6012 58726
rect 6036 58724 6092 58726
rect 6116 58724 6172 58726
rect 6196 58724 6252 58726
rect 5956 57690 6012 57692
rect 6036 57690 6092 57692
rect 6116 57690 6172 57692
rect 6196 57690 6252 57692
rect 5956 57638 5982 57690
rect 5982 57638 6012 57690
rect 6036 57638 6046 57690
rect 6046 57638 6092 57690
rect 6116 57638 6162 57690
rect 6162 57638 6172 57690
rect 6196 57638 6226 57690
rect 6226 57638 6252 57690
rect 5956 57636 6012 57638
rect 6036 57636 6092 57638
rect 6116 57636 6172 57638
rect 6196 57636 6252 57638
rect 5956 56602 6012 56604
rect 6036 56602 6092 56604
rect 6116 56602 6172 56604
rect 6196 56602 6252 56604
rect 5956 56550 5982 56602
rect 5982 56550 6012 56602
rect 6036 56550 6046 56602
rect 6046 56550 6092 56602
rect 6116 56550 6162 56602
rect 6162 56550 6172 56602
rect 6196 56550 6226 56602
rect 6226 56550 6252 56602
rect 5956 56548 6012 56550
rect 6036 56548 6092 56550
rect 6116 56548 6172 56550
rect 6196 56548 6252 56550
rect 5956 55514 6012 55516
rect 6036 55514 6092 55516
rect 6116 55514 6172 55516
rect 6196 55514 6252 55516
rect 5956 55462 5982 55514
rect 5982 55462 6012 55514
rect 6036 55462 6046 55514
rect 6046 55462 6092 55514
rect 6116 55462 6162 55514
rect 6162 55462 6172 55514
rect 6196 55462 6226 55514
rect 6226 55462 6252 55514
rect 5956 55460 6012 55462
rect 6036 55460 6092 55462
rect 6116 55460 6172 55462
rect 6196 55460 6252 55462
rect 5956 54426 6012 54428
rect 6036 54426 6092 54428
rect 6116 54426 6172 54428
rect 6196 54426 6252 54428
rect 5956 54374 5982 54426
rect 5982 54374 6012 54426
rect 6036 54374 6046 54426
rect 6046 54374 6092 54426
rect 6116 54374 6162 54426
rect 6162 54374 6172 54426
rect 6196 54374 6226 54426
rect 6226 54374 6252 54426
rect 5956 54372 6012 54374
rect 6036 54372 6092 54374
rect 6116 54372 6172 54374
rect 6196 54372 6252 54374
rect 5956 53338 6012 53340
rect 6036 53338 6092 53340
rect 6116 53338 6172 53340
rect 6196 53338 6252 53340
rect 5956 53286 5982 53338
rect 5982 53286 6012 53338
rect 6036 53286 6046 53338
rect 6046 53286 6092 53338
rect 6116 53286 6162 53338
rect 6162 53286 6172 53338
rect 6196 53286 6226 53338
rect 6226 53286 6252 53338
rect 5956 53284 6012 53286
rect 6036 53284 6092 53286
rect 6116 53284 6172 53286
rect 6196 53284 6252 53286
rect 5956 52250 6012 52252
rect 6036 52250 6092 52252
rect 6116 52250 6172 52252
rect 6196 52250 6252 52252
rect 5956 52198 5982 52250
rect 5982 52198 6012 52250
rect 6036 52198 6046 52250
rect 6046 52198 6092 52250
rect 6116 52198 6162 52250
rect 6162 52198 6172 52250
rect 6196 52198 6226 52250
rect 6226 52198 6252 52250
rect 5956 52196 6012 52198
rect 6036 52196 6092 52198
rect 6116 52196 6172 52198
rect 6196 52196 6252 52198
rect 5956 51162 6012 51164
rect 6036 51162 6092 51164
rect 6116 51162 6172 51164
rect 6196 51162 6252 51164
rect 5956 51110 5982 51162
rect 5982 51110 6012 51162
rect 6036 51110 6046 51162
rect 6046 51110 6092 51162
rect 6116 51110 6162 51162
rect 6162 51110 6172 51162
rect 6196 51110 6226 51162
rect 6226 51110 6252 51162
rect 5956 51108 6012 51110
rect 6036 51108 6092 51110
rect 6116 51108 6172 51110
rect 6196 51108 6252 51110
rect 7622 171386 7678 171388
rect 7702 171386 7758 171388
rect 7782 171386 7838 171388
rect 7862 171386 7918 171388
rect 7622 171334 7648 171386
rect 7648 171334 7678 171386
rect 7702 171334 7712 171386
rect 7712 171334 7758 171386
rect 7782 171334 7828 171386
rect 7828 171334 7838 171386
rect 7862 171334 7892 171386
rect 7892 171334 7918 171386
rect 7622 171332 7678 171334
rect 7702 171332 7758 171334
rect 7782 171332 7838 171334
rect 7862 171332 7918 171334
rect 7622 170298 7678 170300
rect 7702 170298 7758 170300
rect 7782 170298 7838 170300
rect 7862 170298 7918 170300
rect 7622 170246 7648 170298
rect 7648 170246 7678 170298
rect 7702 170246 7712 170298
rect 7712 170246 7758 170298
rect 7782 170246 7828 170298
rect 7828 170246 7838 170298
rect 7862 170246 7892 170298
rect 7892 170246 7918 170298
rect 7622 170244 7678 170246
rect 7702 170244 7758 170246
rect 7782 170244 7838 170246
rect 7862 170244 7918 170246
rect 7622 169210 7678 169212
rect 7702 169210 7758 169212
rect 7782 169210 7838 169212
rect 7862 169210 7918 169212
rect 7622 169158 7648 169210
rect 7648 169158 7678 169210
rect 7702 169158 7712 169210
rect 7712 169158 7758 169210
rect 7782 169158 7828 169210
rect 7828 169158 7838 169210
rect 7862 169158 7892 169210
rect 7892 169158 7918 169210
rect 7622 169156 7678 169158
rect 7702 169156 7758 169158
rect 7782 169156 7838 169158
rect 7862 169156 7918 169158
rect 7622 168122 7678 168124
rect 7702 168122 7758 168124
rect 7782 168122 7838 168124
rect 7862 168122 7918 168124
rect 7622 168070 7648 168122
rect 7648 168070 7678 168122
rect 7702 168070 7712 168122
rect 7712 168070 7758 168122
rect 7782 168070 7828 168122
rect 7828 168070 7838 168122
rect 7862 168070 7892 168122
rect 7892 168070 7918 168122
rect 7622 168068 7678 168070
rect 7702 168068 7758 168070
rect 7782 168068 7838 168070
rect 7862 168068 7918 168070
rect 7622 167034 7678 167036
rect 7702 167034 7758 167036
rect 7782 167034 7838 167036
rect 7862 167034 7918 167036
rect 7622 166982 7648 167034
rect 7648 166982 7678 167034
rect 7702 166982 7712 167034
rect 7712 166982 7758 167034
rect 7782 166982 7828 167034
rect 7828 166982 7838 167034
rect 7862 166982 7892 167034
rect 7892 166982 7918 167034
rect 7622 166980 7678 166982
rect 7702 166980 7758 166982
rect 7782 166980 7838 166982
rect 7862 166980 7918 166982
rect 7622 165946 7678 165948
rect 7702 165946 7758 165948
rect 7782 165946 7838 165948
rect 7862 165946 7918 165948
rect 7622 165894 7648 165946
rect 7648 165894 7678 165946
rect 7702 165894 7712 165946
rect 7712 165894 7758 165946
rect 7782 165894 7828 165946
rect 7828 165894 7838 165946
rect 7862 165894 7892 165946
rect 7892 165894 7918 165946
rect 7622 165892 7678 165894
rect 7702 165892 7758 165894
rect 7782 165892 7838 165894
rect 7862 165892 7918 165894
rect 7622 164858 7678 164860
rect 7702 164858 7758 164860
rect 7782 164858 7838 164860
rect 7862 164858 7918 164860
rect 7622 164806 7648 164858
rect 7648 164806 7678 164858
rect 7702 164806 7712 164858
rect 7712 164806 7758 164858
rect 7782 164806 7828 164858
rect 7828 164806 7838 164858
rect 7862 164806 7892 164858
rect 7892 164806 7918 164858
rect 7622 164804 7678 164806
rect 7702 164804 7758 164806
rect 7782 164804 7838 164806
rect 7862 164804 7918 164806
rect 7622 163770 7678 163772
rect 7702 163770 7758 163772
rect 7782 163770 7838 163772
rect 7862 163770 7918 163772
rect 7622 163718 7648 163770
rect 7648 163718 7678 163770
rect 7702 163718 7712 163770
rect 7712 163718 7758 163770
rect 7782 163718 7828 163770
rect 7828 163718 7838 163770
rect 7862 163718 7892 163770
rect 7892 163718 7918 163770
rect 7622 163716 7678 163718
rect 7702 163716 7758 163718
rect 7782 163716 7838 163718
rect 7862 163716 7918 163718
rect 7622 162682 7678 162684
rect 7702 162682 7758 162684
rect 7782 162682 7838 162684
rect 7862 162682 7918 162684
rect 7622 162630 7648 162682
rect 7648 162630 7678 162682
rect 7702 162630 7712 162682
rect 7712 162630 7758 162682
rect 7782 162630 7828 162682
rect 7828 162630 7838 162682
rect 7862 162630 7892 162682
rect 7892 162630 7918 162682
rect 7622 162628 7678 162630
rect 7702 162628 7758 162630
rect 7782 162628 7838 162630
rect 7862 162628 7918 162630
rect 7622 161594 7678 161596
rect 7702 161594 7758 161596
rect 7782 161594 7838 161596
rect 7862 161594 7918 161596
rect 7622 161542 7648 161594
rect 7648 161542 7678 161594
rect 7702 161542 7712 161594
rect 7712 161542 7758 161594
rect 7782 161542 7828 161594
rect 7828 161542 7838 161594
rect 7862 161542 7892 161594
rect 7892 161542 7918 161594
rect 7622 161540 7678 161542
rect 7702 161540 7758 161542
rect 7782 161540 7838 161542
rect 7862 161540 7918 161542
rect 7622 160506 7678 160508
rect 7702 160506 7758 160508
rect 7782 160506 7838 160508
rect 7862 160506 7918 160508
rect 7622 160454 7648 160506
rect 7648 160454 7678 160506
rect 7702 160454 7712 160506
rect 7712 160454 7758 160506
rect 7782 160454 7828 160506
rect 7828 160454 7838 160506
rect 7862 160454 7892 160506
rect 7892 160454 7918 160506
rect 7622 160452 7678 160454
rect 7702 160452 7758 160454
rect 7782 160452 7838 160454
rect 7862 160452 7918 160454
rect 7622 159418 7678 159420
rect 7702 159418 7758 159420
rect 7782 159418 7838 159420
rect 7862 159418 7918 159420
rect 7622 159366 7648 159418
rect 7648 159366 7678 159418
rect 7702 159366 7712 159418
rect 7712 159366 7758 159418
rect 7782 159366 7828 159418
rect 7828 159366 7838 159418
rect 7862 159366 7892 159418
rect 7892 159366 7918 159418
rect 7622 159364 7678 159366
rect 7702 159364 7758 159366
rect 7782 159364 7838 159366
rect 7862 159364 7918 159366
rect 7622 158330 7678 158332
rect 7702 158330 7758 158332
rect 7782 158330 7838 158332
rect 7862 158330 7918 158332
rect 7622 158278 7648 158330
rect 7648 158278 7678 158330
rect 7702 158278 7712 158330
rect 7712 158278 7758 158330
rect 7782 158278 7828 158330
rect 7828 158278 7838 158330
rect 7862 158278 7892 158330
rect 7892 158278 7918 158330
rect 7622 158276 7678 158278
rect 7702 158276 7758 158278
rect 7782 158276 7838 158278
rect 7862 158276 7918 158278
rect 6826 50360 6882 50416
rect 5956 50074 6012 50076
rect 6036 50074 6092 50076
rect 6116 50074 6172 50076
rect 6196 50074 6252 50076
rect 5956 50022 5982 50074
rect 5982 50022 6012 50074
rect 6036 50022 6046 50074
rect 6046 50022 6092 50074
rect 6116 50022 6162 50074
rect 6162 50022 6172 50074
rect 6196 50022 6226 50074
rect 6226 50022 6252 50074
rect 5956 50020 6012 50022
rect 6036 50020 6092 50022
rect 6116 50020 6172 50022
rect 6196 50020 6252 50022
rect 5956 48986 6012 48988
rect 6036 48986 6092 48988
rect 6116 48986 6172 48988
rect 6196 48986 6252 48988
rect 5956 48934 5982 48986
rect 5982 48934 6012 48986
rect 6036 48934 6046 48986
rect 6046 48934 6092 48986
rect 6116 48934 6162 48986
rect 6162 48934 6172 48986
rect 6196 48934 6226 48986
rect 6226 48934 6252 48986
rect 5956 48932 6012 48934
rect 6036 48932 6092 48934
rect 6116 48932 6172 48934
rect 6196 48932 6252 48934
rect 5956 47898 6012 47900
rect 6036 47898 6092 47900
rect 6116 47898 6172 47900
rect 6196 47898 6252 47900
rect 5956 47846 5982 47898
rect 5982 47846 6012 47898
rect 6036 47846 6046 47898
rect 6046 47846 6092 47898
rect 6116 47846 6162 47898
rect 6162 47846 6172 47898
rect 6196 47846 6226 47898
rect 6226 47846 6252 47898
rect 5956 47844 6012 47846
rect 6036 47844 6092 47846
rect 6116 47844 6172 47846
rect 6196 47844 6252 47846
rect 5956 46810 6012 46812
rect 6036 46810 6092 46812
rect 6116 46810 6172 46812
rect 6196 46810 6252 46812
rect 5956 46758 5982 46810
rect 5982 46758 6012 46810
rect 6036 46758 6046 46810
rect 6046 46758 6092 46810
rect 6116 46758 6162 46810
rect 6162 46758 6172 46810
rect 6196 46758 6226 46810
rect 6226 46758 6252 46810
rect 5956 46756 6012 46758
rect 6036 46756 6092 46758
rect 6116 46756 6172 46758
rect 6196 46756 6252 46758
rect 5956 45722 6012 45724
rect 6036 45722 6092 45724
rect 6116 45722 6172 45724
rect 6196 45722 6252 45724
rect 5956 45670 5982 45722
rect 5982 45670 6012 45722
rect 6036 45670 6046 45722
rect 6046 45670 6092 45722
rect 6116 45670 6162 45722
rect 6162 45670 6172 45722
rect 6196 45670 6226 45722
rect 6226 45670 6252 45722
rect 5956 45668 6012 45670
rect 6036 45668 6092 45670
rect 6116 45668 6172 45670
rect 6196 45668 6252 45670
rect 5956 44634 6012 44636
rect 6036 44634 6092 44636
rect 6116 44634 6172 44636
rect 6196 44634 6252 44636
rect 5956 44582 5982 44634
rect 5982 44582 6012 44634
rect 6036 44582 6046 44634
rect 6046 44582 6092 44634
rect 6116 44582 6162 44634
rect 6162 44582 6172 44634
rect 6196 44582 6226 44634
rect 6226 44582 6252 44634
rect 5956 44580 6012 44582
rect 6036 44580 6092 44582
rect 6116 44580 6172 44582
rect 6196 44580 6252 44582
rect 5956 43546 6012 43548
rect 6036 43546 6092 43548
rect 6116 43546 6172 43548
rect 6196 43546 6252 43548
rect 5956 43494 5982 43546
rect 5982 43494 6012 43546
rect 6036 43494 6046 43546
rect 6046 43494 6092 43546
rect 6116 43494 6162 43546
rect 6162 43494 6172 43546
rect 6196 43494 6226 43546
rect 6226 43494 6252 43546
rect 5956 43492 6012 43494
rect 6036 43492 6092 43494
rect 6116 43492 6172 43494
rect 6196 43492 6252 43494
rect 5956 42458 6012 42460
rect 6036 42458 6092 42460
rect 6116 42458 6172 42460
rect 6196 42458 6252 42460
rect 5956 42406 5982 42458
rect 5982 42406 6012 42458
rect 6036 42406 6046 42458
rect 6046 42406 6092 42458
rect 6116 42406 6162 42458
rect 6162 42406 6172 42458
rect 6196 42406 6226 42458
rect 6226 42406 6252 42458
rect 5956 42404 6012 42406
rect 6036 42404 6092 42406
rect 6116 42404 6172 42406
rect 6196 42404 6252 42406
rect 5956 41370 6012 41372
rect 6036 41370 6092 41372
rect 6116 41370 6172 41372
rect 6196 41370 6252 41372
rect 5956 41318 5982 41370
rect 5982 41318 6012 41370
rect 6036 41318 6046 41370
rect 6046 41318 6092 41370
rect 6116 41318 6162 41370
rect 6162 41318 6172 41370
rect 6196 41318 6226 41370
rect 6226 41318 6252 41370
rect 5956 41316 6012 41318
rect 6036 41316 6092 41318
rect 6116 41316 6172 41318
rect 6196 41316 6252 41318
rect 5956 40282 6012 40284
rect 6036 40282 6092 40284
rect 6116 40282 6172 40284
rect 6196 40282 6252 40284
rect 5956 40230 5982 40282
rect 5982 40230 6012 40282
rect 6036 40230 6046 40282
rect 6046 40230 6092 40282
rect 6116 40230 6162 40282
rect 6162 40230 6172 40282
rect 6196 40230 6226 40282
rect 6226 40230 6252 40282
rect 5956 40228 6012 40230
rect 6036 40228 6092 40230
rect 6116 40228 6172 40230
rect 6196 40228 6252 40230
rect 5956 39194 6012 39196
rect 6036 39194 6092 39196
rect 6116 39194 6172 39196
rect 6196 39194 6252 39196
rect 5956 39142 5982 39194
rect 5982 39142 6012 39194
rect 6036 39142 6046 39194
rect 6046 39142 6092 39194
rect 6116 39142 6162 39194
rect 6162 39142 6172 39194
rect 6196 39142 6226 39194
rect 6226 39142 6252 39194
rect 5956 39140 6012 39142
rect 6036 39140 6092 39142
rect 6116 39140 6172 39142
rect 6196 39140 6252 39142
rect 5956 38106 6012 38108
rect 6036 38106 6092 38108
rect 6116 38106 6172 38108
rect 6196 38106 6252 38108
rect 5956 38054 5982 38106
rect 5982 38054 6012 38106
rect 6036 38054 6046 38106
rect 6046 38054 6092 38106
rect 6116 38054 6162 38106
rect 6162 38054 6172 38106
rect 6196 38054 6226 38106
rect 6226 38054 6252 38106
rect 5956 38052 6012 38054
rect 6036 38052 6092 38054
rect 6116 38052 6172 38054
rect 6196 38052 6252 38054
rect 5956 37018 6012 37020
rect 6036 37018 6092 37020
rect 6116 37018 6172 37020
rect 6196 37018 6252 37020
rect 5956 36966 5982 37018
rect 5982 36966 6012 37018
rect 6036 36966 6046 37018
rect 6046 36966 6092 37018
rect 6116 36966 6162 37018
rect 6162 36966 6172 37018
rect 6196 36966 6226 37018
rect 6226 36966 6252 37018
rect 5956 36964 6012 36966
rect 6036 36964 6092 36966
rect 6116 36964 6172 36966
rect 6196 36964 6252 36966
rect 5956 35930 6012 35932
rect 6036 35930 6092 35932
rect 6116 35930 6172 35932
rect 6196 35930 6252 35932
rect 5956 35878 5982 35930
rect 5982 35878 6012 35930
rect 6036 35878 6046 35930
rect 6046 35878 6092 35930
rect 6116 35878 6162 35930
rect 6162 35878 6172 35930
rect 6196 35878 6226 35930
rect 6226 35878 6252 35930
rect 5956 35876 6012 35878
rect 6036 35876 6092 35878
rect 6116 35876 6172 35878
rect 6196 35876 6252 35878
rect 5956 34842 6012 34844
rect 6036 34842 6092 34844
rect 6116 34842 6172 34844
rect 6196 34842 6252 34844
rect 5956 34790 5982 34842
rect 5982 34790 6012 34842
rect 6036 34790 6046 34842
rect 6046 34790 6092 34842
rect 6116 34790 6162 34842
rect 6162 34790 6172 34842
rect 6196 34790 6226 34842
rect 6226 34790 6252 34842
rect 5956 34788 6012 34790
rect 6036 34788 6092 34790
rect 6116 34788 6172 34790
rect 6196 34788 6252 34790
rect 5956 33754 6012 33756
rect 6036 33754 6092 33756
rect 6116 33754 6172 33756
rect 6196 33754 6252 33756
rect 5956 33702 5982 33754
rect 5982 33702 6012 33754
rect 6036 33702 6046 33754
rect 6046 33702 6092 33754
rect 6116 33702 6162 33754
rect 6162 33702 6172 33754
rect 6196 33702 6226 33754
rect 6226 33702 6252 33754
rect 5956 33700 6012 33702
rect 6036 33700 6092 33702
rect 6116 33700 6172 33702
rect 6196 33700 6252 33702
rect 5956 32666 6012 32668
rect 6036 32666 6092 32668
rect 6116 32666 6172 32668
rect 6196 32666 6252 32668
rect 5956 32614 5982 32666
rect 5982 32614 6012 32666
rect 6036 32614 6046 32666
rect 6046 32614 6092 32666
rect 6116 32614 6162 32666
rect 6162 32614 6172 32666
rect 6196 32614 6226 32666
rect 6226 32614 6252 32666
rect 5956 32612 6012 32614
rect 6036 32612 6092 32614
rect 6116 32612 6172 32614
rect 6196 32612 6252 32614
rect 5956 31578 6012 31580
rect 6036 31578 6092 31580
rect 6116 31578 6172 31580
rect 6196 31578 6252 31580
rect 5956 31526 5982 31578
rect 5982 31526 6012 31578
rect 6036 31526 6046 31578
rect 6046 31526 6092 31578
rect 6116 31526 6162 31578
rect 6162 31526 6172 31578
rect 6196 31526 6226 31578
rect 6226 31526 6252 31578
rect 5956 31524 6012 31526
rect 6036 31524 6092 31526
rect 6116 31524 6172 31526
rect 6196 31524 6252 31526
rect 5956 30490 6012 30492
rect 6036 30490 6092 30492
rect 6116 30490 6172 30492
rect 6196 30490 6252 30492
rect 5956 30438 5982 30490
rect 5982 30438 6012 30490
rect 6036 30438 6046 30490
rect 6046 30438 6092 30490
rect 6116 30438 6162 30490
rect 6162 30438 6172 30490
rect 6196 30438 6226 30490
rect 6226 30438 6252 30490
rect 5956 30436 6012 30438
rect 6036 30436 6092 30438
rect 6116 30436 6172 30438
rect 6196 30436 6252 30438
rect 5956 29402 6012 29404
rect 6036 29402 6092 29404
rect 6116 29402 6172 29404
rect 6196 29402 6252 29404
rect 5956 29350 5982 29402
rect 5982 29350 6012 29402
rect 6036 29350 6046 29402
rect 6046 29350 6092 29402
rect 6116 29350 6162 29402
rect 6162 29350 6172 29402
rect 6196 29350 6226 29402
rect 6226 29350 6252 29402
rect 5956 29348 6012 29350
rect 6036 29348 6092 29350
rect 6116 29348 6172 29350
rect 6196 29348 6252 29350
rect 5956 28314 6012 28316
rect 6036 28314 6092 28316
rect 6116 28314 6172 28316
rect 6196 28314 6252 28316
rect 5956 28262 5982 28314
rect 5982 28262 6012 28314
rect 6036 28262 6046 28314
rect 6046 28262 6092 28314
rect 6116 28262 6162 28314
rect 6162 28262 6172 28314
rect 6196 28262 6226 28314
rect 6226 28262 6252 28314
rect 5956 28260 6012 28262
rect 6036 28260 6092 28262
rect 6116 28260 6172 28262
rect 6196 28260 6252 28262
rect 5956 27226 6012 27228
rect 6036 27226 6092 27228
rect 6116 27226 6172 27228
rect 6196 27226 6252 27228
rect 5956 27174 5982 27226
rect 5982 27174 6012 27226
rect 6036 27174 6046 27226
rect 6046 27174 6092 27226
rect 6116 27174 6162 27226
rect 6162 27174 6172 27226
rect 6196 27174 6226 27226
rect 6226 27174 6252 27226
rect 5956 27172 6012 27174
rect 6036 27172 6092 27174
rect 6116 27172 6172 27174
rect 6196 27172 6252 27174
rect 5956 26138 6012 26140
rect 6036 26138 6092 26140
rect 6116 26138 6172 26140
rect 6196 26138 6252 26140
rect 5956 26086 5982 26138
rect 5982 26086 6012 26138
rect 6036 26086 6046 26138
rect 6046 26086 6092 26138
rect 6116 26086 6162 26138
rect 6162 26086 6172 26138
rect 6196 26086 6226 26138
rect 6226 26086 6252 26138
rect 5956 26084 6012 26086
rect 6036 26084 6092 26086
rect 6116 26084 6172 26086
rect 6196 26084 6252 26086
rect 5956 25050 6012 25052
rect 6036 25050 6092 25052
rect 6116 25050 6172 25052
rect 6196 25050 6252 25052
rect 5956 24998 5982 25050
rect 5982 24998 6012 25050
rect 6036 24998 6046 25050
rect 6046 24998 6092 25050
rect 6116 24998 6162 25050
rect 6162 24998 6172 25050
rect 6196 24998 6226 25050
rect 6226 24998 6252 25050
rect 5956 24996 6012 24998
rect 6036 24996 6092 24998
rect 6116 24996 6172 24998
rect 6196 24996 6252 24998
rect 5956 23962 6012 23964
rect 6036 23962 6092 23964
rect 6116 23962 6172 23964
rect 6196 23962 6252 23964
rect 5956 23910 5982 23962
rect 5982 23910 6012 23962
rect 6036 23910 6046 23962
rect 6046 23910 6092 23962
rect 6116 23910 6162 23962
rect 6162 23910 6172 23962
rect 6196 23910 6226 23962
rect 6226 23910 6252 23962
rect 5956 23908 6012 23910
rect 6036 23908 6092 23910
rect 6116 23908 6172 23910
rect 6196 23908 6252 23910
rect 5956 22874 6012 22876
rect 6036 22874 6092 22876
rect 6116 22874 6172 22876
rect 6196 22874 6252 22876
rect 5956 22822 5982 22874
rect 5982 22822 6012 22874
rect 6036 22822 6046 22874
rect 6046 22822 6092 22874
rect 6116 22822 6162 22874
rect 6162 22822 6172 22874
rect 6196 22822 6226 22874
rect 6226 22822 6252 22874
rect 5956 22820 6012 22822
rect 6036 22820 6092 22822
rect 6116 22820 6172 22822
rect 6196 22820 6252 22822
rect 5956 21786 6012 21788
rect 6036 21786 6092 21788
rect 6116 21786 6172 21788
rect 6196 21786 6252 21788
rect 5956 21734 5982 21786
rect 5982 21734 6012 21786
rect 6036 21734 6046 21786
rect 6046 21734 6092 21786
rect 6116 21734 6162 21786
rect 6162 21734 6172 21786
rect 6196 21734 6226 21786
rect 6226 21734 6252 21786
rect 5956 21732 6012 21734
rect 6036 21732 6092 21734
rect 6116 21732 6172 21734
rect 6196 21732 6252 21734
rect 5956 20698 6012 20700
rect 6036 20698 6092 20700
rect 6116 20698 6172 20700
rect 6196 20698 6252 20700
rect 5956 20646 5982 20698
rect 5982 20646 6012 20698
rect 6036 20646 6046 20698
rect 6046 20646 6092 20698
rect 6116 20646 6162 20698
rect 6162 20646 6172 20698
rect 6196 20646 6226 20698
rect 6226 20646 6252 20698
rect 5956 20644 6012 20646
rect 6036 20644 6092 20646
rect 6116 20644 6172 20646
rect 6196 20644 6252 20646
rect 5956 19610 6012 19612
rect 6036 19610 6092 19612
rect 6116 19610 6172 19612
rect 6196 19610 6252 19612
rect 5956 19558 5982 19610
rect 5982 19558 6012 19610
rect 6036 19558 6046 19610
rect 6046 19558 6092 19610
rect 6116 19558 6162 19610
rect 6162 19558 6172 19610
rect 6196 19558 6226 19610
rect 6226 19558 6252 19610
rect 5956 19556 6012 19558
rect 6036 19556 6092 19558
rect 6116 19556 6172 19558
rect 6196 19556 6252 19558
rect 5956 18522 6012 18524
rect 6036 18522 6092 18524
rect 6116 18522 6172 18524
rect 6196 18522 6252 18524
rect 5956 18470 5982 18522
rect 5982 18470 6012 18522
rect 6036 18470 6046 18522
rect 6046 18470 6092 18522
rect 6116 18470 6162 18522
rect 6162 18470 6172 18522
rect 6196 18470 6226 18522
rect 6226 18470 6252 18522
rect 5956 18468 6012 18470
rect 6036 18468 6092 18470
rect 6116 18468 6172 18470
rect 6196 18468 6252 18470
rect 5956 17434 6012 17436
rect 6036 17434 6092 17436
rect 6116 17434 6172 17436
rect 6196 17434 6252 17436
rect 5956 17382 5982 17434
rect 5982 17382 6012 17434
rect 6036 17382 6046 17434
rect 6046 17382 6092 17434
rect 6116 17382 6162 17434
rect 6162 17382 6172 17434
rect 6196 17382 6226 17434
rect 6226 17382 6252 17434
rect 5956 17380 6012 17382
rect 6036 17380 6092 17382
rect 6116 17380 6172 17382
rect 6196 17380 6252 17382
rect 4802 17176 4858 17232
rect 4289 16890 4345 16892
rect 4369 16890 4425 16892
rect 4449 16890 4505 16892
rect 4529 16890 4585 16892
rect 4289 16838 4315 16890
rect 4315 16838 4345 16890
rect 4369 16838 4379 16890
rect 4379 16838 4425 16890
rect 4449 16838 4495 16890
rect 4495 16838 4505 16890
rect 4529 16838 4559 16890
rect 4559 16838 4585 16890
rect 4289 16836 4345 16838
rect 4369 16836 4425 16838
rect 4449 16836 4505 16838
rect 4529 16836 4585 16838
rect 5956 16346 6012 16348
rect 6036 16346 6092 16348
rect 6116 16346 6172 16348
rect 6196 16346 6252 16348
rect 5956 16294 5982 16346
rect 5982 16294 6012 16346
rect 6036 16294 6046 16346
rect 6046 16294 6092 16346
rect 6116 16294 6162 16346
rect 6162 16294 6172 16346
rect 6196 16294 6226 16346
rect 6226 16294 6252 16346
rect 5956 16292 6012 16294
rect 6036 16292 6092 16294
rect 6116 16292 6172 16294
rect 6196 16292 6252 16294
rect 4289 15802 4345 15804
rect 4369 15802 4425 15804
rect 4449 15802 4505 15804
rect 4529 15802 4585 15804
rect 4289 15750 4315 15802
rect 4315 15750 4345 15802
rect 4369 15750 4379 15802
rect 4379 15750 4425 15802
rect 4449 15750 4495 15802
rect 4495 15750 4505 15802
rect 4529 15750 4559 15802
rect 4559 15750 4585 15802
rect 4289 15748 4345 15750
rect 4369 15748 4425 15750
rect 4449 15748 4505 15750
rect 4529 15748 4585 15750
rect 5956 15258 6012 15260
rect 6036 15258 6092 15260
rect 6116 15258 6172 15260
rect 6196 15258 6252 15260
rect 5956 15206 5982 15258
rect 5982 15206 6012 15258
rect 6036 15206 6046 15258
rect 6046 15206 6092 15258
rect 6116 15206 6162 15258
rect 6162 15206 6172 15258
rect 6196 15206 6226 15258
rect 6226 15206 6252 15258
rect 5956 15204 6012 15206
rect 6036 15204 6092 15206
rect 6116 15204 6172 15206
rect 6196 15204 6252 15206
rect 4289 14714 4345 14716
rect 4369 14714 4425 14716
rect 4449 14714 4505 14716
rect 4529 14714 4585 14716
rect 4289 14662 4315 14714
rect 4315 14662 4345 14714
rect 4369 14662 4379 14714
rect 4379 14662 4425 14714
rect 4449 14662 4495 14714
rect 4495 14662 4505 14714
rect 4529 14662 4559 14714
rect 4559 14662 4585 14714
rect 4289 14660 4345 14662
rect 4369 14660 4425 14662
rect 4449 14660 4505 14662
rect 4529 14660 4585 14662
rect 5956 14170 6012 14172
rect 6036 14170 6092 14172
rect 6116 14170 6172 14172
rect 6196 14170 6252 14172
rect 5956 14118 5982 14170
rect 5982 14118 6012 14170
rect 6036 14118 6046 14170
rect 6046 14118 6092 14170
rect 6116 14118 6162 14170
rect 6162 14118 6172 14170
rect 6196 14118 6226 14170
rect 6226 14118 6252 14170
rect 5956 14116 6012 14118
rect 6036 14116 6092 14118
rect 6116 14116 6172 14118
rect 6196 14116 6252 14118
rect 4289 13626 4345 13628
rect 4369 13626 4425 13628
rect 4449 13626 4505 13628
rect 4529 13626 4585 13628
rect 4289 13574 4315 13626
rect 4315 13574 4345 13626
rect 4369 13574 4379 13626
rect 4379 13574 4425 13626
rect 4449 13574 4495 13626
rect 4495 13574 4505 13626
rect 4529 13574 4559 13626
rect 4559 13574 4585 13626
rect 4289 13572 4345 13574
rect 4369 13572 4425 13574
rect 4449 13572 4505 13574
rect 4529 13572 4585 13574
rect 5956 13082 6012 13084
rect 6036 13082 6092 13084
rect 6116 13082 6172 13084
rect 6196 13082 6252 13084
rect 5956 13030 5982 13082
rect 5982 13030 6012 13082
rect 6036 13030 6046 13082
rect 6046 13030 6092 13082
rect 6116 13030 6162 13082
rect 6162 13030 6172 13082
rect 6196 13030 6226 13082
rect 6226 13030 6252 13082
rect 5956 13028 6012 13030
rect 6036 13028 6092 13030
rect 6116 13028 6172 13030
rect 6196 13028 6252 13030
rect 4289 12538 4345 12540
rect 4369 12538 4425 12540
rect 4449 12538 4505 12540
rect 4529 12538 4585 12540
rect 4289 12486 4315 12538
rect 4315 12486 4345 12538
rect 4369 12486 4379 12538
rect 4379 12486 4425 12538
rect 4449 12486 4495 12538
rect 4495 12486 4505 12538
rect 4529 12486 4559 12538
rect 4559 12486 4585 12538
rect 4289 12484 4345 12486
rect 4369 12484 4425 12486
rect 4449 12484 4505 12486
rect 4529 12484 4585 12486
rect 5956 11994 6012 11996
rect 6036 11994 6092 11996
rect 6116 11994 6172 11996
rect 6196 11994 6252 11996
rect 5956 11942 5982 11994
rect 5982 11942 6012 11994
rect 6036 11942 6046 11994
rect 6046 11942 6092 11994
rect 6116 11942 6162 11994
rect 6162 11942 6172 11994
rect 6196 11942 6226 11994
rect 6226 11942 6252 11994
rect 5956 11940 6012 11942
rect 6036 11940 6092 11942
rect 6116 11940 6172 11942
rect 6196 11940 6252 11942
rect 4289 11450 4345 11452
rect 4369 11450 4425 11452
rect 4449 11450 4505 11452
rect 4529 11450 4585 11452
rect 4289 11398 4315 11450
rect 4315 11398 4345 11450
rect 4369 11398 4379 11450
rect 4379 11398 4425 11450
rect 4449 11398 4495 11450
rect 4495 11398 4505 11450
rect 4529 11398 4559 11450
rect 4559 11398 4585 11450
rect 4289 11396 4345 11398
rect 4369 11396 4425 11398
rect 4449 11396 4505 11398
rect 4529 11396 4585 11398
rect 5956 10906 6012 10908
rect 6036 10906 6092 10908
rect 6116 10906 6172 10908
rect 6196 10906 6252 10908
rect 5956 10854 5982 10906
rect 5982 10854 6012 10906
rect 6036 10854 6046 10906
rect 6046 10854 6092 10906
rect 6116 10854 6162 10906
rect 6162 10854 6172 10906
rect 6196 10854 6226 10906
rect 6226 10854 6252 10906
rect 5956 10852 6012 10854
rect 6036 10852 6092 10854
rect 6116 10852 6172 10854
rect 6196 10852 6252 10854
rect 4289 10362 4345 10364
rect 4369 10362 4425 10364
rect 4449 10362 4505 10364
rect 4529 10362 4585 10364
rect 4289 10310 4315 10362
rect 4315 10310 4345 10362
rect 4369 10310 4379 10362
rect 4379 10310 4425 10362
rect 4449 10310 4495 10362
rect 4495 10310 4505 10362
rect 4529 10310 4559 10362
rect 4559 10310 4585 10362
rect 4289 10308 4345 10310
rect 4369 10308 4425 10310
rect 4449 10308 4505 10310
rect 4529 10308 4585 10310
rect 5956 9818 6012 9820
rect 6036 9818 6092 9820
rect 6116 9818 6172 9820
rect 6196 9818 6252 9820
rect 5956 9766 5982 9818
rect 5982 9766 6012 9818
rect 6036 9766 6046 9818
rect 6046 9766 6092 9818
rect 6116 9766 6162 9818
rect 6162 9766 6172 9818
rect 6196 9766 6226 9818
rect 6226 9766 6252 9818
rect 5956 9764 6012 9766
rect 6036 9764 6092 9766
rect 6116 9764 6172 9766
rect 6196 9764 6252 9766
rect 4289 9274 4345 9276
rect 4369 9274 4425 9276
rect 4449 9274 4505 9276
rect 4529 9274 4585 9276
rect 4289 9222 4315 9274
rect 4315 9222 4345 9274
rect 4369 9222 4379 9274
rect 4379 9222 4425 9274
rect 4449 9222 4495 9274
rect 4495 9222 4505 9274
rect 4529 9222 4559 9274
rect 4559 9222 4585 9274
rect 4289 9220 4345 9222
rect 4369 9220 4425 9222
rect 4449 9220 4505 9222
rect 4529 9220 4585 9222
rect 5956 8730 6012 8732
rect 6036 8730 6092 8732
rect 6116 8730 6172 8732
rect 6196 8730 6252 8732
rect 5956 8678 5982 8730
rect 5982 8678 6012 8730
rect 6036 8678 6046 8730
rect 6046 8678 6092 8730
rect 6116 8678 6162 8730
rect 6162 8678 6172 8730
rect 6196 8678 6226 8730
rect 6226 8678 6252 8730
rect 5956 8676 6012 8678
rect 6036 8676 6092 8678
rect 6116 8676 6172 8678
rect 6196 8676 6252 8678
rect 4289 8186 4345 8188
rect 4369 8186 4425 8188
rect 4449 8186 4505 8188
rect 4529 8186 4585 8188
rect 4289 8134 4315 8186
rect 4315 8134 4345 8186
rect 4369 8134 4379 8186
rect 4379 8134 4425 8186
rect 4449 8134 4495 8186
rect 4495 8134 4505 8186
rect 4529 8134 4559 8186
rect 4559 8134 4585 8186
rect 4289 8132 4345 8134
rect 4369 8132 4425 8134
rect 4449 8132 4505 8134
rect 4529 8132 4585 8134
rect 5956 7642 6012 7644
rect 6036 7642 6092 7644
rect 6116 7642 6172 7644
rect 6196 7642 6252 7644
rect 5956 7590 5982 7642
rect 5982 7590 6012 7642
rect 6036 7590 6046 7642
rect 6046 7590 6092 7642
rect 6116 7590 6162 7642
rect 6162 7590 6172 7642
rect 6196 7590 6226 7642
rect 6226 7590 6252 7642
rect 5956 7588 6012 7590
rect 6036 7588 6092 7590
rect 6116 7588 6172 7590
rect 6196 7588 6252 7590
rect 4289 7098 4345 7100
rect 4369 7098 4425 7100
rect 4449 7098 4505 7100
rect 4529 7098 4585 7100
rect 4289 7046 4315 7098
rect 4315 7046 4345 7098
rect 4369 7046 4379 7098
rect 4379 7046 4425 7098
rect 4449 7046 4495 7098
rect 4495 7046 4505 7098
rect 4529 7046 4559 7098
rect 4559 7046 4585 7098
rect 4289 7044 4345 7046
rect 4369 7044 4425 7046
rect 4449 7044 4505 7046
rect 4529 7044 4585 7046
rect 5956 6554 6012 6556
rect 6036 6554 6092 6556
rect 6116 6554 6172 6556
rect 6196 6554 6252 6556
rect 5956 6502 5982 6554
rect 5982 6502 6012 6554
rect 6036 6502 6046 6554
rect 6046 6502 6092 6554
rect 6116 6502 6162 6554
rect 6162 6502 6172 6554
rect 6196 6502 6226 6554
rect 6226 6502 6252 6554
rect 5956 6500 6012 6502
rect 6036 6500 6092 6502
rect 6116 6500 6172 6502
rect 6196 6500 6252 6502
rect 4289 6010 4345 6012
rect 4369 6010 4425 6012
rect 4449 6010 4505 6012
rect 4529 6010 4585 6012
rect 4289 5958 4315 6010
rect 4315 5958 4345 6010
rect 4369 5958 4379 6010
rect 4379 5958 4425 6010
rect 4449 5958 4495 6010
rect 4495 5958 4505 6010
rect 4529 5958 4559 6010
rect 4559 5958 4585 6010
rect 4289 5956 4345 5958
rect 4369 5956 4425 5958
rect 4449 5956 4505 5958
rect 4529 5956 4585 5958
rect 5956 5466 6012 5468
rect 6036 5466 6092 5468
rect 6116 5466 6172 5468
rect 6196 5466 6252 5468
rect 5956 5414 5982 5466
rect 5982 5414 6012 5466
rect 6036 5414 6046 5466
rect 6046 5414 6092 5466
rect 6116 5414 6162 5466
rect 6162 5414 6172 5466
rect 6196 5414 6226 5466
rect 6226 5414 6252 5466
rect 5956 5412 6012 5414
rect 6036 5412 6092 5414
rect 6116 5412 6172 5414
rect 6196 5412 6252 5414
rect 4289 4922 4345 4924
rect 4369 4922 4425 4924
rect 4449 4922 4505 4924
rect 4529 4922 4585 4924
rect 4289 4870 4315 4922
rect 4315 4870 4345 4922
rect 4369 4870 4379 4922
rect 4379 4870 4425 4922
rect 4449 4870 4495 4922
rect 4495 4870 4505 4922
rect 4529 4870 4559 4922
rect 4559 4870 4585 4922
rect 4289 4868 4345 4870
rect 4369 4868 4425 4870
rect 4449 4868 4505 4870
rect 4529 4868 4585 4870
rect 5956 4378 6012 4380
rect 6036 4378 6092 4380
rect 6116 4378 6172 4380
rect 6196 4378 6252 4380
rect 5956 4326 5982 4378
rect 5982 4326 6012 4378
rect 6036 4326 6046 4378
rect 6046 4326 6092 4378
rect 6116 4326 6162 4378
rect 6162 4326 6172 4378
rect 6196 4326 6226 4378
rect 6226 4326 6252 4378
rect 5956 4324 6012 4326
rect 6036 4324 6092 4326
rect 6116 4324 6172 4326
rect 6196 4324 6252 4326
rect 7622 157242 7678 157244
rect 7702 157242 7758 157244
rect 7782 157242 7838 157244
rect 7862 157242 7918 157244
rect 7622 157190 7648 157242
rect 7648 157190 7678 157242
rect 7702 157190 7712 157242
rect 7712 157190 7758 157242
rect 7782 157190 7828 157242
rect 7828 157190 7838 157242
rect 7862 157190 7892 157242
rect 7892 157190 7918 157242
rect 7622 157188 7678 157190
rect 7702 157188 7758 157190
rect 7782 157188 7838 157190
rect 7862 157188 7918 157190
rect 7622 156154 7678 156156
rect 7702 156154 7758 156156
rect 7782 156154 7838 156156
rect 7862 156154 7918 156156
rect 7622 156102 7648 156154
rect 7648 156102 7678 156154
rect 7702 156102 7712 156154
rect 7712 156102 7758 156154
rect 7782 156102 7828 156154
rect 7828 156102 7838 156154
rect 7862 156102 7892 156154
rect 7892 156102 7918 156154
rect 7622 156100 7678 156102
rect 7702 156100 7758 156102
rect 7782 156100 7838 156102
rect 7862 156100 7918 156102
rect 7622 155066 7678 155068
rect 7702 155066 7758 155068
rect 7782 155066 7838 155068
rect 7862 155066 7918 155068
rect 7622 155014 7648 155066
rect 7648 155014 7678 155066
rect 7702 155014 7712 155066
rect 7712 155014 7758 155066
rect 7782 155014 7828 155066
rect 7828 155014 7838 155066
rect 7862 155014 7892 155066
rect 7892 155014 7918 155066
rect 7622 155012 7678 155014
rect 7702 155012 7758 155014
rect 7782 155012 7838 155014
rect 7862 155012 7918 155014
rect 7622 153978 7678 153980
rect 7702 153978 7758 153980
rect 7782 153978 7838 153980
rect 7862 153978 7918 153980
rect 7622 153926 7648 153978
rect 7648 153926 7678 153978
rect 7702 153926 7712 153978
rect 7712 153926 7758 153978
rect 7782 153926 7828 153978
rect 7828 153926 7838 153978
rect 7862 153926 7892 153978
rect 7892 153926 7918 153978
rect 7622 153924 7678 153926
rect 7702 153924 7758 153926
rect 7782 153924 7838 153926
rect 7862 153924 7918 153926
rect 7622 152890 7678 152892
rect 7702 152890 7758 152892
rect 7782 152890 7838 152892
rect 7862 152890 7918 152892
rect 7622 152838 7648 152890
rect 7648 152838 7678 152890
rect 7702 152838 7712 152890
rect 7712 152838 7758 152890
rect 7782 152838 7828 152890
rect 7828 152838 7838 152890
rect 7862 152838 7892 152890
rect 7892 152838 7918 152890
rect 7622 152836 7678 152838
rect 7702 152836 7758 152838
rect 7782 152836 7838 152838
rect 7862 152836 7918 152838
rect 7622 151802 7678 151804
rect 7702 151802 7758 151804
rect 7782 151802 7838 151804
rect 7862 151802 7918 151804
rect 7622 151750 7648 151802
rect 7648 151750 7678 151802
rect 7702 151750 7712 151802
rect 7712 151750 7758 151802
rect 7782 151750 7828 151802
rect 7828 151750 7838 151802
rect 7862 151750 7892 151802
rect 7892 151750 7918 151802
rect 7622 151748 7678 151750
rect 7702 151748 7758 151750
rect 7782 151748 7838 151750
rect 7862 151748 7918 151750
rect 7622 150714 7678 150716
rect 7702 150714 7758 150716
rect 7782 150714 7838 150716
rect 7862 150714 7918 150716
rect 7622 150662 7648 150714
rect 7648 150662 7678 150714
rect 7702 150662 7712 150714
rect 7712 150662 7758 150714
rect 7782 150662 7828 150714
rect 7828 150662 7838 150714
rect 7862 150662 7892 150714
rect 7892 150662 7918 150714
rect 7622 150660 7678 150662
rect 7702 150660 7758 150662
rect 7782 150660 7838 150662
rect 7862 150660 7918 150662
rect 7622 149626 7678 149628
rect 7702 149626 7758 149628
rect 7782 149626 7838 149628
rect 7862 149626 7918 149628
rect 7622 149574 7648 149626
rect 7648 149574 7678 149626
rect 7702 149574 7712 149626
rect 7712 149574 7758 149626
rect 7782 149574 7828 149626
rect 7828 149574 7838 149626
rect 7862 149574 7892 149626
rect 7892 149574 7918 149626
rect 7622 149572 7678 149574
rect 7702 149572 7758 149574
rect 7782 149572 7838 149574
rect 7862 149572 7918 149574
rect 7622 148538 7678 148540
rect 7702 148538 7758 148540
rect 7782 148538 7838 148540
rect 7862 148538 7918 148540
rect 7622 148486 7648 148538
rect 7648 148486 7678 148538
rect 7702 148486 7712 148538
rect 7712 148486 7758 148538
rect 7782 148486 7828 148538
rect 7828 148486 7838 148538
rect 7862 148486 7892 148538
rect 7892 148486 7918 148538
rect 7622 148484 7678 148486
rect 7702 148484 7758 148486
rect 7782 148484 7838 148486
rect 7862 148484 7918 148486
rect 7622 147450 7678 147452
rect 7702 147450 7758 147452
rect 7782 147450 7838 147452
rect 7862 147450 7918 147452
rect 7622 147398 7648 147450
rect 7648 147398 7678 147450
rect 7702 147398 7712 147450
rect 7712 147398 7758 147450
rect 7782 147398 7828 147450
rect 7828 147398 7838 147450
rect 7862 147398 7892 147450
rect 7892 147398 7918 147450
rect 7622 147396 7678 147398
rect 7702 147396 7758 147398
rect 7782 147396 7838 147398
rect 7862 147396 7918 147398
rect 7622 146362 7678 146364
rect 7702 146362 7758 146364
rect 7782 146362 7838 146364
rect 7862 146362 7918 146364
rect 7622 146310 7648 146362
rect 7648 146310 7678 146362
rect 7702 146310 7712 146362
rect 7712 146310 7758 146362
rect 7782 146310 7828 146362
rect 7828 146310 7838 146362
rect 7862 146310 7892 146362
rect 7892 146310 7918 146362
rect 7622 146308 7678 146310
rect 7702 146308 7758 146310
rect 7782 146308 7838 146310
rect 7862 146308 7918 146310
rect 7622 145274 7678 145276
rect 7702 145274 7758 145276
rect 7782 145274 7838 145276
rect 7862 145274 7918 145276
rect 7622 145222 7648 145274
rect 7648 145222 7678 145274
rect 7702 145222 7712 145274
rect 7712 145222 7758 145274
rect 7782 145222 7828 145274
rect 7828 145222 7838 145274
rect 7862 145222 7892 145274
rect 7892 145222 7918 145274
rect 7622 145220 7678 145222
rect 7702 145220 7758 145222
rect 7782 145220 7838 145222
rect 7862 145220 7918 145222
rect 7622 144186 7678 144188
rect 7702 144186 7758 144188
rect 7782 144186 7838 144188
rect 7862 144186 7918 144188
rect 7622 144134 7648 144186
rect 7648 144134 7678 144186
rect 7702 144134 7712 144186
rect 7712 144134 7758 144186
rect 7782 144134 7828 144186
rect 7828 144134 7838 144186
rect 7862 144134 7892 144186
rect 7892 144134 7918 144186
rect 7622 144132 7678 144134
rect 7702 144132 7758 144134
rect 7782 144132 7838 144134
rect 7862 144132 7918 144134
rect 7622 143098 7678 143100
rect 7702 143098 7758 143100
rect 7782 143098 7838 143100
rect 7862 143098 7918 143100
rect 7622 143046 7648 143098
rect 7648 143046 7678 143098
rect 7702 143046 7712 143098
rect 7712 143046 7758 143098
rect 7782 143046 7828 143098
rect 7828 143046 7838 143098
rect 7862 143046 7892 143098
rect 7892 143046 7918 143098
rect 7622 143044 7678 143046
rect 7702 143044 7758 143046
rect 7782 143044 7838 143046
rect 7862 143044 7918 143046
rect 7622 142010 7678 142012
rect 7702 142010 7758 142012
rect 7782 142010 7838 142012
rect 7862 142010 7918 142012
rect 7622 141958 7648 142010
rect 7648 141958 7678 142010
rect 7702 141958 7712 142010
rect 7712 141958 7758 142010
rect 7782 141958 7828 142010
rect 7828 141958 7838 142010
rect 7862 141958 7892 142010
rect 7892 141958 7918 142010
rect 7622 141956 7678 141958
rect 7702 141956 7758 141958
rect 7782 141956 7838 141958
rect 7862 141956 7918 141958
rect 7622 140922 7678 140924
rect 7702 140922 7758 140924
rect 7782 140922 7838 140924
rect 7862 140922 7918 140924
rect 7622 140870 7648 140922
rect 7648 140870 7678 140922
rect 7702 140870 7712 140922
rect 7712 140870 7758 140922
rect 7782 140870 7828 140922
rect 7828 140870 7838 140922
rect 7862 140870 7892 140922
rect 7892 140870 7918 140922
rect 7622 140868 7678 140870
rect 7702 140868 7758 140870
rect 7782 140868 7838 140870
rect 7862 140868 7918 140870
rect 7622 139834 7678 139836
rect 7702 139834 7758 139836
rect 7782 139834 7838 139836
rect 7862 139834 7918 139836
rect 7622 139782 7648 139834
rect 7648 139782 7678 139834
rect 7702 139782 7712 139834
rect 7712 139782 7758 139834
rect 7782 139782 7828 139834
rect 7828 139782 7838 139834
rect 7862 139782 7892 139834
rect 7892 139782 7918 139834
rect 7622 139780 7678 139782
rect 7702 139780 7758 139782
rect 7782 139780 7838 139782
rect 7862 139780 7918 139782
rect 7622 138746 7678 138748
rect 7702 138746 7758 138748
rect 7782 138746 7838 138748
rect 7862 138746 7918 138748
rect 7622 138694 7648 138746
rect 7648 138694 7678 138746
rect 7702 138694 7712 138746
rect 7712 138694 7758 138746
rect 7782 138694 7828 138746
rect 7828 138694 7838 138746
rect 7862 138694 7892 138746
rect 7892 138694 7918 138746
rect 7622 138692 7678 138694
rect 7702 138692 7758 138694
rect 7782 138692 7838 138694
rect 7862 138692 7918 138694
rect 7622 137658 7678 137660
rect 7702 137658 7758 137660
rect 7782 137658 7838 137660
rect 7862 137658 7918 137660
rect 7622 137606 7648 137658
rect 7648 137606 7678 137658
rect 7702 137606 7712 137658
rect 7712 137606 7758 137658
rect 7782 137606 7828 137658
rect 7828 137606 7838 137658
rect 7862 137606 7892 137658
rect 7892 137606 7918 137658
rect 7622 137604 7678 137606
rect 7702 137604 7758 137606
rect 7782 137604 7838 137606
rect 7862 137604 7918 137606
rect 7622 136570 7678 136572
rect 7702 136570 7758 136572
rect 7782 136570 7838 136572
rect 7862 136570 7918 136572
rect 7622 136518 7648 136570
rect 7648 136518 7678 136570
rect 7702 136518 7712 136570
rect 7712 136518 7758 136570
rect 7782 136518 7828 136570
rect 7828 136518 7838 136570
rect 7862 136518 7892 136570
rect 7892 136518 7918 136570
rect 7622 136516 7678 136518
rect 7702 136516 7758 136518
rect 7782 136516 7838 136518
rect 7862 136516 7918 136518
rect 7622 135482 7678 135484
rect 7702 135482 7758 135484
rect 7782 135482 7838 135484
rect 7862 135482 7918 135484
rect 7622 135430 7648 135482
rect 7648 135430 7678 135482
rect 7702 135430 7712 135482
rect 7712 135430 7758 135482
rect 7782 135430 7828 135482
rect 7828 135430 7838 135482
rect 7862 135430 7892 135482
rect 7892 135430 7918 135482
rect 7622 135428 7678 135430
rect 7702 135428 7758 135430
rect 7782 135428 7838 135430
rect 7862 135428 7918 135430
rect 7622 134394 7678 134396
rect 7702 134394 7758 134396
rect 7782 134394 7838 134396
rect 7862 134394 7918 134396
rect 7622 134342 7648 134394
rect 7648 134342 7678 134394
rect 7702 134342 7712 134394
rect 7712 134342 7758 134394
rect 7782 134342 7828 134394
rect 7828 134342 7838 134394
rect 7862 134342 7892 134394
rect 7892 134342 7918 134394
rect 7622 134340 7678 134342
rect 7702 134340 7758 134342
rect 7782 134340 7838 134342
rect 7862 134340 7918 134342
rect 7622 133306 7678 133308
rect 7702 133306 7758 133308
rect 7782 133306 7838 133308
rect 7862 133306 7918 133308
rect 7622 133254 7648 133306
rect 7648 133254 7678 133306
rect 7702 133254 7712 133306
rect 7712 133254 7758 133306
rect 7782 133254 7828 133306
rect 7828 133254 7838 133306
rect 7862 133254 7892 133306
rect 7892 133254 7918 133306
rect 7622 133252 7678 133254
rect 7702 133252 7758 133254
rect 7782 133252 7838 133254
rect 7862 133252 7918 133254
rect 7622 132218 7678 132220
rect 7702 132218 7758 132220
rect 7782 132218 7838 132220
rect 7862 132218 7918 132220
rect 7622 132166 7648 132218
rect 7648 132166 7678 132218
rect 7702 132166 7712 132218
rect 7712 132166 7758 132218
rect 7782 132166 7828 132218
rect 7828 132166 7838 132218
rect 7862 132166 7892 132218
rect 7892 132166 7918 132218
rect 7622 132164 7678 132166
rect 7702 132164 7758 132166
rect 7782 132164 7838 132166
rect 7862 132164 7918 132166
rect 7622 131130 7678 131132
rect 7702 131130 7758 131132
rect 7782 131130 7838 131132
rect 7862 131130 7918 131132
rect 7622 131078 7648 131130
rect 7648 131078 7678 131130
rect 7702 131078 7712 131130
rect 7712 131078 7758 131130
rect 7782 131078 7828 131130
rect 7828 131078 7838 131130
rect 7862 131078 7892 131130
rect 7892 131078 7918 131130
rect 7622 131076 7678 131078
rect 7702 131076 7758 131078
rect 7782 131076 7838 131078
rect 7862 131076 7918 131078
rect 7622 130042 7678 130044
rect 7702 130042 7758 130044
rect 7782 130042 7838 130044
rect 7862 130042 7918 130044
rect 7622 129990 7648 130042
rect 7648 129990 7678 130042
rect 7702 129990 7712 130042
rect 7712 129990 7758 130042
rect 7782 129990 7828 130042
rect 7828 129990 7838 130042
rect 7862 129990 7892 130042
rect 7892 129990 7918 130042
rect 7622 129988 7678 129990
rect 7702 129988 7758 129990
rect 7782 129988 7838 129990
rect 7862 129988 7918 129990
rect 7622 128954 7678 128956
rect 7702 128954 7758 128956
rect 7782 128954 7838 128956
rect 7862 128954 7918 128956
rect 7622 128902 7648 128954
rect 7648 128902 7678 128954
rect 7702 128902 7712 128954
rect 7712 128902 7758 128954
rect 7782 128902 7828 128954
rect 7828 128902 7838 128954
rect 7862 128902 7892 128954
rect 7892 128902 7918 128954
rect 7622 128900 7678 128902
rect 7702 128900 7758 128902
rect 7782 128900 7838 128902
rect 7862 128900 7918 128902
rect 7622 127866 7678 127868
rect 7702 127866 7758 127868
rect 7782 127866 7838 127868
rect 7862 127866 7918 127868
rect 7622 127814 7648 127866
rect 7648 127814 7678 127866
rect 7702 127814 7712 127866
rect 7712 127814 7758 127866
rect 7782 127814 7828 127866
rect 7828 127814 7838 127866
rect 7862 127814 7892 127866
rect 7892 127814 7918 127866
rect 7622 127812 7678 127814
rect 7702 127812 7758 127814
rect 7782 127812 7838 127814
rect 7862 127812 7918 127814
rect 7622 126778 7678 126780
rect 7702 126778 7758 126780
rect 7782 126778 7838 126780
rect 7862 126778 7918 126780
rect 7622 126726 7648 126778
rect 7648 126726 7678 126778
rect 7702 126726 7712 126778
rect 7712 126726 7758 126778
rect 7782 126726 7828 126778
rect 7828 126726 7838 126778
rect 7862 126726 7892 126778
rect 7892 126726 7918 126778
rect 7622 126724 7678 126726
rect 7702 126724 7758 126726
rect 7782 126724 7838 126726
rect 7862 126724 7918 126726
rect 7622 125690 7678 125692
rect 7702 125690 7758 125692
rect 7782 125690 7838 125692
rect 7862 125690 7918 125692
rect 7622 125638 7648 125690
rect 7648 125638 7678 125690
rect 7702 125638 7712 125690
rect 7712 125638 7758 125690
rect 7782 125638 7828 125690
rect 7828 125638 7838 125690
rect 7862 125638 7892 125690
rect 7892 125638 7918 125690
rect 7622 125636 7678 125638
rect 7702 125636 7758 125638
rect 7782 125636 7838 125638
rect 7862 125636 7918 125638
rect 7622 124602 7678 124604
rect 7702 124602 7758 124604
rect 7782 124602 7838 124604
rect 7862 124602 7918 124604
rect 7622 124550 7648 124602
rect 7648 124550 7678 124602
rect 7702 124550 7712 124602
rect 7712 124550 7758 124602
rect 7782 124550 7828 124602
rect 7828 124550 7838 124602
rect 7862 124550 7892 124602
rect 7892 124550 7918 124602
rect 7622 124548 7678 124550
rect 7702 124548 7758 124550
rect 7782 124548 7838 124550
rect 7862 124548 7918 124550
rect 7622 123514 7678 123516
rect 7702 123514 7758 123516
rect 7782 123514 7838 123516
rect 7862 123514 7918 123516
rect 7622 123462 7648 123514
rect 7648 123462 7678 123514
rect 7702 123462 7712 123514
rect 7712 123462 7758 123514
rect 7782 123462 7828 123514
rect 7828 123462 7838 123514
rect 7862 123462 7892 123514
rect 7892 123462 7918 123514
rect 7622 123460 7678 123462
rect 7702 123460 7758 123462
rect 7782 123460 7838 123462
rect 7862 123460 7918 123462
rect 7622 122426 7678 122428
rect 7702 122426 7758 122428
rect 7782 122426 7838 122428
rect 7862 122426 7918 122428
rect 7622 122374 7648 122426
rect 7648 122374 7678 122426
rect 7702 122374 7712 122426
rect 7712 122374 7758 122426
rect 7782 122374 7828 122426
rect 7828 122374 7838 122426
rect 7862 122374 7892 122426
rect 7892 122374 7918 122426
rect 7622 122372 7678 122374
rect 7702 122372 7758 122374
rect 7782 122372 7838 122374
rect 7862 122372 7918 122374
rect 7622 121338 7678 121340
rect 7702 121338 7758 121340
rect 7782 121338 7838 121340
rect 7862 121338 7918 121340
rect 7622 121286 7648 121338
rect 7648 121286 7678 121338
rect 7702 121286 7712 121338
rect 7712 121286 7758 121338
rect 7782 121286 7828 121338
rect 7828 121286 7838 121338
rect 7862 121286 7892 121338
rect 7892 121286 7918 121338
rect 7622 121284 7678 121286
rect 7702 121284 7758 121286
rect 7782 121284 7838 121286
rect 7862 121284 7918 121286
rect 7622 120250 7678 120252
rect 7702 120250 7758 120252
rect 7782 120250 7838 120252
rect 7862 120250 7918 120252
rect 7622 120198 7648 120250
rect 7648 120198 7678 120250
rect 7702 120198 7712 120250
rect 7712 120198 7758 120250
rect 7782 120198 7828 120250
rect 7828 120198 7838 120250
rect 7862 120198 7892 120250
rect 7892 120198 7918 120250
rect 7622 120196 7678 120198
rect 7702 120196 7758 120198
rect 7782 120196 7838 120198
rect 7862 120196 7918 120198
rect 7622 119162 7678 119164
rect 7702 119162 7758 119164
rect 7782 119162 7838 119164
rect 7862 119162 7918 119164
rect 7622 119110 7648 119162
rect 7648 119110 7678 119162
rect 7702 119110 7712 119162
rect 7712 119110 7758 119162
rect 7782 119110 7828 119162
rect 7828 119110 7838 119162
rect 7862 119110 7892 119162
rect 7892 119110 7918 119162
rect 7622 119108 7678 119110
rect 7702 119108 7758 119110
rect 7782 119108 7838 119110
rect 7862 119108 7918 119110
rect 7622 118074 7678 118076
rect 7702 118074 7758 118076
rect 7782 118074 7838 118076
rect 7862 118074 7918 118076
rect 7622 118022 7648 118074
rect 7648 118022 7678 118074
rect 7702 118022 7712 118074
rect 7712 118022 7758 118074
rect 7782 118022 7828 118074
rect 7828 118022 7838 118074
rect 7862 118022 7892 118074
rect 7892 118022 7918 118074
rect 7622 118020 7678 118022
rect 7702 118020 7758 118022
rect 7782 118020 7838 118022
rect 7862 118020 7918 118022
rect 7622 116986 7678 116988
rect 7702 116986 7758 116988
rect 7782 116986 7838 116988
rect 7862 116986 7918 116988
rect 7622 116934 7648 116986
rect 7648 116934 7678 116986
rect 7702 116934 7712 116986
rect 7712 116934 7758 116986
rect 7782 116934 7828 116986
rect 7828 116934 7838 116986
rect 7862 116934 7892 116986
rect 7892 116934 7918 116986
rect 7622 116932 7678 116934
rect 7702 116932 7758 116934
rect 7782 116932 7838 116934
rect 7862 116932 7918 116934
rect 7622 115898 7678 115900
rect 7702 115898 7758 115900
rect 7782 115898 7838 115900
rect 7862 115898 7918 115900
rect 7622 115846 7648 115898
rect 7648 115846 7678 115898
rect 7702 115846 7712 115898
rect 7712 115846 7758 115898
rect 7782 115846 7828 115898
rect 7828 115846 7838 115898
rect 7862 115846 7892 115898
rect 7892 115846 7918 115898
rect 7622 115844 7678 115846
rect 7702 115844 7758 115846
rect 7782 115844 7838 115846
rect 7862 115844 7918 115846
rect 7622 114810 7678 114812
rect 7702 114810 7758 114812
rect 7782 114810 7838 114812
rect 7862 114810 7918 114812
rect 7622 114758 7648 114810
rect 7648 114758 7678 114810
rect 7702 114758 7712 114810
rect 7712 114758 7758 114810
rect 7782 114758 7828 114810
rect 7828 114758 7838 114810
rect 7862 114758 7892 114810
rect 7892 114758 7918 114810
rect 7622 114756 7678 114758
rect 7702 114756 7758 114758
rect 7782 114756 7838 114758
rect 7862 114756 7918 114758
rect 7622 113722 7678 113724
rect 7702 113722 7758 113724
rect 7782 113722 7838 113724
rect 7862 113722 7918 113724
rect 7622 113670 7648 113722
rect 7648 113670 7678 113722
rect 7702 113670 7712 113722
rect 7712 113670 7758 113722
rect 7782 113670 7828 113722
rect 7828 113670 7838 113722
rect 7862 113670 7892 113722
rect 7892 113670 7918 113722
rect 7622 113668 7678 113670
rect 7702 113668 7758 113670
rect 7782 113668 7838 113670
rect 7862 113668 7918 113670
rect 7622 112634 7678 112636
rect 7702 112634 7758 112636
rect 7782 112634 7838 112636
rect 7862 112634 7918 112636
rect 7622 112582 7648 112634
rect 7648 112582 7678 112634
rect 7702 112582 7712 112634
rect 7712 112582 7758 112634
rect 7782 112582 7828 112634
rect 7828 112582 7838 112634
rect 7862 112582 7892 112634
rect 7892 112582 7918 112634
rect 7622 112580 7678 112582
rect 7702 112580 7758 112582
rect 7782 112580 7838 112582
rect 7862 112580 7918 112582
rect 7622 111546 7678 111548
rect 7702 111546 7758 111548
rect 7782 111546 7838 111548
rect 7862 111546 7918 111548
rect 7622 111494 7648 111546
rect 7648 111494 7678 111546
rect 7702 111494 7712 111546
rect 7712 111494 7758 111546
rect 7782 111494 7828 111546
rect 7828 111494 7838 111546
rect 7862 111494 7892 111546
rect 7892 111494 7918 111546
rect 7622 111492 7678 111494
rect 7702 111492 7758 111494
rect 7782 111492 7838 111494
rect 7862 111492 7918 111494
rect 7622 110458 7678 110460
rect 7702 110458 7758 110460
rect 7782 110458 7838 110460
rect 7862 110458 7918 110460
rect 7622 110406 7648 110458
rect 7648 110406 7678 110458
rect 7702 110406 7712 110458
rect 7712 110406 7758 110458
rect 7782 110406 7828 110458
rect 7828 110406 7838 110458
rect 7862 110406 7892 110458
rect 7892 110406 7918 110458
rect 7622 110404 7678 110406
rect 7702 110404 7758 110406
rect 7782 110404 7838 110406
rect 7862 110404 7918 110406
rect 7622 109370 7678 109372
rect 7702 109370 7758 109372
rect 7782 109370 7838 109372
rect 7862 109370 7918 109372
rect 7622 109318 7648 109370
rect 7648 109318 7678 109370
rect 7702 109318 7712 109370
rect 7712 109318 7758 109370
rect 7782 109318 7828 109370
rect 7828 109318 7838 109370
rect 7862 109318 7892 109370
rect 7892 109318 7918 109370
rect 7622 109316 7678 109318
rect 7702 109316 7758 109318
rect 7782 109316 7838 109318
rect 7862 109316 7918 109318
rect 7622 108282 7678 108284
rect 7702 108282 7758 108284
rect 7782 108282 7838 108284
rect 7862 108282 7918 108284
rect 7622 108230 7648 108282
rect 7648 108230 7678 108282
rect 7702 108230 7712 108282
rect 7712 108230 7758 108282
rect 7782 108230 7828 108282
rect 7828 108230 7838 108282
rect 7862 108230 7892 108282
rect 7892 108230 7918 108282
rect 7622 108228 7678 108230
rect 7702 108228 7758 108230
rect 7782 108228 7838 108230
rect 7862 108228 7918 108230
rect 7622 107194 7678 107196
rect 7702 107194 7758 107196
rect 7782 107194 7838 107196
rect 7862 107194 7918 107196
rect 7622 107142 7648 107194
rect 7648 107142 7678 107194
rect 7702 107142 7712 107194
rect 7712 107142 7758 107194
rect 7782 107142 7828 107194
rect 7828 107142 7838 107194
rect 7862 107142 7892 107194
rect 7892 107142 7918 107194
rect 7622 107140 7678 107142
rect 7702 107140 7758 107142
rect 7782 107140 7838 107142
rect 7862 107140 7918 107142
rect 7622 106106 7678 106108
rect 7702 106106 7758 106108
rect 7782 106106 7838 106108
rect 7862 106106 7918 106108
rect 7622 106054 7648 106106
rect 7648 106054 7678 106106
rect 7702 106054 7712 106106
rect 7712 106054 7758 106106
rect 7782 106054 7828 106106
rect 7828 106054 7838 106106
rect 7862 106054 7892 106106
rect 7892 106054 7918 106106
rect 7622 106052 7678 106054
rect 7702 106052 7758 106054
rect 7782 106052 7838 106054
rect 7862 106052 7918 106054
rect 7622 105018 7678 105020
rect 7702 105018 7758 105020
rect 7782 105018 7838 105020
rect 7862 105018 7918 105020
rect 7622 104966 7648 105018
rect 7648 104966 7678 105018
rect 7702 104966 7712 105018
rect 7712 104966 7758 105018
rect 7782 104966 7828 105018
rect 7828 104966 7838 105018
rect 7862 104966 7892 105018
rect 7892 104966 7918 105018
rect 7622 104964 7678 104966
rect 7702 104964 7758 104966
rect 7782 104964 7838 104966
rect 7862 104964 7918 104966
rect 7622 103930 7678 103932
rect 7702 103930 7758 103932
rect 7782 103930 7838 103932
rect 7862 103930 7918 103932
rect 7622 103878 7648 103930
rect 7648 103878 7678 103930
rect 7702 103878 7712 103930
rect 7712 103878 7758 103930
rect 7782 103878 7828 103930
rect 7828 103878 7838 103930
rect 7862 103878 7892 103930
rect 7892 103878 7918 103930
rect 7622 103876 7678 103878
rect 7702 103876 7758 103878
rect 7782 103876 7838 103878
rect 7862 103876 7918 103878
rect 7622 102842 7678 102844
rect 7702 102842 7758 102844
rect 7782 102842 7838 102844
rect 7862 102842 7918 102844
rect 7622 102790 7648 102842
rect 7648 102790 7678 102842
rect 7702 102790 7712 102842
rect 7712 102790 7758 102842
rect 7782 102790 7828 102842
rect 7828 102790 7838 102842
rect 7862 102790 7892 102842
rect 7892 102790 7918 102842
rect 7622 102788 7678 102790
rect 7702 102788 7758 102790
rect 7782 102788 7838 102790
rect 7862 102788 7918 102790
rect 7622 101754 7678 101756
rect 7702 101754 7758 101756
rect 7782 101754 7838 101756
rect 7862 101754 7918 101756
rect 7622 101702 7648 101754
rect 7648 101702 7678 101754
rect 7702 101702 7712 101754
rect 7712 101702 7758 101754
rect 7782 101702 7828 101754
rect 7828 101702 7838 101754
rect 7862 101702 7892 101754
rect 7892 101702 7918 101754
rect 7622 101700 7678 101702
rect 7702 101700 7758 101702
rect 7782 101700 7838 101702
rect 7862 101700 7918 101702
rect 7622 100666 7678 100668
rect 7702 100666 7758 100668
rect 7782 100666 7838 100668
rect 7862 100666 7918 100668
rect 7622 100614 7648 100666
rect 7648 100614 7678 100666
rect 7702 100614 7712 100666
rect 7712 100614 7758 100666
rect 7782 100614 7828 100666
rect 7828 100614 7838 100666
rect 7862 100614 7892 100666
rect 7892 100614 7918 100666
rect 7622 100612 7678 100614
rect 7702 100612 7758 100614
rect 7782 100612 7838 100614
rect 7862 100612 7918 100614
rect 7622 99578 7678 99580
rect 7702 99578 7758 99580
rect 7782 99578 7838 99580
rect 7862 99578 7918 99580
rect 7622 99526 7648 99578
rect 7648 99526 7678 99578
rect 7702 99526 7712 99578
rect 7712 99526 7758 99578
rect 7782 99526 7828 99578
rect 7828 99526 7838 99578
rect 7862 99526 7892 99578
rect 7892 99526 7918 99578
rect 7622 99524 7678 99526
rect 7702 99524 7758 99526
rect 7782 99524 7838 99526
rect 7862 99524 7918 99526
rect 7622 98490 7678 98492
rect 7702 98490 7758 98492
rect 7782 98490 7838 98492
rect 7862 98490 7918 98492
rect 7622 98438 7648 98490
rect 7648 98438 7678 98490
rect 7702 98438 7712 98490
rect 7712 98438 7758 98490
rect 7782 98438 7828 98490
rect 7828 98438 7838 98490
rect 7862 98438 7892 98490
rect 7892 98438 7918 98490
rect 7622 98436 7678 98438
rect 7702 98436 7758 98438
rect 7782 98436 7838 98438
rect 7862 98436 7918 98438
rect 7622 97402 7678 97404
rect 7702 97402 7758 97404
rect 7782 97402 7838 97404
rect 7862 97402 7918 97404
rect 7622 97350 7648 97402
rect 7648 97350 7678 97402
rect 7702 97350 7712 97402
rect 7712 97350 7758 97402
rect 7782 97350 7828 97402
rect 7828 97350 7838 97402
rect 7862 97350 7892 97402
rect 7892 97350 7918 97402
rect 7622 97348 7678 97350
rect 7702 97348 7758 97350
rect 7782 97348 7838 97350
rect 7862 97348 7918 97350
rect 7622 96314 7678 96316
rect 7702 96314 7758 96316
rect 7782 96314 7838 96316
rect 7862 96314 7918 96316
rect 7622 96262 7648 96314
rect 7648 96262 7678 96314
rect 7702 96262 7712 96314
rect 7712 96262 7758 96314
rect 7782 96262 7828 96314
rect 7828 96262 7838 96314
rect 7862 96262 7892 96314
rect 7892 96262 7918 96314
rect 7622 96260 7678 96262
rect 7702 96260 7758 96262
rect 7782 96260 7838 96262
rect 7862 96260 7918 96262
rect 7622 95226 7678 95228
rect 7702 95226 7758 95228
rect 7782 95226 7838 95228
rect 7862 95226 7918 95228
rect 7622 95174 7648 95226
rect 7648 95174 7678 95226
rect 7702 95174 7712 95226
rect 7712 95174 7758 95226
rect 7782 95174 7828 95226
rect 7828 95174 7838 95226
rect 7862 95174 7892 95226
rect 7892 95174 7918 95226
rect 7622 95172 7678 95174
rect 7702 95172 7758 95174
rect 7782 95172 7838 95174
rect 7862 95172 7918 95174
rect 7622 94138 7678 94140
rect 7702 94138 7758 94140
rect 7782 94138 7838 94140
rect 7862 94138 7918 94140
rect 7622 94086 7648 94138
rect 7648 94086 7678 94138
rect 7702 94086 7712 94138
rect 7712 94086 7758 94138
rect 7782 94086 7828 94138
rect 7828 94086 7838 94138
rect 7862 94086 7892 94138
rect 7892 94086 7918 94138
rect 7622 94084 7678 94086
rect 7702 94084 7758 94086
rect 7782 94084 7838 94086
rect 7862 94084 7918 94086
rect 7622 93050 7678 93052
rect 7702 93050 7758 93052
rect 7782 93050 7838 93052
rect 7862 93050 7918 93052
rect 7622 92998 7648 93050
rect 7648 92998 7678 93050
rect 7702 92998 7712 93050
rect 7712 92998 7758 93050
rect 7782 92998 7828 93050
rect 7828 92998 7838 93050
rect 7862 92998 7892 93050
rect 7892 92998 7918 93050
rect 7622 92996 7678 92998
rect 7702 92996 7758 92998
rect 7782 92996 7838 92998
rect 7862 92996 7918 92998
rect 7622 91962 7678 91964
rect 7702 91962 7758 91964
rect 7782 91962 7838 91964
rect 7862 91962 7918 91964
rect 7622 91910 7648 91962
rect 7648 91910 7678 91962
rect 7702 91910 7712 91962
rect 7712 91910 7758 91962
rect 7782 91910 7828 91962
rect 7828 91910 7838 91962
rect 7862 91910 7892 91962
rect 7892 91910 7918 91962
rect 7622 91908 7678 91910
rect 7702 91908 7758 91910
rect 7782 91908 7838 91910
rect 7862 91908 7918 91910
rect 7622 90874 7678 90876
rect 7702 90874 7758 90876
rect 7782 90874 7838 90876
rect 7862 90874 7918 90876
rect 7622 90822 7648 90874
rect 7648 90822 7678 90874
rect 7702 90822 7712 90874
rect 7712 90822 7758 90874
rect 7782 90822 7828 90874
rect 7828 90822 7838 90874
rect 7862 90822 7892 90874
rect 7892 90822 7918 90874
rect 7622 90820 7678 90822
rect 7702 90820 7758 90822
rect 7782 90820 7838 90822
rect 7862 90820 7918 90822
rect 7622 89786 7678 89788
rect 7702 89786 7758 89788
rect 7782 89786 7838 89788
rect 7862 89786 7918 89788
rect 7622 89734 7648 89786
rect 7648 89734 7678 89786
rect 7702 89734 7712 89786
rect 7712 89734 7758 89786
rect 7782 89734 7828 89786
rect 7828 89734 7838 89786
rect 7862 89734 7892 89786
rect 7892 89734 7918 89786
rect 7622 89732 7678 89734
rect 7702 89732 7758 89734
rect 7782 89732 7838 89734
rect 7862 89732 7918 89734
rect 7622 88698 7678 88700
rect 7702 88698 7758 88700
rect 7782 88698 7838 88700
rect 7862 88698 7918 88700
rect 7622 88646 7648 88698
rect 7648 88646 7678 88698
rect 7702 88646 7712 88698
rect 7712 88646 7758 88698
rect 7782 88646 7828 88698
rect 7828 88646 7838 88698
rect 7862 88646 7892 88698
rect 7892 88646 7918 88698
rect 7622 88644 7678 88646
rect 7702 88644 7758 88646
rect 7782 88644 7838 88646
rect 7862 88644 7918 88646
rect 7622 87610 7678 87612
rect 7702 87610 7758 87612
rect 7782 87610 7838 87612
rect 7862 87610 7918 87612
rect 7622 87558 7648 87610
rect 7648 87558 7678 87610
rect 7702 87558 7712 87610
rect 7712 87558 7758 87610
rect 7782 87558 7828 87610
rect 7828 87558 7838 87610
rect 7862 87558 7892 87610
rect 7892 87558 7918 87610
rect 7622 87556 7678 87558
rect 7702 87556 7758 87558
rect 7782 87556 7838 87558
rect 7862 87556 7918 87558
rect 7622 86522 7678 86524
rect 7702 86522 7758 86524
rect 7782 86522 7838 86524
rect 7862 86522 7918 86524
rect 7622 86470 7648 86522
rect 7648 86470 7678 86522
rect 7702 86470 7712 86522
rect 7712 86470 7758 86522
rect 7782 86470 7828 86522
rect 7828 86470 7838 86522
rect 7862 86470 7892 86522
rect 7892 86470 7918 86522
rect 7622 86468 7678 86470
rect 7702 86468 7758 86470
rect 7782 86468 7838 86470
rect 7862 86468 7918 86470
rect 7622 85434 7678 85436
rect 7702 85434 7758 85436
rect 7782 85434 7838 85436
rect 7862 85434 7918 85436
rect 7622 85382 7648 85434
rect 7648 85382 7678 85434
rect 7702 85382 7712 85434
rect 7712 85382 7758 85434
rect 7782 85382 7828 85434
rect 7828 85382 7838 85434
rect 7862 85382 7892 85434
rect 7892 85382 7918 85434
rect 7622 85380 7678 85382
rect 7702 85380 7758 85382
rect 7782 85380 7838 85382
rect 7862 85380 7918 85382
rect 7622 84346 7678 84348
rect 7702 84346 7758 84348
rect 7782 84346 7838 84348
rect 7862 84346 7918 84348
rect 7622 84294 7648 84346
rect 7648 84294 7678 84346
rect 7702 84294 7712 84346
rect 7712 84294 7758 84346
rect 7782 84294 7828 84346
rect 7828 84294 7838 84346
rect 7862 84294 7892 84346
rect 7892 84294 7918 84346
rect 7622 84292 7678 84294
rect 7702 84292 7758 84294
rect 7782 84292 7838 84294
rect 7862 84292 7918 84294
rect 8206 83680 8262 83736
rect 7622 83258 7678 83260
rect 7702 83258 7758 83260
rect 7782 83258 7838 83260
rect 7862 83258 7918 83260
rect 7622 83206 7648 83258
rect 7648 83206 7678 83258
rect 7702 83206 7712 83258
rect 7712 83206 7758 83258
rect 7782 83206 7828 83258
rect 7828 83206 7838 83258
rect 7862 83206 7892 83258
rect 7892 83206 7918 83258
rect 7622 83204 7678 83206
rect 7702 83204 7758 83206
rect 7782 83204 7838 83206
rect 7862 83204 7918 83206
rect 7622 82170 7678 82172
rect 7702 82170 7758 82172
rect 7782 82170 7838 82172
rect 7862 82170 7918 82172
rect 7622 82118 7648 82170
rect 7648 82118 7678 82170
rect 7702 82118 7712 82170
rect 7712 82118 7758 82170
rect 7782 82118 7828 82170
rect 7828 82118 7838 82170
rect 7862 82118 7892 82170
rect 7892 82118 7918 82170
rect 7622 82116 7678 82118
rect 7702 82116 7758 82118
rect 7782 82116 7838 82118
rect 7862 82116 7918 82118
rect 7622 81082 7678 81084
rect 7702 81082 7758 81084
rect 7782 81082 7838 81084
rect 7862 81082 7918 81084
rect 7622 81030 7648 81082
rect 7648 81030 7678 81082
rect 7702 81030 7712 81082
rect 7712 81030 7758 81082
rect 7782 81030 7828 81082
rect 7828 81030 7838 81082
rect 7862 81030 7892 81082
rect 7892 81030 7918 81082
rect 7622 81028 7678 81030
rect 7702 81028 7758 81030
rect 7782 81028 7838 81030
rect 7862 81028 7918 81030
rect 7622 79994 7678 79996
rect 7702 79994 7758 79996
rect 7782 79994 7838 79996
rect 7862 79994 7918 79996
rect 7622 79942 7648 79994
rect 7648 79942 7678 79994
rect 7702 79942 7712 79994
rect 7712 79942 7758 79994
rect 7782 79942 7828 79994
rect 7828 79942 7838 79994
rect 7862 79942 7892 79994
rect 7892 79942 7918 79994
rect 7622 79940 7678 79942
rect 7702 79940 7758 79942
rect 7782 79940 7838 79942
rect 7862 79940 7918 79942
rect 7622 78906 7678 78908
rect 7702 78906 7758 78908
rect 7782 78906 7838 78908
rect 7862 78906 7918 78908
rect 7622 78854 7648 78906
rect 7648 78854 7678 78906
rect 7702 78854 7712 78906
rect 7712 78854 7758 78906
rect 7782 78854 7828 78906
rect 7828 78854 7838 78906
rect 7862 78854 7892 78906
rect 7892 78854 7918 78906
rect 7622 78852 7678 78854
rect 7702 78852 7758 78854
rect 7782 78852 7838 78854
rect 7862 78852 7918 78854
rect 7622 77818 7678 77820
rect 7702 77818 7758 77820
rect 7782 77818 7838 77820
rect 7862 77818 7918 77820
rect 7622 77766 7648 77818
rect 7648 77766 7678 77818
rect 7702 77766 7712 77818
rect 7712 77766 7758 77818
rect 7782 77766 7828 77818
rect 7828 77766 7838 77818
rect 7862 77766 7892 77818
rect 7892 77766 7918 77818
rect 7622 77764 7678 77766
rect 7702 77764 7758 77766
rect 7782 77764 7838 77766
rect 7862 77764 7918 77766
rect 7622 76730 7678 76732
rect 7702 76730 7758 76732
rect 7782 76730 7838 76732
rect 7862 76730 7918 76732
rect 7622 76678 7648 76730
rect 7648 76678 7678 76730
rect 7702 76678 7712 76730
rect 7712 76678 7758 76730
rect 7782 76678 7828 76730
rect 7828 76678 7838 76730
rect 7862 76678 7892 76730
rect 7892 76678 7918 76730
rect 7622 76676 7678 76678
rect 7702 76676 7758 76678
rect 7782 76676 7838 76678
rect 7862 76676 7918 76678
rect 7622 75642 7678 75644
rect 7702 75642 7758 75644
rect 7782 75642 7838 75644
rect 7862 75642 7918 75644
rect 7622 75590 7648 75642
rect 7648 75590 7678 75642
rect 7702 75590 7712 75642
rect 7712 75590 7758 75642
rect 7782 75590 7828 75642
rect 7828 75590 7838 75642
rect 7862 75590 7892 75642
rect 7892 75590 7918 75642
rect 7622 75588 7678 75590
rect 7702 75588 7758 75590
rect 7782 75588 7838 75590
rect 7862 75588 7918 75590
rect 7622 74554 7678 74556
rect 7702 74554 7758 74556
rect 7782 74554 7838 74556
rect 7862 74554 7918 74556
rect 7622 74502 7648 74554
rect 7648 74502 7678 74554
rect 7702 74502 7712 74554
rect 7712 74502 7758 74554
rect 7782 74502 7828 74554
rect 7828 74502 7838 74554
rect 7862 74502 7892 74554
rect 7892 74502 7918 74554
rect 7622 74500 7678 74502
rect 7702 74500 7758 74502
rect 7782 74500 7838 74502
rect 7862 74500 7918 74502
rect 7622 73466 7678 73468
rect 7702 73466 7758 73468
rect 7782 73466 7838 73468
rect 7862 73466 7918 73468
rect 7622 73414 7648 73466
rect 7648 73414 7678 73466
rect 7702 73414 7712 73466
rect 7712 73414 7758 73466
rect 7782 73414 7828 73466
rect 7828 73414 7838 73466
rect 7862 73414 7892 73466
rect 7892 73414 7918 73466
rect 7622 73412 7678 73414
rect 7702 73412 7758 73414
rect 7782 73412 7838 73414
rect 7862 73412 7918 73414
rect 7622 72378 7678 72380
rect 7702 72378 7758 72380
rect 7782 72378 7838 72380
rect 7862 72378 7918 72380
rect 7622 72326 7648 72378
rect 7648 72326 7678 72378
rect 7702 72326 7712 72378
rect 7712 72326 7758 72378
rect 7782 72326 7828 72378
rect 7828 72326 7838 72378
rect 7862 72326 7892 72378
rect 7892 72326 7918 72378
rect 7622 72324 7678 72326
rect 7702 72324 7758 72326
rect 7782 72324 7838 72326
rect 7862 72324 7918 72326
rect 7622 71290 7678 71292
rect 7702 71290 7758 71292
rect 7782 71290 7838 71292
rect 7862 71290 7918 71292
rect 7622 71238 7648 71290
rect 7648 71238 7678 71290
rect 7702 71238 7712 71290
rect 7712 71238 7758 71290
rect 7782 71238 7828 71290
rect 7828 71238 7838 71290
rect 7862 71238 7892 71290
rect 7892 71238 7918 71290
rect 7622 71236 7678 71238
rect 7702 71236 7758 71238
rect 7782 71236 7838 71238
rect 7862 71236 7918 71238
rect 7622 70202 7678 70204
rect 7702 70202 7758 70204
rect 7782 70202 7838 70204
rect 7862 70202 7918 70204
rect 7622 70150 7648 70202
rect 7648 70150 7678 70202
rect 7702 70150 7712 70202
rect 7712 70150 7758 70202
rect 7782 70150 7828 70202
rect 7828 70150 7838 70202
rect 7862 70150 7892 70202
rect 7892 70150 7918 70202
rect 7622 70148 7678 70150
rect 7702 70148 7758 70150
rect 7782 70148 7838 70150
rect 7862 70148 7918 70150
rect 7622 69114 7678 69116
rect 7702 69114 7758 69116
rect 7782 69114 7838 69116
rect 7862 69114 7918 69116
rect 7622 69062 7648 69114
rect 7648 69062 7678 69114
rect 7702 69062 7712 69114
rect 7712 69062 7758 69114
rect 7782 69062 7828 69114
rect 7828 69062 7838 69114
rect 7862 69062 7892 69114
rect 7892 69062 7918 69114
rect 7622 69060 7678 69062
rect 7702 69060 7758 69062
rect 7782 69060 7838 69062
rect 7862 69060 7918 69062
rect 7622 68026 7678 68028
rect 7702 68026 7758 68028
rect 7782 68026 7838 68028
rect 7862 68026 7918 68028
rect 7622 67974 7648 68026
rect 7648 67974 7678 68026
rect 7702 67974 7712 68026
rect 7712 67974 7758 68026
rect 7782 67974 7828 68026
rect 7828 67974 7838 68026
rect 7862 67974 7892 68026
rect 7892 67974 7918 68026
rect 7622 67972 7678 67974
rect 7702 67972 7758 67974
rect 7782 67972 7838 67974
rect 7862 67972 7918 67974
rect 7622 66938 7678 66940
rect 7702 66938 7758 66940
rect 7782 66938 7838 66940
rect 7862 66938 7918 66940
rect 7622 66886 7648 66938
rect 7648 66886 7678 66938
rect 7702 66886 7712 66938
rect 7712 66886 7758 66938
rect 7782 66886 7828 66938
rect 7828 66886 7838 66938
rect 7862 66886 7892 66938
rect 7892 66886 7918 66938
rect 7622 66884 7678 66886
rect 7702 66884 7758 66886
rect 7782 66884 7838 66886
rect 7862 66884 7918 66886
rect 7622 65850 7678 65852
rect 7702 65850 7758 65852
rect 7782 65850 7838 65852
rect 7862 65850 7918 65852
rect 7622 65798 7648 65850
rect 7648 65798 7678 65850
rect 7702 65798 7712 65850
rect 7712 65798 7758 65850
rect 7782 65798 7828 65850
rect 7828 65798 7838 65850
rect 7862 65798 7892 65850
rect 7892 65798 7918 65850
rect 7622 65796 7678 65798
rect 7702 65796 7758 65798
rect 7782 65796 7838 65798
rect 7862 65796 7918 65798
rect 7622 64762 7678 64764
rect 7702 64762 7758 64764
rect 7782 64762 7838 64764
rect 7862 64762 7918 64764
rect 7622 64710 7648 64762
rect 7648 64710 7678 64762
rect 7702 64710 7712 64762
rect 7712 64710 7758 64762
rect 7782 64710 7828 64762
rect 7828 64710 7838 64762
rect 7862 64710 7892 64762
rect 7892 64710 7918 64762
rect 7622 64708 7678 64710
rect 7702 64708 7758 64710
rect 7782 64708 7838 64710
rect 7862 64708 7918 64710
rect 7622 63674 7678 63676
rect 7702 63674 7758 63676
rect 7782 63674 7838 63676
rect 7862 63674 7918 63676
rect 7622 63622 7648 63674
rect 7648 63622 7678 63674
rect 7702 63622 7712 63674
rect 7712 63622 7758 63674
rect 7782 63622 7828 63674
rect 7828 63622 7838 63674
rect 7862 63622 7892 63674
rect 7892 63622 7918 63674
rect 7622 63620 7678 63622
rect 7702 63620 7758 63622
rect 7782 63620 7838 63622
rect 7862 63620 7918 63622
rect 7622 62586 7678 62588
rect 7702 62586 7758 62588
rect 7782 62586 7838 62588
rect 7862 62586 7918 62588
rect 7622 62534 7648 62586
rect 7648 62534 7678 62586
rect 7702 62534 7712 62586
rect 7712 62534 7758 62586
rect 7782 62534 7828 62586
rect 7828 62534 7838 62586
rect 7862 62534 7892 62586
rect 7892 62534 7918 62586
rect 7622 62532 7678 62534
rect 7702 62532 7758 62534
rect 7782 62532 7838 62534
rect 7862 62532 7918 62534
rect 7622 61498 7678 61500
rect 7702 61498 7758 61500
rect 7782 61498 7838 61500
rect 7862 61498 7918 61500
rect 7622 61446 7648 61498
rect 7648 61446 7678 61498
rect 7702 61446 7712 61498
rect 7712 61446 7758 61498
rect 7782 61446 7828 61498
rect 7828 61446 7838 61498
rect 7862 61446 7892 61498
rect 7892 61446 7918 61498
rect 7622 61444 7678 61446
rect 7702 61444 7758 61446
rect 7782 61444 7838 61446
rect 7862 61444 7918 61446
rect 7622 60410 7678 60412
rect 7702 60410 7758 60412
rect 7782 60410 7838 60412
rect 7862 60410 7918 60412
rect 7622 60358 7648 60410
rect 7648 60358 7678 60410
rect 7702 60358 7712 60410
rect 7712 60358 7758 60410
rect 7782 60358 7828 60410
rect 7828 60358 7838 60410
rect 7862 60358 7892 60410
rect 7892 60358 7918 60410
rect 7622 60356 7678 60358
rect 7702 60356 7758 60358
rect 7782 60356 7838 60358
rect 7862 60356 7918 60358
rect 7622 59322 7678 59324
rect 7702 59322 7758 59324
rect 7782 59322 7838 59324
rect 7862 59322 7918 59324
rect 7622 59270 7648 59322
rect 7648 59270 7678 59322
rect 7702 59270 7712 59322
rect 7712 59270 7758 59322
rect 7782 59270 7828 59322
rect 7828 59270 7838 59322
rect 7862 59270 7892 59322
rect 7892 59270 7918 59322
rect 7622 59268 7678 59270
rect 7702 59268 7758 59270
rect 7782 59268 7838 59270
rect 7862 59268 7918 59270
rect 7622 58234 7678 58236
rect 7702 58234 7758 58236
rect 7782 58234 7838 58236
rect 7862 58234 7918 58236
rect 7622 58182 7648 58234
rect 7648 58182 7678 58234
rect 7702 58182 7712 58234
rect 7712 58182 7758 58234
rect 7782 58182 7828 58234
rect 7828 58182 7838 58234
rect 7862 58182 7892 58234
rect 7892 58182 7918 58234
rect 7622 58180 7678 58182
rect 7702 58180 7758 58182
rect 7782 58180 7838 58182
rect 7862 58180 7918 58182
rect 7622 57146 7678 57148
rect 7702 57146 7758 57148
rect 7782 57146 7838 57148
rect 7862 57146 7918 57148
rect 7622 57094 7648 57146
rect 7648 57094 7678 57146
rect 7702 57094 7712 57146
rect 7712 57094 7758 57146
rect 7782 57094 7828 57146
rect 7828 57094 7838 57146
rect 7862 57094 7892 57146
rect 7892 57094 7918 57146
rect 7622 57092 7678 57094
rect 7702 57092 7758 57094
rect 7782 57092 7838 57094
rect 7862 57092 7918 57094
rect 7622 56058 7678 56060
rect 7702 56058 7758 56060
rect 7782 56058 7838 56060
rect 7862 56058 7918 56060
rect 7622 56006 7648 56058
rect 7648 56006 7678 56058
rect 7702 56006 7712 56058
rect 7712 56006 7758 56058
rect 7782 56006 7828 56058
rect 7828 56006 7838 56058
rect 7862 56006 7892 56058
rect 7892 56006 7918 56058
rect 7622 56004 7678 56006
rect 7702 56004 7758 56006
rect 7782 56004 7838 56006
rect 7862 56004 7918 56006
rect 7622 54970 7678 54972
rect 7702 54970 7758 54972
rect 7782 54970 7838 54972
rect 7862 54970 7918 54972
rect 7622 54918 7648 54970
rect 7648 54918 7678 54970
rect 7702 54918 7712 54970
rect 7712 54918 7758 54970
rect 7782 54918 7828 54970
rect 7828 54918 7838 54970
rect 7862 54918 7892 54970
rect 7892 54918 7918 54970
rect 7622 54916 7678 54918
rect 7702 54916 7758 54918
rect 7782 54916 7838 54918
rect 7862 54916 7918 54918
rect 7622 53882 7678 53884
rect 7702 53882 7758 53884
rect 7782 53882 7838 53884
rect 7862 53882 7918 53884
rect 7622 53830 7648 53882
rect 7648 53830 7678 53882
rect 7702 53830 7712 53882
rect 7712 53830 7758 53882
rect 7782 53830 7828 53882
rect 7828 53830 7838 53882
rect 7862 53830 7892 53882
rect 7892 53830 7918 53882
rect 7622 53828 7678 53830
rect 7702 53828 7758 53830
rect 7782 53828 7838 53830
rect 7862 53828 7918 53830
rect 7622 52794 7678 52796
rect 7702 52794 7758 52796
rect 7782 52794 7838 52796
rect 7862 52794 7918 52796
rect 7622 52742 7648 52794
rect 7648 52742 7678 52794
rect 7702 52742 7712 52794
rect 7712 52742 7758 52794
rect 7782 52742 7828 52794
rect 7828 52742 7838 52794
rect 7862 52742 7892 52794
rect 7892 52742 7918 52794
rect 7622 52740 7678 52742
rect 7702 52740 7758 52742
rect 7782 52740 7838 52742
rect 7862 52740 7918 52742
rect 7622 51706 7678 51708
rect 7702 51706 7758 51708
rect 7782 51706 7838 51708
rect 7862 51706 7918 51708
rect 7622 51654 7648 51706
rect 7648 51654 7678 51706
rect 7702 51654 7712 51706
rect 7712 51654 7758 51706
rect 7782 51654 7828 51706
rect 7828 51654 7838 51706
rect 7862 51654 7892 51706
rect 7892 51654 7918 51706
rect 7622 51652 7678 51654
rect 7702 51652 7758 51654
rect 7782 51652 7838 51654
rect 7862 51652 7918 51654
rect 7622 50618 7678 50620
rect 7702 50618 7758 50620
rect 7782 50618 7838 50620
rect 7862 50618 7918 50620
rect 7622 50566 7648 50618
rect 7648 50566 7678 50618
rect 7702 50566 7712 50618
rect 7712 50566 7758 50618
rect 7782 50566 7828 50618
rect 7828 50566 7838 50618
rect 7862 50566 7892 50618
rect 7892 50566 7918 50618
rect 7622 50564 7678 50566
rect 7702 50564 7758 50566
rect 7782 50564 7838 50566
rect 7862 50564 7918 50566
rect 7622 49530 7678 49532
rect 7702 49530 7758 49532
rect 7782 49530 7838 49532
rect 7862 49530 7918 49532
rect 7622 49478 7648 49530
rect 7648 49478 7678 49530
rect 7702 49478 7712 49530
rect 7712 49478 7758 49530
rect 7782 49478 7828 49530
rect 7828 49478 7838 49530
rect 7862 49478 7892 49530
rect 7892 49478 7918 49530
rect 7622 49476 7678 49478
rect 7702 49476 7758 49478
rect 7782 49476 7838 49478
rect 7862 49476 7918 49478
rect 7622 48442 7678 48444
rect 7702 48442 7758 48444
rect 7782 48442 7838 48444
rect 7862 48442 7918 48444
rect 7622 48390 7648 48442
rect 7648 48390 7678 48442
rect 7702 48390 7712 48442
rect 7712 48390 7758 48442
rect 7782 48390 7828 48442
rect 7828 48390 7838 48442
rect 7862 48390 7892 48442
rect 7892 48390 7918 48442
rect 7622 48388 7678 48390
rect 7702 48388 7758 48390
rect 7782 48388 7838 48390
rect 7862 48388 7918 48390
rect 7622 47354 7678 47356
rect 7702 47354 7758 47356
rect 7782 47354 7838 47356
rect 7862 47354 7918 47356
rect 7622 47302 7648 47354
rect 7648 47302 7678 47354
rect 7702 47302 7712 47354
rect 7712 47302 7758 47354
rect 7782 47302 7828 47354
rect 7828 47302 7838 47354
rect 7862 47302 7892 47354
rect 7892 47302 7918 47354
rect 7622 47300 7678 47302
rect 7702 47300 7758 47302
rect 7782 47300 7838 47302
rect 7862 47300 7918 47302
rect 7622 46266 7678 46268
rect 7702 46266 7758 46268
rect 7782 46266 7838 46268
rect 7862 46266 7918 46268
rect 7622 46214 7648 46266
rect 7648 46214 7678 46266
rect 7702 46214 7712 46266
rect 7712 46214 7758 46266
rect 7782 46214 7828 46266
rect 7828 46214 7838 46266
rect 7862 46214 7892 46266
rect 7892 46214 7918 46266
rect 7622 46212 7678 46214
rect 7702 46212 7758 46214
rect 7782 46212 7838 46214
rect 7862 46212 7918 46214
rect 7622 45178 7678 45180
rect 7702 45178 7758 45180
rect 7782 45178 7838 45180
rect 7862 45178 7918 45180
rect 7622 45126 7648 45178
rect 7648 45126 7678 45178
rect 7702 45126 7712 45178
rect 7712 45126 7758 45178
rect 7782 45126 7828 45178
rect 7828 45126 7838 45178
rect 7862 45126 7892 45178
rect 7892 45126 7918 45178
rect 7622 45124 7678 45126
rect 7702 45124 7758 45126
rect 7782 45124 7838 45126
rect 7862 45124 7918 45126
rect 7622 44090 7678 44092
rect 7702 44090 7758 44092
rect 7782 44090 7838 44092
rect 7862 44090 7918 44092
rect 7622 44038 7648 44090
rect 7648 44038 7678 44090
rect 7702 44038 7712 44090
rect 7712 44038 7758 44090
rect 7782 44038 7828 44090
rect 7828 44038 7838 44090
rect 7862 44038 7892 44090
rect 7892 44038 7918 44090
rect 7622 44036 7678 44038
rect 7702 44036 7758 44038
rect 7782 44036 7838 44038
rect 7862 44036 7918 44038
rect 7622 43002 7678 43004
rect 7702 43002 7758 43004
rect 7782 43002 7838 43004
rect 7862 43002 7918 43004
rect 7622 42950 7648 43002
rect 7648 42950 7678 43002
rect 7702 42950 7712 43002
rect 7712 42950 7758 43002
rect 7782 42950 7828 43002
rect 7828 42950 7838 43002
rect 7862 42950 7892 43002
rect 7892 42950 7918 43002
rect 7622 42948 7678 42950
rect 7702 42948 7758 42950
rect 7782 42948 7838 42950
rect 7862 42948 7918 42950
rect 7622 41914 7678 41916
rect 7702 41914 7758 41916
rect 7782 41914 7838 41916
rect 7862 41914 7918 41916
rect 7622 41862 7648 41914
rect 7648 41862 7678 41914
rect 7702 41862 7712 41914
rect 7712 41862 7758 41914
rect 7782 41862 7828 41914
rect 7828 41862 7838 41914
rect 7862 41862 7892 41914
rect 7892 41862 7918 41914
rect 7622 41860 7678 41862
rect 7702 41860 7758 41862
rect 7782 41860 7838 41862
rect 7862 41860 7918 41862
rect 7622 40826 7678 40828
rect 7702 40826 7758 40828
rect 7782 40826 7838 40828
rect 7862 40826 7918 40828
rect 7622 40774 7648 40826
rect 7648 40774 7678 40826
rect 7702 40774 7712 40826
rect 7712 40774 7758 40826
rect 7782 40774 7828 40826
rect 7828 40774 7838 40826
rect 7862 40774 7892 40826
rect 7892 40774 7918 40826
rect 7622 40772 7678 40774
rect 7702 40772 7758 40774
rect 7782 40772 7838 40774
rect 7862 40772 7918 40774
rect 7622 39738 7678 39740
rect 7702 39738 7758 39740
rect 7782 39738 7838 39740
rect 7862 39738 7918 39740
rect 7622 39686 7648 39738
rect 7648 39686 7678 39738
rect 7702 39686 7712 39738
rect 7712 39686 7758 39738
rect 7782 39686 7828 39738
rect 7828 39686 7838 39738
rect 7862 39686 7892 39738
rect 7892 39686 7918 39738
rect 7622 39684 7678 39686
rect 7702 39684 7758 39686
rect 7782 39684 7838 39686
rect 7862 39684 7918 39686
rect 7622 38650 7678 38652
rect 7702 38650 7758 38652
rect 7782 38650 7838 38652
rect 7862 38650 7918 38652
rect 7622 38598 7648 38650
rect 7648 38598 7678 38650
rect 7702 38598 7712 38650
rect 7712 38598 7758 38650
rect 7782 38598 7828 38650
rect 7828 38598 7838 38650
rect 7862 38598 7892 38650
rect 7892 38598 7918 38650
rect 7622 38596 7678 38598
rect 7702 38596 7758 38598
rect 7782 38596 7838 38598
rect 7862 38596 7918 38598
rect 7622 37562 7678 37564
rect 7702 37562 7758 37564
rect 7782 37562 7838 37564
rect 7862 37562 7918 37564
rect 7622 37510 7648 37562
rect 7648 37510 7678 37562
rect 7702 37510 7712 37562
rect 7712 37510 7758 37562
rect 7782 37510 7828 37562
rect 7828 37510 7838 37562
rect 7862 37510 7892 37562
rect 7892 37510 7918 37562
rect 7622 37508 7678 37510
rect 7702 37508 7758 37510
rect 7782 37508 7838 37510
rect 7862 37508 7918 37510
rect 7622 36474 7678 36476
rect 7702 36474 7758 36476
rect 7782 36474 7838 36476
rect 7862 36474 7918 36476
rect 7622 36422 7648 36474
rect 7648 36422 7678 36474
rect 7702 36422 7712 36474
rect 7712 36422 7758 36474
rect 7782 36422 7828 36474
rect 7828 36422 7838 36474
rect 7862 36422 7892 36474
rect 7892 36422 7918 36474
rect 7622 36420 7678 36422
rect 7702 36420 7758 36422
rect 7782 36420 7838 36422
rect 7862 36420 7918 36422
rect 7622 35386 7678 35388
rect 7702 35386 7758 35388
rect 7782 35386 7838 35388
rect 7862 35386 7918 35388
rect 7622 35334 7648 35386
rect 7648 35334 7678 35386
rect 7702 35334 7712 35386
rect 7712 35334 7758 35386
rect 7782 35334 7828 35386
rect 7828 35334 7838 35386
rect 7862 35334 7892 35386
rect 7892 35334 7918 35386
rect 7622 35332 7678 35334
rect 7702 35332 7758 35334
rect 7782 35332 7838 35334
rect 7862 35332 7918 35334
rect 7622 34298 7678 34300
rect 7702 34298 7758 34300
rect 7782 34298 7838 34300
rect 7862 34298 7918 34300
rect 7622 34246 7648 34298
rect 7648 34246 7678 34298
rect 7702 34246 7712 34298
rect 7712 34246 7758 34298
rect 7782 34246 7828 34298
rect 7828 34246 7838 34298
rect 7862 34246 7892 34298
rect 7892 34246 7918 34298
rect 7622 34244 7678 34246
rect 7702 34244 7758 34246
rect 7782 34244 7838 34246
rect 7862 34244 7918 34246
rect 7622 33210 7678 33212
rect 7702 33210 7758 33212
rect 7782 33210 7838 33212
rect 7862 33210 7918 33212
rect 7622 33158 7648 33210
rect 7648 33158 7678 33210
rect 7702 33158 7712 33210
rect 7712 33158 7758 33210
rect 7782 33158 7828 33210
rect 7828 33158 7838 33210
rect 7862 33158 7892 33210
rect 7892 33158 7918 33210
rect 7622 33156 7678 33158
rect 7702 33156 7758 33158
rect 7782 33156 7838 33158
rect 7862 33156 7918 33158
rect 7622 32122 7678 32124
rect 7702 32122 7758 32124
rect 7782 32122 7838 32124
rect 7862 32122 7918 32124
rect 7622 32070 7648 32122
rect 7648 32070 7678 32122
rect 7702 32070 7712 32122
rect 7712 32070 7758 32122
rect 7782 32070 7828 32122
rect 7828 32070 7838 32122
rect 7862 32070 7892 32122
rect 7892 32070 7918 32122
rect 7622 32068 7678 32070
rect 7702 32068 7758 32070
rect 7782 32068 7838 32070
rect 7862 32068 7918 32070
rect 7622 31034 7678 31036
rect 7702 31034 7758 31036
rect 7782 31034 7838 31036
rect 7862 31034 7918 31036
rect 7622 30982 7648 31034
rect 7648 30982 7678 31034
rect 7702 30982 7712 31034
rect 7712 30982 7758 31034
rect 7782 30982 7828 31034
rect 7828 30982 7838 31034
rect 7862 30982 7892 31034
rect 7892 30982 7918 31034
rect 7622 30980 7678 30982
rect 7702 30980 7758 30982
rect 7782 30980 7838 30982
rect 7862 30980 7918 30982
rect 7622 29946 7678 29948
rect 7702 29946 7758 29948
rect 7782 29946 7838 29948
rect 7862 29946 7918 29948
rect 7622 29894 7648 29946
rect 7648 29894 7678 29946
rect 7702 29894 7712 29946
rect 7712 29894 7758 29946
rect 7782 29894 7828 29946
rect 7828 29894 7838 29946
rect 7862 29894 7892 29946
rect 7892 29894 7918 29946
rect 7622 29892 7678 29894
rect 7702 29892 7758 29894
rect 7782 29892 7838 29894
rect 7862 29892 7918 29894
rect 7622 28858 7678 28860
rect 7702 28858 7758 28860
rect 7782 28858 7838 28860
rect 7862 28858 7918 28860
rect 7622 28806 7648 28858
rect 7648 28806 7678 28858
rect 7702 28806 7712 28858
rect 7712 28806 7758 28858
rect 7782 28806 7828 28858
rect 7828 28806 7838 28858
rect 7862 28806 7892 28858
rect 7892 28806 7918 28858
rect 7622 28804 7678 28806
rect 7702 28804 7758 28806
rect 7782 28804 7838 28806
rect 7862 28804 7918 28806
rect 7622 27770 7678 27772
rect 7702 27770 7758 27772
rect 7782 27770 7838 27772
rect 7862 27770 7918 27772
rect 7622 27718 7648 27770
rect 7648 27718 7678 27770
rect 7702 27718 7712 27770
rect 7712 27718 7758 27770
rect 7782 27718 7828 27770
rect 7828 27718 7838 27770
rect 7862 27718 7892 27770
rect 7892 27718 7918 27770
rect 7622 27716 7678 27718
rect 7702 27716 7758 27718
rect 7782 27716 7838 27718
rect 7862 27716 7918 27718
rect 7622 26682 7678 26684
rect 7702 26682 7758 26684
rect 7782 26682 7838 26684
rect 7862 26682 7918 26684
rect 7622 26630 7648 26682
rect 7648 26630 7678 26682
rect 7702 26630 7712 26682
rect 7712 26630 7758 26682
rect 7782 26630 7828 26682
rect 7828 26630 7838 26682
rect 7862 26630 7892 26682
rect 7892 26630 7918 26682
rect 7622 26628 7678 26630
rect 7702 26628 7758 26630
rect 7782 26628 7838 26630
rect 7862 26628 7918 26630
rect 7622 25594 7678 25596
rect 7702 25594 7758 25596
rect 7782 25594 7838 25596
rect 7862 25594 7918 25596
rect 7622 25542 7648 25594
rect 7648 25542 7678 25594
rect 7702 25542 7712 25594
rect 7712 25542 7758 25594
rect 7782 25542 7828 25594
rect 7828 25542 7838 25594
rect 7862 25542 7892 25594
rect 7892 25542 7918 25594
rect 7622 25540 7678 25542
rect 7702 25540 7758 25542
rect 7782 25540 7838 25542
rect 7862 25540 7918 25542
rect 7622 24506 7678 24508
rect 7702 24506 7758 24508
rect 7782 24506 7838 24508
rect 7862 24506 7918 24508
rect 7622 24454 7648 24506
rect 7648 24454 7678 24506
rect 7702 24454 7712 24506
rect 7712 24454 7758 24506
rect 7782 24454 7828 24506
rect 7828 24454 7838 24506
rect 7862 24454 7892 24506
rect 7892 24454 7918 24506
rect 7622 24452 7678 24454
rect 7702 24452 7758 24454
rect 7782 24452 7838 24454
rect 7862 24452 7918 24454
rect 7622 23418 7678 23420
rect 7702 23418 7758 23420
rect 7782 23418 7838 23420
rect 7862 23418 7918 23420
rect 7622 23366 7648 23418
rect 7648 23366 7678 23418
rect 7702 23366 7712 23418
rect 7712 23366 7758 23418
rect 7782 23366 7828 23418
rect 7828 23366 7838 23418
rect 7862 23366 7892 23418
rect 7892 23366 7918 23418
rect 7622 23364 7678 23366
rect 7702 23364 7758 23366
rect 7782 23364 7838 23366
rect 7862 23364 7918 23366
rect 7622 22330 7678 22332
rect 7702 22330 7758 22332
rect 7782 22330 7838 22332
rect 7862 22330 7918 22332
rect 7622 22278 7648 22330
rect 7648 22278 7678 22330
rect 7702 22278 7712 22330
rect 7712 22278 7758 22330
rect 7782 22278 7828 22330
rect 7828 22278 7838 22330
rect 7862 22278 7892 22330
rect 7892 22278 7918 22330
rect 7622 22276 7678 22278
rect 7702 22276 7758 22278
rect 7782 22276 7838 22278
rect 7862 22276 7918 22278
rect 7622 21242 7678 21244
rect 7702 21242 7758 21244
rect 7782 21242 7838 21244
rect 7862 21242 7918 21244
rect 7622 21190 7648 21242
rect 7648 21190 7678 21242
rect 7702 21190 7712 21242
rect 7712 21190 7758 21242
rect 7782 21190 7828 21242
rect 7828 21190 7838 21242
rect 7862 21190 7892 21242
rect 7892 21190 7918 21242
rect 7622 21188 7678 21190
rect 7702 21188 7758 21190
rect 7782 21188 7838 21190
rect 7862 21188 7918 21190
rect 7622 20154 7678 20156
rect 7702 20154 7758 20156
rect 7782 20154 7838 20156
rect 7862 20154 7918 20156
rect 7622 20102 7648 20154
rect 7648 20102 7678 20154
rect 7702 20102 7712 20154
rect 7712 20102 7758 20154
rect 7782 20102 7828 20154
rect 7828 20102 7838 20154
rect 7862 20102 7892 20154
rect 7892 20102 7918 20154
rect 7622 20100 7678 20102
rect 7702 20100 7758 20102
rect 7782 20100 7838 20102
rect 7862 20100 7918 20102
rect 7622 19066 7678 19068
rect 7702 19066 7758 19068
rect 7782 19066 7838 19068
rect 7862 19066 7918 19068
rect 7622 19014 7648 19066
rect 7648 19014 7678 19066
rect 7702 19014 7712 19066
rect 7712 19014 7758 19066
rect 7782 19014 7828 19066
rect 7828 19014 7838 19066
rect 7862 19014 7892 19066
rect 7892 19014 7918 19066
rect 7622 19012 7678 19014
rect 7702 19012 7758 19014
rect 7782 19012 7838 19014
rect 7862 19012 7918 19014
rect 7622 17978 7678 17980
rect 7702 17978 7758 17980
rect 7782 17978 7838 17980
rect 7862 17978 7918 17980
rect 7622 17926 7648 17978
rect 7648 17926 7678 17978
rect 7702 17926 7712 17978
rect 7712 17926 7758 17978
rect 7782 17926 7828 17978
rect 7828 17926 7838 17978
rect 7862 17926 7892 17978
rect 7892 17926 7918 17978
rect 7622 17924 7678 17926
rect 7702 17924 7758 17926
rect 7782 17924 7838 17926
rect 7862 17924 7918 17926
rect 7622 16890 7678 16892
rect 7702 16890 7758 16892
rect 7782 16890 7838 16892
rect 7862 16890 7918 16892
rect 7622 16838 7648 16890
rect 7648 16838 7678 16890
rect 7702 16838 7712 16890
rect 7712 16838 7758 16890
rect 7782 16838 7828 16890
rect 7828 16838 7838 16890
rect 7862 16838 7892 16890
rect 7892 16838 7918 16890
rect 7622 16836 7678 16838
rect 7702 16836 7758 16838
rect 7782 16836 7838 16838
rect 7862 16836 7918 16838
rect 7622 15802 7678 15804
rect 7702 15802 7758 15804
rect 7782 15802 7838 15804
rect 7862 15802 7918 15804
rect 7622 15750 7648 15802
rect 7648 15750 7678 15802
rect 7702 15750 7712 15802
rect 7712 15750 7758 15802
rect 7782 15750 7828 15802
rect 7828 15750 7838 15802
rect 7862 15750 7892 15802
rect 7892 15750 7918 15802
rect 7622 15748 7678 15750
rect 7702 15748 7758 15750
rect 7782 15748 7838 15750
rect 7862 15748 7918 15750
rect 7622 14714 7678 14716
rect 7702 14714 7758 14716
rect 7782 14714 7838 14716
rect 7862 14714 7918 14716
rect 7622 14662 7648 14714
rect 7648 14662 7678 14714
rect 7702 14662 7712 14714
rect 7712 14662 7758 14714
rect 7782 14662 7828 14714
rect 7828 14662 7838 14714
rect 7862 14662 7892 14714
rect 7892 14662 7918 14714
rect 7622 14660 7678 14662
rect 7702 14660 7758 14662
rect 7782 14660 7838 14662
rect 7862 14660 7918 14662
rect 7622 13626 7678 13628
rect 7702 13626 7758 13628
rect 7782 13626 7838 13628
rect 7862 13626 7918 13628
rect 7622 13574 7648 13626
rect 7648 13574 7678 13626
rect 7702 13574 7712 13626
rect 7712 13574 7758 13626
rect 7782 13574 7828 13626
rect 7828 13574 7838 13626
rect 7862 13574 7892 13626
rect 7892 13574 7918 13626
rect 7622 13572 7678 13574
rect 7702 13572 7758 13574
rect 7782 13572 7838 13574
rect 7862 13572 7918 13574
rect 7622 12538 7678 12540
rect 7702 12538 7758 12540
rect 7782 12538 7838 12540
rect 7862 12538 7918 12540
rect 7622 12486 7648 12538
rect 7648 12486 7678 12538
rect 7702 12486 7712 12538
rect 7712 12486 7758 12538
rect 7782 12486 7828 12538
rect 7828 12486 7838 12538
rect 7862 12486 7892 12538
rect 7892 12486 7918 12538
rect 7622 12484 7678 12486
rect 7702 12484 7758 12486
rect 7782 12484 7838 12486
rect 7862 12484 7918 12486
rect 7622 11450 7678 11452
rect 7702 11450 7758 11452
rect 7782 11450 7838 11452
rect 7862 11450 7918 11452
rect 7622 11398 7648 11450
rect 7648 11398 7678 11450
rect 7702 11398 7712 11450
rect 7712 11398 7758 11450
rect 7782 11398 7828 11450
rect 7828 11398 7838 11450
rect 7862 11398 7892 11450
rect 7892 11398 7918 11450
rect 7622 11396 7678 11398
rect 7702 11396 7758 11398
rect 7782 11396 7838 11398
rect 7862 11396 7918 11398
rect 7622 10362 7678 10364
rect 7702 10362 7758 10364
rect 7782 10362 7838 10364
rect 7862 10362 7918 10364
rect 7622 10310 7648 10362
rect 7648 10310 7678 10362
rect 7702 10310 7712 10362
rect 7712 10310 7758 10362
rect 7782 10310 7828 10362
rect 7828 10310 7838 10362
rect 7862 10310 7892 10362
rect 7892 10310 7918 10362
rect 7622 10308 7678 10310
rect 7702 10308 7758 10310
rect 7782 10308 7838 10310
rect 7862 10308 7918 10310
rect 7622 9274 7678 9276
rect 7702 9274 7758 9276
rect 7782 9274 7838 9276
rect 7862 9274 7918 9276
rect 7622 9222 7648 9274
rect 7648 9222 7678 9274
rect 7702 9222 7712 9274
rect 7712 9222 7758 9274
rect 7782 9222 7828 9274
rect 7828 9222 7838 9274
rect 7862 9222 7892 9274
rect 7892 9222 7918 9274
rect 7622 9220 7678 9222
rect 7702 9220 7758 9222
rect 7782 9220 7838 9222
rect 7862 9220 7918 9222
rect 7622 8186 7678 8188
rect 7702 8186 7758 8188
rect 7782 8186 7838 8188
rect 7862 8186 7918 8188
rect 7622 8134 7648 8186
rect 7648 8134 7678 8186
rect 7702 8134 7712 8186
rect 7712 8134 7758 8186
rect 7782 8134 7828 8186
rect 7828 8134 7838 8186
rect 7862 8134 7892 8186
rect 7892 8134 7918 8186
rect 7622 8132 7678 8134
rect 7702 8132 7758 8134
rect 7782 8132 7838 8134
rect 7862 8132 7918 8134
rect 7622 7098 7678 7100
rect 7702 7098 7758 7100
rect 7782 7098 7838 7100
rect 7862 7098 7918 7100
rect 7622 7046 7648 7098
rect 7648 7046 7678 7098
rect 7702 7046 7712 7098
rect 7712 7046 7758 7098
rect 7782 7046 7828 7098
rect 7828 7046 7838 7098
rect 7862 7046 7892 7098
rect 7892 7046 7918 7098
rect 7622 7044 7678 7046
rect 7702 7044 7758 7046
rect 7782 7044 7838 7046
rect 7862 7044 7918 7046
rect 7622 6010 7678 6012
rect 7702 6010 7758 6012
rect 7782 6010 7838 6012
rect 7862 6010 7918 6012
rect 7622 5958 7648 6010
rect 7648 5958 7678 6010
rect 7702 5958 7712 6010
rect 7712 5958 7758 6010
rect 7782 5958 7828 6010
rect 7828 5958 7838 6010
rect 7862 5958 7892 6010
rect 7892 5958 7918 6010
rect 7622 5956 7678 5958
rect 7702 5956 7758 5958
rect 7782 5956 7838 5958
rect 7862 5956 7918 5958
rect 7622 4922 7678 4924
rect 7702 4922 7758 4924
rect 7782 4922 7838 4924
rect 7862 4922 7918 4924
rect 7622 4870 7648 4922
rect 7648 4870 7678 4922
rect 7702 4870 7712 4922
rect 7712 4870 7758 4922
rect 7782 4870 7828 4922
rect 7828 4870 7838 4922
rect 7862 4870 7892 4922
rect 7892 4870 7918 4922
rect 7622 4868 7678 4870
rect 7702 4868 7758 4870
rect 7782 4868 7838 4870
rect 7862 4868 7918 4870
rect 4289 3834 4345 3836
rect 4369 3834 4425 3836
rect 4449 3834 4505 3836
rect 4529 3834 4585 3836
rect 4289 3782 4315 3834
rect 4315 3782 4345 3834
rect 4369 3782 4379 3834
rect 4379 3782 4425 3834
rect 4449 3782 4495 3834
rect 4495 3782 4505 3834
rect 4529 3782 4559 3834
rect 4559 3782 4585 3834
rect 4289 3780 4345 3782
rect 4369 3780 4425 3782
rect 4449 3780 4505 3782
rect 4529 3780 4585 3782
rect 5956 3290 6012 3292
rect 6036 3290 6092 3292
rect 6116 3290 6172 3292
rect 6196 3290 6252 3292
rect 5956 3238 5982 3290
rect 5982 3238 6012 3290
rect 6036 3238 6046 3290
rect 6046 3238 6092 3290
rect 6116 3238 6162 3290
rect 6162 3238 6172 3290
rect 6196 3238 6226 3290
rect 6226 3238 6252 3290
rect 5956 3236 6012 3238
rect 6036 3236 6092 3238
rect 6116 3236 6172 3238
rect 6196 3236 6252 3238
rect 4289 2746 4345 2748
rect 4369 2746 4425 2748
rect 4449 2746 4505 2748
rect 4529 2746 4585 2748
rect 4289 2694 4315 2746
rect 4315 2694 4345 2746
rect 4369 2694 4379 2746
rect 4379 2694 4425 2746
rect 4449 2694 4495 2746
rect 4495 2694 4505 2746
rect 4529 2694 4559 2746
rect 4559 2694 4585 2746
rect 4289 2692 4345 2694
rect 4369 2692 4425 2694
rect 4449 2692 4505 2694
rect 4529 2692 4585 2694
rect 5956 2202 6012 2204
rect 6036 2202 6092 2204
rect 6116 2202 6172 2204
rect 6196 2202 6252 2204
rect 5956 2150 5982 2202
rect 5982 2150 6012 2202
rect 6036 2150 6046 2202
rect 6046 2150 6092 2202
rect 6116 2150 6162 2202
rect 6162 2150 6172 2202
rect 6196 2150 6226 2202
rect 6226 2150 6252 2202
rect 5956 2148 6012 2150
rect 6036 2148 6092 2150
rect 6116 2148 6172 2150
rect 6196 2148 6252 2150
rect 7622 3834 7678 3836
rect 7702 3834 7758 3836
rect 7782 3834 7838 3836
rect 7862 3834 7918 3836
rect 7622 3782 7648 3834
rect 7648 3782 7678 3834
rect 7702 3782 7712 3834
rect 7712 3782 7758 3834
rect 7782 3782 7828 3834
rect 7828 3782 7838 3834
rect 7862 3782 7892 3834
rect 7892 3782 7918 3834
rect 7622 3780 7678 3782
rect 7702 3780 7758 3782
rect 7782 3780 7838 3782
rect 7862 3780 7918 3782
rect 7622 2746 7678 2748
rect 7702 2746 7758 2748
rect 7782 2746 7838 2748
rect 7862 2746 7918 2748
rect 7622 2694 7648 2746
rect 7648 2694 7678 2746
rect 7702 2694 7712 2746
rect 7712 2694 7758 2746
rect 7782 2694 7828 2746
rect 7828 2694 7838 2746
rect 7862 2694 7892 2746
rect 7892 2694 7918 2746
rect 7622 2692 7678 2694
rect 7702 2692 7758 2694
rect 7782 2692 7838 2694
rect 7862 2692 7918 2694
<< metal3 >>
rect 2610 330784 2930 330785
rect 2610 330720 2618 330784
rect 2682 330720 2698 330784
rect 2762 330720 2778 330784
rect 2842 330720 2858 330784
rect 2922 330720 2930 330784
rect 2610 330719 2930 330720
rect 5944 330784 6264 330785
rect 5944 330720 5952 330784
rect 6016 330720 6032 330784
rect 6096 330720 6112 330784
rect 6176 330720 6192 330784
rect 6256 330720 6264 330784
rect 5944 330719 6264 330720
rect 4277 330240 4597 330241
rect 4277 330176 4285 330240
rect 4349 330176 4365 330240
rect 4429 330176 4445 330240
rect 4509 330176 4525 330240
rect 4589 330176 4597 330240
rect 4277 330175 4597 330176
rect 7610 330240 7930 330241
rect 7610 330176 7618 330240
rect 7682 330176 7698 330240
rect 7762 330176 7778 330240
rect 7842 330176 7858 330240
rect 7922 330176 7930 330240
rect 7610 330175 7930 330176
rect 2610 329696 2930 329697
rect 2610 329632 2618 329696
rect 2682 329632 2698 329696
rect 2762 329632 2778 329696
rect 2842 329632 2858 329696
rect 2922 329632 2930 329696
rect 2610 329631 2930 329632
rect 5944 329696 6264 329697
rect 5944 329632 5952 329696
rect 6016 329632 6032 329696
rect 6096 329632 6112 329696
rect 6176 329632 6192 329696
rect 6256 329632 6264 329696
rect 5944 329631 6264 329632
rect 4277 329152 4597 329153
rect 4277 329088 4285 329152
rect 4349 329088 4365 329152
rect 4429 329088 4445 329152
rect 4509 329088 4525 329152
rect 4589 329088 4597 329152
rect 4277 329087 4597 329088
rect 7610 329152 7930 329153
rect 7610 329088 7618 329152
rect 7682 329088 7698 329152
rect 7762 329088 7778 329152
rect 7842 329088 7858 329152
rect 7922 329088 7930 329152
rect 7610 329087 7930 329088
rect 2610 328608 2930 328609
rect 2610 328544 2618 328608
rect 2682 328544 2698 328608
rect 2762 328544 2778 328608
rect 2842 328544 2858 328608
rect 2922 328544 2930 328608
rect 2610 328543 2930 328544
rect 5944 328608 6264 328609
rect 5944 328544 5952 328608
rect 6016 328544 6032 328608
rect 6096 328544 6112 328608
rect 6176 328544 6192 328608
rect 6256 328544 6264 328608
rect 5944 328543 6264 328544
rect 4277 328064 4597 328065
rect 4277 328000 4285 328064
rect 4349 328000 4365 328064
rect 4429 328000 4445 328064
rect 4509 328000 4525 328064
rect 4589 328000 4597 328064
rect 4277 327999 4597 328000
rect 7610 328064 7930 328065
rect 7610 328000 7618 328064
rect 7682 328000 7698 328064
rect 7762 328000 7778 328064
rect 7842 328000 7858 328064
rect 7922 328000 7930 328064
rect 7610 327999 7930 328000
rect 2610 327520 2930 327521
rect 2610 327456 2618 327520
rect 2682 327456 2698 327520
rect 2762 327456 2778 327520
rect 2842 327456 2858 327520
rect 2922 327456 2930 327520
rect 2610 327455 2930 327456
rect 5944 327520 6264 327521
rect 5944 327456 5952 327520
rect 6016 327456 6032 327520
rect 6096 327456 6112 327520
rect 6176 327456 6192 327520
rect 6256 327456 6264 327520
rect 5944 327455 6264 327456
rect 4277 326976 4597 326977
rect 4277 326912 4285 326976
rect 4349 326912 4365 326976
rect 4429 326912 4445 326976
rect 4509 326912 4525 326976
rect 4589 326912 4597 326976
rect 4277 326911 4597 326912
rect 7610 326976 7930 326977
rect 7610 326912 7618 326976
rect 7682 326912 7698 326976
rect 7762 326912 7778 326976
rect 7842 326912 7858 326976
rect 7922 326912 7930 326976
rect 7610 326911 7930 326912
rect 2610 326432 2930 326433
rect 2610 326368 2618 326432
rect 2682 326368 2698 326432
rect 2762 326368 2778 326432
rect 2842 326368 2858 326432
rect 2922 326368 2930 326432
rect 2610 326367 2930 326368
rect 5944 326432 6264 326433
rect 5944 326368 5952 326432
rect 6016 326368 6032 326432
rect 6096 326368 6112 326432
rect 6176 326368 6192 326432
rect 6256 326368 6264 326432
rect 5944 326367 6264 326368
rect 4277 325888 4597 325889
rect 4277 325824 4285 325888
rect 4349 325824 4365 325888
rect 4429 325824 4445 325888
rect 4509 325824 4525 325888
rect 4589 325824 4597 325888
rect 4277 325823 4597 325824
rect 7610 325888 7930 325889
rect 7610 325824 7618 325888
rect 7682 325824 7698 325888
rect 7762 325824 7778 325888
rect 7842 325824 7858 325888
rect 7922 325824 7930 325888
rect 7610 325823 7930 325824
rect 2610 325344 2930 325345
rect 2610 325280 2618 325344
rect 2682 325280 2698 325344
rect 2762 325280 2778 325344
rect 2842 325280 2858 325344
rect 2922 325280 2930 325344
rect 2610 325279 2930 325280
rect 5944 325344 6264 325345
rect 5944 325280 5952 325344
rect 6016 325280 6032 325344
rect 6096 325280 6112 325344
rect 6176 325280 6192 325344
rect 6256 325280 6264 325344
rect 5944 325279 6264 325280
rect 4277 324800 4597 324801
rect 4277 324736 4285 324800
rect 4349 324736 4365 324800
rect 4429 324736 4445 324800
rect 4509 324736 4525 324800
rect 4589 324736 4597 324800
rect 4277 324735 4597 324736
rect 7610 324800 7930 324801
rect 7610 324736 7618 324800
rect 7682 324736 7698 324800
rect 7762 324736 7778 324800
rect 7842 324736 7858 324800
rect 7922 324736 7930 324800
rect 7610 324735 7930 324736
rect 2610 324256 2930 324257
rect 2610 324192 2618 324256
rect 2682 324192 2698 324256
rect 2762 324192 2778 324256
rect 2842 324192 2858 324256
rect 2922 324192 2930 324256
rect 2610 324191 2930 324192
rect 5944 324256 6264 324257
rect 5944 324192 5952 324256
rect 6016 324192 6032 324256
rect 6096 324192 6112 324256
rect 6176 324192 6192 324256
rect 6256 324192 6264 324256
rect 5944 324191 6264 324192
rect 4277 323712 4597 323713
rect 4277 323648 4285 323712
rect 4349 323648 4365 323712
rect 4429 323648 4445 323712
rect 4509 323648 4525 323712
rect 4589 323648 4597 323712
rect 4277 323647 4597 323648
rect 7610 323712 7930 323713
rect 7610 323648 7618 323712
rect 7682 323648 7698 323712
rect 7762 323648 7778 323712
rect 7842 323648 7858 323712
rect 7922 323648 7930 323712
rect 7610 323647 7930 323648
rect 2610 323168 2930 323169
rect 2610 323104 2618 323168
rect 2682 323104 2698 323168
rect 2762 323104 2778 323168
rect 2842 323104 2858 323168
rect 2922 323104 2930 323168
rect 2610 323103 2930 323104
rect 5944 323168 6264 323169
rect 5944 323104 5952 323168
rect 6016 323104 6032 323168
rect 6096 323104 6112 323168
rect 6176 323104 6192 323168
rect 6256 323104 6264 323168
rect 5944 323103 6264 323104
rect 4277 322624 4597 322625
rect 4277 322560 4285 322624
rect 4349 322560 4365 322624
rect 4429 322560 4445 322624
rect 4509 322560 4525 322624
rect 4589 322560 4597 322624
rect 4277 322559 4597 322560
rect 7610 322624 7930 322625
rect 7610 322560 7618 322624
rect 7682 322560 7698 322624
rect 7762 322560 7778 322624
rect 7842 322560 7858 322624
rect 7922 322560 7930 322624
rect 7610 322559 7930 322560
rect 2610 322080 2930 322081
rect 2610 322016 2618 322080
rect 2682 322016 2698 322080
rect 2762 322016 2778 322080
rect 2842 322016 2858 322080
rect 2922 322016 2930 322080
rect 2610 322015 2930 322016
rect 5944 322080 6264 322081
rect 5944 322016 5952 322080
rect 6016 322016 6032 322080
rect 6096 322016 6112 322080
rect 6176 322016 6192 322080
rect 6256 322016 6264 322080
rect 5944 322015 6264 322016
rect 4277 321536 4597 321537
rect 4277 321472 4285 321536
rect 4349 321472 4365 321536
rect 4429 321472 4445 321536
rect 4509 321472 4525 321536
rect 4589 321472 4597 321536
rect 4277 321471 4597 321472
rect 7610 321536 7930 321537
rect 7610 321472 7618 321536
rect 7682 321472 7698 321536
rect 7762 321472 7778 321536
rect 7842 321472 7858 321536
rect 7922 321472 7930 321536
rect 7610 321471 7930 321472
rect 2610 320992 2930 320993
rect 2610 320928 2618 320992
rect 2682 320928 2698 320992
rect 2762 320928 2778 320992
rect 2842 320928 2858 320992
rect 2922 320928 2930 320992
rect 2610 320927 2930 320928
rect 5944 320992 6264 320993
rect 5944 320928 5952 320992
rect 6016 320928 6032 320992
rect 6096 320928 6112 320992
rect 6176 320928 6192 320992
rect 6256 320928 6264 320992
rect 5944 320927 6264 320928
rect 4277 320448 4597 320449
rect 4277 320384 4285 320448
rect 4349 320384 4365 320448
rect 4429 320384 4445 320448
rect 4509 320384 4525 320448
rect 4589 320384 4597 320448
rect 4277 320383 4597 320384
rect 7610 320448 7930 320449
rect 7610 320384 7618 320448
rect 7682 320384 7698 320448
rect 7762 320384 7778 320448
rect 7842 320384 7858 320448
rect 7922 320384 7930 320448
rect 7610 320383 7930 320384
rect 2610 319904 2930 319905
rect 2610 319840 2618 319904
rect 2682 319840 2698 319904
rect 2762 319840 2778 319904
rect 2842 319840 2858 319904
rect 2922 319840 2930 319904
rect 2610 319839 2930 319840
rect 5944 319904 6264 319905
rect 5944 319840 5952 319904
rect 6016 319840 6032 319904
rect 6096 319840 6112 319904
rect 6176 319840 6192 319904
rect 6256 319840 6264 319904
rect 5944 319839 6264 319840
rect 4277 319360 4597 319361
rect 4277 319296 4285 319360
rect 4349 319296 4365 319360
rect 4429 319296 4445 319360
rect 4509 319296 4525 319360
rect 4589 319296 4597 319360
rect 4277 319295 4597 319296
rect 7610 319360 7930 319361
rect 7610 319296 7618 319360
rect 7682 319296 7698 319360
rect 7762 319296 7778 319360
rect 7842 319296 7858 319360
rect 7922 319296 7930 319360
rect 7610 319295 7930 319296
rect 2610 318816 2930 318817
rect 2610 318752 2618 318816
rect 2682 318752 2698 318816
rect 2762 318752 2778 318816
rect 2842 318752 2858 318816
rect 2922 318752 2930 318816
rect 2610 318751 2930 318752
rect 5944 318816 6264 318817
rect 5944 318752 5952 318816
rect 6016 318752 6032 318816
rect 6096 318752 6112 318816
rect 6176 318752 6192 318816
rect 6256 318752 6264 318816
rect 5944 318751 6264 318752
rect 4277 318272 4597 318273
rect 4277 318208 4285 318272
rect 4349 318208 4365 318272
rect 4429 318208 4445 318272
rect 4509 318208 4525 318272
rect 4589 318208 4597 318272
rect 4277 318207 4597 318208
rect 7610 318272 7930 318273
rect 7610 318208 7618 318272
rect 7682 318208 7698 318272
rect 7762 318208 7778 318272
rect 7842 318208 7858 318272
rect 7922 318208 7930 318272
rect 7610 318207 7930 318208
rect 2610 317728 2930 317729
rect 2610 317664 2618 317728
rect 2682 317664 2698 317728
rect 2762 317664 2778 317728
rect 2842 317664 2858 317728
rect 2922 317664 2930 317728
rect 2610 317663 2930 317664
rect 5944 317728 6264 317729
rect 5944 317664 5952 317728
rect 6016 317664 6032 317728
rect 6096 317664 6112 317728
rect 6176 317664 6192 317728
rect 6256 317664 6264 317728
rect 5944 317663 6264 317664
rect 4277 317184 4597 317185
rect 4277 317120 4285 317184
rect 4349 317120 4365 317184
rect 4429 317120 4445 317184
rect 4509 317120 4525 317184
rect 4589 317120 4597 317184
rect 4277 317119 4597 317120
rect 7610 317184 7930 317185
rect 7610 317120 7618 317184
rect 7682 317120 7698 317184
rect 7762 317120 7778 317184
rect 7842 317120 7858 317184
rect 7922 317120 7930 317184
rect 7610 317119 7930 317120
rect 2610 316640 2930 316641
rect 2610 316576 2618 316640
rect 2682 316576 2698 316640
rect 2762 316576 2778 316640
rect 2842 316576 2858 316640
rect 2922 316576 2930 316640
rect 2610 316575 2930 316576
rect 5944 316640 6264 316641
rect 5944 316576 5952 316640
rect 6016 316576 6032 316640
rect 6096 316576 6112 316640
rect 6176 316576 6192 316640
rect 6256 316576 6264 316640
rect 5944 316575 6264 316576
rect 9520 316344 10000 316464
rect 4277 316096 4597 316097
rect 4277 316032 4285 316096
rect 4349 316032 4365 316096
rect 4429 316032 4445 316096
rect 4509 316032 4525 316096
rect 4589 316032 4597 316096
rect 4277 316031 4597 316032
rect 7610 316096 7930 316097
rect 7610 316032 7618 316096
rect 7682 316032 7698 316096
rect 7762 316032 7778 316096
rect 7842 316032 7858 316096
rect 7922 316032 7930 316096
rect 7610 316031 7930 316032
rect 7281 315890 7347 315893
rect 9630 315890 9690 316344
rect 7281 315888 9690 315890
rect 7281 315832 7286 315888
rect 7342 315832 9690 315888
rect 7281 315830 9690 315832
rect 7281 315827 7347 315830
rect 2610 315552 2930 315553
rect 2610 315488 2618 315552
rect 2682 315488 2698 315552
rect 2762 315488 2778 315552
rect 2842 315488 2858 315552
rect 2922 315488 2930 315552
rect 2610 315487 2930 315488
rect 5944 315552 6264 315553
rect 5944 315488 5952 315552
rect 6016 315488 6032 315552
rect 6096 315488 6112 315552
rect 6176 315488 6192 315552
rect 6256 315488 6264 315552
rect 5944 315487 6264 315488
rect 4277 315008 4597 315009
rect 4277 314944 4285 315008
rect 4349 314944 4365 315008
rect 4429 314944 4445 315008
rect 4509 314944 4525 315008
rect 4589 314944 4597 315008
rect 4277 314943 4597 314944
rect 7610 315008 7930 315009
rect 7610 314944 7618 315008
rect 7682 314944 7698 315008
rect 7762 314944 7778 315008
rect 7842 314944 7858 315008
rect 7922 314944 7930 315008
rect 7610 314943 7930 314944
rect 2610 314464 2930 314465
rect 2610 314400 2618 314464
rect 2682 314400 2698 314464
rect 2762 314400 2778 314464
rect 2842 314400 2858 314464
rect 2922 314400 2930 314464
rect 2610 314399 2930 314400
rect 5944 314464 6264 314465
rect 5944 314400 5952 314464
rect 6016 314400 6032 314464
rect 6096 314400 6112 314464
rect 6176 314400 6192 314464
rect 6256 314400 6264 314464
rect 5944 314399 6264 314400
rect 4277 313920 4597 313921
rect 4277 313856 4285 313920
rect 4349 313856 4365 313920
rect 4429 313856 4445 313920
rect 4509 313856 4525 313920
rect 4589 313856 4597 313920
rect 4277 313855 4597 313856
rect 7610 313920 7930 313921
rect 7610 313856 7618 313920
rect 7682 313856 7698 313920
rect 7762 313856 7778 313920
rect 7842 313856 7858 313920
rect 7922 313856 7930 313920
rect 7610 313855 7930 313856
rect 2610 313376 2930 313377
rect 2610 313312 2618 313376
rect 2682 313312 2698 313376
rect 2762 313312 2778 313376
rect 2842 313312 2858 313376
rect 2922 313312 2930 313376
rect 2610 313311 2930 313312
rect 5944 313376 6264 313377
rect 5944 313312 5952 313376
rect 6016 313312 6032 313376
rect 6096 313312 6112 313376
rect 6176 313312 6192 313376
rect 6256 313312 6264 313376
rect 5944 313311 6264 313312
rect 4277 312832 4597 312833
rect 4277 312768 4285 312832
rect 4349 312768 4365 312832
rect 4429 312768 4445 312832
rect 4509 312768 4525 312832
rect 4589 312768 4597 312832
rect 4277 312767 4597 312768
rect 7610 312832 7930 312833
rect 7610 312768 7618 312832
rect 7682 312768 7698 312832
rect 7762 312768 7778 312832
rect 7842 312768 7858 312832
rect 7922 312768 7930 312832
rect 7610 312767 7930 312768
rect 2610 312288 2930 312289
rect 2610 312224 2618 312288
rect 2682 312224 2698 312288
rect 2762 312224 2778 312288
rect 2842 312224 2858 312288
rect 2922 312224 2930 312288
rect 2610 312223 2930 312224
rect 5944 312288 6264 312289
rect 5944 312224 5952 312288
rect 6016 312224 6032 312288
rect 6096 312224 6112 312288
rect 6176 312224 6192 312288
rect 6256 312224 6264 312288
rect 5944 312223 6264 312224
rect 4277 311744 4597 311745
rect 4277 311680 4285 311744
rect 4349 311680 4365 311744
rect 4429 311680 4445 311744
rect 4509 311680 4525 311744
rect 4589 311680 4597 311744
rect 4277 311679 4597 311680
rect 7610 311744 7930 311745
rect 7610 311680 7618 311744
rect 7682 311680 7698 311744
rect 7762 311680 7778 311744
rect 7842 311680 7858 311744
rect 7922 311680 7930 311744
rect 7610 311679 7930 311680
rect 2610 311200 2930 311201
rect 2610 311136 2618 311200
rect 2682 311136 2698 311200
rect 2762 311136 2778 311200
rect 2842 311136 2858 311200
rect 2922 311136 2930 311200
rect 2610 311135 2930 311136
rect 5944 311200 6264 311201
rect 5944 311136 5952 311200
rect 6016 311136 6032 311200
rect 6096 311136 6112 311200
rect 6176 311136 6192 311200
rect 6256 311136 6264 311200
rect 5944 311135 6264 311136
rect 4277 310656 4597 310657
rect 4277 310592 4285 310656
rect 4349 310592 4365 310656
rect 4429 310592 4445 310656
rect 4509 310592 4525 310656
rect 4589 310592 4597 310656
rect 4277 310591 4597 310592
rect 7610 310656 7930 310657
rect 7610 310592 7618 310656
rect 7682 310592 7698 310656
rect 7762 310592 7778 310656
rect 7842 310592 7858 310656
rect 7922 310592 7930 310656
rect 7610 310591 7930 310592
rect 2610 310112 2930 310113
rect 2610 310048 2618 310112
rect 2682 310048 2698 310112
rect 2762 310048 2778 310112
rect 2842 310048 2858 310112
rect 2922 310048 2930 310112
rect 2610 310047 2930 310048
rect 5944 310112 6264 310113
rect 5944 310048 5952 310112
rect 6016 310048 6032 310112
rect 6096 310048 6112 310112
rect 6176 310048 6192 310112
rect 6256 310048 6264 310112
rect 5944 310047 6264 310048
rect 4277 309568 4597 309569
rect 4277 309504 4285 309568
rect 4349 309504 4365 309568
rect 4429 309504 4445 309568
rect 4509 309504 4525 309568
rect 4589 309504 4597 309568
rect 4277 309503 4597 309504
rect 7610 309568 7930 309569
rect 7610 309504 7618 309568
rect 7682 309504 7698 309568
rect 7762 309504 7778 309568
rect 7842 309504 7858 309568
rect 7922 309504 7930 309568
rect 7610 309503 7930 309504
rect 0 309136 480 309256
rect 62 308682 122 309136
rect 2610 309024 2930 309025
rect 2610 308960 2618 309024
rect 2682 308960 2698 309024
rect 2762 308960 2778 309024
rect 2842 308960 2858 309024
rect 2922 308960 2930 309024
rect 2610 308959 2930 308960
rect 5944 309024 6264 309025
rect 5944 308960 5952 309024
rect 6016 308960 6032 309024
rect 6096 308960 6112 309024
rect 6176 308960 6192 309024
rect 6256 308960 6264 309024
rect 5944 308959 6264 308960
rect 2221 308682 2287 308685
rect 62 308680 2287 308682
rect 62 308624 2226 308680
rect 2282 308624 2287 308680
rect 62 308622 2287 308624
rect 2221 308619 2287 308622
rect 4277 308480 4597 308481
rect 4277 308416 4285 308480
rect 4349 308416 4365 308480
rect 4429 308416 4445 308480
rect 4509 308416 4525 308480
rect 4589 308416 4597 308480
rect 4277 308415 4597 308416
rect 7610 308480 7930 308481
rect 7610 308416 7618 308480
rect 7682 308416 7698 308480
rect 7762 308416 7778 308480
rect 7842 308416 7858 308480
rect 7922 308416 7930 308480
rect 7610 308415 7930 308416
rect 2610 307936 2930 307937
rect 2610 307872 2618 307936
rect 2682 307872 2698 307936
rect 2762 307872 2778 307936
rect 2842 307872 2858 307936
rect 2922 307872 2930 307936
rect 2610 307871 2930 307872
rect 5944 307936 6264 307937
rect 5944 307872 5952 307936
rect 6016 307872 6032 307936
rect 6096 307872 6112 307936
rect 6176 307872 6192 307936
rect 6256 307872 6264 307936
rect 5944 307871 6264 307872
rect 4277 307392 4597 307393
rect 4277 307328 4285 307392
rect 4349 307328 4365 307392
rect 4429 307328 4445 307392
rect 4509 307328 4525 307392
rect 4589 307328 4597 307392
rect 4277 307327 4597 307328
rect 7610 307392 7930 307393
rect 7610 307328 7618 307392
rect 7682 307328 7698 307392
rect 7762 307328 7778 307392
rect 7842 307328 7858 307392
rect 7922 307328 7930 307392
rect 7610 307327 7930 307328
rect 2610 306848 2930 306849
rect 2610 306784 2618 306848
rect 2682 306784 2698 306848
rect 2762 306784 2778 306848
rect 2842 306784 2858 306848
rect 2922 306784 2930 306848
rect 2610 306783 2930 306784
rect 5944 306848 6264 306849
rect 5944 306784 5952 306848
rect 6016 306784 6032 306848
rect 6096 306784 6112 306848
rect 6176 306784 6192 306848
rect 6256 306784 6264 306848
rect 5944 306783 6264 306784
rect 4277 306304 4597 306305
rect 4277 306240 4285 306304
rect 4349 306240 4365 306304
rect 4429 306240 4445 306304
rect 4509 306240 4525 306304
rect 4589 306240 4597 306304
rect 4277 306239 4597 306240
rect 7610 306304 7930 306305
rect 7610 306240 7618 306304
rect 7682 306240 7698 306304
rect 7762 306240 7778 306304
rect 7842 306240 7858 306304
rect 7922 306240 7930 306304
rect 7610 306239 7930 306240
rect 2610 305760 2930 305761
rect 2610 305696 2618 305760
rect 2682 305696 2698 305760
rect 2762 305696 2778 305760
rect 2842 305696 2858 305760
rect 2922 305696 2930 305760
rect 2610 305695 2930 305696
rect 5944 305760 6264 305761
rect 5944 305696 5952 305760
rect 6016 305696 6032 305760
rect 6096 305696 6112 305760
rect 6176 305696 6192 305760
rect 6256 305696 6264 305760
rect 5944 305695 6264 305696
rect 4277 305216 4597 305217
rect 4277 305152 4285 305216
rect 4349 305152 4365 305216
rect 4429 305152 4445 305216
rect 4509 305152 4525 305216
rect 4589 305152 4597 305216
rect 4277 305151 4597 305152
rect 7610 305216 7930 305217
rect 7610 305152 7618 305216
rect 7682 305152 7698 305216
rect 7762 305152 7778 305216
rect 7842 305152 7858 305216
rect 7922 305152 7930 305216
rect 7610 305151 7930 305152
rect 2610 304672 2930 304673
rect 2610 304608 2618 304672
rect 2682 304608 2698 304672
rect 2762 304608 2778 304672
rect 2842 304608 2858 304672
rect 2922 304608 2930 304672
rect 2610 304607 2930 304608
rect 5944 304672 6264 304673
rect 5944 304608 5952 304672
rect 6016 304608 6032 304672
rect 6096 304608 6112 304672
rect 6176 304608 6192 304672
rect 6256 304608 6264 304672
rect 5944 304607 6264 304608
rect 4277 304128 4597 304129
rect 4277 304064 4285 304128
rect 4349 304064 4365 304128
rect 4429 304064 4445 304128
rect 4509 304064 4525 304128
rect 4589 304064 4597 304128
rect 4277 304063 4597 304064
rect 7610 304128 7930 304129
rect 7610 304064 7618 304128
rect 7682 304064 7698 304128
rect 7762 304064 7778 304128
rect 7842 304064 7858 304128
rect 7922 304064 7930 304128
rect 7610 304063 7930 304064
rect 2610 303584 2930 303585
rect 2610 303520 2618 303584
rect 2682 303520 2698 303584
rect 2762 303520 2778 303584
rect 2842 303520 2858 303584
rect 2922 303520 2930 303584
rect 2610 303519 2930 303520
rect 5944 303584 6264 303585
rect 5944 303520 5952 303584
rect 6016 303520 6032 303584
rect 6096 303520 6112 303584
rect 6176 303520 6192 303584
rect 6256 303520 6264 303584
rect 5944 303519 6264 303520
rect 4277 303040 4597 303041
rect 4277 302976 4285 303040
rect 4349 302976 4365 303040
rect 4429 302976 4445 303040
rect 4509 302976 4525 303040
rect 4589 302976 4597 303040
rect 4277 302975 4597 302976
rect 7610 303040 7930 303041
rect 7610 302976 7618 303040
rect 7682 302976 7698 303040
rect 7762 302976 7778 303040
rect 7842 302976 7858 303040
rect 7922 302976 7930 303040
rect 7610 302975 7930 302976
rect 2610 302496 2930 302497
rect 2610 302432 2618 302496
rect 2682 302432 2698 302496
rect 2762 302432 2778 302496
rect 2842 302432 2858 302496
rect 2922 302432 2930 302496
rect 2610 302431 2930 302432
rect 5944 302496 6264 302497
rect 5944 302432 5952 302496
rect 6016 302432 6032 302496
rect 6096 302432 6112 302496
rect 6176 302432 6192 302496
rect 6256 302432 6264 302496
rect 5944 302431 6264 302432
rect 4277 301952 4597 301953
rect 4277 301888 4285 301952
rect 4349 301888 4365 301952
rect 4429 301888 4445 301952
rect 4509 301888 4525 301952
rect 4589 301888 4597 301952
rect 4277 301887 4597 301888
rect 7610 301952 7930 301953
rect 7610 301888 7618 301952
rect 7682 301888 7698 301952
rect 7762 301888 7778 301952
rect 7842 301888 7858 301952
rect 7922 301888 7930 301952
rect 7610 301887 7930 301888
rect 2610 301408 2930 301409
rect 2610 301344 2618 301408
rect 2682 301344 2698 301408
rect 2762 301344 2778 301408
rect 2842 301344 2858 301408
rect 2922 301344 2930 301408
rect 2610 301343 2930 301344
rect 5944 301408 6264 301409
rect 5944 301344 5952 301408
rect 6016 301344 6032 301408
rect 6096 301344 6112 301408
rect 6176 301344 6192 301408
rect 6256 301344 6264 301408
rect 5944 301343 6264 301344
rect 4277 300864 4597 300865
rect 4277 300800 4285 300864
rect 4349 300800 4365 300864
rect 4429 300800 4445 300864
rect 4509 300800 4525 300864
rect 4589 300800 4597 300864
rect 4277 300799 4597 300800
rect 7610 300864 7930 300865
rect 7610 300800 7618 300864
rect 7682 300800 7698 300864
rect 7762 300800 7778 300864
rect 7842 300800 7858 300864
rect 7922 300800 7930 300864
rect 7610 300799 7930 300800
rect 2610 300320 2930 300321
rect 2610 300256 2618 300320
rect 2682 300256 2698 300320
rect 2762 300256 2778 300320
rect 2842 300256 2858 300320
rect 2922 300256 2930 300320
rect 2610 300255 2930 300256
rect 5944 300320 6264 300321
rect 5944 300256 5952 300320
rect 6016 300256 6032 300320
rect 6096 300256 6112 300320
rect 6176 300256 6192 300320
rect 6256 300256 6264 300320
rect 5944 300255 6264 300256
rect 4277 299776 4597 299777
rect 4277 299712 4285 299776
rect 4349 299712 4365 299776
rect 4429 299712 4445 299776
rect 4509 299712 4525 299776
rect 4589 299712 4597 299776
rect 4277 299711 4597 299712
rect 7610 299776 7930 299777
rect 7610 299712 7618 299776
rect 7682 299712 7698 299776
rect 7762 299712 7778 299776
rect 7842 299712 7858 299776
rect 7922 299712 7930 299776
rect 7610 299711 7930 299712
rect 2610 299232 2930 299233
rect 2610 299168 2618 299232
rect 2682 299168 2698 299232
rect 2762 299168 2778 299232
rect 2842 299168 2858 299232
rect 2922 299168 2930 299232
rect 2610 299167 2930 299168
rect 5944 299232 6264 299233
rect 5944 299168 5952 299232
rect 6016 299168 6032 299232
rect 6096 299168 6112 299232
rect 6176 299168 6192 299232
rect 6256 299168 6264 299232
rect 5944 299167 6264 299168
rect 4277 298688 4597 298689
rect 4277 298624 4285 298688
rect 4349 298624 4365 298688
rect 4429 298624 4445 298688
rect 4509 298624 4525 298688
rect 4589 298624 4597 298688
rect 4277 298623 4597 298624
rect 7610 298688 7930 298689
rect 7610 298624 7618 298688
rect 7682 298624 7698 298688
rect 7762 298624 7778 298688
rect 7842 298624 7858 298688
rect 7922 298624 7930 298688
rect 7610 298623 7930 298624
rect 2610 298144 2930 298145
rect 2610 298080 2618 298144
rect 2682 298080 2698 298144
rect 2762 298080 2778 298144
rect 2842 298080 2858 298144
rect 2922 298080 2930 298144
rect 2610 298079 2930 298080
rect 5944 298144 6264 298145
rect 5944 298080 5952 298144
rect 6016 298080 6032 298144
rect 6096 298080 6112 298144
rect 6176 298080 6192 298144
rect 6256 298080 6264 298144
rect 5944 298079 6264 298080
rect 4277 297600 4597 297601
rect 4277 297536 4285 297600
rect 4349 297536 4365 297600
rect 4429 297536 4445 297600
rect 4509 297536 4525 297600
rect 4589 297536 4597 297600
rect 4277 297535 4597 297536
rect 7610 297600 7930 297601
rect 7610 297536 7618 297600
rect 7682 297536 7698 297600
rect 7762 297536 7778 297600
rect 7842 297536 7858 297600
rect 7922 297536 7930 297600
rect 7610 297535 7930 297536
rect 2610 297056 2930 297057
rect 2610 296992 2618 297056
rect 2682 296992 2698 297056
rect 2762 296992 2778 297056
rect 2842 296992 2858 297056
rect 2922 296992 2930 297056
rect 2610 296991 2930 296992
rect 5944 297056 6264 297057
rect 5944 296992 5952 297056
rect 6016 296992 6032 297056
rect 6096 296992 6112 297056
rect 6176 296992 6192 297056
rect 6256 296992 6264 297056
rect 5944 296991 6264 296992
rect 4277 296512 4597 296513
rect 4277 296448 4285 296512
rect 4349 296448 4365 296512
rect 4429 296448 4445 296512
rect 4509 296448 4525 296512
rect 4589 296448 4597 296512
rect 4277 296447 4597 296448
rect 7610 296512 7930 296513
rect 7610 296448 7618 296512
rect 7682 296448 7698 296512
rect 7762 296448 7778 296512
rect 7842 296448 7858 296512
rect 7922 296448 7930 296512
rect 7610 296447 7930 296448
rect 2610 295968 2930 295969
rect 2610 295904 2618 295968
rect 2682 295904 2698 295968
rect 2762 295904 2778 295968
rect 2842 295904 2858 295968
rect 2922 295904 2930 295968
rect 2610 295903 2930 295904
rect 5944 295968 6264 295969
rect 5944 295904 5952 295968
rect 6016 295904 6032 295968
rect 6096 295904 6112 295968
rect 6176 295904 6192 295968
rect 6256 295904 6264 295968
rect 5944 295903 6264 295904
rect 4277 295424 4597 295425
rect 4277 295360 4285 295424
rect 4349 295360 4365 295424
rect 4429 295360 4445 295424
rect 4509 295360 4525 295424
rect 4589 295360 4597 295424
rect 4277 295359 4597 295360
rect 7610 295424 7930 295425
rect 7610 295360 7618 295424
rect 7682 295360 7698 295424
rect 7762 295360 7778 295424
rect 7842 295360 7858 295424
rect 7922 295360 7930 295424
rect 7610 295359 7930 295360
rect 2610 294880 2930 294881
rect 2610 294816 2618 294880
rect 2682 294816 2698 294880
rect 2762 294816 2778 294880
rect 2842 294816 2858 294880
rect 2922 294816 2930 294880
rect 2610 294815 2930 294816
rect 5944 294880 6264 294881
rect 5944 294816 5952 294880
rect 6016 294816 6032 294880
rect 6096 294816 6112 294880
rect 6176 294816 6192 294880
rect 6256 294816 6264 294880
rect 5944 294815 6264 294816
rect 4277 294336 4597 294337
rect 4277 294272 4285 294336
rect 4349 294272 4365 294336
rect 4429 294272 4445 294336
rect 4509 294272 4525 294336
rect 4589 294272 4597 294336
rect 4277 294271 4597 294272
rect 7610 294336 7930 294337
rect 7610 294272 7618 294336
rect 7682 294272 7698 294336
rect 7762 294272 7778 294336
rect 7842 294272 7858 294336
rect 7922 294272 7930 294336
rect 7610 294271 7930 294272
rect 2610 293792 2930 293793
rect 2610 293728 2618 293792
rect 2682 293728 2698 293792
rect 2762 293728 2778 293792
rect 2842 293728 2858 293792
rect 2922 293728 2930 293792
rect 2610 293727 2930 293728
rect 5944 293792 6264 293793
rect 5944 293728 5952 293792
rect 6016 293728 6032 293792
rect 6096 293728 6112 293792
rect 6176 293728 6192 293792
rect 6256 293728 6264 293792
rect 5944 293727 6264 293728
rect 4277 293248 4597 293249
rect 4277 293184 4285 293248
rect 4349 293184 4365 293248
rect 4429 293184 4445 293248
rect 4509 293184 4525 293248
rect 4589 293184 4597 293248
rect 4277 293183 4597 293184
rect 7610 293248 7930 293249
rect 7610 293184 7618 293248
rect 7682 293184 7698 293248
rect 7762 293184 7778 293248
rect 7842 293184 7858 293248
rect 7922 293184 7930 293248
rect 7610 293183 7930 293184
rect 2610 292704 2930 292705
rect 2610 292640 2618 292704
rect 2682 292640 2698 292704
rect 2762 292640 2778 292704
rect 2842 292640 2858 292704
rect 2922 292640 2930 292704
rect 2610 292639 2930 292640
rect 5944 292704 6264 292705
rect 5944 292640 5952 292704
rect 6016 292640 6032 292704
rect 6096 292640 6112 292704
rect 6176 292640 6192 292704
rect 6256 292640 6264 292704
rect 5944 292639 6264 292640
rect 4277 292160 4597 292161
rect 4277 292096 4285 292160
rect 4349 292096 4365 292160
rect 4429 292096 4445 292160
rect 4509 292096 4525 292160
rect 4589 292096 4597 292160
rect 4277 292095 4597 292096
rect 7610 292160 7930 292161
rect 7610 292096 7618 292160
rect 7682 292096 7698 292160
rect 7762 292096 7778 292160
rect 7842 292096 7858 292160
rect 7922 292096 7930 292160
rect 7610 292095 7930 292096
rect 2610 291616 2930 291617
rect 2610 291552 2618 291616
rect 2682 291552 2698 291616
rect 2762 291552 2778 291616
rect 2842 291552 2858 291616
rect 2922 291552 2930 291616
rect 2610 291551 2930 291552
rect 5944 291616 6264 291617
rect 5944 291552 5952 291616
rect 6016 291552 6032 291616
rect 6096 291552 6112 291616
rect 6176 291552 6192 291616
rect 6256 291552 6264 291616
rect 5944 291551 6264 291552
rect 4277 291072 4597 291073
rect 4277 291008 4285 291072
rect 4349 291008 4365 291072
rect 4429 291008 4445 291072
rect 4509 291008 4525 291072
rect 4589 291008 4597 291072
rect 4277 291007 4597 291008
rect 7610 291072 7930 291073
rect 7610 291008 7618 291072
rect 7682 291008 7698 291072
rect 7762 291008 7778 291072
rect 7842 291008 7858 291072
rect 7922 291008 7930 291072
rect 7610 291007 7930 291008
rect 2610 290528 2930 290529
rect 2610 290464 2618 290528
rect 2682 290464 2698 290528
rect 2762 290464 2778 290528
rect 2842 290464 2858 290528
rect 2922 290464 2930 290528
rect 2610 290463 2930 290464
rect 5944 290528 6264 290529
rect 5944 290464 5952 290528
rect 6016 290464 6032 290528
rect 6096 290464 6112 290528
rect 6176 290464 6192 290528
rect 6256 290464 6264 290528
rect 5944 290463 6264 290464
rect 4277 289984 4597 289985
rect 4277 289920 4285 289984
rect 4349 289920 4365 289984
rect 4429 289920 4445 289984
rect 4509 289920 4525 289984
rect 4589 289920 4597 289984
rect 4277 289919 4597 289920
rect 7610 289984 7930 289985
rect 7610 289920 7618 289984
rect 7682 289920 7698 289984
rect 7762 289920 7778 289984
rect 7842 289920 7858 289984
rect 7922 289920 7930 289984
rect 7610 289919 7930 289920
rect 2610 289440 2930 289441
rect 2610 289376 2618 289440
rect 2682 289376 2698 289440
rect 2762 289376 2778 289440
rect 2842 289376 2858 289440
rect 2922 289376 2930 289440
rect 2610 289375 2930 289376
rect 5944 289440 6264 289441
rect 5944 289376 5952 289440
rect 6016 289376 6032 289440
rect 6096 289376 6112 289440
rect 6176 289376 6192 289440
rect 6256 289376 6264 289440
rect 5944 289375 6264 289376
rect 4277 288896 4597 288897
rect 4277 288832 4285 288896
rect 4349 288832 4365 288896
rect 4429 288832 4445 288896
rect 4509 288832 4525 288896
rect 4589 288832 4597 288896
rect 4277 288831 4597 288832
rect 7610 288896 7930 288897
rect 7610 288832 7618 288896
rect 7682 288832 7698 288896
rect 7762 288832 7778 288896
rect 7842 288832 7858 288896
rect 7922 288832 7930 288896
rect 7610 288831 7930 288832
rect 2610 288352 2930 288353
rect 2610 288288 2618 288352
rect 2682 288288 2698 288352
rect 2762 288288 2778 288352
rect 2842 288288 2858 288352
rect 2922 288288 2930 288352
rect 2610 288287 2930 288288
rect 5944 288352 6264 288353
rect 5944 288288 5952 288352
rect 6016 288288 6032 288352
rect 6096 288288 6112 288352
rect 6176 288288 6192 288352
rect 6256 288288 6264 288352
rect 5944 288287 6264 288288
rect 4277 287808 4597 287809
rect 4277 287744 4285 287808
rect 4349 287744 4365 287808
rect 4429 287744 4445 287808
rect 4509 287744 4525 287808
rect 4589 287744 4597 287808
rect 4277 287743 4597 287744
rect 7610 287808 7930 287809
rect 7610 287744 7618 287808
rect 7682 287744 7698 287808
rect 7762 287744 7778 287808
rect 7842 287744 7858 287808
rect 7922 287744 7930 287808
rect 7610 287743 7930 287744
rect 2610 287264 2930 287265
rect 2610 287200 2618 287264
rect 2682 287200 2698 287264
rect 2762 287200 2778 287264
rect 2842 287200 2858 287264
rect 2922 287200 2930 287264
rect 2610 287199 2930 287200
rect 5944 287264 6264 287265
rect 5944 287200 5952 287264
rect 6016 287200 6032 287264
rect 6096 287200 6112 287264
rect 6176 287200 6192 287264
rect 6256 287200 6264 287264
rect 5944 287199 6264 287200
rect 4277 286720 4597 286721
rect 4277 286656 4285 286720
rect 4349 286656 4365 286720
rect 4429 286656 4445 286720
rect 4509 286656 4525 286720
rect 4589 286656 4597 286720
rect 4277 286655 4597 286656
rect 7610 286720 7930 286721
rect 7610 286656 7618 286720
rect 7682 286656 7698 286720
rect 7762 286656 7778 286720
rect 7842 286656 7858 286720
rect 7922 286656 7930 286720
rect 7610 286655 7930 286656
rect 2610 286176 2930 286177
rect 2610 286112 2618 286176
rect 2682 286112 2698 286176
rect 2762 286112 2778 286176
rect 2842 286112 2858 286176
rect 2922 286112 2930 286176
rect 2610 286111 2930 286112
rect 5944 286176 6264 286177
rect 5944 286112 5952 286176
rect 6016 286112 6032 286176
rect 6096 286112 6112 286176
rect 6176 286112 6192 286176
rect 6256 286112 6264 286176
rect 5944 286111 6264 286112
rect 4277 285632 4597 285633
rect 4277 285568 4285 285632
rect 4349 285568 4365 285632
rect 4429 285568 4445 285632
rect 4509 285568 4525 285632
rect 4589 285568 4597 285632
rect 4277 285567 4597 285568
rect 7610 285632 7930 285633
rect 7610 285568 7618 285632
rect 7682 285568 7698 285632
rect 7762 285568 7778 285632
rect 7842 285568 7858 285632
rect 7922 285568 7930 285632
rect 7610 285567 7930 285568
rect 2610 285088 2930 285089
rect 2610 285024 2618 285088
rect 2682 285024 2698 285088
rect 2762 285024 2778 285088
rect 2842 285024 2858 285088
rect 2922 285024 2930 285088
rect 2610 285023 2930 285024
rect 5944 285088 6264 285089
rect 5944 285024 5952 285088
rect 6016 285024 6032 285088
rect 6096 285024 6112 285088
rect 6176 285024 6192 285088
rect 6256 285024 6264 285088
rect 5944 285023 6264 285024
rect 4277 284544 4597 284545
rect 4277 284480 4285 284544
rect 4349 284480 4365 284544
rect 4429 284480 4445 284544
rect 4509 284480 4525 284544
rect 4589 284480 4597 284544
rect 4277 284479 4597 284480
rect 7610 284544 7930 284545
rect 7610 284480 7618 284544
rect 7682 284480 7698 284544
rect 7762 284480 7778 284544
rect 7842 284480 7858 284544
rect 7922 284480 7930 284544
rect 7610 284479 7930 284480
rect 2610 284000 2930 284001
rect 2610 283936 2618 284000
rect 2682 283936 2698 284000
rect 2762 283936 2778 284000
rect 2842 283936 2858 284000
rect 2922 283936 2930 284000
rect 2610 283935 2930 283936
rect 5944 284000 6264 284001
rect 5944 283936 5952 284000
rect 6016 283936 6032 284000
rect 6096 283936 6112 284000
rect 6176 283936 6192 284000
rect 6256 283936 6264 284000
rect 5944 283935 6264 283936
rect 4277 283456 4597 283457
rect 4277 283392 4285 283456
rect 4349 283392 4365 283456
rect 4429 283392 4445 283456
rect 4509 283392 4525 283456
rect 4589 283392 4597 283456
rect 4277 283391 4597 283392
rect 7610 283456 7930 283457
rect 7610 283392 7618 283456
rect 7682 283392 7698 283456
rect 7762 283392 7778 283456
rect 7842 283392 7858 283456
rect 7922 283392 7930 283456
rect 7610 283391 7930 283392
rect 9520 283024 10000 283144
rect 2610 282912 2930 282913
rect 2610 282848 2618 282912
rect 2682 282848 2698 282912
rect 2762 282848 2778 282912
rect 2842 282848 2858 282912
rect 2922 282848 2930 282912
rect 2610 282847 2930 282848
rect 5944 282912 6264 282913
rect 5944 282848 5952 282912
rect 6016 282848 6032 282912
rect 6096 282848 6112 282912
rect 6176 282848 6192 282912
rect 6256 282848 6264 282912
rect 5944 282847 6264 282848
rect 6269 282570 6335 282573
rect 9630 282570 9690 283024
rect 6269 282568 9690 282570
rect 6269 282512 6274 282568
rect 6330 282512 9690 282568
rect 6269 282510 9690 282512
rect 6269 282507 6335 282510
rect 4277 282368 4597 282369
rect 4277 282304 4285 282368
rect 4349 282304 4365 282368
rect 4429 282304 4445 282368
rect 4509 282304 4525 282368
rect 4589 282304 4597 282368
rect 4277 282303 4597 282304
rect 7610 282368 7930 282369
rect 7610 282304 7618 282368
rect 7682 282304 7698 282368
rect 7762 282304 7778 282368
rect 7842 282304 7858 282368
rect 7922 282304 7930 282368
rect 7610 282303 7930 282304
rect 2610 281824 2930 281825
rect 2610 281760 2618 281824
rect 2682 281760 2698 281824
rect 2762 281760 2778 281824
rect 2842 281760 2858 281824
rect 2922 281760 2930 281824
rect 2610 281759 2930 281760
rect 5944 281824 6264 281825
rect 5944 281760 5952 281824
rect 6016 281760 6032 281824
rect 6096 281760 6112 281824
rect 6176 281760 6192 281824
rect 6256 281760 6264 281824
rect 5944 281759 6264 281760
rect 4277 281280 4597 281281
rect 4277 281216 4285 281280
rect 4349 281216 4365 281280
rect 4429 281216 4445 281280
rect 4509 281216 4525 281280
rect 4589 281216 4597 281280
rect 4277 281215 4597 281216
rect 7610 281280 7930 281281
rect 7610 281216 7618 281280
rect 7682 281216 7698 281280
rect 7762 281216 7778 281280
rect 7842 281216 7858 281280
rect 7922 281216 7930 281280
rect 7610 281215 7930 281216
rect 2610 280736 2930 280737
rect 2610 280672 2618 280736
rect 2682 280672 2698 280736
rect 2762 280672 2778 280736
rect 2842 280672 2858 280736
rect 2922 280672 2930 280736
rect 2610 280671 2930 280672
rect 5944 280736 6264 280737
rect 5944 280672 5952 280736
rect 6016 280672 6032 280736
rect 6096 280672 6112 280736
rect 6176 280672 6192 280736
rect 6256 280672 6264 280736
rect 5944 280671 6264 280672
rect 4277 280192 4597 280193
rect 4277 280128 4285 280192
rect 4349 280128 4365 280192
rect 4429 280128 4445 280192
rect 4509 280128 4525 280192
rect 4589 280128 4597 280192
rect 4277 280127 4597 280128
rect 7610 280192 7930 280193
rect 7610 280128 7618 280192
rect 7682 280128 7698 280192
rect 7762 280128 7778 280192
rect 7842 280128 7858 280192
rect 7922 280128 7930 280192
rect 7610 280127 7930 280128
rect 2610 279648 2930 279649
rect 2610 279584 2618 279648
rect 2682 279584 2698 279648
rect 2762 279584 2778 279648
rect 2842 279584 2858 279648
rect 2922 279584 2930 279648
rect 2610 279583 2930 279584
rect 5944 279648 6264 279649
rect 5944 279584 5952 279648
rect 6016 279584 6032 279648
rect 6096 279584 6112 279648
rect 6176 279584 6192 279648
rect 6256 279584 6264 279648
rect 5944 279583 6264 279584
rect 4277 279104 4597 279105
rect 4277 279040 4285 279104
rect 4349 279040 4365 279104
rect 4429 279040 4445 279104
rect 4509 279040 4525 279104
rect 4589 279040 4597 279104
rect 4277 279039 4597 279040
rect 7610 279104 7930 279105
rect 7610 279040 7618 279104
rect 7682 279040 7698 279104
rect 7762 279040 7778 279104
rect 7842 279040 7858 279104
rect 7922 279040 7930 279104
rect 7610 279039 7930 279040
rect 2610 278560 2930 278561
rect 2610 278496 2618 278560
rect 2682 278496 2698 278560
rect 2762 278496 2778 278560
rect 2842 278496 2858 278560
rect 2922 278496 2930 278560
rect 2610 278495 2930 278496
rect 5944 278560 6264 278561
rect 5944 278496 5952 278560
rect 6016 278496 6032 278560
rect 6096 278496 6112 278560
rect 6176 278496 6192 278560
rect 6256 278496 6264 278560
rect 5944 278495 6264 278496
rect 4277 278016 4597 278017
rect 4277 277952 4285 278016
rect 4349 277952 4365 278016
rect 4429 277952 4445 278016
rect 4509 277952 4525 278016
rect 4589 277952 4597 278016
rect 4277 277951 4597 277952
rect 7610 278016 7930 278017
rect 7610 277952 7618 278016
rect 7682 277952 7698 278016
rect 7762 277952 7778 278016
rect 7842 277952 7858 278016
rect 7922 277952 7930 278016
rect 7610 277951 7930 277952
rect 2610 277472 2930 277473
rect 2610 277408 2618 277472
rect 2682 277408 2698 277472
rect 2762 277408 2778 277472
rect 2842 277408 2858 277472
rect 2922 277408 2930 277472
rect 2610 277407 2930 277408
rect 5944 277472 6264 277473
rect 5944 277408 5952 277472
rect 6016 277408 6032 277472
rect 6096 277408 6112 277472
rect 6176 277408 6192 277472
rect 6256 277408 6264 277472
rect 5944 277407 6264 277408
rect 4277 276928 4597 276929
rect 4277 276864 4285 276928
rect 4349 276864 4365 276928
rect 4429 276864 4445 276928
rect 4509 276864 4525 276928
rect 4589 276864 4597 276928
rect 4277 276863 4597 276864
rect 7610 276928 7930 276929
rect 7610 276864 7618 276928
rect 7682 276864 7698 276928
rect 7762 276864 7778 276928
rect 7842 276864 7858 276928
rect 7922 276864 7930 276928
rect 7610 276863 7930 276864
rect 2610 276384 2930 276385
rect 2610 276320 2618 276384
rect 2682 276320 2698 276384
rect 2762 276320 2778 276384
rect 2842 276320 2858 276384
rect 2922 276320 2930 276384
rect 2610 276319 2930 276320
rect 5944 276384 6264 276385
rect 5944 276320 5952 276384
rect 6016 276320 6032 276384
rect 6096 276320 6112 276384
rect 6176 276320 6192 276384
rect 6256 276320 6264 276384
rect 5944 276319 6264 276320
rect 4277 275840 4597 275841
rect 4277 275776 4285 275840
rect 4349 275776 4365 275840
rect 4429 275776 4445 275840
rect 4509 275776 4525 275840
rect 4589 275776 4597 275840
rect 4277 275775 4597 275776
rect 7610 275840 7930 275841
rect 7610 275776 7618 275840
rect 7682 275776 7698 275840
rect 7762 275776 7778 275840
rect 7842 275776 7858 275840
rect 7922 275776 7930 275840
rect 7610 275775 7930 275776
rect 2610 275296 2930 275297
rect 2610 275232 2618 275296
rect 2682 275232 2698 275296
rect 2762 275232 2778 275296
rect 2842 275232 2858 275296
rect 2922 275232 2930 275296
rect 2610 275231 2930 275232
rect 5944 275296 6264 275297
rect 5944 275232 5952 275296
rect 6016 275232 6032 275296
rect 6096 275232 6112 275296
rect 6176 275232 6192 275296
rect 6256 275232 6264 275296
rect 5944 275231 6264 275232
rect 4277 274752 4597 274753
rect 4277 274688 4285 274752
rect 4349 274688 4365 274752
rect 4429 274688 4445 274752
rect 4509 274688 4525 274752
rect 4589 274688 4597 274752
rect 4277 274687 4597 274688
rect 7610 274752 7930 274753
rect 7610 274688 7618 274752
rect 7682 274688 7698 274752
rect 7762 274688 7778 274752
rect 7842 274688 7858 274752
rect 7922 274688 7930 274752
rect 7610 274687 7930 274688
rect 2610 274208 2930 274209
rect 2610 274144 2618 274208
rect 2682 274144 2698 274208
rect 2762 274144 2778 274208
rect 2842 274144 2858 274208
rect 2922 274144 2930 274208
rect 2610 274143 2930 274144
rect 5944 274208 6264 274209
rect 5944 274144 5952 274208
rect 6016 274144 6032 274208
rect 6096 274144 6112 274208
rect 6176 274144 6192 274208
rect 6256 274144 6264 274208
rect 5944 274143 6264 274144
rect 4277 273664 4597 273665
rect 4277 273600 4285 273664
rect 4349 273600 4365 273664
rect 4429 273600 4445 273664
rect 4509 273600 4525 273664
rect 4589 273600 4597 273664
rect 4277 273599 4597 273600
rect 7610 273664 7930 273665
rect 7610 273600 7618 273664
rect 7682 273600 7698 273664
rect 7762 273600 7778 273664
rect 7842 273600 7858 273664
rect 7922 273600 7930 273664
rect 7610 273599 7930 273600
rect 2610 273120 2930 273121
rect 2610 273056 2618 273120
rect 2682 273056 2698 273120
rect 2762 273056 2778 273120
rect 2842 273056 2858 273120
rect 2922 273056 2930 273120
rect 2610 273055 2930 273056
rect 5944 273120 6264 273121
rect 5944 273056 5952 273120
rect 6016 273056 6032 273120
rect 6096 273056 6112 273120
rect 6176 273056 6192 273120
rect 6256 273056 6264 273120
rect 5944 273055 6264 273056
rect 4277 272576 4597 272577
rect 4277 272512 4285 272576
rect 4349 272512 4365 272576
rect 4429 272512 4445 272576
rect 4509 272512 4525 272576
rect 4589 272512 4597 272576
rect 4277 272511 4597 272512
rect 7610 272576 7930 272577
rect 7610 272512 7618 272576
rect 7682 272512 7698 272576
rect 7762 272512 7778 272576
rect 7842 272512 7858 272576
rect 7922 272512 7930 272576
rect 7610 272511 7930 272512
rect 2610 272032 2930 272033
rect 2610 271968 2618 272032
rect 2682 271968 2698 272032
rect 2762 271968 2778 272032
rect 2842 271968 2858 272032
rect 2922 271968 2930 272032
rect 2610 271967 2930 271968
rect 5944 272032 6264 272033
rect 5944 271968 5952 272032
rect 6016 271968 6032 272032
rect 6096 271968 6112 272032
rect 6176 271968 6192 272032
rect 6256 271968 6264 272032
rect 5944 271967 6264 271968
rect 4277 271488 4597 271489
rect 4277 271424 4285 271488
rect 4349 271424 4365 271488
rect 4429 271424 4445 271488
rect 4509 271424 4525 271488
rect 4589 271424 4597 271488
rect 4277 271423 4597 271424
rect 7610 271488 7930 271489
rect 7610 271424 7618 271488
rect 7682 271424 7698 271488
rect 7762 271424 7778 271488
rect 7842 271424 7858 271488
rect 7922 271424 7930 271488
rect 7610 271423 7930 271424
rect 2610 270944 2930 270945
rect 2610 270880 2618 270944
rect 2682 270880 2698 270944
rect 2762 270880 2778 270944
rect 2842 270880 2858 270944
rect 2922 270880 2930 270944
rect 2610 270879 2930 270880
rect 5944 270944 6264 270945
rect 5944 270880 5952 270944
rect 6016 270880 6032 270944
rect 6096 270880 6112 270944
rect 6176 270880 6192 270944
rect 6256 270880 6264 270944
rect 5944 270879 6264 270880
rect 4277 270400 4597 270401
rect 4277 270336 4285 270400
rect 4349 270336 4365 270400
rect 4429 270336 4445 270400
rect 4509 270336 4525 270400
rect 4589 270336 4597 270400
rect 4277 270335 4597 270336
rect 7610 270400 7930 270401
rect 7610 270336 7618 270400
rect 7682 270336 7698 270400
rect 7762 270336 7778 270400
rect 7842 270336 7858 270400
rect 7922 270336 7930 270400
rect 7610 270335 7930 270336
rect 2610 269856 2930 269857
rect 2610 269792 2618 269856
rect 2682 269792 2698 269856
rect 2762 269792 2778 269856
rect 2842 269792 2858 269856
rect 2922 269792 2930 269856
rect 2610 269791 2930 269792
rect 5944 269856 6264 269857
rect 5944 269792 5952 269856
rect 6016 269792 6032 269856
rect 6096 269792 6112 269856
rect 6176 269792 6192 269856
rect 6256 269792 6264 269856
rect 5944 269791 6264 269792
rect 4277 269312 4597 269313
rect 4277 269248 4285 269312
rect 4349 269248 4365 269312
rect 4429 269248 4445 269312
rect 4509 269248 4525 269312
rect 4589 269248 4597 269312
rect 4277 269247 4597 269248
rect 7610 269312 7930 269313
rect 7610 269248 7618 269312
rect 7682 269248 7698 269312
rect 7762 269248 7778 269312
rect 7842 269248 7858 269312
rect 7922 269248 7930 269312
rect 7610 269247 7930 269248
rect 2610 268768 2930 268769
rect 2610 268704 2618 268768
rect 2682 268704 2698 268768
rect 2762 268704 2778 268768
rect 2842 268704 2858 268768
rect 2922 268704 2930 268768
rect 2610 268703 2930 268704
rect 5944 268768 6264 268769
rect 5944 268704 5952 268768
rect 6016 268704 6032 268768
rect 6096 268704 6112 268768
rect 6176 268704 6192 268768
rect 6256 268704 6264 268768
rect 5944 268703 6264 268704
rect 4277 268224 4597 268225
rect 4277 268160 4285 268224
rect 4349 268160 4365 268224
rect 4429 268160 4445 268224
rect 4509 268160 4525 268224
rect 4589 268160 4597 268224
rect 4277 268159 4597 268160
rect 7610 268224 7930 268225
rect 7610 268160 7618 268224
rect 7682 268160 7698 268224
rect 7762 268160 7778 268224
rect 7842 268160 7858 268224
rect 7922 268160 7930 268224
rect 7610 268159 7930 268160
rect 2610 267680 2930 267681
rect 2610 267616 2618 267680
rect 2682 267616 2698 267680
rect 2762 267616 2778 267680
rect 2842 267616 2858 267680
rect 2922 267616 2930 267680
rect 2610 267615 2930 267616
rect 5944 267680 6264 267681
rect 5944 267616 5952 267680
rect 6016 267616 6032 267680
rect 6096 267616 6112 267680
rect 6176 267616 6192 267680
rect 6256 267616 6264 267680
rect 5944 267615 6264 267616
rect 4277 267136 4597 267137
rect 4277 267072 4285 267136
rect 4349 267072 4365 267136
rect 4429 267072 4445 267136
rect 4509 267072 4525 267136
rect 4589 267072 4597 267136
rect 4277 267071 4597 267072
rect 7610 267136 7930 267137
rect 7610 267072 7618 267136
rect 7682 267072 7698 267136
rect 7762 267072 7778 267136
rect 7842 267072 7858 267136
rect 7922 267072 7930 267136
rect 7610 267071 7930 267072
rect 2610 266592 2930 266593
rect 2610 266528 2618 266592
rect 2682 266528 2698 266592
rect 2762 266528 2778 266592
rect 2842 266528 2858 266592
rect 2922 266528 2930 266592
rect 2610 266527 2930 266528
rect 5944 266592 6264 266593
rect 5944 266528 5952 266592
rect 6016 266528 6032 266592
rect 6096 266528 6112 266592
rect 6176 266528 6192 266592
rect 6256 266528 6264 266592
rect 5944 266527 6264 266528
rect 4277 266048 4597 266049
rect 4277 265984 4285 266048
rect 4349 265984 4365 266048
rect 4429 265984 4445 266048
rect 4509 265984 4525 266048
rect 4589 265984 4597 266048
rect 4277 265983 4597 265984
rect 7610 266048 7930 266049
rect 7610 265984 7618 266048
rect 7682 265984 7698 266048
rect 7762 265984 7778 266048
rect 7842 265984 7858 266048
rect 7922 265984 7930 266048
rect 7610 265983 7930 265984
rect 2610 265504 2930 265505
rect 2610 265440 2618 265504
rect 2682 265440 2698 265504
rect 2762 265440 2778 265504
rect 2842 265440 2858 265504
rect 2922 265440 2930 265504
rect 2610 265439 2930 265440
rect 5944 265504 6264 265505
rect 5944 265440 5952 265504
rect 6016 265440 6032 265504
rect 6096 265440 6112 265504
rect 6176 265440 6192 265504
rect 6256 265440 6264 265504
rect 5944 265439 6264 265440
rect 4277 264960 4597 264961
rect 4277 264896 4285 264960
rect 4349 264896 4365 264960
rect 4429 264896 4445 264960
rect 4509 264896 4525 264960
rect 4589 264896 4597 264960
rect 4277 264895 4597 264896
rect 7610 264960 7930 264961
rect 7610 264896 7618 264960
rect 7682 264896 7698 264960
rect 7762 264896 7778 264960
rect 7842 264896 7858 264960
rect 7922 264896 7930 264960
rect 7610 264895 7930 264896
rect 2610 264416 2930 264417
rect 2610 264352 2618 264416
rect 2682 264352 2698 264416
rect 2762 264352 2778 264416
rect 2842 264352 2858 264416
rect 2922 264352 2930 264416
rect 2610 264351 2930 264352
rect 5944 264416 6264 264417
rect 5944 264352 5952 264416
rect 6016 264352 6032 264416
rect 6096 264352 6112 264416
rect 6176 264352 6192 264416
rect 6256 264352 6264 264416
rect 5944 264351 6264 264352
rect 4277 263872 4597 263873
rect 4277 263808 4285 263872
rect 4349 263808 4365 263872
rect 4429 263808 4445 263872
rect 4509 263808 4525 263872
rect 4589 263808 4597 263872
rect 4277 263807 4597 263808
rect 7610 263872 7930 263873
rect 7610 263808 7618 263872
rect 7682 263808 7698 263872
rect 7762 263808 7778 263872
rect 7842 263808 7858 263872
rect 7922 263808 7930 263872
rect 7610 263807 7930 263808
rect 2610 263328 2930 263329
rect 2610 263264 2618 263328
rect 2682 263264 2698 263328
rect 2762 263264 2778 263328
rect 2842 263264 2858 263328
rect 2922 263264 2930 263328
rect 2610 263263 2930 263264
rect 5944 263328 6264 263329
rect 5944 263264 5952 263328
rect 6016 263264 6032 263328
rect 6096 263264 6112 263328
rect 6176 263264 6192 263328
rect 6256 263264 6264 263328
rect 5944 263263 6264 263264
rect 4277 262784 4597 262785
rect 4277 262720 4285 262784
rect 4349 262720 4365 262784
rect 4429 262720 4445 262784
rect 4509 262720 4525 262784
rect 4589 262720 4597 262784
rect 4277 262719 4597 262720
rect 7610 262784 7930 262785
rect 7610 262720 7618 262784
rect 7682 262720 7698 262784
rect 7762 262720 7778 262784
rect 7842 262720 7858 262784
rect 7922 262720 7930 262784
rect 7610 262719 7930 262720
rect 2610 262240 2930 262241
rect 2610 262176 2618 262240
rect 2682 262176 2698 262240
rect 2762 262176 2778 262240
rect 2842 262176 2858 262240
rect 2922 262176 2930 262240
rect 2610 262175 2930 262176
rect 5944 262240 6264 262241
rect 5944 262176 5952 262240
rect 6016 262176 6032 262240
rect 6096 262176 6112 262240
rect 6176 262176 6192 262240
rect 6256 262176 6264 262240
rect 5944 262175 6264 262176
rect 4277 261696 4597 261697
rect 0 261536 480 261656
rect 4277 261632 4285 261696
rect 4349 261632 4365 261696
rect 4429 261632 4445 261696
rect 4509 261632 4525 261696
rect 4589 261632 4597 261696
rect 4277 261631 4597 261632
rect 7610 261696 7930 261697
rect 7610 261632 7618 261696
rect 7682 261632 7698 261696
rect 7762 261632 7778 261696
rect 7842 261632 7858 261696
rect 7922 261632 7930 261696
rect 7610 261631 7930 261632
rect 62 261354 122 261536
rect 2497 261354 2563 261357
rect 62 261352 2563 261354
rect 62 261296 2502 261352
rect 2558 261296 2563 261352
rect 62 261294 2563 261296
rect 2497 261291 2563 261294
rect 2610 261152 2930 261153
rect 2610 261088 2618 261152
rect 2682 261088 2698 261152
rect 2762 261088 2778 261152
rect 2842 261088 2858 261152
rect 2922 261088 2930 261152
rect 2610 261087 2930 261088
rect 5944 261152 6264 261153
rect 5944 261088 5952 261152
rect 6016 261088 6032 261152
rect 6096 261088 6112 261152
rect 6176 261088 6192 261152
rect 6256 261088 6264 261152
rect 5944 261087 6264 261088
rect 4277 260608 4597 260609
rect 4277 260544 4285 260608
rect 4349 260544 4365 260608
rect 4429 260544 4445 260608
rect 4509 260544 4525 260608
rect 4589 260544 4597 260608
rect 4277 260543 4597 260544
rect 7610 260608 7930 260609
rect 7610 260544 7618 260608
rect 7682 260544 7698 260608
rect 7762 260544 7778 260608
rect 7842 260544 7858 260608
rect 7922 260544 7930 260608
rect 7610 260543 7930 260544
rect 2610 260064 2930 260065
rect 2610 260000 2618 260064
rect 2682 260000 2698 260064
rect 2762 260000 2778 260064
rect 2842 260000 2858 260064
rect 2922 260000 2930 260064
rect 2610 259999 2930 260000
rect 5944 260064 6264 260065
rect 5944 260000 5952 260064
rect 6016 260000 6032 260064
rect 6096 260000 6112 260064
rect 6176 260000 6192 260064
rect 6256 260000 6264 260064
rect 5944 259999 6264 260000
rect 4277 259520 4597 259521
rect 4277 259456 4285 259520
rect 4349 259456 4365 259520
rect 4429 259456 4445 259520
rect 4509 259456 4525 259520
rect 4589 259456 4597 259520
rect 4277 259455 4597 259456
rect 7610 259520 7930 259521
rect 7610 259456 7618 259520
rect 7682 259456 7698 259520
rect 7762 259456 7778 259520
rect 7842 259456 7858 259520
rect 7922 259456 7930 259520
rect 7610 259455 7930 259456
rect 2610 258976 2930 258977
rect 2610 258912 2618 258976
rect 2682 258912 2698 258976
rect 2762 258912 2778 258976
rect 2842 258912 2858 258976
rect 2922 258912 2930 258976
rect 2610 258911 2930 258912
rect 5944 258976 6264 258977
rect 5944 258912 5952 258976
rect 6016 258912 6032 258976
rect 6096 258912 6112 258976
rect 6176 258912 6192 258976
rect 6256 258912 6264 258976
rect 5944 258911 6264 258912
rect 4277 258432 4597 258433
rect 4277 258368 4285 258432
rect 4349 258368 4365 258432
rect 4429 258368 4445 258432
rect 4509 258368 4525 258432
rect 4589 258368 4597 258432
rect 4277 258367 4597 258368
rect 7610 258432 7930 258433
rect 7610 258368 7618 258432
rect 7682 258368 7698 258432
rect 7762 258368 7778 258432
rect 7842 258368 7858 258432
rect 7922 258368 7930 258432
rect 7610 258367 7930 258368
rect 2610 257888 2930 257889
rect 2610 257824 2618 257888
rect 2682 257824 2698 257888
rect 2762 257824 2778 257888
rect 2842 257824 2858 257888
rect 2922 257824 2930 257888
rect 2610 257823 2930 257824
rect 5944 257888 6264 257889
rect 5944 257824 5952 257888
rect 6016 257824 6032 257888
rect 6096 257824 6112 257888
rect 6176 257824 6192 257888
rect 6256 257824 6264 257888
rect 5944 257823 6264 257824
rect 4277 257344 4597 257345
rect 4277 257280 4285 257344
rect 4349 257280 4365 257344
rect 4429 257280 4445 257344
rect 4509 257280 4525 257344
rect 4589 257280 4597 257344
rect 4277 257279 4597 257280
rect 7610 257344 7930 257345
rect 7610 257280 7618 257344
rect 7682 257280 7698 257344
rect 7762 257280 7778 257344
rect 7842 257280 7858 257344
rect 7922 257280 7930 257344
rect 7610 257279 7930 257280
rect 2610 256800 2930 256801
rect 2610 256736 2618 256800
rect 2682 256736 2698 256800
rect 2762 256736 2778 256800
rect 2842 256736 2858 256800
rect 2922 256736 2930 256800
rect 2610 256735 2930 256736
rect 5944 256800 6264 256801
rect 5944 256736 5952 256800
rect 6016 256736 6032 256800
rect 6096 256736 6112 256800
rect 6176 256736 6192 256800
rect 6256 256736 6264 256800
rect 5944 256735 6264 256736
rect 4277 256256 4597 256257
rect 4277 256192 4285 256256
rect 4349 256192 4365 256256
rect 4429 256192 4445 256256
rect 4509 256192 4525 256256
rect 4589 256192 4597 256256
rect 4277 256191 4597 256192
rect 7610 256256 7930 256257
rect 7610 256192 7618 256256
rect 7682 256192 7698 256256
rect 7762 256192 7778 256256
rect 7842 256192 7858 256256
rect 7922 256192 7930 256256
rect 7610 256191 7930 256192
rect 2610 255712 2930 255713
rect 2610 255648 2618 255712
rect 2682 255648 2698 255712
rect 2762 255648 2778 255712
rect 2842 255648 2858 255712
rect 2922 255648 2930 255712
rect 2610 255647 2930 255648
rect 5944 255712 6264 255713
rect 5944 255648 5952 255712
rect 6016 255648 6032 255712
rect 6096 255648 6112 255712
rect 6176 255648 6192 255712
rect 6256 255648 6264 255712
rect 5944 255647 6264 255648
rect 4277 255168 4597 255169
rect 4277 255104 4285 255168
rect 4349 255104 4365 255168
rect 4429 255104 4445 255168
rect 4509 255104 4525 255168
rect 4589 255104 4597 255168
rect 4277 255103 4597 255104
rect 7610 255168 7930 255169
rect 7610 255104 7618 255168
rect 7682 255104 7698 255168
rect 7762 255104 7778 255168
rect 7842 255104 7858 255168
rect 7922 255104 7930 255168
rect 7610 255103 7930 255104
rect 2610 254624 2930 254625
rect 2610 254560 2618 254624
rect 2682 254560 2698 254624
rect 2762 254560 2778 254624
rect 2842 254560 2858 254624
rect 2922 254560 2930 254624
rect 2610 254559 2930 254560
rect 5944 254624 6264 254625
rect 5944 254560 5952 254624
rect 6016 254560 6032 254624
rect 6096 254560 6112 254624
rect 6176 254560 6192 254624
rect 6256 254560 6264 254624
rect 5944 254559 6264 254560
rect 4277 254080 4597 254081
rect 4277 254016 4285 254080
rect 4349 254016 4365 254080
rect 4429 254016 4445 254080
rect 4509 254016 4525 254080
rect 4589 254016 4597 254080
rect 4277 254015 4597 254016
rect 7610 254080 7930 254081
rect 7610 254016 7618 254080
rect 7682 254016 7698 254080
rect 7762 254016 7778 254080
rect 7842 254016 7858 254080
rect 7922 254016 7930 254080
rect 7610 254015 7930 254016
rect 2610 253536 2930 253537
rect 2610 253472 2618 253536
rect 2682 253472 2698 253536
rect 2762 253472 2778 253536
rect 2842 253472 2858 253536
rect 2922 253472 2930 253536
rect 2610 253471 2930 253472
rect 5944 253536 6264 253537
rect 5944 253472 5952 253536
rect 6016 253472 6032 253536
rect 6096 253472 6112 253536
rect 6176 253472 6192 253536
rect 6256 253472 6264 253536
rect 5944 253471 6264 253472
rect 4277 252992 4597 252993
rect 4277 252928 4285 252992
rect 4349 252928 4365 252992
rect 4429 252928 4445 252992
rect 4509 252928 4525 252992
rect 4589 252928 4597 252992
rect 4277 252927 4597 252928
rect 7610 252992 7930 252993
rect 7610 252928 7618 252992
rect 7682 252928 7698 252992
rect 7762 252928 7778 252992
rect 7842 252928 7858 252992
rect 7922 252928 7930 252992
rect 7610 252927 7930 252928
rect 2610 252448 2930 252449
rect 2610 252384 2618 252448
rect 2682 252384 2698 252448
rect 2762 252384 2778 252448
rect 2842 252384 2858 252448
rect 2922 252384 2930 252448
rect 2610 252383 2930 252384
rect 5944 252448 6264 252449
rect 5944 252384 5952 252448
rect 6016 252384 6032 252448
rect 6096 252384 6112 252448
rect 6176 252384 6192 252448
rect 6256 252384 6264 252448
rect 5944 252383 6264 252384
rect 4277 251904 4597 251905
rect 4277 251840 4285 251904
rect 4349 251840 4365 251904
rect 4429 251840 4445 251904
rect 4509 251840 4525 251904
rect 4589 251840 4597 251904
rect 4277 251839 4597 251840
rect 7610 251904 7930 251905
rect 7610 251840 7618 251904
rect 7682 251840 7698 251904
rect 7762 251840 7778 251904
rect 7842 251840 7858 251904
rect 7922 251840 7930 251904
rect 7610 251839 7930 251840
rect 2610 251360 2930 251361
rect 2610 251296 2618 251360
rect 2682 251296 2698 251360
rect 2762 251296 2778 251360
rect 2842 251296 2858 251360
rect 2922 251296 2930 251360
rect 2610 251295 2930 251296
rect 5944 251360 6264 251361
rect 5944 251296 5952 251360
rect 6016 251296 6032 251360
rect 6096 251296 6112 251360
rect 6176 251296 6192 251360
rect 6256 251296 6264 251360
rect 5944 251295 6264 251296
rect 4277 250816 4597 250817
rect 4277 250752 4285 250816
rect 4349 250752 4365 250816
rect 4429 250752 4445 250816
rect 4509 250752 4525 250816
rect 4589 250752 4597 250816
rect 4277 250751 4597 250752
rect 7610 250816 7930 250817
rect 7610 250752 7618 250816
rect 7682 250752 7698 250816
rect 7762 250752 7778 250816
rect 7842 250752 7858 250816
rect 7922 250752 7930 250816
rect 7610 250751 7930 250752
rect 2610 250272 2930 250273
rect 2610 250208 2618 250272
rect 2682 250208 2698 250272
rect 2762 250208 2778 250272
rect 2842 250208 2858 250272
rect 2922 250208 2930 250272
rect 2610 250207 2930 250208
rect 5944 250272 6264 250273
rect 5944 250208 5952 250272
rect 6016 250208 6032 250272
rect 6096 250208 6112 250272
rect 6176 250208 6192 250272
rect 6256 250208 6264 250272
rect 5944 250207 6264 250208
rect 4277 249728 4597 249729
rect 4277 249664 4285 249728
rect 4349 249664 4365 249728
rect 4429 249664 4445 249728
rect 4509 249664 4525 249728
rect 4589 249664 4597 249728
rect 4277 249663 4597 249664
rect 7610 249728 7930 249729
rect 7610 249664 7618 249728
rect 7682 249664 7698 249728
rect 7762 249664 7778 249728
rect 7842 249664 7858 249728
rect 7922 249664 7930 249728
rect 9520 249704 10000 249824
rect 7610 249663 7930 249664
rect 6361 249250 6427 249253
rect 9630 249250 9690 249704
rect 6361 249248 9690 249250
rect 6361 249192 6366 249248
rect 6422 249192 9690 249248
rect 6361 249190 9690 249192
rect 6361 249187 6427 249190
rect 2610 249184 2930 249185
rect 2610 249120 2618 249184
rect 2682 249120 2698 249184
rect 2762 249120 2778 249184
rect 2842 249120 2858 249184
rect 2922 249120 2930 249184
rect 2610 249119 2930 249120
rect 5944 249184 6264 249185
rect 5944 249120 5952 249184
rect 6016 249120 6032 249184
rect 6096 249120 6112 249184
rect 6176 249120 6192 249184
rect 6256 249120 6264 249184
rect 5944 249119 6264 249120
rect 4277 248640 4597 248641
rect 4277 248576 4285 248640
rect 4349 248576 4365 248640
rect 4429 248576 4445 248640
rect 4509 248576 4525 248640
rect 4589 248576 4597 248640
rect 4277 248575 4597 248576
rect 7610 248640 7930 248641
rect 7610 248576 7618 248640
rect 7682 248576 7698 248640
rect 7762 248576 7778 248640
rect 7842 248576 7858 248640
rect 7922 248576 7930 248640
rect 7610 248575 7930 248576
rect 2610 248096 2930 248097
rect 2610 248032 2618 248096
rect 2682 248032 2698 248096
rect 2762 248032 2778 248096
rect 2842 248032 2858 248096
rect 2922 248032 2930 248096
rect 2610 248031 2930 248032
rect 5944 248096 6264 248097
rect 5944 248032 5952 248096
rect 6016 248032 6032 248096
rect 6096 248032 6112 248096
rect 6176 248032 6192 248096
rect 6256 248032 6264 248096
rect 5944 248031 6264 248032
rect 4277 247552 4597 247553
rect 4277 247488 4285 247552
rect 4349 247488 4365 247552
rect 4429 247488 4445 247552
rect 4509 247488 4525 247552
rect 4589 247488 4597 247552
rect 4277 247487 4597 247488
rect 7610 247552 7930 247553
rect 7610 247488 7618 247552
rect 7682 247488 7698 247552
rect 7762 247488 7778 247552
rect 7842 247488 7858 247552
rect 7922 247488 7930 247552
rect 7610 247487 7930 247488
rect 2610 247008 2930 247009
rect 2610 246944 2618 247008
rect 2682 246944 2698 247008
rect 2762 246944 2778 247008
rect 2842 246944 2858 247008
rect 2922 246944 2930 247008
rect 2610 246943 2930 246944
rect 5944 247008 6264 247009
rect 5944 246944 5952 247008
rect 6016 246944 6032 247008
rect 6096 246944 6112 247008
rect 6176 246944 6192 247008
rect 6256 246944 6264 247008
rect 5944 246943 6264 246944
rect 4277 246464 4597 246465
rect 4277 246400 4285 246464
rect 4349 246400 4365 246464
rect 4429 246400 4445 246464
rect 4509 246400 4525 246464
rect 4589 246400 4597 246464
rect 4277 246399 4597 246400
rect 7610 246464 7930 246465
rect 7610 246400 7618 246464
rect 7682 246400 7698 246464
rect 7762 246400 7778 246464
rect 7842 246400 7858 246464
rect 7922 246400 7930 246464
rect 7610 246399 7930 246400
rect 2610 245920 2930 245921
rect 2610 245856 2618 245920
rect 2682 245856 2698 245920
rect 2762 245856 2778 245920
rect 2842 245856 2858 245920
rect 2922 245856 2930 245920
rect 2610 245855 2930 245856
rect 5944 245920 6264 245921
rect 5944 245856 5952 245920
rect 6016 245856 6032 245920
rect 6096 245856 6112 245920
rect 6176 245856 6192 245920
rect 6256 245856 6264 245920
rect 5944 245855 6264 245856
rect 4277 245376 4597 245377
rect 4277 245312 4285 245376
rect 4349 245312 4365 245376
rect 4429 245312 4445 245376
rect 4509 245312 4525 245376
rect 4589 245312 4597 245376
rect 4277 245311 4597 245312
rect 7610 245376 7930 245377
rect 7610 245312 7618 245376
rect 7682 245312 7698 245376
rect 7762 245312 7778 245376
rect 7842 245312 7858 245376
rect 7922 245312 7930 245376
rect 7610 245311 7930 245312
rect 2610 244832 2930 244833
rect 2610 244768 2618 244832
rect 2682 244768 2698 244832
rect 2762 244768 2778 244832
rect 2842 244768 2858 244832
rect 2922 244768 2930 244832
rect 2610 244767 2930 244768
rect 5944 244832 6264 244833
rect 5944 244768 5952 244832
rect 6016 244768 6032 244832
rect 6096 244768 6112 244832
rect 6176 244768 6192 244832
rect 6256 244768 6264 244832
rect 5944 244767 6264 244768
rect 4277 244288 4597 244289
rect 4277 244224 4285 244288
rect 4349 244224 4365 244288
rect 4429 244224 4445 244288
rect 4509 244224 4525 244288
rect 4589 244224 4597 244288
rect 4277 244223 4597 244224
rect 7610 244288 7930 244289
rect 7610 244224 7618 244288
rect 7682 244224 7698 244288
rect 7762 244224 7778 244288
rect 7842 244224 7858 244288
rect 7922 244224 7930 244288
rect 7610 244223 7930 244224
rect 2610 243744 2930 243745
rect 2610 243680 2618 243744
rect 2682 243680 2698 243744
rect 2762 243680 2778 243744
rect 2842 243680 2858 243744
rect 2922 243680 2930 243744
rect 2610 243679 2930 243680
rect 5944 243744 6264 243745
rect 5944 243680 5952 243744
rect 6016 243680 6032 243744
rect 6096 243680 6112 243744
rect 6176 243680 6192 243744
rect 6256 243680 6264 243744
rect 5944 243679 6264 243680
rect 4277 243200 4597 243201
rect 4277 243136 4285 243200
rect 4349 243136 4365 243200
rect 4429 243136 4445 243200
rect 4509 243136 4525 243200
rect 4589 243136 4597 243200
rect 4277 243135 4597 243136
rect 7610 243200 7930 243201
rect 7610 243136 7618 243200
rect 7682 243136 7698 243200
rect 7762 243136 7778 243200
rect 7842 243136 7858 243200
rect 7922 243136 7930 243200
rect 7610 243135 7930 243136
rect 2610 242656 2930 242657
rect 2610 242592 2618 242656
rect 2682 242592 2698 242656
rect 2762 242592 2778 242656
rect 2842 242592 2858 242656
rect 2922 242592 2930 242656
rect 2610 242591 2930 242592
rect 5944 242656 6264 242657
rect 5944 242592 5952 242656
rect 6016 242592 6032 242656
rect 6096 242592 6112 242656
rect 6176 242592 6192 242656
rect 6256 242592 6264 242656
rect 5944 242591 6264 242592
rect 4277 242112 4597 242113
rect 4277 242048 4285 242112
rect 4349 242048 4365 242112
rect 4429 242048 4445 242112
rect 4509 242048 4525 242112
rect 4589 242048 4597 242112
rect 4277 242047 4597 242048
rect 7610 242112 7930 242113
rect 7610 242048 7618 242112
rect 7682 242048 7698 242112
rect 7762 242048 7778 242112
rect 7842 242048 7858 242112
rect 7922 242048 7930 242112
rect 7610 242047 7930 242048
rect 2610 241568 2930 241569
rect 2610 241504 2618 241568
rect 2682 241504 2698 241568
rect 2762 241504 2778 241568
rect 2842 241504 2858 241568
rect 2922 241504 2930 241568
rect 2610 241503 2930 241504
rect 5944 241568 6264 241569
rect 5944 241504 5952 241568
rect 6016 241504 6032 241568
rect 6096 241504 6112 241568
rect 6176 241504 6192 241568
rect 6256 241504 6264 241568
rect 5944 241503 6264 241504
rect 4277 241024 4597 241025
rect 4277 240960 4285 241024
rect 4349 240960 4365 241024
rect 4429 240960 4445 241024
rect 4509 240960 4525 241024
rect 4589 240960 4597 241024
rect 4277 240959 4597 240960
rect 7610 241024 7930 241025
rect 7610 240960 7618 241024
rect 7682 240960 7698 241024
rect 7762 240960 7778 241024
rect 7842 240960 7858 241024
rect 7922 240960 7930 241024
rect 7610 240959 7930 240960
rect 2610 240480 2930 240481
rect 2610 240416 2618 240480
rect 2682 240416 2698 240480
rect 2762 240416 2778 240480
rect 2842 240416 2858 240480
rect 2922 240416 2930 240480
rect 2610 240415 2930 240416
rect 5944 240480 6264 240481
rect 5944 240416 5952 240480
rect 6016 240416 6032 240480
rect 6096 240416 6112 240480
rect 6176 240416 6192 240480
rect 6256 240416 6264 240480
rect 5944 240415 6264 240416
rect 4277 239936 4597 239937
rect 4277 239872 4285 239936
rect 4349 239872 4365 239936
rect 4429 239872 4445 239936
rect 4509 239872 4525 239936
rect 4589 239872 4597 239936
rect 4277 239871 4597 239872
rect 7610 239936 7930 239937
rect 7610 239872 7618 239936
rect 7682 239872 7698 239936
rect 7762 239872 7778 239936
rect 7842 239872 7858 239936
rect 7922 239872 7930 239936
rect 7610 239871 7930 239872
rect 2610 239392 2930 239393
rect 2610 239328 2618 239392
rect 2682 239328 2698 239392
rect 2762 239328 2778 239392
rect 2842 239328 2858 239392
rect 2922 239328 2930 239392
rect 2610 239327 2930 239328
rect 5944 239392 6264 239393
rect 5944 239328 5952 239392
rect 6016 239328 6032 239392
rect 6096 239328 6112 239392
rect 6176 239328 6192 239392
rect 6256 239328 6264 239392
rect 5944 239327 6264 239328
rect 4277 238848 4597 238849
rect 4277 238784 4285 238848
rect 4349 238784 4365 238848
rect 4429 238784 4445 238848
rect 4509 238784 4525 238848
rect 4589 238784 4597 238848
rect 4277 238783 4597 238784
rect 7610 238848 7930 238849
rect 7610 238784 7618 238848
rect 7682 238784 7698 238848
rect 7762 238784 7778 238848
rect 7842 238784 7858 238848
rect 7922 238784 7930 238848
rect 7610 238783 7930 238784
rect 2610 238304 2930 238305
rect 2610 238240 2618 238304
rect 2682 238240 2698 238304
rect 2762 238240 2778 238304
rect 2842 238240 2858 238304
rect 2922 238240 2930 238304
rect 2610 238239 2930 238240
rect 5944 238304 6264 238305
rect 5944 238240 5952 238304
rect 6016 238240 6032 238304
rect 6096 238240 6112 238304
rect 6176 238240 6192 238304
rect 6256 238240 6264 238304
rect 5944 238239 6264 238240
rect 4277 237760 4597 237761
rect 4277 237696 4285 237760
rect 4349 237696 4365 237760
rect 4429 237696 4445 237760
rect 4509 237696 4525 237760
rect 4589 237696 4597 237760
rect 4277 237695 4597 237696
rect 7610 237760 7930 237761
rect 7610 237696 7618 237760
rect 7682 237696 7698 237760
rect 7762 237696 7778 237760
rect 7842 237696 7858 237760
rect 7922 237696 7930 237760
rect 7610 237695 7930 237696
rect 2610 237216 2930 237217
rect 2610 237152 2618 237216
rect 2682 237152 2698 237216
rect 2762 237152 2778 237216
rect 2842 237152 2858 237216
rect 2922 237152 2930 237216
rect 2610 237151 2930 237152
rect 5944 237216 6264 237217
rect 5944 237152 5952 237216
rect 6016 237152 6032 237216
rect 6096 237152 6112 237216
rect 6176 237152 6192 237216
rect 6256 237152 6264 237216
rect 5944 237151 6264 237152
rect 4277 236672 4597 236673
rect 4277 236608 4285 236672
rect 4349 236608 4365 236672
rect 4429 236608 4445 236672
rect 4509 236608 4525 236672
rect 4589 236608 4597 236672
rect 4277 236607 4597 236608
rect 7610 236672 7930 236673
rect 7610 236608 7618 236672
rect 7682 236608 7698 236672
rect 7762 236608 7778 236672
rect 7842 236608 7858 236672
rect 7922 236608 7930 236672
rect 7610 236607 7930 236608
rect 2610 236128 2930 236129
rect 2610 236064 2618 236128
rect 2682 236064 2698 236128
rect 2762 236064 2778 236128
rect 2842 236064 2858 236128
rect 2922 236064 2930 236128
rect 2610 236063 2930 236064
rect 5944 236128 6264 236129
rect 5944 236064 5952 236128
rect 6016 236064 6032 236128
rect 6096 236064 6112 236128
rect 6176 236064 6192 236128
rect 6256 236064 6264 236128
rect 5944 236063 6264 236064
rect 4277 235584 4597 235585
rect 4277 235520 4285 235584
rect 4349 235520 4365 235584
rect 4429 235520 4445 235584
rect 4509 235520 4525 235584
rect 4589 235520 4597 235584
rect 4277 235519 4597 235520
rect 7610 235584 7930 235585
rect 7610 235520 7618 235584
rect 7682 235520 7698 235584
rect 7762 235520 7778 235584
rect 7842 235520 7858 235584
rect 7922 235520 7930 235584
rect 7610 235519 7930 235520
rect 2610 235040 2930 235041
rect 2610 234976 2618 235040
rect 2682 234976 2698 235040
rect 2762 234976 2778 235040
rect 2842 234976 2858 235040
rect 2922 234976 2930 235040
rect 2610 234975 2930 234976
rect 5944 235040 6264 235041
rect 5944 234976 5952 235040
rect 6016 234976 6032 235040
rect 6096 234976 6112 235040
rect 6176 234976 6192 235040
rect 6256 234976 6264 235040
rect 5944 234975 6264 234976
rect 4277 234496 4597 234497
rect 4277 234432 4285 234496
rect 4349 234432 4365 234496
rect 4429 234432 4445 234496
rect 4509 234432 4525 234496
rect 4589 234432 4597 234496
rect 4277 234431 4597 234432
rect 7610 234496 7930 234497
rect 7610 234432 7618 234496
rect 7682 234432 7698 234496
rect 7762 234432 7778 234496
rect 7842 234432 7858 234496
rect 7922 234432 7930 234496
rect 7610 234431 7930 234432
rect 2610 233952 2930 233953
rect 2610 233888 2618 233952
rect 2682 233888 2698 233952
rect 2762 233888 2778 233952
rect 2842 233888 2858 233952
rect 2922 233888 2930 233952
rect 2610 233887 2930 233888
rect 5944 233952 6264 233953
rect 5944 233888 5952 233952
rect 6016 233888 6032 233952
rect 6096 233888 6112 233952
rect 6176 233888 6192 233952
rect 6256 233888 6264 233952
rect 5944 233887 6264 233888
rect 4277 233408 4597 233409
rect 4277 233344 4285 233408
rect 4349 233344 4365 233408
rect 4429 233344 4445 233408
rect 4509 233344 4525 233408
rect 4589 233344 4597 233408
rect 4277 233343 4597 233344
rect 7610 233408 7930 233409
rect 7610 233344 7618 233408
rect 7682 233344 7698 233408
rect 7762 233344 7778 233408
rect 7842 233344 7858 233408
rect 7922 233344 7930 233408
rect 7610 233343 7930 233344
rect 2610 232864 2930 232865
rect 2610 232800 2618 232864
rect 2682 232800 2698 232864
rect 2762 232800 2778 232864
rect 2842 232800 2858 232864
rect 2922 232800 2930 232864
rect 2610 232799 2930 232800
rect 5944 232864 6264 232865
rect 5944 232800 5952 232864
rect 6016 232800 6032 232864
rect 6096 232800 6112 232864
rect 6176 232800 6192 232864
rect 6256 232800 6264 232864
rect 5944 232799 6264 232800
rect 4277 232320 4597 232321
rect 4277 232256 4285 232320
rect 4349 232256 4365 232320
rect 4429 232256 4445 232320
rect 4509 232256 4525 232320
rect 4589 232256 4597 232320
rect 4277 232255 4597 232256
rect 7610 232320 7930 232321
rect 7610 232256 7618 232320
rect 7682 232256 7698 232320
rect 7762 232256 7778 232320
rect 7842 232256 7858 232320
rect 7922 232256 7930 232320
rect 7610 232255 7930 232256
rect 2610 231776 2930 231777
rect 2610 231712 2618 231776
rect 2682 231712 2698 231776
rect 2762 231712 2778 231776
rect 2842 231712 2858 231776
rect 2922 231712 2930 231776
rect 2610 231711 2930 231712
rect 5944 231776 6264 231777
rect 5944 231712 5952 231776
rect 6016 231712 6032 231776
rect 6096 231712 6112 231776
rect 6176 231712 6192 231776
rect 6256 231712 6264 231776
rect 5944 231711 6264 231712
rect 4277 231232 4597 231233
rect 4277 231168 4285 231232
rect 4349 231168 4365 231232
rect 4429 231168 4445 231232
rect 4509 231168 4525 231232
rect 4589 231168 4597 231232
rect 4277 231167 4597 231168
rect 7610 231232 7930 231233
rect 7610 231168 7618 231232
rect 7682 231168 7698 231232
rect 7762 231168 7778 231232
rect 7842 231168 7858 231232
rect 7922 231168 7930 231232
rect 7610 231167 7930 231168
rect 2610 230688 2930 230689
rect 2610 230624 2618 230688
rect 2682 230624 2698 230688
rect 2762 230624 2778 230688
rect 2842 230624 2858 230688
rect 2922 230624 2930 230688
rect 2610 230623 2930 230624
rect 5944 230688 6264 230689
rect 5944 230624 5952 230688
rect 6016 230624 6032 230688
rect 6096 230624 6112 230688
rect 6176 230624 6192 230688
rect 6256 230624 6264 230688
rect 5944 230623 6264 230624
rect 4277 230144 4597 230145
rect 4277 230080 4285 230144
rect 4349 230080 4365 230144
rect 4429 230080 4445 230144
rect 4509 230080 4525 230144
rect 4589 230080 4597 230144
rect 4277 230079 4597 230080
rect 7610 230144 7930 230145
rect 7610 230080 7618 230144
rect 7682 230080 7698 230144
rect 7762 230080 7778 230144
rect 7842 230080 7858 230144
rect 7922 230080 7930 230144
rect 7610 230079 7930 230080
rect 2610 229600 2930 229601
rect 2610 229536 2618 229600
rect 2682 229536 2698 229600
rect 2762 229536 2778 229600
rect 2842 229536 2858 229600
rect 2922 229536 2930 229600
rect 2610 229535 2930 229536
rect 5944 229600 6264 229601
rect 5944 229536 5952 229600
rect 6016 229536 6032 229600
rect 6096 229536 6112 229600
rect 6176 229536 6192 229600
rect 6256 229536 6264 229600
rect 5944 229535 6264 229536
rect 4277 229056 4597 229057
rect 4277 228992 4285 229056
rect 4349 228992 4365 229056
rect 4429 228992 4445 229056
rect 4509 228992 4525 229056
rect 4589 228992 4597 229056
rect 4277 228991 4597 228992
rect 7610 229056 7930 229057
rect 7610 228992 7618 229056
rect 7682 228992 7698 229056
rect 7762 228992 7778 229056
rect 7842 228992 7858 229056
rect 7922 228992 7930 229056
rect 7610 228991 7930 228992
rect 2610 228512 2930 228513
rect 2610 228448 2618 228512
rect 2682 228448 2698 228512
rect 2762 228448 2778 228512
rect 2842 228448 2858 228512
rect 2922 228448 2930 228512
rect 2610 228447 2930 228448
rect 5944 228512 6264 228513
rect 5944 228448 5952 228512
rect 6016 228448 6032 228512
rect 6096 228448 6112 228512
rect 6176 228448 6192 228512
rect 6256 228448 6264 228512
rect 5944 228447 6264 228448
rect 4277 227968 4597 227969
rect 4277 227904 4285 227968
rect 4349 227904 4365 227968
rect 4429 227904 4445 227968
rect 4509 227904 4525 227968
rect 4589 227904 4597 227968
rect 4277 227903 4597 227904
rect 7610 227968 7930 227969
rect 7610 227904 7618 227968
rect 7682 227904 7698 227968
rect 7762 227904 7778 227968
rect 7842 227904 7858 227968
rect 7922 227904 7930 227968
rect 7610 227903 7930 227904
rect 2610 227424 2930 227425
rect 2610 227360 2618 227424
rect 2682 227360 2698 227424
rect 2762 227360 2778 227424
rect 2842 227360 2858 227424
rect 2922 227360 2930 227424
rect 2610 227359 2930 227360
rect 5944 227424 6264 227425
rect 5944 227360 5952 227424
rect 6016 227360 6032 227424
rect 6096 227360 6112 227424
rect 6176 227360 6192 227424
rect 6256 227360 6264 227424
rect 5944 227359 6264 227360
rect 4277 226880 4597 226881
rect 4277 226816 4285 226880
rect 4349 226816 4365 226880
rect 4429 226816 4445 226880
rect 4509 226816 4525 226880
rect 4589 226816 4597 226880
rect 4277 226815 4597 226816
rect 7610 226880 7930 226881
rect 7610 226816 7618 226880
rect 7682 226816 7698 226880
rect 7762 226816 7778 226880
rect 7842 226816 7858 226880
rect 7922 226816 7930 226880
rect 7610 226815 7930 226816
rect 2610 226336 2930 226337
rect 2610 226272 2618 226336
rect 2682 226272 2698 226336
rect 2762 226272 2778 226336
rect 2842 226272 2858 226336
rect 2922 226272 2930 226336
rect 2610 226271 2930 226272
rect 5944 226336 6264 226337
rect 5944 226272 5952 226336
rect 6016 226272 6032 226336
rect 6096 226272 6112 226336
rect 6176 226272 6192 226336
rect 6256 226272 6264 226336
rect 5944 226271 6264 226272
rect 4277 225792 4597 225793
rect 4277 225728 4285 225792
rect 4349 225728 4365 225792
rect 4429 225728 4445 225792
rect 4509 225728 4525 225792
rect 4589 225728 4597 225792
rect 4277 225727 4597 225728
rect 7610 225792 7930 225793
rect 7610 225728 7618 225792
rect 7682 225728 7698 225792
rect 7762 225728 7778 225792
rect 7842 225728 7858 225792
rect 7922 225728 7930 225792
rect 7610 225727 7930 225728
rect 2610 225248 2930 225249
rect 2610 225184 2618 225248
rect 2682 225184 2698 225248
rect 2762 225184 2778 225248
rect 2842 225184 2858 225248
rect 2922 225184 2930 225248
rect 2610 225183 2930 225184
rect 5944 225248 6264 225249
rect 5944 225184 5952 225248
rect 6016 225184 6032 225248
rect 6096 225184 6112 225248
rect 6176 225184 6192 225248
rect 6256 225184 6264 225248
rect 5944 225183 6264 225184
rect 4277 224704 4597 224705
rect 4277 224640 4285 224704
rect 4349 224640 4365 224704
rect 4429 224640 4445 224704
rect 4509 224640 4525 224704
rect 4589 224640 4597 224704
rect 4277 224639 4597 224640
rect 7610 224704 7930 224705
rect 7610 224640 7618 224704
rect 7682 224640 7698 224704
rect 7762 224640 7778 224704
rect 7842 224640 7858 224704
rect 7922 224640 7930 224704
rect 7610 224639 7930 224640
rect 2610 224160 2930 224161
rect 2610 224096 2618 224160
rect 2682 224096 2698 224160
rect 2762 224096 2778 224160
rect 2842 224096 2858 224160
rect 2922 224096 2930 224160
rect 2610 224095 2930 224096
rect 5944 224160 6264 224161
rect 5944 224096 5952 224160
rect 6016 224096 6032 224160
rect 6096 224096 6112 224160
rect 6176 224096 6192 224160
rect 6256 224096 6264 224160
rect 5944 224095 6264 224096
rect 4277 223616 4597 223617
rect 4277 223552 4285 223616
rect 4349 223552 4365 223616
rect 4429 223552 4445 223616
rect 4509 223552 4525 223616
rect 4589 223552 4597 223616
rect 4277 223551 4597 223552
rect 7610 223616 7930 223617
rect 7610 223552 7618 223616
rect 7682 223552 7698 223616
rect 7762 223552 7778 223616
rect 7842 223552 7858 223616
rect 7922 223552 7930 223616
rect 7610 223551 7930 223552
rect 2610 223072 2930 223073
rect 2610 223008 2618 223072
rect 2682 223008 2698 223072
rect 2762 223008 2778 223072
rect 2842 223008 2858 223072
rect 2922 223008 2930 223072
rect 2610 223007 2930 223008
rect 5944 223072 6264 223073
rect 5944 223008 5952 223072
rect 6016 223008 6032 223072
rect 6096 223008 6112 223072
rect 6176 223008 6192 223072
rect 6256 223008 6264 223072
rect 5944 223007 6264 223008
rect 4277 222528 4597 222529
rect 4277 222464 4285 222528
rect 4349 222464 4365 222528
rect 4429 222464 4445 222528
rect 4509 222464 4525 222528
rect 4589 222464 4597 222528
rect 4277 222463 4597 222464
rect 7610 222528 7930 222529
rect 7610 222464 7618 222528
rect 7682 222464 7698 222528
rect 7762 222464 7778 222528
rect 7842 222464 7858 222528
rect 7922 222464 7930 222528
rect 7610 222463 7930 222464
rect 2610 221984 2930 221985
rect 2610 221920 2618 221984
rect 2682 221920 2698 221984
rect 2762 221920 2778 221984
rect 2842 221920 2858 221984
rect 2922 221920 2930 221984
rect 2610 221919 2930 221920
rect 5944 221984 6264 221985
rect 5944 221920 5952 221984
rect 6016 221920 6032 221984
rect 6096 221920 6112 221984
rect 6176 221920 6192 221984
rect 6256 221920 6264 221984
rect 5944 221919 6264 221920
rect 4277 221440 4597 221441
rect 4277 221376 4285 221440
rect 4349 221376 4365 221440
rect 4429 221376 4445 221440
rect 4509 221376 4525 221440
rect 4589 221376 4597 221440
rect 4277 221375 4597 221376
rect 7610 221440 7930 221441
rect 7610 221376 7618 221440
rect 7682 221376 7698 221440
rect 7762 221376 7778 221440
rect 7842 221376 7858 221440
rect 7922 221376 7930 221440
rect 7610 221375 7930 221376
rect 2610 220896 2930 220897
rect 2610 220832 2618 220896
rect 2682 220832 2698 220896
rect 2762 220832 2778 220896
rect 2842 220832 2858 220896
rect 2922 220832 2930 220896
rect 2610 220831 2930 220832
rect 5944 220896 6264 220897
rect 5944 220832 5952 220896
rect 6016 220832 6032 220896
rect 6096 220832 6112 220896
rect 6176 220832 6192 220896
rect 6256 220832 6264 220896
rect 5944 220831 6264 220832
rect 4277 220352 4597 220353
rect 4277 220288 4285 220352
rect 4349 220288 4365 220352
rect 4429 220288 4445 220352
rect 4509 220288 4525 220352
rect 4589 220288 4597 220352
rect 4277 220287 4597 220288
rect 7610 220352 7930 220353
rect 7610 220288 7618 220352
rect 7682 220288 7698 220352
rect 7762 220288 7778 220352
rect 7842 220288 7858 220352
rect 7922 220288 7930 220352
rect 7610 220287 7930 220288
rect 2610 219808 2930 219809
rect 2610 219744 2618 219808
rect 2682 219744 2698 219808
rect 2762 219744 2778 219808
rect 2842 219744 2858 219808
rect 2922 219744 2930 219808
rect 2610 219743 2930 219744
rect 5944 219808 6264 219809
rect 5944 219744 5952 219808
rect 6016 219744 6032 219808
rect 6096 219744 6112 219808
rect 6176 219744 6192 219808
rect 6256 219744 6264 219808
rect 5944 219743 6264 219744
rect 4277 219264 4597 219265
rect 4277 219200 4285 219264
rect 4349 219200 4365 219264
rect 4429 219200 4445 219264
rect 4509 219200 4525 219264
rect 4589 219200 4597 219264
rect 4277 219199 4597 219200
rect 7610 219264 7930 219265
rect 7610 219200 7618 219264
rect 7682 219200 7698 219264
rect 7762 219200 7778 219264
rect 7842 219200 7858 219264
rect 7922 219200 7930 219264
rect 7610 219199 7930 219200
rect 2610 218720 2930 218721
rect 2610 218656 2618 218720
rect 2682 218656 2698 218720
rect 2762 218656 2778 218720
rect 2842 218656 2858 218720
rect 2922 218656 2930 218720
rect 2610 218655 2930 218656
rect 5944 218720 6264 218721
rect 5944 218656 5952 218720
rect 6016 218656 6032 218720
rect 6096 218656 6112 218720
rect 6176 218656 6192 218720
rect 6256 218656 6264 218720
rect 5944 218655 6264 218656
rect 4277 218176 4597 218177
rect 4277 218112 4285 218176
rect 4349 218112 4365 218176
rect 4429 218112 4445 218176
rect 4509 218112 4525 218176
rect 4589 218112 4597 218176
rect 4277 218111 4597 218112
rect 7610 218176 7930 218177
rect 7610 218112 7618 218176
rect 7682 218112 7698 218176
rect 7762 218112 7778 218176
rect 7842 218112 7858 218176
rect 7922 218112 7930 218176
rect 7610 218111 7930 218112
rect 2610 217632 2930 217633
rect 2610 217568 2618 217632
rect 2682 217568 2698 217632
rect 2762 217568 2778 217632
rect 2842 217568 2858 217632
rect 2922 217568 2930 217632
rect 2610 217567 2930 217568
rect 5944 217632 6264 217633
rect 5944 217568 5952 217632
rect 6016 217568 6032 217632
rect 6096 217568 6112 217632
rect 6176 217568 6192 217632
rect 6256 217568 6264 217632
rect 5944 217567 6264 217568
rect 4277 217088 4597 217089
rect 4277 217024 4285 217088
rect 4349 217024 4365 217088
rect 4429 217024 4445 217088
rect 4509 217024 4525 217088
rect 4589 217024 4597 217088
rect 4277 217023 4597 217024
rect 7610 217088 7930 217089
rect 7610 217024 7618 217088
rect 7682 217024 7698 217088
rect 7762 217024 7778 217088
rect 7842 217024 7858 217088
rect 7922 217024 7930 217088
rect 7610 217023 7930 217024
rect 2610 216544 2930 216545
rect 2610 216480 2618 216544
rect 2682 216480 2698 216544
rect 2762 216480 2778 216544
rect 2842 216480 2858 216544
rect 2922 216480 2930 216544
rect 2610 216479 2930 216480
rect 5944 216544 6264 216545
rect 5944 216480 5952 216544
rect 6016 216480 6032 216544
rect 6096 216480 6112 216544
rect 6176 216480 6192 216544
rect 6256 216480 6264 216544
rect 5944 216479 6264 216480
rect 9520 216384 10000 216504
rect 7005 216202 7071 216205
rect 9630 216202 9690 216384
rect 7005 216200 9690 216202
rect 7005 216144 7010 216200
rect 7066 216144 9690 216200
rect 7005 216142 9690 216144
rect 7005 216139 7071 216142
rect 4277 216000 4597 216001
rect 4277 215936 4285 216000
rect 4349 215936 4365 216000
rect 4429 215936 4445 216000
rect 4509 215936 4525 216000
rect 4589 215936 4597 216000
rect 4277 215935 4597 215936
rect 7610 216000 7930 216001
rect 7610 215936 7618 216000
rect 7682 215936 7698 216000
rect 7762 215936 7778 216000
rect 7842 215936 7858 216000
rect 7922 215936 7930 216000
rect 7610 215935 7930 215936
rect 2610 215456 2930 215457
rect 2610 215392 2618 215456
rect 2682 215392 2698 215456
rect 2762 215392 2778 215456
rect 2842 215392 2858 215456
rect 2922 215392 2930 215456
rect 2610 215391 2930 215392
rect 5944 215456 6264 215457
rect 5944 215392 5952 215456
rect 6016 215392 6032 215456
rect 6096 215392 6112 215456
rect 6176 215392 6192 215456
rect 6256 215392 6264 215456
rect 5944 215391 6264 215392
rect 4277 214912 4597 214913
rect 4277 214848 4285 214912
rect 4349 214848 4365 214912
rect 4429 214848 4445 214912
rect 4509 214848 4525 214912
rect 4589 214848 4597 214912
rect 4277 214847 4597 214848
rect 7610 214912 7930 214913
rect 7610 214848 7618 214912
rect 7682 214848 7698 214912
rect 7762 214848 7778 214912
rect 7842 214848 7858 214912
rect 7922 214848 7930 214912
rect 7610 214847 7930 214848
rect 2610 214368 2930 214369
rect 2610 214304 2618 214368
rect 2682 214304 2698 214368
rect 2762 214304 2778 214368
rect 2842 214304 2858 214368
rect 2922 214304 2930 214368
rect 2610 214303 2930 214304
rect 5944 214368 6264 214369
rect 5944 214304 5952 214368
rect 6016 214304 6032 214368
rect 6096 214304 6112 214368
rect 6176 214304 6192 214368
rect 6256 214304 6264 214368
rect 5944 214303 6264 214304
rect 0 214024 480 214056
rect 0 213968 110 214024
rect 166 213968 480 214024
rect 0 213936 480 213968
rect 4277 213824 4597 213825
rect 4277 213760 4285 213824
rect 4349 213760 4365 213824
rect 4429 213760 4445 213824
rect 4509 213760 4525 213824
rect 4589 213760 4597 213824
rect 4277 213759 4597 213760
rect 7610 213824 7930 213825
rect 7610 213760 7618 213824
rect 7682 213760 7698 213824
rect 7762 213760 7778 213824
rect 7842 213760 7858 213824
rect 7922 213760 7930 213824
rect 7610 213759 7930 213760
rect 2610 213280 2930 213281
rect 2610 213216 2618 213280
rect 2682 213216 2698 213280
rect 2762 213216 2778 213280
rect 2842 213216 2858 213280
rect 2922 213216 2930 213280
rect 2610 213215 2930 213216
rect 5944 213280 6264 213281
rect 5944 213216 5952 213280
rect 6016 213216 6032 213280
rect 6096 213216 6112 213280
rect 6176 213216 6192 213280
rect 6256 213216 6264 213280
rect 5944 213215 6264 213216
rect 4277 212736 4597 212737
rect 4277 212672 4285 212736
rect 4349 212672 4365 212736
rect 4429 212672 4445 212736
rect 4509 212672 4525 212736
rect 4589 212672 4597 212736
rect 4277 212671 4597 212672
rect 7610 212736 7930 212737
rect 7610 212672 7618 212736
rect 7682 212672 7698 212736
rect 7762 212672 7778 212736
rect 7842 212672 7858 212736
rect 7922 212672 7930 212736
rect 7610 212671 7930 212672
rect 2610 212192 2930 212193
rect 2610 212128 2618 212192
rect 2682 212128 2698 212192
rect 2762 212128 2778 212192
rect 2842 212128 2858 212192
rect 2922 212128 2930 212192
rect 2610 212127 2930 212128
rect 5944 212192 6264 212193
rect 5944 212128 5952 212192
rect 6016 212128 6032 212192
rect 6096 212128 6112 212192
rect 6176 212128 6192 212192
rect 6256 212128 6264 212192
rect 5944 212127 6264 212128
rect 4277 211648 4597 211649
rect 4277 211584 4285 211648
rect 4349 211584 4365 211648
rect 4429 211584 4445 211648
rect 4509 211584 4525 211648
rect 4589 211584 4597 211648
rect 4277 211583 4597 211584
rect 7610 211648 7930 211649
rect 7610 211584 7618 211648
rect 7682 211584 7698 211648
rect 7762 211584 7778 211648
rect 7842 211584 7858 211648
rect 7922 211584 7930 211648
rect 7610 211583 7930 211584
rect 2610 211104 2930 211105
rect 2610 211040 2618 211104
rect 2682 211040 2698 211104
rect 2762 211040 2778 211104
rect 2842 211040 2858 211104
rect 2922 211040 2930 211104
rect 2610 211039 2930 211040
rect 5944 211104 6264 211105
rect 5944 211040 5952 211104
rect 6016 211040 6032 211104
rect 6096 211040 6112 211104
rect 6176 211040 6192 211104
rect 6256 211040 6264 211104
rect 5944 211039 6264 211040
rect 4277 210560 4597 210561
rect 4277 210496 4285 210560
rect 4349 210496 4365 210560
rect 4429 210496 4445 210560
rect 4509 210496 4525 210560
rect 4589 210496 4597 210560
rect 4277 210495 4597 210496
rect 7610 210560 7930 210561
rect 7610 210496 7618 210560
rect 7682 210496 7698 210560
rect 7762 210496 7778 210560
rect 7842 210496 7858 210560
rect 7922 210496 7930 210560
rect 7610 210495 7930 210496
rect 2610 210016 2930 210017
rect 2610 209952 2618 210016
rect 2682 209952 2698 210016
rect 2762 209952 2778 210016
rect 2842 209952 2858 210016
rect 2922 209952 2930 210016
rect 2610 209951 2930 209952
rect 5944 210016 6264 210017
rect 5944 209952 5952 210016
rect 6016 209952 6032 210016
rect 6096 209952 6112 210016
rect 6176 209952 6192 210016
rect 6256 209952 6264 210016
rect 5944 209951 6264 209952
rect 4277 209472 4597 209473
rect 4277 209408 4285 209472
rect 4349 209408 4365 209472
rect 4429 209408 4445 209472
rect 4509 209408 4525 209472
rect 4589 209408 4597 209472
rect 4277 209407 4597 209408
rect 7610 209472 7930 209473
rect 7610 209408 7618 209472
rect 7682 209408 7698 209472
rect 7762 209408 7778 209472
rect 7842 209408 7858 209472
rect 7922 209408 7930 209472
rect 7610 209407 7930 209408
rect 2610 208928 2930 208929
rect 2610 208864 2618 208928
rect 2682 208864 2698 208928
rect 2762 208864 2778 208928
rect 2842 208864 2858 208928
rect 2922 208864 2930 208928
rect 2610 208863 2930 208864
rect 5944 208928 6264 208929
rect 5944 208864 5952 208928
rect 6016 208864 6032 208928
rect 6096 208864 6112 208928
rect 6176 208864 6192 208928
rect 6256 208864 6264 208928
rect 5944 208863 6264 208864
rect 4277 208384 4597 208385
rect 4277 208320 4285 208384
rect 4349 208320 4365 208384
rect 4429 208320 4445 208384
rect 4509 208320 4525 208384
rect 4589 208320 4597 208384
rect 4277 208319 4597 208320
rect 7610 208384 7930 208385
rect 7610 208320 7618 208384
rect 7682 208320 7698 208384
rect 7762 208320 7778 208384
rect 7842 208320 7858 208384
rect 7922 208320 7930 208384
rect 7610 208319 7930 208320
rect 2610 207840 2930 207841
rect 2610 207776 2618 207840
rect 2682 207776 2698 207840
rect 2762 207776 2778 207840
rect 2842 207776 2858 207840
rect 2922 207776 2930 207840
rect 2610 207775 2930 207776
rect 5944 207840 6264 207841
rect 5944 207776 5952 207840
rect 6016 207776 6032 207840
rect 6096 207776 6112 207840
rect 6176 207776 6192 207840
rect 6256 207776 6264 207840
rect 5944 207775 6264 207776
rect 4277 207296 4597 207297
rect 4277 207232 4285 207296
rect 4349 207232 4365 207296
rect 4429 207232 4445 207296
rect 4509 207232 4525 207296
rect 4589 207232 4597 207296
rect 4277 207231 4597 207232
rect 7610 207296 7930 207297
rect 7610 207232 7618 207296
rect 7682 207232 7698 207296
rect 7762 207232 7778 207296
rect 7842 207232 7858 207296
rect 7922 207232 7930 207296
rect 7610 207231 7930 207232
rect 2610 206752 2930 206753
rect 2610 206688 2618 206752
rect 2682 206688 2698 206752
rect 2762 206688 2778 206752
rect 2842 206688 2858 206752
rect 2922 206688 2930 206752
rect 2610 206687 2930 206688
rect 5944 206752 6264 206753
rect 5944 206688 5952 206752
rect 6016 206688 6032 206752
rect 6096 206688 6112 206752
rect 6176 206688 6192 206752
rect 6256 206688 6264 206752
rect 5944 206687 6264 206688
rect 4277 206208 4597 206209
rect 4277 206144 4285 206208
rect 4349 206144 4365 206208
rect 4429 206144 4445 206208
rect 4509 206144 4525 206208
rect 4589 206144 4597 206208
rect 4277 206143 4597 206144
rect 7610 206208 7930 206209
rect 7610 206144 7618 206208
rect 7682 206144 7698 206208
rect 7762 206144 7778 206208
rect 7842 206144 7858 206208
rect 7922 206144 7930 206208
rect 7610 206143 7930 206144
rect 2610 205664 2930 205665
rect 2610 205600 2618 205664
rect 2682 205600 2698 205664
rect 2762 205600 2778 205664
rect 2842 205600 2858 205664
rect 2922 205600 2930 205664
rect 2610 205599 2930 205600
rect 5944 205664 6264 205665
rect 5944 205600 5952 205664
rect 6016 205600 6032 205664
rect 6096 205600 6112 205664
rect 6176 205600 6192 205664
rect 6256 205600 6264 205664
rect 5944 205599 6264 205600
rect 4277 205120 4597 205121
rect 4277 205056 4285 205120
rect 4349 205056 4365 205120
rect 4429 205056 4445 205120
rect 4509 205056 4525 205120
rect 4589 205056 4597 205120
rect 4277 205055 4597 205056
rect 7610 205120 7930 205121
rect 7610 205056 7618 205120
rect 7682 205056 7698 205120
rect 7762 205056 7778 205120
rect 7842 205056 7858 205120
rect 7922 205056 7930 205120
rect 7610 205055 7930 205056
rect 2610 204576 2930 204577
rect 2610 204512 2618 204576
rect 2682 204512 2698 204576
rect 2762 204512 2778 204576
rect 2842 204512 2858 204576
rect 2922 204512 2930 204576
rect 2610 204511 2930 204512
rect 5944 204576 6264 204577
rect 5944 204512 5952 204576
rect 6016 204512 6032 204576
rect 6096 204512 6112 204576
rect 6176 204512 6192 204576
rect 6256 204512 6264 204576
rect 5944 204511 6264 204512
rect 4277 204032 4597 204033
rect 4277 203968 4285 204032
rect 4349 203968 4365 204032
rect 4429 203968 4445 204032
rect 4509 203968 4525 204032
rect 4589 203968 4597 204032
rect 4277 203967 4597 203968
rect 7610 204032 7930 204033
rect 7610 203968 7618 204032
rect 7682 203968 7698 204032
rect 7762 203968 7778 204032
rect 7842 203968 7858 204032
rect 7922 203968 7930 204032
rect 7610 203967 7930 203968
rect 2610 203488 2930 203489
rect 2610 203424 2618 203488
rect 2682 203424 2698 203488
rect 2762 203424 2778 203488
rect 2842 203424 2858 203488
rect 2922 203424 2930 203488
rect 2610 203423 2930 203424
rect 5944 203488 6264 203489
rect 5944 203424 5952 203488
rect 6016 203424 6032 203488
rect 6096 203424 6112 203488
rect 6176 203424 6192 203488
rect 6256 203424 6264 203488
rect 5944 203423 6264 203424
rect 4277 202944 4597 202945
rect 4277 202880 4285 202944
rect 4349 202880 4365 202944
rect 4429 202880 4445 202944
rect 4509 202880 4525 202944
rect 4589 202880 4597 202944
rect 4277 202879 4597 202880
rect 7610 202944 7930 202945
rect 7610 202880 7618 202944
rect 7682 202880 7698 202944
rect 7762 202880 7778 202944
rect 7842 202880 7858 202944
rect 7922 202880 7930 202944
rect 7610 202879 7930 202880
rect 2610 202400 2930 202401
rect 2610 202336 2618 202400
rect 2682 202336 2698 202400
rect 2762 202336 2778 202400
rect 2842 202336 2858 202400
rect 2922 202336 2930 202400
rect 2610 202335 2930 202336
rect 5944 202400 6264 202401
rect 5944 202336 5952 202400
rect 6016 202336 6032 202400
rect 6096 202336 6112 202400
rect 6176 202336 6192 202400
rect 6256 202336 6264 202400
rect 5944 202335 6264 202336
rect 4277 201856 4597 201857
rect 4277 201792 4285 201856
rect 4349 201792 4365 201856
rect 4429 201792 4445 201856
rect 4509 201792 4525 201856
rect 4589 201792 4597 201856
rect 4277 201791 4597 201792
rect 7610 201856 7930 201857
rect 7610 201792 7618 201856
rect 7682 201792 7698 201856
rect 7762 201792 7778 201856
rect 7842 201792 7858 201856
rect 7922 201792 7930 201856
rect 7610 201791 7930 201792
rect 2610 201312 2930 201313
rect 2610 201248 2618 201312
rect 2682 201248 2698 201312
rect 2762 201248 2778 201312
rect 2842 201248 2858 201312
rect 2922 201248 2930 201312
rect 2610 201247 2930 201248
rect 5944 201312 6264 201313
rect 5944 201248 5952 201312
rect 6016 201248 6032 201312
rect 6096 201248 6112 201312
rect 6176 201248 6192 201312
rect 6256 201248 6264 201312
rect 5944 201247 6264 201248
rect 4277 200768 4597 200769
rect 4277 200704 4285 200768
rect 4349 200704 4365 200768
rect 4429 200704 4445 200768
rect 4509 200704 4525 200768
rect 4589 200704 4597 200768
rect 4277 200703 4597 200704
rect 7610 200768 7930 200769
rect 7610 200704 7618 200768
rect 7682 200704 7698 200768
rect 7762 200704 7778 200768
rect 7842 200704 7858 200768
rect 7922 200704 7930 200768
rect 7610 200703 7930 200704
rect 2610 200224 2930 200225
rect 2610 200160 2618 200224
rect 2682 200160 2698 200224
rect 2762 200160 2778 200224
rect 2842 200160 2858 200224
rect 2922 200160 2930 200224
rect 2610 200159 2930 200160
rect 5944 200224 6264 200225
rect 5944 200160 5952 200224
rect 6016 200160 6032 200224
rect 6096 200160 6112 200224
rect 6176 200160 6192 200224
rect 6256 200160 6264 200224
rect 5944 200159 6264 200160
rect 4277 199680 4597 199681
rect 4277 199616 4285 199680
rect 4349 199616 4365 199680
rect 4429 199616 4445 199680
rect 4509 199616 4525 199680
rect 4589 199616 4597 199680
rect 4277 199615 4597 199616
rect 7610 199680 7930 199681
rect 7610 199616 7618 199680
rect 7682 199616 7698 199680
rect 7762 199616 7778 199680
rect 7842 199616 7858 199680
rect 7922 199616 7930 199680
rect 7610 199615 7930 199616
rect 2610 199136 2930 199137
rect 2610 199072 2618 199136
rect 2682 199072 2698 199136
rect 2762 199072 2778 199136
rect 2842 199072 2858 199136
rect 2922 199072 2930 199136
rect 2610 199071 2930 199072
rect 5944 199136 6264 199137
rect 5944 199072 5952 199136
rect 6016 199072 6032 199136
rect 6096 199072 6112 199136
rect 6176 199072 6192 199136
rect 6256 199072 6264 199136
rect 5944 199071 6264 199072
rect 4277 198592 4597 198593
rect 4277 198528 4285 198592
rect 4349 198528 4365 198592
rect 4429 198528 4445 198592
rect 4509 198528 4525 198592
rect 4589 198528 4597 198592
rect 4277 198527 4597 198528
rect 7610 198592 7930 198593
rect 7610 198528 7618 198592
rect 7682 198528 7698 198592
rect 7762 198528 7778 198592
rect 7842 198528 7858 198592
rect 7922 198528 7930 198592
rect 7610 198527 7930 198528
rect 2610 198048 2930 198049
rect 2610 197984 2618 198048
rect 2682 197984 2698 198048
rect 2762 197984 2778 198048
rect 2842 197984 2858 198048
rect 2922 197984 2930 198048
rect 2610 197983 2930 197984
rect 5944 198048 6264 198049
rect 5944 197984 5952 198048
rect 6016 197984 6032 198048
rect 6096 197984 6112 198048
rect 6176 197984 6192 198048
rect 6256 197984 6264 198048
rect 5944 197983 6264 197984
rect 4277 197504 4597 197505
rect 4277 197440 4285 197504
rect 4349 197440 4365 197504
rect 4429 197440 4445 197504
rect 4509 197440 4525 197504
rect 4589 197440 4597 197504
rect 4277 197439 4597 197440
rect 7610 197504 7930 197505
rect 7610 197440 7618 197504
rect 7682 197440 7698 197504
rect 7762 197440 7778 197504
rect 7842 197440 7858 197504
rect 7922 197440 7930 197504
rect 7610 197439 7930 197440
rect 2610 196960 2930 196961
rect 2610 196896 2618 196960
rect 2682 196896 2698 196960
rect 2762 196896 2778 196960
rect 2842 196896 2858 196960
rect 2922 196896 2930 196960
rect 2610 196895 2930 196896
rect 5944 196960 6264 196961
rect 5944 196896 5952 196960
rect 6016 196896 6032 196960
rect 6096 196896 6112 196960
rect 6176 196896 6192 196960
rect 6256 196896 6264 196960
rect 5944 196895 6264 196896
rect 4277 196416 4597 196417
rect 4277 196352 4285 196416
rect 4349 196352 4365 196416
rect 4429 196352 4445 196416
rect 4509 196352 4525 196416
rect 4589 196352 4597 196416
rect 4277 196351 4597 196352
rect 7610 196416 7930 196417
rect 7610 196352 7618 196416
rect 7682 196352 7698 196416
rect 7762 196352 7778 196416
rect 7842 196352 7858 196416
rect 7922 196352 7930 196416
rect 7610 196351 7930 196352
rect 2610 195872 2930 195873
rect 2610 195808 2618 195872
rect 2682 195808 2698 195872
rect 2762 195808 2778 195872
rect 2842 195808 2858 195872
rect 2922 195808 2930 195872
rect 2610 195807 2930 195808
rect 5944 195872 6264 195873
rect 5944 195808 5952 195872
rect 6016 195808 6032 195872
rect 6096 195808 6112 195872
rect 6176 195808 6192 195872
rect 6256 195808 6264 195872
rect 5944 195807 6264 195808
rect 4277 195328 4597 195329
rect 4277 195264 4285 195328
rect 4349 195264 4365 195328
rect 4429 195264 4445 195328
rect 4509 195264 4525 195328
rect 4589 195264 4597 195328
rect 4277 195263 4597 195264
rect 7610 195328 7930 195329
rect 7610 195264 7618 195328
rect 7682 195264 7698 195328
rect 7762 195264 7778 195328
rect 7842 195264 7858 195328
rect 7922 195264 7930 195328
rect 7610 195263 7930 195264
rect 2610 194784 2930 194785
rect 2610 194720 2618 194784
rect 2682 194720 2698 194784
rect 2762 194720 2778 194784
rect 2842 194720 2858 194784
rect 2922 194720 2930 194784
rect 2610 194719 2930 194720
rect 5944 194784 6264 194785
rect 5944 194720 5952 194784
rect 6016 194720 6032 194784
rect 6096 194720 6112 194784
rect 6176 194720 6192 194784
rect 6256 194720 6264 194784
rect 5944 194719 6264 194720
rect 4277 194240 4597 194241
rect 4277 194176 4285 194240
rect 4349 194176 4365 194240
rect 4429 194176 4445 194240
rect 4509 194176 4525 194240
rect 4589 194176 4597 194240
rect 4277 194175 4597 194176
rect 7610 194240 7930 194241
rect 7610 194176 7618 194240
rect 7682 194176 7698 194240
rect 7762 194176 7778 194240
rect 7842 194176 7858 194240
rect 7922 194176 7930 194240
rect 7610 194175 7930 194176
rect 2610 193696 2930 193697
rect 2610 193632 2618 193696
rect 2682 193632 2698 193696
rect 2762 193632 2778 193696
rect 2842 193632 2858 193696
rect 2922 193632 2930 193696
rect 2610 193631 2930 193632
rect 5944 193696 6264 193697
rect 5944 193632 5952 193696
rect 6016 193632 6032 193696
rect 6096 193632 6112 193696
rect 6176 193632 6192 193696
rect 6256 193632 6264 193696
rect 5944 193631 6264 193632
rect 4277 193152 4597 193153
rect 4277 193088 4285 193152
rect 4349 193088 4365 193152
rect 4429 193088 4445 193152
rect 4509 193088 4525 193152
rect 4589 193088 4597 193152
rect 4277 193087 4597 193088
rect 7610 193152 7930 193153
rect 7610 193088 7618 193152
rect 7682 193088 7698 193152
rect 7762 193088 7778 193152
rect 7842 193088 7858 193152
rect 7922 193088 7930 193152
rect 7610 193087 7930 193088
rect 2610 192608 2930 192609
rect 2610 192544 2618 192608
rect 2682 192544 2698 192608
rect 2762 192544 2778 192608
rect 2842 192544 2858 192608
rect 2922 192544 2930 192608
rect 2610 192543 2930 192544
rect 5944 192608 6264 192609
rect 5944 192544 5952 192608
rect 6016 192544 6032 192608
rect 6096 192544 6112 192608
rect 6176 192544 6192 192608
rect 6256 192544 6264 192608
rect 5944 192543 6264 192544
rect 4277 192064 4597 192065
rect 4277 192000 4285 192064
rect 4349 192000 4365 192064
rect 4429 192000 4445 192064
rect 4509 192000 4525 192064
rect 4589 192000 4597 192064
rect 4277 191999 4597 192000
rect 7610 192064 7930 192065
rect 7610 192000 7618 192064
rect 7682 192000 7698 192064
rect 7762 192000 7778 192064
rect 7842 192000 7858 192064
rect 7922 192000 7930 192064
rect 7610 191999 7930 192000
rect 2610 191520 2930 191521
rect 2610 191456 2618 191520
rect 2682 191456 2698 191520
rect 2762 191456 2778 191520
rect 2842 191456 2858 191520
rect 2922 191456 2930 191520
rect 2610 191455 2930 191456
rect 5944 191520 6264 191521
rect 5944 191456 5952 191520
rect 6016 191456 6032 191520
rect 6096 191456 6112 191520
rect 6176 191456 6192 191520
rect 6256 191456 6264 191520
rect 5944 191455 6264 191456
rect 4277 190976 4597 190977
rect 4277 190912 4285 190976
rect 4349 190912 4365 190976
rect 4429 190912 4445 190976
rect 4509 190912 4525 190976
rect 4589 190912 4597 190976
rect 4277 190911 4597 190912
rect 7610 190976 7930 190977
rect 7610 190912 7618 190976
rect 7682 190912 7698 190976
rect 7762 190912 7778 190976
rect 7842 190912 7858 190976
rect 7922 190912 7930 190976
rect 7610 190911 7930 190912
rect 2610 190432 2930 190433
rect 2610 190368 2618 190432
rect 2682 190368 2698 190432
rect 2762 190368 2778 190432
rect 2842 190368 2858 190432
rect 2922 190368 2930 190432
rect 2610 190367 2930 190368
rect 5944 190432 6264 190433
rect 5944 190368 5952 190432
rect 6016 190368 6032 190432
rect 6096 190368 6112 190432
rect 6176 190368 6192 190432
rect 6256 190368 6264 190432
rect 5944 190367 6264 190368
rect 4277 189888 4597 189889
rect 4277 189824 4285 189888
rect 4349 189824 4365 189888
rect 4429 189824 4445 189888
rect 4509 189824 4525 189888
rect 4589 189824 4597 189888
rect 4277 189823 4597 189824
rect 7610 189888 7930 189889
rect 7610 189824 7618 189888
rect 7682 189824 7698 189888
rect 7762 189824 7778 189888
rect 7842 189824 7858 189888
rect 7922 189824 7930 189888
rect 7610 189823 7930 189824
rect 2610 189344 2930 189345
rect 2610 189280 2618 189344
rect 2682 189280 2698 189344
rect 2762 189280 2778 189344
rect 2842 189280 2858 189344
rect 2922 189280 2930 189344
rect 2610 189279 2930 189280
rect 5944 189344 6264 189345
rect 5944 189280 5952 189344
rect 6016 189280 6032 189344
rect 6096 189280 6112 189344
rect 6176 189280 6192 189344
rect 6256 189280 6264 189344
rect 5944 189279 6264 189280
rect 4277 188800 4597 188801
rect 4277 188736 4285 188800
rect 4349 188736 4365 188800
rect 4429 188736 4445 188800
rect 4509 188736 4525 188800
rect 4589 188736 4597 188800
rect 4277 188735 4597 188736
rect 7610 188800 7930 188801
rect 7610 188736 7618 188800
rect 7682 188736 7698 188800
rect 7762 188736 7778 188800
rect 7842 188736 7858 188800
rect 7922 188736 7930 188800
rect 7610 188735 7930 188736
rect 2610 188256 2930 188257
rect 2610 188192 2618 188256
rect 2682 188192 2698 188256
rect 2762 188192 2778 188256
rect 2842 188192 2858 188256
rect 2922 188192 2930 188256
rect 2610 188191 2930 188192
rect 5944 188256 6264 188257
rect 5944 188192 5952 188256
rect 6016 188192 6032 188256
rect 6096 188192 6112 188256
rect 6176 188192 6192 188256
rect 6256 188192 6264 188256
rect 5944 188191 6264 188192
rect 4277 187712 4597 187713
rect 4277 187648 4285 187712
rect 4349 187648 4365 187712
rect 4429 187648 4445 187712
rect 4509 187648 4525 187712
rect 4589 187648 4597 187712
rect 4277 187647 4597 187648
rect 7610 187712 7930 187713
rect 7610 187648 7618 187712
rect 7682 187648 7698 187712
rect 7762 187648 7778 187712
rect 7842 187648 7858 187712
rect 7922 187648 7930 187712
rect 7610 187647 7930 187648
rect 2610 187168 2930 187169
rect 2610 187104 2618 187168
rect 2682 187104 2698 187168
rect 2762 187104 2778 187168
rect 2842 187104 2858 187168
rect 2922 187104 2930 187168
rect 2610 187103 2930 187104
rect 5944 187168 6264 187169
rect 5944 187104 5952 187168
rect 6016 187104 6032 187168
rect 6096 187104 6112 187168
rect 6176 187104 6192 187168
rect 6256 187104 6264 187168
rect 5944 187103 6264 187104
rect 4277 186624 4597 186625
rect 4277 186560 4285 186624
rect 4349 186560 4365 186624
rect 4429 186560 4445 186624
rect 4509 186560 4525 186624
rect 4589 186560 4597 186624
rect 4277 186559 4597 186560
rect 7610 186624 7930 186625
rect 7610 186560 7618 186624
rect 7682 186560 7698 186624
rect 7762 186560 7778 186624
rect 7842 186560 7858 186624
rect 7922 186560 7930 186624
rect 7610 186559 7930 186560
rect 2610 186080 2930 186081
rect 2610 186016 2618 186080
rect 2682 186016 2698 186080
rect 2762 186016 2778 186080
rect 2842 186016 2858 186080
rect 2922 186016 2930 186080
rect 2610 186015 2930 186016
rect 5944 186080 6264 186081
rect 5944 186016 5952 186080
rect 6016 186016 6032 186080
rect 6096 186016 6112 186080
rect 6176 186016 6192 186080
rect 6256 186016 6264 186080
rect 5944 186015 6264 186016
rect 4277 185536 4597 185537
rect 4277 185472 4285 185536
rect 4349 185472 4365 185536
rect 4429 185472 4445 185536
rect 4509 185472 4525 185536
rect 4589 185472 4597 185536
rect 4277 185471 4597 185472
rect 7610 185536 7930 185537
rect 7610 185472 7618 185536
rect 7682 185472 7698 185536
rect 7762 185472 7778 185536
rect 7842 185472 7858 185536
rect 7922 185472 7930 185536
rect 7610 185471 7930 185472
rect 2610 184992 2930 184993
rect 2610 184928 2618 184992
rect 2682 184928 2698 184992
rect 2762 184928 2778 184992
rect 2842 184928 2858 184992
rect 2922 184928 2930 184992
rect 2610 184927 2930 184928
rect 5944 184992 6264 184993
rect 5944 184928 5952 184992
rect 6016 184928 6032 184992
rect 6096 184928 6112 184992
rect 6176 184928 6192 184992
rect 6256 184928 6264 184992
rect 5944 184927 6264 184928
rect 4277 184448 4597 184449
rect 4277 184384 4285 184448
rect 4349 184384 4365 184448
rect 4429 184384 4445 184448
rect 4509 184384 4525 184448
rect 4589 184384 4597 184448
rect 4277 184383 4597 184384
rect 7610 184448 7930 184449
rect 7610 184384 7618 184448
rect 7682 184384 7698 184448
rect 7762 184384 7778 184448
rect 7842 184384 7858 184448
rect 7922 184384 7930 184448
rect 7610 184383 7930 184384
rect 2610 183904 2930 183905
rect 2610 183840 2618 183904
rect 2682 183840 2698 183904
rect 2762 183840 2778 183904
rect 2842 183840 2858 183904
rect 2922 183840 2930 183904
rect 2610 183839 2930 183840
rect 5944 183904 6264 183905
rect 5944 183840 5952 183904
rect 6016 183840 6032 183904
rect 6096 183840 6112 183904
rect 6176 183840 6192 183904
rect 6256 183840 6264 183904
rect 5944 183839 6264 183840
rect 4277 183360 4597 183361
rect 4277 183296 4285 183360
rect 4349 183296 4365 183360
rect 4429 183296 4445 183360
rect 4509 183296 4525 183360
rect 4589 183296 4597 183360
rect 4277 183295 4597 183296
rect 7610 183360 7930 183361
rect 7610 183296 7618 183360
rect 7682 183296 7698 183360
rect 7762 183296 7778 183360
rect 7842 183296 7858 183360
rect 7922 183296 7930 183360
rect 7610 183295 7930 183296
rect 9520 183064 10000 183184
rect 2610 182816 2930 182817
rect 2610 182752 2618 182816
rect 2682 182752 2698 182816
rect 2762 182752 2778 182816
rect 2842 182752 2858 182816
rect 2922 182752 2930 182816
rect 2610 182751 2930 182752
rect 5944 182816 6264 182817
rect 5944 182752 5952 182816
rect 6016 182752 6032 182816
rect 6096 182752 6112 182816
rect 6176 182752 6192 182816
rect 6256 182752 6264 182816
rect 5944 182751 6264 182752
rect 6637 182610 6703 182613
rect 9630 182610 9690 183064
rect 6637 182608 9690 182610
rect 6637 182552 6642 182608
rect 6698 182552 9690 182608
rect 6637 182550 9690 182552
rect 6637 182547 6703 182550
rect 4277 182272 4597 182273
rect 4277 182208 4285 182272
rect 4349 182208 4365 182272
rect 4429 182208 4445 182272
rect 4509 182208 4525 182272
rect 4589 182208 4597 182272
rect 4277 182207 4597 182208
rect 7610 182272 7930 182273
rect 7610 182208 7618 182272
rect 7682 182208 7698 182272
rect 7762 182208 7778 182272
rect 7842 182208 7858 182272
rect 7922 182208 7930 182272
rect 7610 182207 7930 182208
rect 2610 181728 2930 181729
rect 2610 181664 2618 181728
rect 2682 181664 2698 181728
rect 2762 181664 2778 181728
rect 2842 181664 2858 181728
rect 2922 181664 2930 181728
rect 2610 181663 2930 181664
rect 5944 181728 6264 181729
rect 5944 181664 5952 181728
rect 6016 181664 6032 181728
rect 6096 181664 6112 181728
rect 6176 181664 6192 181728
rect 6256 181664 6264 181728
rect 5944 181663 6264 181664
rect 4277 181184 4597 181185
rect 4277 181120 4285 181184
rect 4349 181120 4365 181184
rect 4429 181120 4445 181184
rect 4509 181120 4525 181184
rect 4589 181120 4597 181184
rect 4277 181119 4597 181120
rect 7610 181184 7930 181185
rect 7610 181120 7618 181184
rect 7682 181120 7698 181184
rect 7762 181120 7778 181184
rect 7842 181120 7858 181184
rect 7922 181120 7930 181184
rect 7610 181119 7930 181120
rect 2610 180640 2930 180641
rect 2610 180576 2618 180640
rect 2682 180576 2698 180640
rect 2762 180576 2778 180640
rect 2842 180576 2858 180640
rect 2922 180576 2930 180640
rect 2610 180575 2930 180576
rect 5944 180640 6264 180641
rect 5944 180576 5952 180640
rect 6016 180576 6032 180640
rect 6096 180576 6112 180640
rect 6176 180576 6192 180640
rect 6256 180576 6264 180640
rect 5944 180575 6264 180576
rect 4277 180096 4597 180097
rect 4277 180032 4285 180096
rect 4349 180032 4365 180096
rect 4429 180032 4445 180096
rect 4509 180032 4525 180096
rect 4589 180032 4597 180096
rect 4277 180031 4597 180032
rect 7610 180096 7930 180097
rect 7610 180032 7618 180096
rect 7682 180032 7698 180096
rect 7762 180032 7778 180096
rect 7842 180032 7858 180096
rect 7922 180032 7930 180096
rect 7610 180031 7930 180032
rect 2610 179552 2930 179553
rect 2610 179488 2618 179552
rect 2682 179488 2698 179552
rect 2762 179488 2778 179552
rect 2842 179488 2858 179552
rect 2922 179488 2930 179552
rect 2610 179487 2930 179488
rect 5944 179552 6264 179553
rect 5944 179488 5952 179552
rect 6016 179488 6032 179552
rect 6096 179488 6112 179552
rect 6176 179488 6192 179552
rect 6256 179488 6264 179552
rect 5944 179487 6264 179488
rect 4277 179008 4597 179009
rect 4277 178944 4285 179008
rect 4349 178944 4365 179008
rect 4429 178944 4445 179008
rect 4509 178944 4525 179008
rect 4589 178944 4597 179008
rect 4277 178943 4597 178944
rect 7610 179008 7930 179009
rect 7610 178944 7618 179008
rect 7682 178944 7698 179008
rect 7762 178944 7778 179008
rect 7842 178944 7858 179008
rect 7922 178944 7930 179008
rect 7610 178943 7930 178944
rect 2610 178464 2930 178465
rect 2610 178400 2618 178464
rect 2682 178400 2698 178464
rect 2762 178400 2778 178464
rect 2842 178400 2858 178464
rect 2922 178400 2930 178464
rect 2610 178399 2930 178400
rect 5944 178464 6264 178465
rect 5944 178400 5952 178464
rect 6016 178400 6032 178464
rect 6096 178400 6112 178464
rect 6176 178400 6192 178464
rect 6256 178400 6264 178464
rect 5944 178399 6264 178400
rect 4277 177920 4597 177921
rect 4277 177856 4285 177920
rect 4349 177856 4365 177920
rect 4429 177856 4445 177920
rect 4509 177856 4525 177920
rect 4589 177856 4597 177920
rect 4277 177855 4597 177856
rect 7610 177920 7930 177921
rect 7610 177856 7618 177920
rect 7682 177856 7698 177920
rect 7762 177856 7778 177920
rect 7842 177856 7858 177920
rect 7922 177856 7930 177920
rect 7610 177855 7930 177856
rect 2610 177376 2930 177377
rect 2610 177312 2618 177376
rect 2682 177312 2698 177376
rect 2762 177312 2778 177376
rect 2842 177312 2858 177376
rect 2922 177312 2930 177376
rect 2610 177311 2930 177312
rect 5944 177376 6264 177377
rect 5944 177312 5952 177376
rect 6016 177312 6032 177376
rect 6096 177312 6112 177376
rect 6176 177312 6192 177376
rect 6256 177312 6264 177376
rect 5944 177311 6264 177312
rect 4277 176832 4597 176833
rect 4277 176768 4285 176832
rect 4349 176768 4365 176832
rect 4429 176768 4445 176832
rect 4509 176768 4525 176832
rect 4589 176768 4597 176832
rect 4277 176767 4597 176768
rect 7610 176832 7930 176833
rect 7610 176768 7618 176832
rect 7682 176768 7698 176832
rect 7762 176768 7778 176832
rect 7842 176768 7858 176832
rect 7922 176768 7930 176832
rect 7610 176767 7930 176768
rect 2610 176288 2930 176289
rect 2610 176224 2618 176288
rect 2682 176224 2698 176288
rect 2762 176224 2778 176288
rect 2842 176224 2858 176288
rect 2922 176224 2930 176288
rect 2610 176223 2930 176224
rect 5944 176288 6264 176289
rect 5944 176224 5952 176288
rect 6016 176224 6032 176288
rect 6096 176224 6112 176288
rect 6176 176224 6192 176288
rect 6256 176224 6264 176288
rect 5944 176223 6264 176224
rect 4277 175744 4597 175745
rect 4277 175680 4285 175744
rect 4349 175680 4365 175744
rect 4429 175680 4445 175744
rect 4509 175680 4525 175744
rect 4589 175680 4597 175744
rect 4277 175679 4597 175680
rect 7610 175744 7930 175745
rect 7610 175680 7618 175744
rect 7682 175680 7698 175744
rect 7762 175680 7778 175744
rect 7842 175680 7858 175744
rect 7922 175680 7930 175744
rect 7610 175679 7930 175680
rect 2610 175200 2930 175201
rect 2610 175136 2618 175200
rect 2682 175136 2698 175200
rect 2762 175136 2778 175200
rect 2842 175136 2858 175200
rect 2922 175136 2930 175200
rect 2610 175135 2930 175136
rect 5944 175200 6264 175201
rect 5944 175136 5952 175200
rect 6016 175136 6032 175200
rect 6096 175136 6112 175200
rect 6176 175136 6192 175200
rect 6256 175136 6264 175200
rect 5944 175135 6264 175136
rect 4277 174656 4597 174657
rect 4277 174592 4285 174656
rect 4349 174592 4365 174656
rect 4429 174592 4445 174656
rect 4509 174592 4525 174656
rect 4589 174592 4597 174656
rect 4277 174591 4597 174592
rect 7610 174656 7930 174657
rect 7610 174592 7618 174656
rect 7682 174592 7698 174656
rect 7762 174592 7778 174656
rect 7842 174592 7858 174656
rect 7922 174592 7930 174656
rect 7610 174591 7930 174592
rect 2610 174112 2930 174113
rect 2610 174048 2618 174112
rect 2682 174048 2698 174112
rect 2762 174048 2778 174112
rect 2842 174048 2858 174112
rect 2922 174048 2930 174112
rect 2610 174047 2930 174048
rect 5944 174112 6264 174113
rect 5944 174048 5952 174112
rect 6016 174048 6032 174112
rect 6096 174048 6112 174112
rect 6176 174048 6192 174112
rect 6256 174048 6264 174112
rect 5944 174047 6264 174048
rect 4277 173568 4597 173569
rect 4277 173504 4285 173568
rect 4349 173504 4365 173568
rect 4429 173504 4445 173568
rect 4509 173504 4525 173568
rect 4589 173504 4597 173568
rect 4277 173503 4597 173504
rect 7610 173568 7930 173569
rect 7610 173504 7618 173568
rect 7682 173504 7698 173568
rect 7762 173504 7778 173568
rect 7842 173504 7858 173568
rect 7922 173504 7930 173568
rect 7610 173503 7930 173504
rect 2610 173024 2930 173025
rect 2610 172960 2618 173024
rect 2682 172960 2698 173024
rect 2762 172960 2778 173024
rect 2842 172960 2858 173024
rect 2922 172960 2930 173024
rect 2610 172959 2930 172960
rect 5944 173024 6264 173025
rect 5944 172960 5952 173024
rect 6016 172960 6032 173024
rect 6096 172960 6112 173024
rect 6176 172960 6192 173024
rect 6256 172960 6264 173024
rect 5944 172959 6264 172960
rect 4277 172480 4597 172481
rect 4277 172416 4285 172480
rect 4349 172416 4365 172480
rect 4429 172416 4445 172480
rect 4509 172416 4525 172480
rect 4589 172416 4597 172480
rect 4277 172415 4597 172416
rect 7610 172480 7930 172481
rect 7610 172416 7618 172480
rect 7682 172416 7698 172480
rect 7762 172416 7778 172480
rect 7842 172416 7858 172480
rect 7922 172416 7930 172480
rect 7610 172415 7930 172416
rect 2610 171936 2930 171937
rect 2610 171872 2618 171936
rect 2682 171872 2698 171936
rect 2762 171872 2778 171936
rect 2842 171872 2858 171936
rect 2922 171872 2930 171936
rect 2610 171871 2930 171872
rect 5944 171936 6264 171937
rect 5944 171872 5952 171936
rect 6016 171872 6032 171936
rect 6096 171872 6112 171936
rect 6176 171872 6192 171936
rect 6256 171872 6264 171936
rect 5944 171871 6264 171872
rect 4277 171392 4597 171393
rect 4277 171328 4285 171392
rect 4349 171328 4365 171392
rect 4429 171328 4445 171392
rect 4509 171328 4525 171392
rect 4589 171328 4597 171392
rect 4277 171327 4597 171328
rect 7610 171392 7930 171393
rect 7610 171328 7618 171392
rect 7682 171328 7698 171392
rect 7762 171328 7778 171392
rect 7842 171328 7858 171392
rect 7922 171328 7930 171392
rect 7610 171327 7930 171328
rect 2610 170848 2930 170849
rect 2610 170784 2618 170848
rect 2682 170784 2698 170848
rect 2762 170784 2778 170848
rect 2842 170784 2858 170848
rect 2922 170784 2930 170848
rect 2610 170783 2930 170784
rect 5944 170848 6264 170849
rect 5944 170784 5952 170848
rect 6016 170784 6032 170848
rect 6096 170784 6112 170848
rect 6176 170784 6192 170848
rect 6256 170784 6264 170848
rect 5944 170783 6264 170784
rect 4277 170304 4597 170305
rect 4277 170240 4285 170304
rect 4349 170240 4365 170304
rect 4429 170240 4445 170304
rect 4509 170240 4525 170304
rect 4589 170240 4597 170304
rect 4277 170239 4597 170240
rect 7610 170304 7930 170305
rect 7610 170240 7618 170304
rect 7682 170240 7698 170304
rect 7762 170240 7778 170304
rect 7842 170240 7858 170304
rect 7922 170240 7930 170304
rect 7610 170239 7930 170240
rect 2610 169760 2930 169761
rect 2610 169696 2618 169760
rect 2682 169696 2698 169760
rect 2762 169696 2778 169760
rect 2842 169696 2858 169760
rect 2922 169696 2930 169760
rect 2610 169695 2930 169696
rect 5944 169760 6264 169761
rect 5944 169696 5952 169760
rect 6016 169696 6032 169760
rect 6096 169696 6112 169760
rect 6176 169696 6192 169760
rect 6256 169696 6264 169760
rect 5944 169695 6264 169696
rect 4277 169216 4597 169217
rect 4277 169152 4285 169216
rect 4349 169152 4365 169216
rect 4429 169152 4445 169216
rect 4509 169152 4525 169216
rect 4589 169152 4597 169216
rect 4277 169151 4597 169152
rect 7610 169216 7930 169217
rect 7610 169152 7618 169216
rect 7682 169152 7698 169216
rect 7762 169152 7778 169216
rect 7842 169152 7858 169216
rect 7922 169152 7930 169216
rect 7610 169151 7930 169152
rect 2610 168672 2930 168673
rect 2610 168608 2618 168672
rect 2682 168608 2698 168672
rect 2762 168608 2778 168672
rect 2842 168608 2858 168672
rect 2922 168608 2930 168672
rect 2610 168607 2930 168608
rect 5944 168672 6264 168673
rect 5944 168608 5952 168672
rect 6016 168608 6032 168672
rect 6096 168608 6112 168672
rect 6176 168608 6192 168672
rect 6256 168608 6264 168672
rect 5944 168607 6264 168608
rect 4277 168128 4597 168129
rect 4277 168064 4285 168128
rect 4349 168064 4365 168128
rect 4429 168064 4445 168128
rect 4509 168064 4525 168128
rect 4589 168064 4597 168128
rect 4277 168063 4597 168064
rect 7610 168128 7930 168129
rect 7610 168064 7618 168128
rect 7682 168064 7698 168128
rect 7762 168064 7778 168128
rect 7842 168064 7858 168128
rect 7922 168064 7930 168128
rect 7610 168063 7930 168064
rect 2610 167584 2930 167585
rect 2610 167520 2618 167584
rect 2682 167520 2698 167584
rect 2762 167520 2778 167584
rect 2842 167520 2858 167584
rect 2922 167520 2930 167584
rect 2610 167519 2930 167520
rect 5944 167584 6264 167585
rect 5944 167520 5952 167584
rect 6016 167520 6032 167584
rect 6096 167520 6112 167584
rect 6176 167520 6192 167584
rect 6256 167520 6264 167584
rect 5944 167519 6264 167520
rect 4277 167040 4597 167041
rect 4277 166976 4285 167040
rect 4349 166976 4365 167040
rect 4429 166976 4445 167040
rect 4509 166976 4525 167040
rect 4589 166976 4597 167040
rect 4277 166975 4597 166976
rect 7610 167040 7930 167041
rect 7610 166976 7618 167040
rect 7682 166976 7698 167040
rect 7762 166976 7778 167040
rect 7842 166976 7858 167040
rect 7922 166976 7930 167040
rect 7610 166975 7930 166976
rect 2610 166496 2930 166497
rect 0 166336 480 166456
rect 2610 166432 2618 166496
rect 2682 166432 2698 166496
rect 2762 166432 2778 166496
rect 2842 166432 2858 166496
rect 2922 166432 2930 166496
rect 2610 166431 2930 166432
rect 5944 166496 6264 166497
rect 5944 166432 5952 166496
rect 6016 166432 6032 166496
rect 6096 166432 6112 166496
rect 6176 166432 6192 166496
rect 6256 166432 6264 166496
rect 5944 166431 6264 166432
rect 62 165882 122 166336
rect 4277 165952 4597 165953
rect 4277 165888 4285 165952
rect 4349 165888 4365 165952
rect 4429 165888 4445 165952
rect 4509 165888 4525 165952
rect 4589 165888 4597 165952
rect 4277 165887 4597 165888
rect 7610 165952 7930 165953
rect 7610 165888 7618 165952
rect 7682 165888 7698 165952
rect 7762 165888 7778 165952
rect 7842 165888 7858 165952
rect 7922 165888 7930 165952
rect 7610 165887 7930 165888
rect 3417 165882 3483 165885
rect 62 165880 3483 165882
rect 62 165824 3422 165880
rect 3478 165824 3483 165880
rect 62 165822 3483 165824
rect 3417 165819 3483 165822
rect 2610 165408 2930 165409
rect 2610 165344 2618 165408
rect 2682 165344 2698 165408
rect 2762 165344 2778 165408
rect 2842 165344 2858 165408
rect 2922 165344 2930 165408
rect 2610 165343 2930 165344
rect 5944 165408 6264 165409
rect 5944 165344 5952 165408
rect 6016 165344 6032 165408
rect 6096 165344 6112 165408
rect 6176 165344 6192 165408
rect 6256 165344 6264 165408
rect 5944 165343 6264 165344
rect 4277 164864 4597 164865
rect 4277 164800 4285 164864
rect 4349 164800 4365 164864
rect 4429 164800 4445 164864
rect 4509 164800 4525 164864
rect 4589 164800 4597 164864
rect 4277 164799 4597 164800
rect 7610 164864 7930 164865
rect 7610 164800 7618 164864
rect 7682 164800 7698 164864
rect 7762 164800 7778 164864
rect 7842 164800 7858 164864
rect 7922 164800 7930 164864
rect 7610 164799 7930 164800
rect 2610 164320 2930 164321
rect 2610 164256 2618 164320
rect 2682 164256 2698 164320
rect 2762 164256 2778 164320
rect 2842 164256 2858 164320
rect 2922 164256 2930 164320
rect 2610 164255 2930 164256
rect 5944 164320 6264 164321
rect 5944 164256 5952 164320
rect 6016 164256 6032 164320
rect 6096 164256 6112 164320
rect 6176 164256 6192 164320
rect 6256 164256 6264 164320
rect 5944 164255 6264 164256
rect 4277 163776 4597 163777
rect 4277 163712 4285 163776
rect 4349 163712 4365 163776
rect 4429 163712 4445 163776
rect 4509 163712 4525 163776
rect 4589 163712 4597 163776
rect 4277 163711 4597 163712
rect 7610 163776 7930 163777
rect 7610 163712 7618 163776
rect 7682 163712 7698 163776
rect 7762 163712 7778 163776
rect 7842 163712 7858 163776
rect 7922 163712 7930 163776
rect 7610 163711 7930 163712
rect 2610 163232 2930 163233
rect 2610 163168 2618 163232
rect 2682 163168 2698 163232
rect 2762 163168 2778 163232
rect 2842 163168 2858 163232
rect 2922 163168 2930 163232
rect 2610 163167 2930 163168
rect 5944 163232 6264 163233
rect 5944 163168 5952 163232
rect 6016 163168 6032 163232
rect 6096 163168 6112 163232
rect 6176 163168 6192 163232
rect 6256 163168 6264 163232
rect 5944 163167 6264 163168
rect 4277 162688 4597 162689
rect 4277 162624 4285 162688
rect 4349 162624 4365 162688
rect 4429 162624 4445 162688
rect 4509 162624 4525 162688
rect 4589 162624 4597 162688
rect 4277 162623 4597 162624
rect 7610 162688 7930 162689
rect 7610 162624 7618 162688
rect 7682 162624 7698 162688
rect 7762 162624 7778 162688
rect 7842 162624 7858 162688
rect 7922 162624 7930 162688
rect 7610 162623 7930 162624
rect 2610 162144 2930 162145
rect 2610 162080 2618 162144
rect 2682 162080 2698 162144
rect 2762 162080 2778 162144
rect 2842 162080 2858 162144
rect 2922 162080 2930 162144
rect 2610 162079 2930 162080
rect 5944 162144 6264 162145
rect 5944 162080 5952 162144
rect 6016 162080 6032 162144
rect 6096 162080 6112 162144
rect 6176 162080 6192 162144
rect 6256 162080 6264 162144
rect 5944 162079 6264 162080
rect 4277 161600 4597 161601
rect 4277 161536 4285 161600
rect 4349 161536 4365 161600
rect 4429 161536 4445 161600
rect 4509 161536 4525 161600
rect 4589 161536 4597 161600
rect 4277 161535 4597 161536
rect 7610 161600 7930 161601
rect 7610 161536 7618 161600
rect 7682 161536 7698 161600
rect 7762 161536 7778 161600
rect 7842 161536 7858 161600
rect 7922 161536 7930 161600
rect 7610 161535 7930 161536
rect 2610 161056 2930 161057
rect 2610 160992 2618 161056
rect 2682 160992 2698 161056
rect 2762 160992 2778 161056
rect 2842 160992 2858 161056
rect 2922 160992 2930 161056
rect 2610 160991 2930 160992
rect 5944 161056 6264 161057
rect 5944 160992 5952 161056
rect 6016 160992 6032 161056
rect 6096 160992 6112 161056
rect 6176 160992 6192 161056
rect 6256 160992 6264 161056
rect 5944 160991 6264 160992
rect 4277 160512 4597 160513
rect 4277 160448 4285 160512
rect 4349 160448 4365 160512
rect 4429 160448 4445 160512
rect 4509 160448 4525 160512
rect 4589 160448 4597 160512
rect 4277 160447 4597 160448
rect 7610 160512 7930 160513
rect 7610 160448 7618 160512
rect 7682 160448 7698 160512
rect 7762 160448 7778 160512
rect 7842 160448 7858 160512
rect 7922 160448 7930 160512
rect 7610 160447 7930 160448
rect 2610 159968 2930 159969
rect 2610 159904 2618 159968
rect 2682 159904 2698 159968
rect 2762 159904 2778 159968
rect 2842 159904 2858 159968
rect 2922 159904 2930 159968
rect 2610 159903 2930 159904
rect 5944 159968 6264 159969
rect 5944 159904 5952 159968
rect 6016 159904 6032 159968
rect 6096 159904 6112 159968
rect 6176 159904 6192 159968
rect 6256 159904 6264 159968
rect 5944 159903 6264 159904
rect 4277 159424 4597 159425
rect 4277 159360 4285 159424
rect 4349 159360 4365 159424
rect 4429 159360 4445 159424
rect 4509 159360 4525 159424
rect 4589 159360 4597 159424
rect 4277 159359 4597 159360
rect 7610 159424 7930 159425
rect 7610 159360 7618 159424
rect 7682 159360 7698 159424
rect 7762 159360 7778 159424
rect 7842 159360 7858 159424
rect 7922 159360 7930 159424
rect 7610 159359 7930 159360
rect 2610 158880 2930 158881
rect 2610 158816 2618 158880
rect 2682 158816 2698 158880
rect 2762 158816 2778 158880
rect 2842 158816 2858 158880
rect 2922 158816 2930 158880
rect 2610 158815 2930 158816
rect 5944 158880 6264 158881
rect 5944 158816 5952 158880
rect 6016 158816 6032 158880
rect 6096 158816 6112 158880
rect 6176 158816 6192 158880
rect 6256 158816 6264 158880
rect 5944 158815 6264 158816
rect 4277 158336 4597 158337
rect 4277 158272 4285 158336
rect 4349 158272 4365 158336
rect 4429 158272 4445 158336
rect 4509 158272 4525 158336
rect 4589 158272 4597 158336
rect 4277 158271 4597 158272
rect 7610 158336 7930 158337
rect 7610 158272 7618 158336
rect 7682 158272 7698 158336
rect 7762 158272 7778 158336
rect 7842 158272 7858 158336
rect 7922 158272 7930 158336
rect 7610 158271 7930 158272
rect 2610 157792 2930 157793
rect 2610 157728 2618 157792
rect 2682 157728 2698 157792
rect 2762 157728 2778 157792
rect 2842 157728 2858 157792
rect 2922 157728 2930 157792
rect 2610 157727 2930 157728
rect 5944 157792 6264 157793
rect 5944 157728 5952 157792
rect 6016 157728 6032 157792
rect 6096 157728 6112 157792
rect 6176 157728 6192 157792
rect 6256 157728 6264 157792
rect 5944 157727 6264 157728
rect 4277 157248 4597 157249
rect 4277 157184 4285 157248
rect 4349 157184 4365 157248
rect 4429 157184 4445 157248
rect 4509 157184 4525 157248
rect 4589 157184 4597 157248
rect 4277 157183 4597 157184
rect 7610 157248 7930 157249
rect 7610 157184 7618 157248
rect 7682 157184 7698 157248
rect 7762 157184 7778 157248
rect 7842 157184 7858 157248
rect 7922 157184 7930 157248
rect 7610 157183 7930 157184
rect 2610 156704 2930 156705
rect 2610 156640 2618 156704
rect 2682 156640 2698 156704
rect 2762 156640 2778 156704
rect 2842 156640 2858 156704
rect 2922 156640 2930 156704
rect 2610 156639 2930 156640
rect 5944 156704 6264 156705
rect 5944 156640 5952 156704
rect 6016 156640 6032 156704
rect 6096 156640 6112 156704
rect 6176 156640 6192 156704
rect 6256 156640 6264 156704
rect 5944 156639 6264 156640
rect 4277 156160 4597 156161
rect 4277 156096 4285 156160
rect 4349 156096 4365 156160
rect 4429 156096 4445 156160
rect 4509 156096 4525 156160
rect 4589 156096 4597 156160
rect 4277 156095 4597 156096
rect 7610 156160 7930 156161
rect 7610 156096 7618 156160
rect 7682 156096 7698 156160
rect 7762 156096 7778 156160
rect 7842 156096 7858 156160
rect 7922 156096 7930 156160
rect 7610 156095 7930 156096
rect 2610 155616 2930 155617
rect 2610 155552 2618 155616
rect 2682 155552 2698 155616
rect 2762 155552 2778 155616
rect 2842 155552 2858 155616
rect 2922 155552 2930 155616
rect 2610 155551 2930 155552
rect 5944 155616 6264 155617
rect 5944 155552 5952 155616
rect 6016 155552 6032 155616
rect 6096 155552 6112 155616
rect 6176 155552 6192 155616
rect 6256 155552 6264 155616
rect 5944 155551 6264 155552
rect 4277 155072 4597 155073
rect 4277 155008 4285 155072
rect 4349 155008 4365 155072
rect 4429 155008 4445 155072
rect 4509 155008 4525 155072
rect 4589 155008 4597 155072
rect 4277 155007 4597 155008
rect 7610 155072 7930 155073
rect 7610 155008 7618 155072
rect 7682 155008 7698 155072
rect 7762 155008 7778 155072
rect 7842 155008 7858 155072
rect 7922 155008 7930 155072
rect 7610 155007 7930 155008
rect 2610 154528 2930 154529
rect 2610 154464 2618 154528
rect 2682 154464 2698 154528
rect 2762 154464 2778 154528
rect 2842 154464 2858 154528
rect 2922 154464 2930 154528
rect 2610 154463 2930 154464
rect 5944 154528 6264 154529
rect 5944 154464 5952 154528
rect 6016 154464 6032 154528
rect 6096 154464 6112 154528
rect 6176 154464 6192 154528
rect 6256 154464 6264 154528
rect 5944 154463 6264 154464
rect 4277 153984 4597 153985
rect 4277 153920 4285 153984
rect 4349 153920 4365 153984
rect 4429 153920 4445 153984
rect 4509 153920 4525 153984
rect 4589 153920 4597 153984
rect 4277 153919 4597 153920
rect 7610 153984 7930 153985
rect 7610 153920 7618 153984
rect 7682 153920 7698 153984
rect 7762 153920 7778 153984
rect 7842 153920 7858 153984
rect 7922 153920 7930 153984
rect 7610 153919 7930 153920
rect 2610 153440 2930 153441
rect 2610 153376 2618 153440
rect 2682 153376 2698 153440
rect 2762 153376 2778 153440
rect 2842 153376 2858 153440
rect 2922 153376 2930 153440
rect 2610 153375 2930 153376
rect 5944 153440 6264 153441
rect 5944 153376 5952 153440
rect 6016 153376 6032 153440
rect 6096 153376 6112 153440
rect 6176 153376 6192 153440
rect 6256 153376 6264 153440
rect 5944 153375 6264 153376
rect 4277 152896 4597 152897
rect 4277 152832 4285 152896
rect 4349 152832 4365 152896
rect 4429 152832 4445 152896
rect 4509 152832 4525 152896
rect 4589 152832 4597 152896
rect 4277 152831 4597 152832
rect 7610 152896 7930 152897
rect 7610 152832 7618 152896
rect 7682 152832 7698 152896
rect 7762 152832 7778 152896
rect 7842 152832 7858 152896
rect 7922 152832 7930 152896
rect 7610 152831 7930 152832
rect 2610 152352 2930 152353
rect 2610 152288 2618 152352
rect 2682 152288 2698 152352
rect 2762 152288 2778 152352
rect 2842 152288 2858 152352
rect 2922 152288 2930 152352
rect 2610 152287 2930 152288
rect 5944 152352 6264 152353
rect 5944 152288 5952 152352
rect 6016 152288 6032 152352
rect 6096 152288 6112 152352
rect 6176 152288 6192 152352
rect 6256 152288 6264 152352
rect 5944 152287 6264 152288
rect 4277 151808 4597 151809
rect 4277 151744 4285 151808
rect 4349 151744 4365 151808
rect 4429 151744 4445 151808
rect 4509 151744 4525 151808
rect 4589 151744 4597 151808
rect 4277 151743 4597 151744
rect 7610 151808 7930 151809
rect 7610 151744 7618 151808
rect 7682 151744 7698 151808
rect 7762 151744 7778 151808
rect 7842 151744 7858 151808
rect 7922 151744 7930 151808
rect 7610 151743 7930 151744
rect 2610 151264 2930 151265
rect 2610 151200 2618 151264
rect 2682 151200 2698 151264
rect 2762 151200 2778 151264
rect 2842 151200 2858 151264
rect 2922 151200 2930 151264
rect 2610 151199 2930 151200
rect 5944 151264 6264 151265
rect 5944 151200 5952 151264
rect 6016 151200 6032 151264
rect 6096 151200 6112 151264
rect 6176 151200 6192 151264
rect 6256 151200 6264 151264
rect 5944 151199 6264 151200
rect 4277 150720 4597 150721
rect 4277 150656 4285 150720
rect 4349 150656 4365 150720
rect 4429 150656 4445 150720
rect 4509 150656 4525 150720
rect 4589 150656 4597 150720
rect 4277 150655 4597 150656
rect 7610 150720 7930 150721
rect 7610 150656 7618 150720
rect 7682 150656 7698 150720
rect 7762 150656 7778 150720
rect 7842 150656 7858 150720
rect 7922 150656 7930 150720
rect 7610 150655 7930 150656
rect 3509 150378 3575 150381
rect 3509 150376 9690 150378
rect 3509 150320 3514 150376
rect 3570 150320 9690 150376
rect 3509 150318 9690 150320
rect 3509 150315 3575 150318
rect 2610 150176 2930 150177
rect 2610 150112 2618 150176
rect 2682 150112 2698 150176
rect 2762 150112 2778 150176
rect 2842 150112 2858 150176
rect 2922 150112 2930 150176
rect 2610 150111 2930 150112
rect 5944 150176 6264 150177
rect 5944 150112 5952 150176
rect 6016 150112 6032 150176
rect 6096 150112 6112 150176
rect 6176 150112 6192 150176
rect 6256 150112 6264 150176
rect 5944 150111 6264 150112
rect 9630 149864 9690 150318
rect 9520 149744 10000 149864
rect 4277 149632 4597 149633
rect 4277 149568 4285 149632
rect 4349 149568 4365 149632
rect 4429 149568 4445 149632
rect 4509 149568 4525 149632
rect 4589 149568 4597 149632
rect 4277 149567 4597 149568
rect 7610 149632 7930 149633
rect 7610 149568 7618 149632
rect 7682 149568 7698 149632
rect 7762 149568 7778 149632
rect 7842 149568 7858 149632
rect 7922 149568 7930 149632
rect 7610 149567 7930 149568
rect 2610 149088 2930 149089
rect 2610 149024 2618 149088
rect 2682 149024 2698 149088
rect 2762 149024 2778 149088
rect 2842 149024 2858 149088
rect 2922 149024 2930 149088
rect 2610 149023 2930 149024
rect 5944 149088 6264 149089
rect 5944 149024 5952 149088
rect 6016 149024 6032 149088
rect 6096 149024 6112 149088
rect 6176 149024 6192 149088
rect 6256 149024 6264 149088
rect 5944 149023 6264 149024
rect 4277 148544 4597 148545
rect 4277 148480 4285 148544
rect 4349 148480 4365 148544
rect 4429 148480 4445 148544
rect 4509 148480 4525 148544
rect 4589 148480 4597 148544
rect 4277 148479 4597 148480
rect 7610 148544 7930 148545
rect 7610 148480 7618 148544
rect 7682 148480 7698 148544
rect 7762 148480 7778 148544
rect 7842 148480 7858 148544
rect 7922 148480 7930 148544
rect 7610 148479 7930 148480
rect 2610 148000 2930 148001
rect 2610 147936 2618 148000
rect 2682 147936 2698 148000
rect 2762 147936 2778 148000
rect 2842 147936 2858 148000
rect 2922 147936 2930 148000
rect 2610 147935 2930 147936
rect 5944 148000 6264 148001
rect 5944 147936 5952 148000
rect 6016 147936 6032 148000
rect 6096 147936 6112 148000
rect 6176 147936 6192 148000
rect 6256 147936 6264 148000
rect 5944 147935 6264 147936
rect 4277 147456 4597 147457
rect 4277 147392 4285 147456
rect 4349 147392 4365 147456
rect 4429 147392 4445 147456
rect 4509 147392 4525 147456
rect 4589 147392 4597 147456
rect 4277 147391 4597 147392
rect 7610 147456 7930 147457
rect 7610 147392 7618 147456
rect 7682 147392 7698 147456
rect 7762 147392 7778 147456
rect 7842 147392 7858 147456
rect 7922 147392 7930 147456
rect 7610 147391 7930 147392
rect 2610 146912 2930 146913
rect 2610 146848 2618 146912
rect 2682 146848 2698 146912
rect 2762 146848 2778 146912
rect 2842 146848 2858 146912
rect 2922 146848 2930 146912
rect 2610 146847 2930 146848
rect 5944 146912 6264 146913
rect 5944 146848 5952 146912
rect 6016 146848 6032 146912
rect 6096 146848 6112 146912
rect 6176 146848 6192 146912
rect 6256 146848 6264 146912
rect 5944 146847 6264 146848
rect 4277 146368 4597 146369
rect 4277 146304 4285 146368
rect 4349 146304 4365 146368
rect 4429 146304 4445 146368
rect 4509 146304 4525 146368
rect 4589 146304 4597 146368
rect 4277 146303 4597 146304
rect 7610 146368 7930 146369
rect 7610 146304 7618 146368
rect 7682 146304 7698 146368
rect 7762 146304 7778 146368
rect 7842 146304 7858 146368
rect 7922 146304 7930 146368
rect 7610 146303 7930 146304
rect 2610 145824 2930 145825
rect 2610 145760 2618 145824
rect 2682 145760 2698 145824
rect 2762 145760 2778 145824
rect 2842 145760 2858 145824
rect 2922 145760 2930 145824
rect 2610 145759 2930 145760
rect 5944 145824 6264 145825
rect 5944 145760 5952 145824
rect 6016 145760 6032 145824
rect 6096 145760 6112 145824
rect 6176 145760 6192 145824
rect 6256 145760 6264 145824
rect 5944 145759 6264 145760
rect 4277 145280 4597 145281
rect 4277 145216 4285 145280
rect 4349 145216 4365 145280
rect 4429 145216 4445 145280
rect 4509 145216 4525 145280
rect 4589 145216 4597 145280
rect 4277 145215 4597 145216
rect 7610 145280 7930 145281
rect 7610 145216 7618 145280
rect 7682 145216 7698 145280
rect 7762 145216 7778 145280
rect 7842 145216 7858 145280
rect 7922 145216 7930 145280
rect 7610 145215 7930 145216
rect 2610 144736 2930 144737
rect 2610 144672 2618 144736
rect 2682 144672 2698 144736
rect 2762 144672 2778 144736
rect 2842 144672 2858 144736
rect 2922 144672 2930 144736
rect 2610 144671 2930 144672
rect 5944 144736 6264 144737
rect 5944 144672 5952 144736
rect 6016 144672 6032 144736
rect 6096 144672 6112 144736
rect 6176 144672 6192 144736
rect 6256 144672 6264 144736
rect 5944 144671 6264 144672
rect 4277 144192 4597 144193
rect 4277 144128 4285 144192
rect 4349 144128 4365 144192
rect 4429 144128 4445 144192
rect 4509 144128 4525 144192
rect 4589 144128 4597 144192
rect 4277 144127 4597 144128
rect 7610 144192 7930 144193
rect 7610 144128 7618 144192
rect 7682 144128 7698 144192
rect 7762 144128 7778 144192
rect 7842 144128 7858 144192
rect 7922 144128 7930 144192
rect 7610 144127 7930 144128
rect 2610 143648 2930 143649
rect 2610 143584 2618 143648
rect 2682 143584 2698 143648
rect 2762 143584 2778 143648
rect 2842 143584 2858 143648
rect 2922 143584 2930 143648
rect 2610 143583 2930 143584
rect 5944 143648 6264 143649
rect 5944 143584 5952 143648
rect 6016 143584 6032 143648
rect 6096 143584 6112 143648
rect 6176 143584 6192 143648
rect 6256 143584 6264 143648
rect 5944 143583 6264 143584
rect 4277 143104 4597 143105
rect 4277 143040 4285 143104
rect 4349 143040 4365 143104
rect 4429 143040 4445 143104
rect 4509 143040 4525 143104
rect 4589 143040 4597 143104
rect 4277 143039 4597 143040
rect 7610 143104 7930 143105
rect 7610 143040 7618 143104
rect 7682 143040 7698 143104
rect 7762 143040 7778 143104
rect 7842 143040 7858 143104
rect 7922 143040 7930 143104
rect 7610 143039 7930 143040
rect 2610 142560 2930 142561
rect 2610 142496 2618 142560
rect 2682 142496 2698 142560
rect 2762 142496 2778 142560
rect 2842 142496 2858 142560
rect 2922 142496 2930 142560
rect 2610 142495 2930 142496
rect 5944 142560 6264 142561
rect 5944 142496 5952 142560
rect 6016 142496 6032 142560
rect 6096 142496 6112 142560
rect 6176 142496 6192 142560
rect 6256 142496 6264 142560
rect 5944 142495 6264 142496
rect 4277 142016 4597 142017
rect 4277 141952 4285 142016
rect 4349 141952 4365 142016
rect 4429 141952 4445 142016
rect 4509 141952 4525 142016
rect 4589 141952 4597 142016
rect 4277 141951 4597 141952
rect 7610 142016 7930 142017
rect 7610 141952 7618 142016
rect 7682 141952 7698 142016
rect 7762 141952 7778 142016
rect 7842 141952 7858 142016
rect 7922 141952 7930 142016
rect 7610 141951 7930 141952
rect 2610 141472 2930 141473
rect 2610 141408 2618 141472
rect 2682 141408 2698 141472
rect 2762 141408 2778 141472
rect 2842 141408 2858 141472
rect 2922 141408 2930 141472
rect 2610 141407 2930 141408
rect 5944 141472 6264 141473
rect 5944 141408 5952 141472
rect 6016 141408 6032 141472
rect 6096 141408 6112 141472
rect 6176 141408 6192 141472
rect 6256 141408 6264 141472
rect 5944 141407 6264 141408
rect 4277 140928 4597 140929
rect 4277 140864 4285 140928
rect 4349 140864 4365 140928
rect 4429 140864 4445 140928
rect 4509 140864 4525 140928
rect 4589 140864 4597 140928
rect 4277 140863 4597 140864
rect 7610 140928 7930 140929
rect 7610 140864 7618 140928
rect 7682 140864 7698 140928
rect 7762 140864 7778 140928
rect 7842 140864 7858 140928
rect 7922 140864 7930 140928
rect 7610 140863 7930 140864
rect 2610 140384 2930 140385
rect 2610 140320 2618 140384
rect 2682 140320 2698 140384
rect 2762 140320 2778 140384
rect 2842 140320 2858 140384
rect 2922 140320 2930 140384
rect 2610 140319 2930 140320
rect 5944 140384 6264 140385
rect 5944 140320 5952 140384
rect 6016 140320 6032 140384
rect 6096 140320 6112 140384
rect 6176 140320 6192 140384
rect 6256 140320 6264 140384
rect 5944 140319 6264 140320
rect 4277 139840 4597 139841
rect 4277 139776 4285 139840
rect 4349 139776 4365 139840
rect 4429 139776 4445 139840
rect 4509 139776 4525 139840
rect 4589 139776 4597 139840
rect 4277 139775 4597 139776
rect 7610 139840 7930 139841
rect 7610 139776 7618 139840
rect 7682 139776 7698 139840
rect 7762 139776 7778 139840
rect 7842 139776 7858 139840
rect 7922 139776 7930 139840
rect 7610 139775 7930 139776
rect 2610 139296 2930 139297
rect 2610 139232 2618 139296
rect 2682 139232 2698 139296
rect 2762 139232 2778 139296
rect 2842 139232 2858 139296
rect 2922 139232 2930 139296
rect 2610 139231 2930 139232
rect 5944 139296 6264 139297
rect 5944 139232 5952 139296
rect 6016 139232 6032 139296
rect 6096 139232 6112 139296
rect 6176 139232 6192 139296
rect 6256 139232 6264 139296
rect 5944 139231 6264 139232
rect 4277 138752 4597 138753
rect 4277 138688 4285 138752
rect 4349 138688 4365 138752
rect 4429 138688 4445 138752
rect 4509 138688 4525 138752
rect 4589 138688 4597 138752
rect 4277 138687 4597 138688
rect 7610 138752 7930 138753
rect 7610 138688 7618 138752
rect 7682 138688 7698 138752
rect 7762 138688 7778 138752
rect 7842 138688 7858 138752
rect 7922 138688 7930 138752
rect 7610 138687 7930 138688
rect 2610 138208 2930 138209
rect 2610 138144 2618 138208
rect 2682 138144 2698 138208
rect 2762 138144 2778 138208
rect 2842 138144 2858 138208
rect 2922 138144 2930 138208
rect 2610 138143 2930 138144
rect 5944 138208 6264 138209
rect 5944 138144 5952 138208
rect 6016 138144 6032 138208
rect 6096 138144 6112 138208
rect 6176 138144 6192 138208
rect 6256 138144 6264 138208
rect 5944 138143 6264 138144
rect 4277 137664 4597 137665
rect 4277 137600 4285 137664
rect 4349 137600 4365 137664
rect 4429 137600 4445 137664
rect 4509 137600 4525 137664
rect 4589 137600 4597 137664
rect 4277 137599 4597 137600
rect 7610 137664 7930 137665
rect 7610 137600 7618 137664
rect 7682 137600 7698 137664
rect 7762 137600 7778 137664
rect 7842 137600 7858 137664
rect 7922 137600 7930 137664
rect 7610 137599 7930 137600
rect 2610 137120 2930 137121
rect 2610 137056 2618 137120
rect 2682 137056 2698 137120
rect 2762 137056 2778 137120
rect 2842 137056 2858 137120
rect 2922 137056 2930 137120
rect 2610 137055 2930 137056
rect 5944 137120 6264 137121
rect 5944 137056 5952 137120
rect 6016 137056 6032 137120
rect 6096 137056 6112 137120
rect 6176 137056 6192 137120
rect 6256 137056 6264 137120
rect 5944 137055 6264 137056
rect 4277 136576 4597 136577
rect 4277 136512 4285 136576
rect 4349 136512 4365 136576
rect 4429 136512 4445 136576
rect 4509 136512 4525 136576
rect 4589 136512 4597 136576
rect 4277 136511 4597 136512
rect 7610 136576 7930 136577
rect 7610 136512 7618 136576
rect 7682 136512 7698 136576
rect 7762 136512 7778 136576
rect 7842 136512 7858 136576
rect 7922 136512 7930 136576
rect 7610 136511 7930 136512
rect 2610 136032 2930 136033
rect 2610 135968 2618 136032
rect 2682 135968 2698 136032
rect 2762 135968 2778 136032
rect 2842 135968 2858 136032
rect 2922 135968 2930 136032
rect 2610 135967 2930 135968
rect 5944 136032 6264 136033
rect 5944 135968 5952 136032
rect 6016 135968 6032 136032
rect 6096 135968 6112 136032
rect 6176 135968 6192 136032
rect 6256 135968 6264 136032
rect 5944 135967 6264 135968
rect 4277 135488 4597 135489
rect 4277 135424 4285 135488
rect 4349 135424 4365 135488
rect 4429 135424 4445 135488
rect 4509 135424 4525 135488
rect 4589 135424 4597 135488
rect 4277 135423 4597 135424
rect 7610 135488 7930 135489
rect 7610 135424 7618 135488
rect 7682 135424 7698 135488
rect 7762 135424 7778 135488
rect 7842 135424 7858 135488
rect 7922 135424 7930 135488
rect 7610 135423 7930 135424
rect 2610 134944 2930 134945
rect 2610 134880 2618 134944
rect 2682 134880 2698 134944
rect 2762 134880 2778 134944
rect 2842 134880 2858 134944
rect 2922 134880 2930 134944
rect 2610 134879 2930 134880
rect 5944 134944 6264 134945
rect 5944 134880 5952 134944
rect 6016 134880 6032 134944
rect 6096 134880 6112 134944
rect 6176 134880 6192 134944
rect 6256 134880 6264 134944
rect 5944 134879 6264 134880
rect 4277 134400 4597 134401
rect 4277 134336 4285 134400
rect 4349 134336 4365 134400
rect 4429 134336 4445 134400
rect 4509 134336 4525 134400
rect 4589 134336 4597 134400
rect 4277 134335 4597 134336
rect 7610 134400 7930 134401
rect 7610 134336 7618 134400
rect 7682 134336 7698 134400
rect 7762 134336 7778 134400
rect 7842 134336 7858 134400
rect 7922 134336 7930 134400
rect 7610 134335 7930 134336
rect 2610 133856 2930 133857
rect 2610 133792 2618 133856
rect 2682 133792 2698 133856
rect 2762 133792 2778 133856
rect 2842 133792 2858 133856
rect 2922 133792 2930 133856
rect 2610 133791 2930 133792
rect 5944 133856 6264 133857
rect 5944 133792 5952 133856
rect 6016 133792 6032 133856
rect 6096 133792 6112 133856
rect 6176 133792 6192 133856
rect 6256 133792 6264 133856
rect 5944 133791 6264 133792
rect 4277 133312 4597 133313
rect 4277 133248 4285 133312
rect 4349 133248 4365 133312
rect 4429 133248 4445 133312
rect 4509 133248 4525 133312
rect 4589 133248 4597 133312
rect 4277 133247 4597 133248
rect 7610 133312 7930 133313
rect 7610 133248 7618 133312
rect 7682 133248 7698 133312
rect 7762 133248 7778 133312
rect 7842 133248 7858 133312
rect 7922 133248 7930 133312
rect 7610 133247 7930 133248
rect 2610 132768 2930 132769
rect 2610 132704 2618 132768
rect 2682 132704 2698 132768
rect 2762 132704 2778 132768
rect 2842 132704 2858 132768
rect 2922 132704 2930 132768
rect 2610 132703 2930 132704
rect 5944 132768 6264 132769
rect 5944 132704 5952 132768
rect 6016 132704 6032 132768
rect 6096 132704 6112 132768
rect 6176 132704 6192 132768
rect 6256 132704 6264 132768
rect 5944 132703 6264 132704
rect 4277 132224 4597 132225
rect 4277 132160 4285 132224
rect 4349 132160 4365 132224
rect 4429 132160 4445 132224
rect 4509 132160 4525 132224
rect 4589 132160 4597 132224
rect 4277 132159 4597 132160
rect 7610 132224 7930 132225
rect 7610 132160 7618 132224
rect 7682 132160 7698 132224
rect 7762 132160 7778 132224
rect 7842 132160 7858 132224
rect 7922 132160 7930 132224
rect 7610 132159 7930 132160
rect 2610 131680 2930 131681
rect 2610 131616 2618 131680
rect 2682 131616 2698 131680
rect 2762 131616 2778 131680
rect 2842 131616 2858 131680
rect 2922 131616 2930 131680
rect 2610 131615 2930 131616
rect 5944 131680 6264 131681
rect 5944 131616 5952 131680
rect 6016 131616 6032 131680
rect 6096 131616 6112 131680
rect 6176 131616 6192 131680
rect 6256 131616 6264 131680
rect 5944 131615 6264 131616
rect 4277 131136 4597 131137
rect 4277 131072 4285 131136
rect 4349 131072 4365 131136
rect 4429 131072 4445 131136
rect 4509 131072 4525 131136
rect 4589 131072 4597 131136
rect 4277 131071 4597 131072
rect 7610 131136 7930 131137
rect 7610 131072 7618 131136
rect 7682 131072 7698 131136
rect 7762 131072 7778 131136
rect 7842 131072 7858 131136
rect 7922 131072 7930 131136
rect 7610 131071 7930 131072
rect 2610 130592 2930 130593
rect 2610 130528 2618 130592
rect 2682 130528 2698 130592
rect 2762 130528 2778 130592
rect 2842 130528 2858 130592
rect 2922 130528 2930 130592
rect 2610 130527 2930 130528
rect 5944 130592 6264 130593
rect 5944 130528 5952 130592
rect 6016 130528 6032 130592
rect 6096 130528 6112 130592
rect 6176 130528 6192 130592
rect 6256 130528 6264 130592
rect 5944 130527 6264 130528
rect 4277 130048 4597 130049
rect 4277 129984 4285 130048
rect 4349 129984 4365 130048
rect 4429 129984 4445 130048
rect 4509 129984 4525 130048
rect 4589 129984 4597 130048
rect 4277 129983 4597 129984
rect 7610 130048 7930 130049
rect 7610 129984 7618 130048
rect 7682 129984 7698 130048
rect 7762 129984 7778 130048
rect 7842 129984 7858 130048
rect 7922 129984 7930 130048
rect 7610 129983 7930 129984
rect 2610 129504 2930 129505
rect 2610 129440 2618 129504
rect 2682 129440 2698 129504
rect 2762 129440 2778 129504
rect 2842 129440 2858 129504
rect 2922 129440 2930 129504
rect 2610 129439 2930 129440
rect 5944 129504 6264 129505
rect 5944 129440 5952 129504
rect 6016 129440 6032 129504
rect 6096 129440 6112 129504
rect 6176 129440 6192 129504
rect 6256 129440 6264 129504
rect 5944 129439 6264 129440
rect 4277 128960 4597 128961
rect 4277 128896 4285 128960
rect 4349 128896 4365 128960
rect 4429 128896 4445 128960
rect 4509 128896 4525 128960
rect 4589 128896 4597 128960
rect 4277 128895 4597 128896
rect 7610 128960 7930 128961
rect 7610 128896 7618 128960
rect 7682 128896 7698 128960
rect 7762 128896 7778 128960
rect 7842 128896 7858 128960
rect 7922 128896 7930 128960
rect 7610 128895 7930 128896
rect 2610 128416 2930 128417
rect 2610 128352 2618 128416
rect 2682 128352 2698 128416
rect 2762 128352 2778 128416
rect 2842 128352 2858 128416
rect 2922 128352 2930 128416
rect 2610 128351 2930 128352
rect 5944 128416 6264 128417
rect 5944 128352 5952 128416
rect 6016 128352 6032 128416
rect 6096 128352 6112 128416
rect 6176 128352 6192 128416
rect 6256 128352 6264 128416
rect 5944 128351 6264 128352
rect 4277 127872 4597 127873
rect 4277 127808 4285 127872
rect 4349 127808 4365 127872
rect 4429 127808 4445 127872
rect 4509 127808 4525 127872
rect 4589 127808 4597 127872
rect 4277 127807 4597 127808
rect 7610 127872 7930 127873
rect 7610 127808 7618 127872
rect 7682 127808 7698 127872
rect 7762 127808 7778 127872
rect 7842 127808 7858 127872
rect 7922 127808 7930 127872
rect 7610 127807 7930 127808
rect 2610 127328 2930 127329
rect 2610 127264 2618 127328
rect 2682 127264 2698 127328
rect 2762 127264 2778 127328
rect 2842 127264 2858 127328
rect 2922 127264 2930 127328
rect 2610 127263 2930 127264
rect 5944 127328 6264 127329
rect 5944 127264 5952 127328
rect 6016 127264 6032 127328
rect 6096 127264 6112 127328
rect 6176 127264 6192 127328
rect 6256 127264 6264 127328
rect 5944 127263 6264 127264
rect 4277 126784 4597 126785
rect 4277 126720 4285 126784
rect 4349 126720 4365 126784
rect 4429 126720 4445 126784
rect 4509 126720 4525 126784
rect 4589 126720 4597 126784
rect 4277 126719 4597 126720
rect 7610 126784 7930 126785
rect 7610 126720 7618 126784
rect 7682 126720 7698 126784
rect 7762 126720 7778 126784
rect 7842 126720 7858 126784
rect 7922 126720 7930 126784
rect 7610 126719 7930 126720
rect 2610 126240 2930 126241
rect 2610 126176 2618 126240
rect 2682 126176 2698 126240
rect 2762 126176 2778 126240
rect 2842 126176 2858 126240
rect 2922 126176 2930 126240
rect 2610 126175 2930 126176
rect 5944 126240 6264 126241
rect 5944 126176 5952 126240
rect 6016 126176 6032 126240
rect 6096 126176 6112 126240
rect 6176 126176 6192 126240
rect 6256 126176 6264 126240
rect 5944 126175 6264 126176
rect 4277 125696 4597 125697
rect 4277 125632 4285 125696
rect 4349 125632 4365 125696
rect 4429 125632 4445 125696
rect 4509 125632 4525 125696
rect 4589 125632 4597 125696
rect 4277 125631 4597 125632
rect 7610 125696 7930 125697
rect 7610 125632 7618 125696
rect 7682 125632 7698 125696
rect 7762 125632 7778 125696
rect 7842 125632 7858 125696
rect 7922 125632 7930 125696
rect 7610 125631 7930 125632
rect 2610 125152 2930 125153
rect 2610 125088 2618 125152
rect 2682 125088 2698 125152
rect 2762 125088 2778 125152
rect 2842 125088 2858 125152
rect 2922 125088 2930 125152
rect 2610 125087 2930 125088
rect 5944 125152 6264 125153
rect 5944 125088 5952 125152
rect 6016 125088 6032 125152
rect 6096 125088 6112 125152
rect 6176 125088 6192 125152
rect 6256 125088 6264 125152
rect 5944 125087 6264 125088
rect 4277 124608 4597 124609
rect 4277 124544 4285 124608
rect 4349 124544 4365 124608
rect 4429 124544 4445 124608
rect 4509 124544 4525 124608
rect 4589 124544 4597 124608
rect 4277 124543 4597 124544
rect 7610 124608 7930 124609
rect 7610 124544 7618 124608
rect 7682 124544 7698 124608
rect 7762 124544 7778 124608
rect 7842 124544 7858 124608
rect 7922 124544 7930 124608
rect 7610 124543 7930 124544
rect 2610 124064 2930 124065
rect 2610 124000 2618 124064
rect 2682 124000 2698 124064
rect 2762 124000 2778 124064
rect 2842 124000 2858 124064
rect 2922 124000 2930 124064
rect 2610 123999 2930 124000
rect 5944 124064 6264 124065
rect 5944 124000 5952 124064
rect 6016 124000 6032 124064
rect 6096 124000 6112 124064
rect 6176 124000 6192 124064
rect 6256 124000 6264 124064
rect 5944 123999 6264 124000
rect 4277 123520 4597 123521
rect 4277 123456 4285 123520
rect 4349 123456 4365 123520
rect 4429 123456 4445 123520
rect 4509 123456 4525 123520
rect 4589 123456 4597 123520
rect 4277 123455 4597 123456
rect 7610 123520 7930 123521
rect 7610 123456 7618 123520
rect 7682 123456 7698 123520
rect 7762 123456 7778 123520
rect 7842 123456 7858 123520
rect 7922 123456 7930 123520
rect 7610 123455 7930 123456
rect 2610 122976 2930 122977
rect 2610 122912 2618 122976
rect 2682 122912 2698 122976
rect 2762 122912 2778 122976
rect 2842 122912 2858 122976
rect 2922 122912 2930 122976
rect 2610 122911 2930 122912
rect 5944 122976 6264 122977
rect 5944 122912 5952 122976
rect 6016 122912 6032 122976
rect 6096 122912 6112 122976
rect 6176 122912 6192 122976
rect 6256 122912 6264 122976
rect 5944 122911 6264 122912
rect 4277 122432 4597 122433
rect 4277 122368 4285 122432
rect 4349 122368 4365 122432
rect 4429 122368 4445 122432
rect 4509 122368 4525 122432
rect 4589 122368 4597 122432
rect 4277 122367 4597 122368
rect 7610 122432 7930 122433
rect 7610 122368 7618 122432
rect 7682 122368 7698 122432
rect 7762 122368 7778 122432
rect 7842 122368 7858 122432
rect 7922 122368 7930 122432
rect 7610 122367 7930 122368
rect 2610 121888 2930 121889
rect 2610 121824 2618 121888
rect 2682 121824 2698 121888
rect 2762 121824 2778 121888
rect 2842 121824 2858 121888
rect 2922 121824 2930 121888
rect 2610 121823 2930 121824
rect 5944 121888 6264 121889
rect 5944 121824 5952 121888
rect 6016 121824 6032 121888
rect 6096 121824 6112 121888
rect 6176 121824 6192 121888
rect 6256 121824 6264 121888
rect 5944 121823 6264 121824
rect 4277 121344 4597 121345
rect 4277 121280 4285 121344
rect 4349 121280 4365 121344
rect 4429 121280 4445 121344
rect 4509 121280 4525 121344
rect 4589 121280 4597 121344
rect 4277 121279 4597 121280
rect 7610 121344 7930 121345
rect 7610 121280 7618 121344
rect 7682 121280 7698 121344
rect 7762 121280 7778 121344
rect 7842 121280 7858 121344
rect 7922 121280 7930 121344
rect 7610 121279 7930 121280
rect 2610 120800 2930 120801
rect 2610 120736 2618 120800
rect 2682 120736 2698 120800
rect 2762 120736 2778 120800
rect 2842 120736 2858 120800
rect 2922 120736 2930 120800
rect 2610 120735 2930 120736
rect 5944 120800 6264 120801
rect 5944 120736 5952 120800
rect 6016 120736 6032 120800
rect 6096 120736 6112 120800
rect 6176 120736 6192 120800
rect 6256 120736 6264 120800
rect 5944 120735 6264 120736
rect 4277 120256 4597 120257
rect 4277 120192 4285 120256
rect 4349 120192 4365 120256
rect 4429 120192 4445 120256
rect 4509 120192 4525 120256
rect 4589 120192 4597 120256
rect 4277 120191 4597 120192
rect 7610 120256 7930 120257
rect 7610 120192 7618 120256
rect 7682 120192 7698 120256
rect 7762 120192 7778 120256
rect 7842 120192 7858 120256
rect 7922 120192 7930 120256
rect 7610 120191 7930 120192
rect 2610 119712 2930 119713
rect 2610 119648 2618 119712
rect 2682 119648 2698 119712
rect 2762 119648 2778 119712
rect 2842 119648 2858 119712
rect 2922 119648 2930 119712
rect 2610 119647 2930 119648
rect 5944 119712 6264 119713
rect 5944 119648 5952 119712
rect 6016 119648 6032 119712
rect 6096 119648 6112 119712
rect 6176 119648 6192 119712
rect 6256 119648 6264 119712
rect 5944 119647 6264 119648
rect 4277 119168 4597 119169
rect 4277 119104 4285 119168
rect 4349 119104 4365 119168
rect 4429 119104 4445 119168
rect 4509 119104 4525 119168
rect 4589 119104 4597 119168
rect 4277 119103 4597 119104
rect 7610 119168 7930 119169
rect 7610 119104 7618 119168
rect 7682 119104 7698 119168
rect 7762 119104 7778 119168
rect 7842 119104 7858 119168
rect 7922 119104 7930 119168
rect 7610 119103 7930 119104
rect 0 118824 480 118856
rect 0 118768 18 118824
rect 74 118768 480 118824
rect 0 118736 480 118768
rect 2610 118624 2930 118625
rect 2610 118560 2618 118624
rect 2682 118560 2698 118624
rect 2762 118560 2778 118624
rect 2842 118560 2858 118624
rect 2922 118560 2930 118624
rect 2610 118559 2930 118560
rect 5944 118624 6264 118625
rect 5944 118560 5952 118624
rect 6016 118560 6032 118624
rect 6096 118560 6112 118624
rect 6176 118560 6192 118624
rect 6256 118560 6264 118624
rect 5944 118559 6264 118560
rect 4277 118080 4597 118081
rect 4277 118016 4285 118080
rect 4349 118016 4365 118080
rect 4429 118016 4445 118080
rect 4509 118016 4525 118080
rect 4589 118016 4597 118080
rect 4277 118015 4597 118016
rect 7610 118080 7930 118081
rect 7610 118016 7618 118080
rect 7682 118016 7698 118080
rect 7762 118016 7778 118080
rect 7842 118016 7858 118080
rect 7922 118016 7930 118080
rect 7610 118015 7930 118016
rect 2610 117536 2930 117537
rect 2610 117472 2618 117536
rect 2682 117472 2698 117536
rect 2762 117472 2778 117536
rect 2842 117472 2858 117536
rect 2922 117472 2930 117536
rect 2610 117471 2930 117472
rect 5944 117536 6264 117537
rect 5944 117472 5952 117536
rect 6016 117472 6032 117536
rect 6096 117472 6112 117536
rect 6176 117472 6192 117536
rect 6256 117472 6264 117536
rect 5944 117471 6264 117472
rect 4277 116992 4597 116993
rect 4277 116928 4285 116992
rect 4349 116928 4365 116992
rect 4429 116928 4445 116992
rect 4509 116928 4525 116992
rect 4589 116928 4597 116992
rect 4277 116927 4597 116928
rect 7610 116992 7930 116993
rect 7610 116928 7618 116992
rect 7682 116928 7698 116992
rect 7762 116928 7778 116992
rect 7842 116928 7858 116992
rect 7922 116928 7930 116992
rect 7610 116927 7930 116928
rect 6729 116786 6795 116789
rect 6729 116784 9690 116786
rect 6729 116728 6734 116784
rect 6790 116728 9690 116784
rect 6729 116726 9690 116728
rect 6729 116723 6795 116726
rect 9630 116544 9690 116726
rect 2610 116448 2930 116449
rect 2610 116384 2618 116448
rect 2682 116384 2698 116448
rect 2762 116384 2778 116448
rect 2842 116384 2858 116448
rect 2922 116384 2930 116448
rect 2610 116383 2930 116384
rect 5944 116448 6264 116449
rect 5944 116384 5952 116448
rect 6016 116384 6032 116448
rect 6096 116384 6112 116448
rect 6176 116384 6192 116448
rect 6256 116384 6264 116448
rect 9520 116424 10000 116544
rect 5944 116383 6264 116384
rect 4277 115904 4597 115905
rect 4277 115840 4285 115904
rect 4349 115840 4365 115904
rect 4429 115840 4445 115904
rect 4509 115840 4525 115904
rect 4589 115840 4597 115904
rect 4277 115839 4597 115840
rect 7610 115904 7930 115905
rect 7610 115840 7618 115904
rect 7682 115840 7698 115904
rect 7762 115840 7778 115904
rect 7842 115840 7858 115904
rect 7922 115840 7930 115904
rect 7610 115839 7930 115840
rect 2610 115360 2930 115361
rect 2610 115296 2618 115360
rect 2682 115296 2698 115360
rect 2762 115296 2778 115360
rect 2842 115296 2858 115360
rect 2922 115296 2930 115360
rect 2610 115295 2930 115296
rect 5944 115360 6264 115361
rect 5944 115296 5952 115360
rect 6016 115296 6032 115360
rect 6096 115296 6112 115360
rect 6176 115296 6192 115360
rect 6256 115296 6264 115360
rect 5944 115295 6264 115296
rect 4277 114816 4597 114817
rect 4277 114752 4285 114816
rect 4349 114752 4365 114816
rect 4429 114752 4445 114816
rect 4509 114752 4525 114816
rect 4589 114752 4597 114816
rect 4277 114751 4597 114752
rect 7610 114816 7930 114817
rect 7610 114752 7618 114816
rect 7682 114752 7698 114816
rect 7762 114752 7778 114816
rect 7842 114752 7858 114816
rect 7922 114752 7930 114816
rect 7610 114751 7930 114752
rect 2610 114272 2930 114273
rect 2610 114208 2618 114272
rect 2682 114208 2698 114272
rect 2762 114208 2778 114272
rect 2842 114208 2858 114272
rect 2922 114208 2930 114272
rect 2610 114207 2930 114208
rect 5944 114272 6264 114273
rect 5944 114208 5952 114272
rect 6016 114208 6032 114272
rect 6096 114208 6112 114272
rect 6176 114208 6192 114272
rect 6256 114208 6264 114272
rect 5944 114207 6264 114208
rect 4277 113728 4597 113729
rect 4277 113664 4285 113728
rect 4349 113664 4365 113728
rect 4429 113664 4445 113728
rect 4509 113664 4525 113728
rect 4589 113664 4597 113728
rect 4277 113663 4597 113664
rect 7610 113728 7930 113729
rect 7610 113664 7618 113728
rect 7682 113664 7698 113728
rect 7762 113664 7778 113728
rect 7842 113664 7858 113728
rect 7922 113664 7930 113728
rect 7610 113663 7930 113664
rect 2610 113184 2930 113185
rect 2610 113120 2618 113184
rect 2682 113120 2698 113184
rect 2762 113120 2778 113184
rect 2842 113120 2858 113184
rect 2922 113120 2930 113184
rect 2610 113119 2930 113120
rect 5944 113184 6264 113185
rect 5944 113120 5952 113184
rect 6016 113120 6032 113184
rect 6096 113120 6112 113184
rect 6176 113120 6192 113184
rect 6256 113120 6264 113184
rect 5944 113119 6264 113120
rect 4277 112640 4597 112641
rect 4277 112576 4285 112640
rect 4349 112576 4365 112640
rect 4429 112576 4445 112640
rect 4509 112576 4525 112640
rect 4589 112576 4597 112640
rect 4277 112575 4597 112576
rect 7610 112640 7930 112641
rect 7610 112576 7618 112640
rect 7682 112576 7698 112640
rect 7762 112576 7778 112640
rect 7842 112576 7858 112640
rect 7922 112576 7930 112640
rect 7610 112575 7930 112576
rect 2610 112096 2930 112097
rect 2610 112032 2618 112096
rect 2682 112032 2698 112096
rect 2762 112032 2778 112096
rect 2842 112032 2858 112096
rect 2922 112032 2930 112096
rect 2610 112031 2930 112032
rect 5944 112096 6264 112097
rect 5944 112032 5952 112096
rect 6016 112032 6032 112096
rect 6096 112032 6112 112096
rect 6176 112032 6192 112096
rect 6256 112032 6264 112096
rect 5944 112031 6264 112032
rect 4277 111552 4597 111553
rect 4277 111488 4285 111552
rect 4349 111488 4365 111552
rect 4429 111488 4445 111552
rect 4509 111488 4525 111552
rect 4589 111488 4597 111552
rect 4277 111487 4597 111488
rect 7610 111552 7930 111553
rect 7610 111488 7618 111552
rect 7682 111488 7698 111552
rect 7762 111488 7778 111552
rect 7842 111488 7858 111552
rect 7922 111488 7930 111552
rect 7610 111487 7930 111488
rect 2610 111008 2930 111009
rect 2610 110944 2618 111008
rect 2682 110944 2698 111008
rect 2762 110944 2778 111008
rect 2842 110944 2858 111008
rect 2922 110944 2930 111008
rect 2610 110943 2930 110944
rect 5944 111008 6264 111009
rect 5944 110944 5952 111008
rect 6016 110944 6032 111008
rect 6096 110944 6112 111008
rect 6176 110944 6192 111008
rect 6256 110944 6264 111008
rect 5944 110943 6264 110944
rect 4277 110464 4597 110465
rect 4277 110400 4285 110464
rect 4349 110400 4365 110464
rect 4429 110400 4445 110464
rect 4509 110400 4525 110464
rect 4589 110400 4597 110464
rect 4277 110399 4597 110400
rect 7610 110464 7930 110465
rect 7610 110400 7618 110464
rect 7682 110400 7698 110464
rect 7762 110400 7778 110464
rect 7842 110400 7858 110464
rect 7922 110400 7930 110464
rect 7610 110399 7930 110400
rect 2610 109920 2930 109921
rect 2610 109856 2618 109920
rect 2682 109856 2698 109920
rect 2762 109856 2778 109920
rect 2842 109856 2858 109920
rect 2922 109856 2930 109920
rect 2610 109855 2930 109856
rect 5944 109920 6264 109921
rect 5944 109856 5952 109920
rect 6016 109856 6032 109920
rect 6096 109856 6112 109920
rect 6176 109856 6192 109920
rect 6256 109856 6264 109920
rect 5944 109855 6264 109856
rect 4277 109376 4597 109377
rect 4277 109312 4285 109376
rect 4349 109312 4365 109376
rect 4429 109312 4445 109376
rect 4509 109312 4525 109376
rect 4589 109312 4597 109376
rect 4277 109311 4597 109312
rect 7610 109376 7930 109377
rect 7610 109312 7618 109376
rect 7682 109312 7698 109376
rect 7762 109312 7778 109376
rect 7842 109312 7858 109376
rect 7922 109312 7930 109376
rect 7610 109311 7930 109312
rect 2610 108832 2930 108833
rect 2610 108768 2618 108832
rect 2682 108768 2698 108832
rect 2762 108768 2778 108832
rect 2842 108768 2858 108832
rect 2922 108768 2930 108832
rect 2610 108767 2930 108768
rect 5944 108832 6264 108833
rect 5944 108768 5952 108832
rect 6016 108768 6032 108832
rect 6096 108768 6112 108832
rect 6176 108768 6192 108832
rect 6256 108768 6264 108832
rect 5944 108767 6264 108768
rect 4277 108288 4597 108289
rect 4277 108224 4285 108288
rect 4349 108224 4365 108288
rect 4429 108224 4445 108288
rect 4509 108224 4525 108288
rect 4589 108224 4597 108288
rect 4277 108223 4597 108224
rect 7610 108288 7930 108289
rect 7610 108224 7618 108288
rect 7682 108224 7698 108288
rect 7762 108224 7778 108288
rect 7842 108224 7858 108288
rect 7922 108224 7930 108288
rect 7610 108223 7930 108224
rect 2610 107744 2930 107745
rect 2610 107680 2618 107744
rect 2682 107680 2698 107744
rect 2762 107680 2778 107744
rect 2842 107680 2858 107744
rect 2922 107680 2930 107744
rect 2610 107679 2930 107680
rect 5944 107744 6264 107745
rect 5944 107680 5952 107744
rect 6016 107680 6032 107744
rect 6096 107680 6112 107744
rect 6176 107680 6192 107744
rect 6256 107680 6264 107744
rect 5944 107679 6264 107680
rect 4277 107200 4597 107201
rect 4277 107136 4285 107200
rect 4349 107136 4365 107200
rect 4429 107136 4445 107200
rect 4509 107136 4525 107200
rect 4589 107136 4597 107200
rect 4277 107135 4597 107136
rect 7610 107200 7930 107201
rect 7610 107136 7618 107200
rect 7682 107136 7698 107200
rect 7762 107136 7778 107200
rect 7842 107136 7858 107200
rect 7922 107136 7930 107200
rect 7610 107135 7930 107136
rect 2610 106656 2930 106657
rect 2610 106592 2618 106656
rect 2682 106592 2698 106656
rect 2762 106592 2778 106656
rect 2842 106592 2858 106656
rect 2922 106592 2930 106656
rect 2610 106591 2930 106592
rect 5944 106656 6264 106657
rect 5944 106592 5952 106656
rect 6016 106592 6032 106656
rect 6096 106592 6112 106656
rect 6176 106592 6192 106656
rect 6256 106592 6264 106656
rect 5944 106591 6264 106592
rect 4277 106112 4597 106113
rect 4277 106048 4285 106112
rect 4349 106048 4365 106112
rect 4429 106048 4445 106112
rect 4509 106048 4525 106112
rect 4589 106048 4597 106112
rect 4277 106047 4597 106048
rect 7610 106112 7930 106113
rect 7610 106048 7618 106112
rect 7682 106048 7698 106112
rect 7762 106048 7778 106112
rect 7842 106048 7858 106112
rect 7922 106048 7930 106112
rect 7610 106047 7930 106048
rect 2610 105568 2930 105569
rect 2610 105504 2618 105568
rect 2682 105504 2698 105568
rect 2762 105504 2778 105568
rect 2842 105504 2858 105568
rect 2922 105504 2930 105568
rect 2610 105503 2930 105504
rect 5944 105568 6264 105569
rect 5944 105504 5952 105568
rect 6016 105504 6032 105568
rect 6096 105504 6112 105568
rect 6176 105504 6192 105568
rect 6256 105504 6264 105568
rect 5944 105503 6264 105504
rect 4277 105024 4597 105025
rect 4277 104960 4285 105024
rect 4349 104960 4365 105024
rect 4429 104960 4445 105024
rect 4509 104960 4525 105024
rect 4589 104960 4597 105024
rect 4277 104959 4597 104960
rect 7610 105024 7930 105025
rect 7610 104960 7618 105024
rect 7682 104960 7698 105024
rect 7762 104960 7778 105024
rect 7842 104960 7858 105024
rect 7922 104960 7930 105024
rect 7610 104959 7930 104960
rect 2610 104480 2930 104481
rect 2610 104416 2618 104480
rect 2682 104416 2698 104480
rect 2762 104416 2778 104480
rect 2842 104416 2858 104480
rect 2922 104416 2930 104480
rect 2610 104415 2930 104416
rect 5944 104480 6264 104481
rect 5944 104416 5952 104480
rect 6016 104416 6032 104480
rect 6096 104416 6112 104480
rect 6176 104416 6192 104480
rect 6256 104416 6264 104480
rect 5944 104415 6264 104416
rect 4277 103936 4597 103937
rect 4277 103872 4285 103936
rect 4349 103872 4365 103936
rect 4429 103872 4445 103936
rect 4509 103872 4525 103936
rect 4589 103872 4597 103936
rect 4277 103871 4597 103872
rect 7610 103936 7930 103937
rect 7610 103872 7618 103936
rect 7682 103872 7698 103936
rect 7762 103872 7778 103936
rect 7842 103872 7858 103936
rect 7922 103872 7930 103936
rect 7610 103871 7930 103872
rect 2610 103392 2930 103393
rect 2610 103328 2618 103392
rect 2682 103328 2698 103392
rect 2762 103328 2778 103392
rect 2842 103328 2858 103392
rect 2922 103328 2930 103392
rect 2610 103327 2930 103328
rect 5944 103392 6264 103393
rect 5944 103328 5952 103392
rect 6016 103328 6032 103392
rect 6096 103328 6112 103392
rect 6176 103328 6192 103392
rect 6256 103328 6264 103392
rect 5944 103327 6264 103328
rect 4277 102848 4597 102849
rect 4277 102784 4285 102848
rect 4349 102784 4365 102848
rect 4429 102784 4445 102848
rect 4509 102784 4525 102848
rect 4589 102784 4597 102848
rect 4277 102783 4597 102784
rect 7610 102848 7930 102849
rect 7610 102784 7618 102848
rect 7682 102784 7698 102848
rect 7762 102784 7778 102848
rect 7842 102784 7858 102848
rect 7922 102784 7930 102848
rect 7610 102783 7930 102784
rect 2610 102304 2930 102305
rect 2610 102240 2618 102304
rect 2682 102240 2698 102304
rect 2762 102240 2778 102304
rect 2842 102240 2858 102304
rect 2922 102240 2930 102304
rect 2610 102239 2930 102240
rect 5944 102304 6264 102305
rect 5944 102240 5952 102304
rect 6016 102240 6032 102304
rect 6096 102240 6112 102304
rect 6176 102240 6192 102304
rect 6256 102240 6264 102304
rect 5944 102239 6264 102240
rect 4277 101760 4597 101761
rect 4277 101696 4285 101760
rect 4349 101696 4365 101760
rect 4429 101696 4445 101760
rect 4509 101696 4525 101760
rect 4589 101696 4597 101760
rect 4277 101695 4597 101696
rect 7610 101760 7930 101761
rect 7610 101696 7618 101760
rect 7682 101696 7698 101760
rect 7762 101696 7778 101760
rect 7842 101696 7858 101760
rect 7922 101696 7930 101760
rect 7610 101695 7930 101696
rect 2610 101216 2930 101217
rect 2610 101152 2618 101216
rect 2682 101152 2698 101216
rect 2762 101152 2778 101216
rect 2842 101152 2858 101216
rect 2922 101152 2930 101216
rect 2610 101151 2930 101152
rect 5944 101216 6264 101217
rect 5944 101152 5952 101216
rect 6016 101152 6032 101216
rect 6096 101152 6112 101216
rect 6176 101152 6192 101216
rect 6256 101152 6264 101216
rect 5944 101151 6264 101152
rect 4277 100672 4597 100673
rect 4277 100608 4285 100672
rect 4349 100608 4365 100672
rect 4429 100608 4445 100672
rect 4509 100608 4525 100672
rect 4589 100608 4597 100672
rect 4277 100607 4597 100608
rect 7610 100672 7930 100673
rect 7610 100608 7618 100672
rect 7682 100608 7698 100672
rect 7762 100608 7778 100672
rect 7842 100608 7858 100672
rect 7922 100608 7930 100672
rect 7610 100607 7930 100608
rect 2610 100128 2930 100129
rect 2610 100064 2618 100128
rect 2682 100064 2698 100128
rect 2762 100064 2778 100128
rect 2842 100064 2858 100128
rect 2922 100064 2930 100128
rect 2610 100063 2930 100064
rect 5944 100128 6264 100129
rect 5944 100064 5952 100128
rect 6016 100064 6032 100128
rect 6096 100064 6112 100128
rect 6176 100064 6192 100128
rect 6256 100064 6264 100128
rect 5944 100063 6264 100064
rect 4277 99584 4597 99585
rect 4277 99520 4285 99584
rect 4349 99520 4365 99584
rect 4429 99520 4445 99584
rect 4509 99520 4525 99584
rect 4589 99520 4597 99584
rect 4277 99519 4597 99520
rect 7610 99584 7930 99585
rect 7610 99520 7618 99584
rect 7682 99520 7698 99584
rect 7762 99520 7778 99584
rect 7842 99520 7858 99584
rect 7922 99520 7930 99584
rect 7610 99519 7930 99520
rect 2610 99040 2930 99041
rect 2610 98976 2618 99040
rect 2682 98976 2698 99040
rect 2762 98976 2778 99040
rect 2842 98976 2858 99040
rect 2922 98976 2930 99040
rect 2610 98975 2930 98976
rect 5944 99040 6264 99041
rect 5944 98976 5952 99040
rect 6016 98976 6032 99040
rect 6096 98976 6112 99040
rect 6176 98976 6192 99040
rect 6256 98976 6264 99040
rect 5944 98975 6264 98976
rect 4277 98496 4597 98497
rect 4277 98432 4285 98496
rect 4349 98432 4365 98496
rect 4429 98432 4445 98496
rect 4509 98432 4525 98496
rect 4589 98432 4597 98496
rect 4277 98431 4597 98432
rect 7610 98496 7930 98497
rect 7610 98432 7618 98496
rect 7682 98432 7698 98496
rect 7762 98432 7778 98496
rect 7842 98432 7858 98496
rect 7922 98432 7930 98496
rect 7610 98431 7930 98432
rect 2610 97952 2930 97953
rect 2610 97888 2618 97952
rect 2682 97888 2698 97952
rect 2762 97888 2778 97952
rect 2842 97888 2858 97952
rect 2922 97888 2930 97952
rect 2610 97887 2930 97888
rect 5944 97952 6264 97953
rect 5944 97888 5952 97952
rect 6016 97888 6032 97952
rect 6096 97888 6112 97952
rect 6176 97888 6192 97952
rect 6256 97888 6264 97952
rect 5944 97887 6264 97888
rect 4277 97408 4597 97409
rect 4277 97344 4285 97408
rect 4349 97344 4365 97408
rect 4429 97344 4445 97408
rect 4509 97344 4525 97408
rect 4589 97344 4597 97408
rect 4277 97343 4597 97344
rect 7610 97408 7930 97409
rect 7610 97344 7618 97408
rect 7682 97344 7698 97408
rect 7762 97344 7778 97408
rect 7842 97344 7858 97408
rect 7922 97344 7930 97408
rect 7610 97343 7930 97344
rect 2610 96864 2930 96865
rect 2610 96800 2618 96864
rect 2682 96800 2698 96864
rect 2762 96800 2778 96864
rect 2842 96800 2858 96864
rect 2922 96800 2930 96864
rect 2610 96799 2930 96800
rect 5944 96864 6264 96865
rect 5944 96800 5952 96864
rect 6016 96800 6032 96864
rect 6096 96800 6112 96864
rect 6176 96800 6192 96864
rect 6256 96800 6264 96864
rect 5944 96799 6264 96800
rect 4277 96320 4597 96321
rect 4277 96256 4285 96320
rect 4349 96256 4365 96320
rect 4429 96256 4445 96320
rect 4509 96256 4525 96320
rect 4589 96256 4597 96320
rect 4277 96255 4597 96256
rect 7610 96320 7930 96321
rect 7610 96256 7618 96320
rect 7682 96256 7698 96320
rect 7762 96256 7778 96320
rect 7842 96256 7858 96320
rect 7922 96256 7930 96320
rect 7610 96255 7930 96256
rect 2610 95776 2930 95777
rect 2610 95712 2618 95776
rect 2682 95712 2698 95776
rect 2762 95712 2778 95776
rect 2842 95712 2858 95776
rect 2922 95712 2930 95776
rect 2610 95711 2930 95712
rect 5944 95776 6264 95777
rect 5944 95712 5952 95776
rect 6016 95712 6032 95776
rect 6096 95712 6112 95776
rect 6176 95712 6192 95776
rect 6256 95712 6264 95776
rect 5944 95711 6264 95712
rect 4277 95232 4597 95233
rect 4277 95168 4285 95232
rect 4349 95168 4365 95232
rect 4429 95168 4445 95232
rect 4509 95168 4525 95232
rect 4589 95168 4597 95232
rect 4277 95167 4597 95168
rect 7610 95232 7930 95233
rect 7610 95168 7618 95232
rect 7682 95168 7698 95232
rect 7762 95168 7778 95232
rect 7842 95168 7858 95232
rect 7922 95168 7930 95232
rect 7610 95167 7930 95168
rect 2610 94688 2930 94689
rect 2610 94624 2618 94688
rect 2682 94624 2698 94688
rect 2762 94624 2778 94688
rect 2842 94624 2858 94688
rect 2922 94624 2930 94688
rect 2610 94623 2930 94624
rect 5944 94688 6264 94689
rect 5944 94624 5952 94688
rect 6016 94624 6032 94688
rect 6096 94624 6112 94688
rect 6176 94624 6192 94688
rect 6256 94624 6264 94688
rect 5944 94623 6264 94624
rect 4277 94144 4597 94145
rect 4277 94080 4285 94144
rect 4349 94080 4365 94144
rect 4429 94080 4445 94144
rect 4509 94080 4525 94144
rect 4589 94080 4597 94144
rect 4277 94079 4597 94080
rect 7610 94144 7930 94145
rect 7610 94080 7618 94144
rect 7682 94080 7698 94144
rect 7762 94080 7778 94144
rect 7842 94080 7858 94144
rect 7922 94080 7930 94144
rect 7610 94079 7930 94080
rect 2610 93600 2930 93601
rect 2610 93536 2618 93600
rect 2682 93536 2698 93600
rect 2762 93536 2778 93600
rect 2842 93536 2858 93600
rect 2922 93536 2930 93600
rect 2610 93535 2930 93536
rect 5944 93600 6264 93601
rect 5944 93536 5952 93600
rect 6016 93536 6032 93600
rect 6096 93536 6112 93600
rect 6176 93536 6192 93600
rect 6256 93536 6264 93600
rect 5944 93535 6264 93536
rect 4277 93056 4597 93057
rect 4277 92992 4285 93056
rect 4349 92992 4365 93056
rect 4429 92992 4445 93056
rect 4509 92992 4525 93056
rect 4589 92992 4597 93056
rect 4277 92991 4597 92992
rect 7610 93056 7930 93057
rect 7610 92992 7618 93056
rect 7682 92992 7698 93056
rect 7762 92992 7778 93056
rect 7842 92992 7858 93056
rect 7922 92992 7930 93056
rect 7610 92991 7930 92992
rect 2610 92512 2930 92513
rect 2610 92448 2618 92512
rect 2682 92448 2698 92512
rect 2762 92448 2778 92512
rect 2842 92448 2858 92512
rect 2922 92448 2930 92512
rect 2610 92447 2930 92448
rect 5944 92512 6264 92513
rect 5944 92448 5952 92512
rect 6016 92448 6032 92512
rect 6096 92448 6112 92512
rect 6176 92448 6192 92512
rect 6256 92448 6264 92512
rect 5944 92447 6264 92448
rect 4277 91968 4597 91969
rect 4277 91904 4285 91968
rect 4349 91904 4365 91968
rect 4429 91904 4445 91968
rect 4509 91904 4525 91968
rect 4589 91904 4597 91968
rect 4277 91903 4597 91904
rect 7610 91968 7930 91969
rect 7610 91904 7618 91968
rect 7682 91904 7698 91968
rect 7762 91904 7778 91968
rect 7842 91904 7858 91968
rect 7922 91904 7930 91968
rect 7610 91903 7930 91904
rect 2610 91424 2930 91425
rect 2610 91360 2618 91424
rect 2682 91360 2698 91424
rect 2762 91360 2778 91424
rect 2842 91360 2858 91424
rect 2922 91360 2930 91424
rect 2610 91359 2930 91360
rect 5944 91424 6264 91425
rect 5944 91360 5952 91424
rect 6016 91360 6032 91424
rect 6096 91360 6112 91424
rect 6176 91360 6192 91424
rect 6256 91360 6264 91424
rect 5944 91359 6264 91360
rect 4277 90880 4597 90881
rect 4277 90816 4285 90880
rect 4349 90816 4365 90880
rect 4429 90816 4445 90880
rect 4509 90816 4525 90880
rect 4589 90816 4597 90880
rect 4277 90815 4597 90816
rect 7610 90880 7930 90881
rect 7610 90816 7618 90880
rect 7682 90816 7698 90880
rect 7762 90816 7778 90880
rect 7842 90816 7858 90880
rect 7922 90816 7930 90880
rect 7610 90815 7930 90816
rect 2610 90336 2930 90337
rect 2610 90272 2618 90336
rect 2682 90272 2698 90336
rect 2762 90272 2778 90336
rect 2842 90272 2858 90336
rect 2922 90272 2930 90336
rect 2610 90271 2930 90272
rect 5944 90336 6264 90337
rect 5944 90272 5952 90336
rect 6016 90272 6032 90336
rect 6096 90272 6112 90336
rect 6176 90272 6192 90336
rect 6256 90272 6264 90336
rect 5944 90271 6264 90272
rect 4277 89792 4597 89793
rect 4277 89728 4285 89792
rect 4349 89728 4365 89792
rect 4429 89728 4445 89792
rect 4509 89728 4525 89792
rect 4589 89728 4597 89792
rect 4277 89727 4597 89728
rect 7610 89792 7930 89793
rect 7610 89728 7618 89792
rect 7682 89728 7698 89792
rect 7762 89728 7778 89792
rect 7842 89728 7858 89792
rect 7922 89728 7930 89792
rect 7610 89727 7930 89728
rect 2610 89248 2930 89249
rect 2610 89184 2618 89248
rect 2682 89184 2698 89248
rect 2762 89184 2778 89248
rect 2842 89184 2858 89248
rect 2922 89184 2930 89248
rect 2610 89183 2930 89184
rect 5944 89248 6264 89249
rect 5944 89184 5952 89248
rect 6016 89184 6032 89248
rect 6096 89184 6112 89248
rect 6176 89184 6192 89248
rect 6256 89184 6264 89248
rect 5944 89183 6264 89184
rect 4277 88704 4597 88705
rect 4277 88640 4285 88704
rect 4349 88640 4365 88704
rect 4429 88640 4445 88704
rect 4509 88640 4525 88704
rect 4589 88640 4597 88704
rect 4277 88639 4597 88640
rect 7610 88704 7930 88705
rect 7610 88640 7618 88704
rect 7682 88640 7698 88704
rect 7762 88640 7778 88704
rect 7842 88640 7858 88704
rect 7922 88640 7930 88704
rect 7610 88639 7930 88640
rect 2610 88160 2930 88161
rect 2610 88096 2618 88160
rect 2682 88096 2698 88160
rect 2762 88096 2778 88160
rect 2842 88096 2858 88160
rect 2922 88096 2930 88160
rect 2610 88095 2930 88096
rect 5944 88160 6264 88161
rect 5944 88096 5952 88160
rect 6016 88096 6032 88160
rect 6096 88096 6112 88160
rect 6176 88096 6192 88160
rect 6256 88096 6264 88160
rect 5944 88095 6264 88096
rect 4277 87616 4597 87617
rect 4277 87552 4285 87616
rect 4349 87552 4365 87616
rect 4429 87552 4445 87616
rect 4509 87552 4525 87616
rect 4589 87552 4597 87616
rect 4277 87551 4597 87552
rect 7610 87616 7930 87617
rect 7610 87552 7618 87616
rect 7682 87552 7698 87616
rect 7762 87552 7778 87616
rect 7842 87552 7858 87616
rect 7922 87552 7930 87616
rect 7610 87551 7930 87552
rect 2610 87072 2930 87073
rect 2610 87008 2618 87072
rect 2682 87008 2698 87072
rect 2762 87008 2778 87072
rect 2842 87008 2858 87072
rect 2922 87008 2930 87072
rect 2610 87007 2930 87008
rect 5944 87072 6264 87073
rect 5944 87008 5952 87072
rect 6016 87008 6032 87072
rect 6096 87008 6112 87072
rect 6176 87008 6192 87072
rect 6256 87008 6264 87072
rect 5944 87007 6264 87008
rect 4277 86528 4597 86529
rect 4277 86464 4285 86528
rect 4349 86464 4365 86528
rect 4429 86464 4445 86528
rect 4509 86464 4525 86528
rect 4589 86464 4597 86528
rect 4277 86463 4597 86464
rect 7610 86528 7930 86529
rect 7610 86464 7618 86528
rect 7682 86464 7698 86528
rect 7762 86464 7778 86528
rect 7842 86464 7858 86528
rect 7922 86464 7930 86528
rect 7610 86463 7930 86464
rect 2610 85984 2930 85985
rect 2610 85920 2618 85984
rect 2682 85920 2698 85984
rect 2762 85920 2778 85984
rect 2842 85920 2858 85984
rect 2922 85920 2930 85984
rect 2610 85919 2930 85920
rect 5944 85984 6264 85985
rect 5944 85920 5952 85984
rect 6016 85920 6032 85984
rect 6096 85920 6112 85984
rect 6176 85920 6192 85984
rect 6256 85920 6264 85984
rect 5944 85919 6264 85920
rect 4277 85440 4597 85441
rect 4277 85376 4285 85440
rect 4349 85376 4365 85440
rect 4429 85376 4445 85440
rect 4509 85376 4525 85440
rect 4589 85376 4597 85440
rect 4277 85375 4597 85376
rect 7610 85440 7930 85441
rect 7610 85376 7618 85440
rect 7682 85376 7698 85440
rect 7762 85376 7778 85440
rect 7842 85376 7858 85440
rect 7922 85376 7930 85440
rect 7610 85375 7930 85376
rect 2610 84896 2930 84897
rect 2610 84832 2618 84896
rect 2682 84832 2698 84896
rect 2762 84832 2778 84896
rect 2842 84832 2858 84896
rect 2922 84832 2930 84896
rect 2610 84831 2930 84832
rect 5944 84896 6264 84897
rect 5944 84832 5952 84896
rect 6016 84832 6032 84896
rect 6096 84832 6112 84896
rect 6176 84832 6192 84896
rect 6256 84832 6264 84896
rect 5944 84831 6264 84832
rect 4277 84352 4597 84353
rect 4277 84288 4285 84352
rect 4349 84288 4365 84352
rect 4429 84288 4445 84352
rect 4509 84288 4525 84352
rect 4589 84288 4597 84352
rect 4277 84287 4597 84288
rect 7610 84352 7930 84353
rect 7610 84288 7618 84352
rect 7682 84288 7698 84352
rect 7762 84288 7778 84352
rect 7842 84288 7858 84352
rect 7922 84288 7930 84352
rect 7610 84287 7930 84288
rect 2610 83808 2930 83809
rect 2610 83744 2618 83808
rect 2682 83744 2698 83808
rect 2762 83744 2778 83808
rect 2842 83744 2858 83808
rect 2922 83744 2930 83808
rect 2610 83743 2930 83744
rect 5944 83808 6264 83809
rect 5944 83744 5952 83808
rect 6016 83744 6032 83808
rect 6096 83744 6112 83808
rect 6176 83744 6192 83808
rect 6256 83744 6264 83808
rect 5944 83743 6264 83744
rect 8201 83738 8267 83741
rect 8201 83736 9690 83738
rect 8201 83680 8206 83736
rect 8262 83680 9690 83736
rect 8201 83678 9690 83680
rect 8201 83675 8267 83678
rect 4277 83264 4597 83265
rect 4277 83200 4285 83264
rect 4349 83200 4365 83264
rect 4429 83200 4445 83264
rect 4509 83200 4525 83264
rect 4589 83200 4597 83264
rect 4277 83199 4597 83200
rect 7610 83264 7930 83265
rect 7610 83200 7618 83264
rect 7682 83200 7698 83264
rect 7762 83200 7778 83264
rect 7842 83200 7858 83264
rect 7922 83200 7930 83264
rect 9630 83224 9690 83678
rect 7610 83199 7930 83200
rect 9520 83104 10000 83224
rect 2610 82720 2930 82721
rect 2610 82656 2618 82720
rect 2682 82656 2698 82720
rect 2762 82656 2778 82720
rect 2842 82656 2858 82720
rect 2922 82656 2930 82720
rect 2610 82655 2930 82656
rect 5944 82720 6264 82721
rect 5944 82656 5952 82720
rect 6016 82656 6032 82720
rect 6096 82656 6112 82720
rect 6176 82656 6192 82720
rect 6256 82656 6264 82720
rect 5944 82655 6264 82656
rect 4277 82176 4597 82177
rect 4277 82112 4285 82176
rect 4349 82112 4365 82176
rect 4429 82112 4445 82176
rect 4509 82112 4525 82176
rect 4589 82112 4597 82176
rect 4277 82111 4597 82112
rect 7610 82176 7930 82177
rect 7610 82112 7618 82176
rect 7682 82112 7698 82176
rect 7762 82112 7778 82176
rect 7842 82112 7858 82176
rect 7922 82112 7930 82176
rect 7610 82111 7930 82112
rect 2610 81632 2930 81633
rect 2610 81568 2618 81632
rect 2682 81568 2698 81632
rect 2762 81568 2778 81632
rect 2842 81568 2858 81632
rect 2922 81568 2930 81632
rect 2610 81567 2930 81568
rect 5944 81632 6264 81633
rect 5944 81568 5952 81632
rect 6016 81568 6032 81632
rect 6096 81568 6112 81632
rect 6176 81568 6192 81632
rect 6256 81568 6264 81632
rect 5944 81567 6264 81568
rect 4277 81088 4597 81089
rect 4277 81024 4285 81088
rect 4349 81024 4365 81088
rect 4429 81024 4445 81088
rect 4509 81024 4525 81088
rect 4589 81024 4597 81088
rect 4277 81023 4597 81024
rect 7610 81088 7930 81089
rect 7610 81024 7618 81088
rect 7682 81024 7698 81088
rect 7762 81024 7778 81088
rect 7842 81024 7858 81088
rect 7922 81024 7930 81088
rect 7610 81023 7930 81024
rect 2610 80544 2930 80545
rect 2610 80480 2618 80544
rect 2682 80480 2698 80544
rect 2762 80480 2778 80544
rect 2842 80480 2858 80544
rect 2922 80480 2930 80544
rect 2610 80479 2930 80480
rect 5944 80544 6264 80545
rect 5944 80480 5952 80544
rect 6016 80480 6032 80544
rect 6096 80480 6112 80544
rect 6176 80480 6192 80544
rect 6256 80480 6264 80544
rect 5944 80479 6264 80480
rect 4277 80000 4597 80001
rect 4277 79936 4285 80000
rect 4349 79936 4365 80000
rect 4429 79936 4445 80000
rect 4509 79936 4525 80000
rect 4589 79936 4597 80000
rect 4277 79935 4597 79936
rect 7610 80000 7930 80001
rect 7610 79936 7618 80000
rect 7682 79936 7698 80000
rect 7762 79936 7778 80000
rect 7842 79936 7858 80000
rect 7922 79936 7930 80000
rect 7610 79935 7930 79936
rect 2610 79456 2930 79457
rect 2610 79392 2618 79456
rect 2682 79392 2698 79456
rect 2762 79392 2778 79456
rect 2842 79392 2858 79456
rect 2922 79392 2930 79456
rect 2610 79391 2930 79392
rect 5944 79456 6264 79457
rect 5944 79392 5952 79456
rect 6016 79392 6032 79456
rect 6096 79392 6112 79456
rect 6176 79392 6192 79456
rect 6256 79392 6264 79456
rect 5944 79391 6264 79392
rect 4277 78912 4597 78913
rect 4277 78848 4285 78912
rect 4349 78848 4365 78912
rect 4429 78848 4445 78912
rect 4509 78848 4525 78912
rect 4589 78848 4597 78912
rect 4277 78847 4597 78848
rect 7610 78912 7930 78913
rect 7610 78848 7618 78912
rect 7682 78848 7698 78912
rect 7762 78848 7778 78912
rect 7842 78848 7858 78912
rect 7922 78848 7930 78912
rect 7610 78847 7930 78848
rect 2610 78368 2930 78369
rect 2610 78304 2618 78368
rect 2682 78304 2698 78368
rect 2762 78304 2778 78368
rect 2842 78304 2858 78368
rect 2922 78304 2930 78368
rect 2610 78303 2930 78304
rect 5944 78368 6264 78369
rect 5944 78304 5952 78368
rect 6016 78304 6032 78368
rect 6096 78304 6112 78368
rect 6176 78304 6192 78368
rect 6256 78304 6264 78368
rect 5944 78303 6264 78304
rect 4277 77824 4597 77825
rect 4277 77760 4285 77824
rect 4349 77760 4365 77824
rect 4429 77760 4445 77824
rect 4509 77760 4525 77824
rect 4589 77760 4597 77824
rect 4277 77759 4597 77760
rect 7610 77824 7930 77825
rect 7610 77760 7618 77824
rect 7682 77760 7698 77824
rect 7762 77760 7778 77824
rect 7842 77760 7858 77824
rect 7922 77760 7930 77824
rect 7610 77759 7930 77760
rect 2610 77280 2930 77281
rect 2610 77216 2618 77280
rect 2682 77216 2698 77280
rect 2762 77216 2778 77280
rect 2842 77216 2858 77280
rect 2922 77216 2930 77280
rect 2610 77215 2930 77216
rect 5944 77280 6264 77281
rect 5944 77216 5952 77280
rect 6016 77216 6032 77280
rect 6096 77216 6112 77280
rect 6176 77216 6192 77280
rect 6256 77216 6264 77280
rect 5944 77215 6264 77216
rect 4277 76736 4597 76737
rect 4277 76672 4285 76736
rect 4349 76672 4365 76736
rect 4429 76672 4445 76736
rect 4509 76672 4525 76736
rect 4589 76672 4597 76736
rect 4277 76671 4597 76672
rect 7610 76736 7930 76737
rect 7610 76672 7618 76736
rect 7682 76672 7698 76736
rect 7762 76672 7778 76736
rect 7842 76672 7858 76736
rect 7922 76672 7930 76736
rect 7610 76671 7930 76672
rect 2610 76192 2930 76193
rect 2610 76128 2618 76192
rect 2682 76128 2698 76192
rect 2762 76128 2778 76192
rect 2842 76128 2858 76192
rect 2922 76128 2930 76192
rect 2610 76127 2930 76128
rect 5944 76192 6264 76193
rect 5944 76128 5952 76192
rect 6016 76128 6032 76192
rect 6096 76128 6112 76192
rect 6176 76128 6192 76192
rect 6256 76128 6264 76192
rect 5944 76127 6264 76128
rect 4277 75648 4597 75649
rect 4277 75584 4285 75648
rect 4349 75584 4365 75648
rect 4429 75584 4445 75648
rect 4509 75584 4525 75648
rect 4589 75584 4597 75648
rect 4277 75583 4597 75584
rect 7610 75648 7930 75649
rect 7610 75584 7618 75648
rect 7682 75584 7698 75648
rect 7762 75584 7778 75648
rect 7842 75584 7858 75648
rect 7922 75584 7930 75648
rect 7610 75583 7930 75584
rect 2610 75104 2930 75105
rect 2610 75040 2618 75104
rect 2682 75040 2698 75104
rect 2762 75040 2778 75104
rect 2842 75040 2858 75104
rect 2922 75040 2930 75104
rect 2610 75039 2930 75040
rect 5944 75104 6264 75105
rect 5944 75040 5952 75104
rect 6016 75040 6032 75104
rect 6096 75040 6112 75104
rect 6176 75040 6192 75104
rect 6256 75040 6264 75104
rect 5944 75039 6264 75040
rect 4277 74560 4597 74561
rect 4277 74496 4285 74560
rect 4349 74496 4365 74560
rect 4429 74496 4445 74560
rect 4509 74496 4525 74560
rect 4589 74496 4597 74560
rect 4277 74495 4597 74496
rect 7610 74560 7930 74561
rect 7610 74496 7618 74560
rect 7682 74496 7698 74560
rect 7762 74496 7778 74560
rect 7842 74496 7858 74560
rect 7922 74496 7930 74560
rect 7610 74495 7930 74496
rect 2610 74016 2930 74017
rect 2610 73952 2618 74016
rect 2682 73952 2698 74016
rect 2762 73952 2778 74016
rect 2842 73952 2858 74016
rect 2922 73952 2930 74016
rect 2610 73951 2930 73952
rect 5944 74016 6264 74017
rect 5944 73952 5952 74016
rect 6016 73952 6032 74016
rect 6096 73952 6112 74016
rect 6176 73952 6192 74016
rect 6256 73952 6264 74016
rect 5944 73951 6264 73952
rect 4277 73472 4597 73473
rect 4277 73408 4285 73472
rect 4349 73408 4365 73472
rect 4429 73408 4445 73472
rect 4509 73408 4525 73472
rect 4589 73408 4597 73472
rect 4277 73407 4597 73408
rect 7610 73472 7930 73473
rect 7610 73408 7618 73472
rect 7682 73408 7698 73472
rect 7762 73408 7778 73472
rect 7842 73408 7858 73472
rect 7922 73408 7930 73472
rect 7610 73407 7930 73408
rect 2610 72928 2930 72929
rect 2610 72864 2618 72928
rect 2682 72864 2698 72928
rect 2762 72864 2778 72928
rect 2842 72864 2858 72928
rect 2922 72864 2930 72928
rect 2610 72863 2930 72864
rect 5944 72928 6264 72929
rect 5944 72864 5952 72928
rect 6016 72864 6032 72928
rect 6096 72864 6112 72928
rect 6176 72864 6192 72928
rect 6256 72864 6264 72928
rect 5944 72863 6264 72864
rect 4277 72384 4597 72385
rect 4277 72320 4285 72384
rect 4349 72320 4365 72384
rect 4429 72320 4445 72384
rect 4509 72320 4525 72384
rect 4589 72320 4597 72384
rect 4277 72319 4597 72320
rect 7610 72384 7930 72385
rect 7610 72320 7618 72384
rect 7682 72320 7698 72384
rect 7762 72320 7778 72384
rect 7842 72320 7858 72384
rect 7922 72320 7930 72384
rect 7610 72319 7930 72320
rect 2610 71840 2930 71841
rect 2610 71776 2618 71840
rect 2682 71776 2698 71840
rect 2762 71776 2778 71840
rect 2842 71776 2858 71840
rect 2922 71776 2930 71840
rect 2610 71775 2930 71776
rect 5944 71840 6264 71841
rect 5944 71776 5952 71840
rect 6016 71776 6032 71840
rect 6096 71776 6112 71840
rect 6176 71776 6192 71840
rect 6256 71776 6264 71840
rect 5944 71775 6264 71776
rect 4277 71296 4597 71297
rect 0 71224 480 71256
rect 4277 71232 4285 71296
rect 4349 71232 4365 71296
rect 4429 71232 4445 71296
rect 4509 71232 4525 71296
rect 4589 71232 4597 71296
rect 4277 71231 4597 71232
rect 7610 71296 7930 71297
rect 7610 71232 7618 71296
rect 7682 71232 7698 71296
rect 7762 71232 7778 71296
rect 7842 71232 7858 71296
rect 7922 71232 7930 71296
rect 7610 71231 7930 71232
rect 0 71168 110 71224
rect 166 71168 480 71224
rect 0 71136 480 71168
rect 2610 70752 2930 70753
rect 2610 70688 2618 70752
rect 2682 70688 2698 70752
rect 2762 70688 2778 70752
rect 2842 70688 2858 70752
rect 2922 70688 2930 70752
rect 2610 70687 2930 70688
rect 5944 70752 6264 70753
rect 5944 70688 5952 70752
rect 6016 70688 6032 70752
rect 6096 70688 6112 70752
rect 6176 70688 6192 70752
rect 6256 70688 6264 70752
rect 5944 70687 6264 70688
rect 4277 70208 4597 70209
rect 4277 70144 4285 70208
rect 4349 70144 4365 70208
rect 4429 70144 4445 70208
rect 4509 70144 4525 70208
rect 4589 70144 4597 70208
rect 4277 70143 4597 70144
rect 7610 70208 7930 70209
rect 7610 70144 7618 70208
rect 7682 70144 7698 70208
rect 7762 70144 7778 70208
rect 7842 70144 7858 70208
rect 7922 70144 7930 70208
rect 7610 70143 7930 70144
rect 2610 69664 2930 69665
rect 2610 69600 2618 69664
rect 2682 69600 2698 69664
rect 2762 69600 2778 69664
rect 2842 69600 2858 69664
rect 2922 69600 2930 69664
rect 2610 69599 2930 69600
rect 5944 69664 6264 69665
rect 5944 69600 5952 69664
rect 6016 69600 6032 69664
rect 6096 69600 6112 69664
rect 6176 69600 6192 69664
rect 6256 69600 6264 69664
rect 5944 69599 6264 69600
rect 4277 69120 4597 69121
rect 4277 69056 4285 69120
rect 4349 69056 4365 69120
rect 4429 69056 4445 69120
rect 4509 69056 4525 69120
rect 4589 69056 4597 69120
rect 4277 69055 4597 69056
rect 7610 69120 7930 69121
rect 7610 69056 7618 69120
rect 7682 69056 7698 69120
rect 7762 69056 7778 69120
rect 7842 69056 7858 69120
rect 7922 69056 7930 69120
rect 7610 69055 7930 69056
rect 2610 68576 2930 68577
rect 2610 68512 2618 68576
rect 2682 68512 2698 68576
rect 2762 68512 2778 68576
rect 2842 68512 2858 68576
rect 2922 68512 2930 68576
rect 2610 68511 2930 68512
rect 5944 68576 6264 68577
rect 5944 68512 5952 68576
rect 6016 68512 6032 68576
rect 6096 68512 6112 68576
rect 6176 68512 6192 68576
rect 6256 68512 6264 68576
rect 5944 68511 6264 68512
rect 4277 68032 4597 68033
rect 4277 67968 4285 68032
rect 4349 67968 4365 68032
rect 4429 67968 4445 68032
rect 4509 67968 4525 68032
rect 4589 67968 4597 68032
rect 4277 67967 4597 67968
rect 7610 68032 7930 68033
rect 7610 67968 7618 68032
rect 7682 67968 7698 68032
rect 7762 67968 7778 68032
rect 7842 67968 7858 68032
rect 7922 67968 7930 68032
rect 7610 67967 7930 67968
rect 2610 67488 2930 67489
rect 2610 67424 2618 67488
rect 2682 67424 2698 67488
rect 2762 67424 2778 67488
rect 2842 67424 2858 67488
rect 2922 67424 2930 67488
rect 2610 67423 2930 67424
rect 5944 67488 6264 67489
rect 5944 67424 5952 67488
rect 6016 67424 6032 67488
rect 6096 67424 6112 67488
rect 6176 67424 6192 67488
rect 6256 67424 6264 67488
rect 5944 67423 6264 67424
rect 4277 66944 4597 66945
rect 4277 66880 4285 66944
rect 4349 66880 4365 66944
rect 4429 66880 4445 66944
rect 4509 66880 4525 66944
rect 4589 66880 4597 66944
rect 4277 66879 4597 66880
rect 7610 66944 7930 66945
rect 7610 66880 7618 66944
rect 7682 66880 7698 66944
rect 7762 66880 7778 66944
rect 7842 66880 7858 66944
rect 7922 66880 7930 66944
rect 7610 66879 7930 66880
rect 2610 66400 2930 66401
rect 2610 66336 2618 66400
rect 2682 66336 2698 66400
rect 2762 66336 2778 66400
rect 2842 66336 2858 66400
rect 2922 66336 2930 66400
rect 2610 66335 2930 66336
rect 5944 66400 6264 66401
rect 5944 66336 5952 66400
rect 6016 66336 6032 66400
rect 6096 66336 6112 66400
rect 6176 66336 6192 66400
rect 6256 66336 6264 66400
rect 5944 66335 6264 66336
rect 4277 65856 4597 65857
rect 4277 65792 4285 65856
rect 4349 65792 4365 65856
rect 4429 65792 4445 65856
rect 4509 65792 4525 65856
rect 4589 65792 4597 65856
rect 4277 65791 4597 65792
rect 7610 65856 7930 65857
rect 7610 65792 7618 65856
rect 7682 65792 7698 65856
rect 7762 65792 7778 65856
rect 7842 65792 7858 65856
rect 7922 65792 7930 65856
rect 7610 65791 7930 65792
rect 2610 65312 2930 65313
rect 2610 65248 2618 65312
rect 2682 65248 2698 65312
rect 2762 65248 2778 65312
rect 2842 65248 2858 65312
rect 2922 65248 2930 65312
rect 2610 65247 2930 65248
rect 5944 65312 6264 65313
rect 5944 65248 5952 65312
rect 6016 65248 6032 65312
rect 6096 65248 6112 65312
rect 6176 65248 6192 65312
rect 6256 65248 6264 65312
rect 5944 65247 6264 65248
rect 4277 64768 4597 64769
rect 4277 64704 4285 64768
rect 4349 64704 4365 64768
rect 4429 64704 4445 64768
rect 4509 64704 4525 64768
rect 4589 64704 4597 64768
rect 4277 64703 4597 64704
rect 7610 64768 7930 64769
rect 7610 64704 7618 64768
rect 7682 64704 7698 64768
rect 7762 64704 7778 64768
rect 7842 64704 7858 64768
rect 7922 64704 7930 64768
rect 7610 64703 7930 64704
rect 2610 64224 2930 64225
rect 2610 64160 2618 64224
rect 2682 64160 2698 64224
rect 2762 64160 2778 64224
rect 2842 64160 2858 64224
rect 2922 64160 2930 64224
rect 2610 64159 2930 64160
rect 5944 64224 6264 64225
rect 5944 64160 5952 64224
rect 6016 64160 6032 64224
rect 6096 64160 6112 64224
rect 6176 64160 6192 64224
rect 6256 64160 6264 64224
rect 5944 64159 6264 64160
rect 4277 63680 4597 63681
rect 4277 63616 4285 63680
rect 4349 63616 4365 63680
rect 4429 63616 4445 63680
rect 4509 63616 4525 63680
rect 4589 63616 4597 63680
rect 4277 63615 4597 63616
rect 7610 63680 7930 63681
rect 7610 63616 7618 63680
rect 7682 63616 7698 63680
rect 7762 63616 7778 63680
rect 7842 63616 7858 63680
rect 7922 63616 7930 63680
rect 7610 63615 7930 63616
rect 2610 63136 2930 63137
rect 2610 63072 2618 63136
rect 2682 63072 2698 63136
rect 2762 63072 2778 63136
rect 2842 63072 2858 63136
rect 2922 63072 2930 63136
rect 2610 63071 2930 63072
rect 5944 63136 6264 63137
rect 5944 63072 5952 63136
rect 6016 63072 6032 63136
rect 6096 63072 6112 63136
rect 6176 63072 6192 63136
rect 6256 63072 6264 63136
rect 5944 63071 6264 63072
rect 4277 62592 4597 62593
rect 4277 62528 4285 62592
rect 4349 62528 4365 62592
rect 4429 62528 4445 62592
rect 4509 62528 4525 62592
rect 4589 62528 4597 62592
rect 4277 62527 4597 62528
rect 7610 62592 7930 62593
rect 7610 62528 7618 62592
rect 7682 62528 7698 62592
rect 7762 62528 7778 62592
rect 7842 62528 7858 62592
rect 7922 62528 7930 62592
rect 7610 62527 7930 62528
rect 2610 62048 2930 62049
rect 2610 61984 2618 62048
rect 2682 61984 2698 62048
rect 2762 61984 2778 62048
rect 2842 61984 2858 62048
rect 2922 61984 2930 62048
rect 2610 61983 2930 61984
rect 5944 62048 6264 62049
rect 5944 61984 5952 62048
rect 6016 61984 6032 62048
rect 6096 61984 6112 62048
rect 6176 61984 6192 62048
rect 6256 61984 6264 62048
rect 5944 61983 6264 61984
rect 4277 61504 4597 61505
rect 4277 61440 4285 61504
rect 4349 61440 4365 61504
rect 4429 61440 4445 61504
rect 4509 61440 4525 61504
rect 4589 61440 4597 61504
rect 4277 61439 4597 61440
rect 7610 61504 7930 61505
rect 7610 61440 7618 61504
rect 7682 61440 7698 61504
rect 7762 61440 7778 61504
rect 7842 61440 7858 61504
rect 7922 61440 7930 61504
rect 7610 61439 7930 61440
rect 2610 60960 2930 60961
rect 2610 60896 2618 60960
rect 2682 60896 2698 60960
rect 2762 60896 2778 60960
rect 2842 60896 2858 60960
rect 2922 60896 2930 60960
rect 2610 60895 2930 60896
rect 5944 60960 6264 60961
rect 5944 60896 5952 60960
rect 6016 60896 6032 60960
rect 6096 60896 6112 60960
rect 6176 60896 6192 60960
rect 6256 60896 6264 60960
rect 5944 60895 6264 60896
rect 4277 60416 4597 60417
rect 4277 60352 4285 60416
rect 4349 60352 4365 60416
rect 4429 60352 4445 60416
rect 4509 60352 4525 60416
rect 4589 60352 4597 60416
rect 4277 60351 4597 60352
rect 7610 60416 7930 60417
rect 7610 60352 7618 60416
rect 7682 60352 7698 60416
rect 7762 60352 7778 60416
rect 7842 60352 7858 60416
rect 7922 60352 7930 60416
rect 7610 60351 7930 60352
rect 2610 59872 2930 59873
rect 2610 59808 2618 59872
rect 2682 59808 2698 59872
rect 2762 59808 2778 59872
rect 2842 59808 2858 59872
rect 2922 59808 2930 59872
rect 2610 59807 2930 59808
rect 5944 59872 6264 59873
rect 5944 59808 5952 59872
rect 6016 59808 6032 59872
rect 6096 59808 6112 59872
rect 6176 59808 6192 59872
rect 6256 59808 6264 59872
rect 5944 59807 6264 59808
rect 4277 59328 4597 59329
rect 4277 59264 4285 59328
rect 4349 59264 4365 59328
rect 4429 59264 4445 59328
rect 4509 59264 4525 59328
rect 4589 59264 4597 59328
rect 4277 59263 4597 59264
rect 7610 59328 7930 59329
rect 7610 59264 7618 59328
rect 7682 59264 7698 59328
rect 7762 59264 7778 59328
rect 7842 59264 7858 59328
rect 7922 59264 7930 59328
rect 7610 59263 7930 59264
rect 2610 58784 2930 58785
rect 2610 58720 2618 58784
rect 2682 58720 2698 58784
rect 2762 58720 2778 58784
rect 2842 58720 2858 58784
rect 2922 58720 2930 58784
rect 2610 58719 2930 58720
rect 5944 58784 6264 58785
rect 5944 58720 5952 58784
rect 6016 58720 6032 58784
rect 6096 58720 6112 58784
rect 6176 58720 6192 58784
rect 6256 58720 6264 58784
rect 5944 58719 6264 58720
rect 4277 58240 4597 58241
rect 4277 58176 4285 58240
rect 4349 58176 4365 58240
rect 4429 58176 4445 58240
rect 4509 58176 4525 58240
rect 4589 58176 4597 58240
rect 4277 58175 4597 58176
rect 7610 58240 7930 58241
rect 7610 58176 7618 58240
rect 7682 58176 7698 58240
rect 7762 58176 7778 58240
rect 7842 58176 7858 58240
rect 7922 58176 7930 58240
rect 7610 58175 7930 58176
rect 2610 57696 2930 57697
rect 2610 57632 2618 57696
rect 2682 57632 2698 57696
rect 2762 57632 2778 57696
rect 2842 57632 2858 57696
rect 2922 57632 2930 57696
rect 2610 57631 2930 57632
rect 5944 57696 6264 57697
rect 5944 57632 5952 57696
rect 6016 57632 6032 57696
rect 6096 57632 6112 57696
rect 6176 57632 6192 57696
rect 6256 57632 6264 57696
rect 5944 57631 6264 57632
rect 4277 57152 4597 57153
rect 4277 57088 4285 57152
rect 4349 57088 4365 57152
rect 4429 57088 4445 57152
rect 4509 57088 4525 57152
rect 4589 57088 4597 57152
rect 4277 57087 4597 57088
rect 7610 57152 7930 57153
rect 7610 57088 7618 57152
rect 7682 57088 7698 57152
rect 7762 57088 7778 57152
rect 7842 57088 7858 57152
rect 7922 57088 7930 57152
rect 7610 57087 7930 57088
rect 2610 56608 2930 56609
rect 2610 56544 2618 56608
rect 2682 56544 2698 56608
rect 2762 56544 2778 56608
rect 2842 56544 2858 56608
rect 2922 56544 2930 56608
rect 2610 56543 2930 56544
rect 5944 56608 6264 56609
rect 5944 56544 5952 56608
rect 6016 56544 6032 56608
rect 6096 56544 6112 56608
rect 6176 56544 6192 56608
rect 6256 56544 6264 56608
rect 5944 56543 6264 56544
rect 4277 56064 4597 56065
rect 4277 56000 4285 56064
rect 4349 56000 4365 56064
rect 4429 56000 4445 56064
rect 4509 56000 4525 56064
rect 4589 56000 4597 56064
rect 4277 55999 4597 56000
rect 7610 56064 7930 56065
rect 7610 56000 7618 56064
rect 7682 56000 7698 56064
rect 7762 56000 7778 56064
rect 7842 56000 7858 56064
rect 7922 56000 7930 56064
rect 7610 55999 7930 56000
rect 2610 55520 2930 55521
rect 2610 55456 2618 55520
rect 2682 55456 2698 55520
rect 2762 55456 2778 55520
rect 2842 55456 2858 55520
rect 2922 55456 2930 55520
rect 2610 55455 2930 55456
rect 5944 55520 6264 55521
rect 5944 55456 5952 55520
rect 6016 55456 6032 55520
rect 6096 55456 6112 55520
rect 6176 55456 6192 55520
rect 6256 55456 6264 55520
rect 5944 55455 6264 55456
rect 4277 54976 4597 54977
rect 4277 54912 4285 54976
rect 4349 54912 4365 54976
rect 4429 54912 4445 54976
rect 4509 54912 4525 54976
rect 4589 54912 4597 54976
rect 4277 54911 4597 54912
rect 7610 54976 7930 54977
rect 7610 54912 7618 54976
rect 7682 54912 7698 54976
rect 7762 54912 7778 54976
rect 7842 54912 7858 54976
rect 7922 54912 7930 54976
rect 7610 54911 7930 54912
rect 2610 54432 2930 54433
rect 2610 54368 2618 54432
rect 2682 54368 2698 54432
rect 2762 54368 2778 54432
rect 2842 54368 2858 54432
rect 2922 54368 2930 54432
rect 2610 54367 2930 54368
rect 5944 54432 6264 54433
rect 5944 54368 5952 54432
rect 6016 54368 6032 54432
rect 6096 54368 6112 54432
rect 6176 54368 6192 54432
rect 6256 54368 6264 54432
rect 5944 54367 6264 54368
rect 4277 53888 4597 53889
rect 4277 53824 4285 53888
rect 4349 53824 4365 53888
rect 4429 53824 4445 53888
rect 4509 53824 4525 53888
rect 4589 53824 4597 53888
rect 4277 53823 4597 53824
rect 7610 53888 7930 53889
rect 7610 53824 7618 53888
rect 7682 53824 7698 53888
rect 7762 53824 7778 53888
rect 7842 53824 7858 53888
rect 7922 53824 7930 53888
rect 7610 53823 7930 53824
rect 2610 53344 2930 53345
rect 2610 53280 2618 53344
rect 2682 53280 2698 53344
rect 2762 53280 2778 53344
rect 2842 53280 2858 53344
rect 2922 53280 2930 53344
rect 2610 53279 2930 53280
rect 5944 53344 6264 53345
rect 5944 53280 5952 53344
rect 6016 53280 6032 53344
rect 6096 53280 6112 53344
rect 6176 53280 6192 53344
rect 6256 53280 6264 53344
rect 5944 53279 6264 53280
rect 4277 52800 4597 52801
rect 4277 52736 4285 52800
rect 4349 52736 4365 52800
rect 4429 52736 4445 52800
rect 4509 52736 4525 52800
rect 4589 52736 4597 52800
rect 4277 52735 4597 52736
rect 7610 52800 7930 52801
rect 7610 52736 7618 52800
rect 7682 52736 7698 52800
rect 7762 52736 7778 52800
rect 7842 52736 7858 52800
rect 7922 52736 7930 52800
rect 7610 52735 7930 52736
rect 2610 52256 2930 52257
rect 2610 52192 2618 52256
rect 2682 52192 2698 52256
rect 2762 52192 2778 52256
rect 2842 52192 2858 52256
rect 2922 52192 2930 52256
rect 2610 52191 2930 52192
rect 5944 52256 6264 52257
rect 5944 52192 5952 52256
rect 6016 52192 6032 52256
rect 6096 52192 6112 52256
rect 6176 52192 6192 52256
rect 6256 52192 6264 52256
rect 5944 52191 6264 52192
rect 4277 51712 4597 51713
rect 4277 51648 4285 51712
rect 4349 51648 4365 51712
rect 4429 51648 4445 51712
rect 4509 51648 4525 51712
rect 4589 51648 4597 51712
rect 4277 51647 4597 51648
rect 7610 51712 7930 51713
rect 7610 51648 7618 51712
rect 7682 51648 7698 51712
rect 7762 51648 7778 51712
rect 7842 51648 7858 51712
rect 7922 51648 7930 51712
rect 7610 51647 7930 51648
rect 2610 51168 2930 51169
rect 2610 51104 2618 51168
rect 2682 51104 2698 51168
rect 2762 51104 2778 51168
rect 2842 51104 2858 51168
rect 2922 51104 2930 51168
rect 2610 51103 2930 51104
rect 5944 51168 6264 51169
rect 5944 51104 5952 51168
rect 6016 51104 6032 51168
rect 6096 51104 6112 51168
rect 6176 51104 6192 51168
rect 6256 51104 6264 51168
rect 5944 51103 6264 51104
rect 4277 50624 4597 50625
rect 4277 50560 4285 50624
rect 4349 50560 4365 50624
rect 4429 50560 4445 50624
rect 4509 50560 4525 50624
rect 4589 50560 4597 50624
rect 4277 50559 4597 50560
rect 7610 50624 7930 50625
rect 7610 50560 7618 50624
rect 7682 50560 7698 50624
rect 7762 50560 7778 50624
rect 7842 50560 7858 50624
rect 7922 50560 7930 50624
rect 7610 50559 7930 50560
rect 6821 50418 6887 50421
rect 6821 50416 9690 50418
rect 6821 50360 6826 50416
rect 6882 50360 9690 50416
rect 6821 50358 9690 50360
rect 6821 50355 6887 50358
rect 2610 50080 2930 50081
rect 2610 50016 2618 50080
rect 2682 50016 2698 50080
rect 2762 50016 2778 50080
rect 2842 50016 2858 50080
rect 2922 50016 2930 50080
rect 2610 50015 2930 50016
rect 5944 50080 6264 50081
rect 5944 50016 5952 50080
rect 6016 50016 6032 50080
rect 6096 50016 6112 50080
rect 6176 50016 6192 50080
rect 6256 50016 6264 50080
rect 5944 50015 6264 50016
rect 9630 49904 9690 50358
rect 9520 49784 10000 49904
rect 4277 49536 4597 49537
rect 4277 49472 4285 49536
rect 4349 49472 4365 49536
rect 4429 49472 4445 49536
rect 4509 49472 4525 49536
rect 4589 49472 4597 49536
rect 4277 49471 4597 49472
rect 7610 49536 7930 49537
rect 7610 49472 7618 49536
rect 7682 49472 7698 49536
rect 7762 49472 7778 49536
rect 7842 49472 7858 49536
rect 7922 49472 7930 49536
rect 7610 49471 7930 49472
rect 2610 48992 2930 48993
rect 2610 48928 2618 48992
rect 2682 48928 2698 48992
rect 2762 48928 2778 48992
rect 2842 48928 2858 48992
rect 2922 48928 2930 48992
rect 2610 48927 2930 48928
rect 5944 48992 6264 48993
rect 5944 48928 5952 48992
rect 6016 48928 6032 48992
rect 6096 48928 6112 48992
rect 6176 48928 6192 48992
rect 6256 48928 6264 48992
rect 5944 48927 6264 48928
rect 4277 48448 4597 48449
rect 4277 48384 4285 48448
rect 4349 48384 4365 48448
rect 4429 48384 4445 48448
rect 4509 48384 4525 48448
rect 4589 48384 4597 48448
rect 4277 48383 4597 48384
rect 7610 48448 7930 48449
rect 7610 48384 7618 48448
rect 7682 48384 7698 48448
rect 7762 48384 7778 48448
rect 7842 48384 7858 48448
rect 7922 48384 7930 48448
rect 7610 48383 7930 48384
rect 2610 47904 2930 47905
rect 2610 47840 2618 47904
rect 2682 47840 2698 47904
rect 2762 47840 2778 47904
rect 2842 47840 2858 47904
rect 2922 47840 2930 47904
rect 2610 47839 2930 47840
rect 5944 47904 6264 47905
rect 5944 47840 5952 47904
rect 6016 47840 6032 47904
rect 6096 47840 6112 47904
rect 6176 47840 6192 47904
rect 6256 47840 6264 47904
rect 5944 47839 6264 47840
rect 4277 47360 4597 47361
rect 4277 47296 4285 47360
rect 4349 47296 4365 47360
rect 4429 47296 4445 47360
rect 4509 47296 4525 47360
rect 4589 47296 4597 47360
rect 4277 47295 4597 47296
rect 7610 47360 7930 47361
rect 7610 47296 7618 47360
rect 7682 47296 7698 47360
rect 7762 47296 7778 47360
rect 7842 47296 7858 47360
rect 7922 47296 7930 47360
rect 7610 47295 7930 47296
rect 2610 46816 2930 46817
rect 2610 46752 2618 46816
rect 2682 46752 2698 46816
rect 2762 46752 2778 46816
rect 2842 46752 2858 46816
rect 2922 46752 2930 46816
rect 2610 46751 2930 46752
rect 5944 46816 6264 46817
rect 5944 46752 5952 46816
rect 6016 46752 6032 46816
rect 6096 46752 6112 46816
rect 6176 46752 6192 46816
rect 6256 46752 6264 46816
rect 5944 46751 6264 46752
rect 4277 46272 4597 46273
rect 4277 46208 4285 46272
rect 4349 46208 4365 46272
rect 4429 46208 4445 46272
rect 4509 46208 4525 46272
rect 4589 46208 4597 46272
rect 4277 46207 4597 46208
rect 7610 46272 7930 46273
rect 7610 46208 7618 46272
rect 7682 46208 7698 46272
rect 7762 46208 7778 46272
rect 7842 46208 7858 46272
rect 7922 46208 7930 46272
rect 7610 46207 7930 46208
rect 2610 45728 2930 45729
rect 2610 45664 2618 45728
rect 2682 45664 2698 45728
rect 2762 45664 2778 45728
rect 2842 45664 2858 45728
rect 2922 45664 2930 45728
rect 2610 45663 2930 45664
rect 5944 45728 6264 45729
rect 5944 45664 5952 45728
rect 6016 45664 6032 45728
rect 6096 45664 6112 45728
rect 6176 45664 6192 45728
rect 6256 45664 6264 45728
rect 5944 45663 6264 45664
rect 4277 45184 4597 45185
rect 4277 45120 4285 45184
rect 4349 45120 4365 45184
rect 4429 45120 4445 45184
rect 4509 45120 4525 45184
rect 4589 45120 4597 45184
rect 4277 45119 4597 45120
rect 7610 45184 7930 45185
rect 7610 45120 7618 45184
rect 7682 45120 7698 45184
rect 7762 45120 7778 45184
rect 7842 45120 7858 45184
rect 7922 45120 7930 45184
rect 7610 45119 7930 45120
rect 2610 44640 2930 44641
rect 2610 44576 2618 44640
rect 2682 44576 2698 44640
rect 2762 44576 2778 44640
rect 2842 44576 2858 44640
rect 2922 44576 2930 44640
rect 2610 44575 2930 44576
rect 5944 44640 6264 44641
rect 5944 44576 5952 44640
rect 6016 44576 6032 44640
rect 6096 44576 6112 44640
rect 6176 44576 6192 44640
rect 6256 44576 6264 44640
rect 5944 44575 6264 44576
rect 4277 44096 4597 44097
rect 4277 44032 4285 44096
rect 4349 44032 4365 44096
rect 4429 44032 4445 44096
rect 4509 44032 4525 44096
rect 4589 44032 4597 44096
rect 4277 44031 4597 44032
rect 7610 44096 7930 44097
rect 7610 44032 7618 44096
rect 7682 44032 7698 44096
rect 7762 44032 7778 44096
rect 7842 44032 7858 44096
rect 7922 44032 7930 44096
rect 7610 44031 7930 44032
rect 2610 43552 2930 43553
rect 2610 43488 2618 43552
rect 2682 43488 2698 43552
rect 2762 43488 2778 43552
rect 2842 43488 2858 43552
rect 2922 43488 2930 43552
rect 2610 43487 2930 43488
rect 5944 43552 6264 43553
rect 5944 43488 5952 43552
rect 6016 43488 6032 43552
rect 6096 43488 6112 43552
rect 6176 43488 6192 43552
rect 6256 43488 6264 43552
rect 5944 43487 6264 43488
rect 4277 43008 4597 43009
rect 4277 42944 4285 43008
rect 4349 42944 4365 43008
rect 4429 42944 4445 43008
rect 4509 42944 4525 43008
rect 4589 42944 4597 43008
rect 4277 42943 4597 42944
rect 7610 43008 7930 43009
rect 7610 42944 7618 43008
rect 7682 42944 7698 43008
rect 7762 42944 7778 43008
rect 7842 42944 7858 43008
rect 7922 42944 7930 43008
rect 7610 42943 7930 42944
rect 2610 42464 2930 42465
rect 2610 42400 2618 42464
rect 2682 42400 2698 42464
rect 2762 42400 2778 42464
rect 2842 42400 2858 42464
rect 2922 42400 2930 42464
rect 2610 42399 2930 42400
rect 5944 42464 6264 42465
rect 5944 42400 5952 42464
rect 6016 42400 6032 42464
rect 6096 42400 6112 42464
rect 6176 42400 6192 42464
rect 6256 42400 6264 42464
rect 5944 42399 6264 42400
rect 4277 41920 4597 41921
rect 4277 41856 4285 41920
rect 4349 41856 4365 41920
rect 4429 41856 4445 41920
rect 4509 41856 4525 41920
rect 4589 41856 4597 41920
rect 4277 41855 4597 41856
rect 7610 41920 7930 41921
rect 7610 41856 7618 41920
rect 7682 41856 7698 41920
rect 7762 41856 7778 41920
rect 7842 41856 7858 41920
rect 7922 41856 7930 41920
rect 7610 41855 7930 41856
rect 2610 41376 2930 41377
rect 2610 41312 2618 41376
rect 2682 41312 2698 41376
rect 2762 41312 2778 41376
rect 2842 41312 2858 41376
rect 2922 41312 2930 41376
rect 2610 41311 2930 41312
rect 5944 41376 6264 41377
rect 5944 41312 5952 41376
rect 6016 41312 6032 41376
rect 6096 41312 6112 41376
rect 6176 41312 6192 41376
rect 6256 41312 6264 41376
rect 5944 41311 6264 41312
rect 4277 40832 4597 40833
rect 4277 40768 4285 40832
rect 4349 40768 4365 40832
rect 4429 40768 4445 40832
rect 4509 40768 4525 40832
rect 4589 40768 4597 40832
rect 4277 40767 4597 40768
rect 7610 40832 7930 40833
rect 7610 40768 7618 40832
rect 7682 40768 7698 40832
rect 7762 40768 7778 40832
rect 7842 40768 7858 40832
rect 7922 40768 7930 40832
rect 7610 40767 7930 40768
rect 2610 40288 2930 40289
rect 2610 40224 2618 40288
rect 2682 40224 2698 40288
rect 2762 40224 2778 40288
rect 2842 40224 2858 40288
rect 2922 40224 2930 40288
rect 2610 40223 2930 40224
rect 5944 40288 6264 40289
rect 5944 40224 5952 40288
rect 6016 40224 6032 40288
rect 6096 40224 6112 40288
rect 6176 40224 6192 40288
rect 6256 40224 6264 40288
rect 5944 40223 6264 40224
rect 4277 39744 4597 39745
rect 4277 39680 4285 39744
rect 4349 39680 4365 39744
rect 4429 39680 4445 39744
rect 4509 39680 4525 39744
rect 4589 39680 4597 39744
rect 4277 39679 4597 39680
rect 7610 39744 7930 39745
rect 7610 39680 7618 39744
rect 7682 39680 7698 39744
rect 7762 39680 7778 39744
rect 7842 39680 7858 39744
rect 7922 39680 7930 39744
rect 7610 39679 7930 39680
rect 2610 39200 2930 39201
rect 2610 39136 2618 39200
rect 2682 39136 2698 39200
rect 2762 39136 2778 39200
rect 2842 39136 2858 39200
rect 2922 39136 2930 39200
rect 2610 39135 2930 39136
rect 5944 39200 6264 39201
rect 5944 39136 5952 39200
rect 6016 39136 6032 39200
rect 6096 39136 6112 39200
rect 6176 39136 6192 39200
rect 6256 39136 6264 39200
rect 5944 39135 6264 39136
rect 4277 38656 4597 38657
rect 4277 38592 4285 38656
rect 4349 38592 4365 38656
rect 4429 38592 4445 38656
rect 4509 38592 4525 38656
rect 4589 38592 4597 38656
rect 4277 38591 4597 38592
rect 7610 38656 7930 38657
rect 7610 38592 7618 38656
rect 7682 38592 7698 38656
rect 7762 38592 7778 38656
rect 7842 38592 7858 38656
rect 7922 38592 7930 38656
rect 7610 38591 7930 38592
rect 2610 38112 2930 38113
rect 2610 38048 2618 38112
rect 2682 38048 2698 38112
rect 2762 38048 2778 38112
rect 2842 38048 2858 38112
rect 2922 38048 2930 38112
rect 2610 38047 2930 38048
rect 5944 38112 6264 38113
rect 5944 38048 5952 38112
rect 6016 38048 6032 38112
rect 6096 38048 6112 38112
rect 6176 38048 6192 38112
rect 6256 38048 6264 38112
rect 5944 38047 6264 38048
rect 4277 37568 4597 37569
rect 4277 37504 4285 37568
rect 4349 37504 4365 37568
rect 4429 37504 4445 37568
rect 4509 37504 4525 37568
rect 4589 37504 4597 37568
rect 4277 37503 4597 37504
rect 7610 37568 7930 37569
rect 7610 37504 7618 37568
rect 7682 37504 7698 37568
rect 7762 37504 7778 37568
rect 7842 37504 7858 37568
rect 7922 37504 7930 37568
rect 7610 37503 7930 37504
rect 2610 37024 2930 37025
rect 2610 36960 2618 37024
rect 2682 36960 2698 37024
rect 2762 36960 2778 37024
rect 2842 36960 2858 37024
rect 2922 36960 2930 37024
rect 2610 36959 2930 36960
rect 5944 37024 6264 37025
rect 5944 36960 5952 37024
rect 6016 36960 6032 37024
rect 6096 36960 6112 37024
rect 6176 36960 6192 37024
rect 6256 36960 6264 37024
rect 5944 36959 6264 36960
rect 4277 36480 4597 36481
rect 4277 36416 4285 36480
rect 4349 36416 4365 36480
rect 4429 36416 4445 36480
rect 4509 36416 4525 36480
rect 4589 36416 4597 36480
rect 4277 36415 4597 36416
rect 7610 36480 7930 36481
rect 7610 36416 7618 36480
rect 7682 36416 7698 36480
rect 7762 36416 7778 36480
rect 7842 36416 7858 36480
rect 7922 36416 7930 36480
rect 7610 36415 7930 36416
rect 2610 35936 2930 35937
rect 2610 35872 2618 35936
rect 2682 35872 2698 35936
rect 2762 35872 2778 35936
rect 2842 35872 2858 35936
rect 2922 35872 2930 35936
rect 2610 35871 2930 35872
rect 5944 35936 6264 35937
rect 5944 35872 5952 35936
rect 6016 35872 6032 35936
rect 6096 35872 6112 35936
rect 6176 35872 6192 35936
rect 6256 35872 6264 35936
rect 5944 35871 6264 35872
rect 4277 35392 4597 35393
rect 4277 35328 4285 35392
rect 4349 35328 4365 35392
rect 4429 35328 4445 35392
rect 4509 35328 4525 35392
rect 4589 35328 4597 35392
rect 4277 35327 4597 35328
rect 7610 35392 7930 35393
rect 7610 35328 7618 35392
rect 7682 35328 7698 35392
rect 7762 35328 7778 35392
rect 7842 35328 7858 35392
rect 7922 35328 7930 35392
rect 7610 35327 7930 35328
rect 2610 34848 2930 34849
rect 2610 34784 2618 34848
rect 2682 34784 2698 34848
rect 2762 34784 2778 34848
rect 2842 34784 2858 34848
rect 2922 34784 2930 34848
rect 2610 34783 2930 34784
rect 5944 34848 6264 34849
rect 5944 34784 5952 34848
rect 6016 34784 6032 34848
rect 6096 34784 6112 34848
rect 6176 34784 6192 34848
rect 6256 34784 6264 34848
rect 5944 34783 6264 34784
rect 4277 34304 4597 34305
rect 4277 34240 4285 34304
rect 4349 34240 4365 34304
rect 4429 34240 4445 34304
rect 4509 34240 4525 34304
rect 4589 34240 4597 34304
rect 4277 34239 4597 34240
rect 7610 34304 7930 34305
rect 7610 34240 7618 34304
rect 7682 34240 7698 34304
rect 7762 34240 7778 34304
rect 7842 34240 7858 34304
rect 7922 34240 7930 34304
rect 7610 34239 7930 34240
rect 2610 33760 2930 33761
rect 2610 33696 2618 33760
rect 2682 33696 2698 33760
rect 2762 33696 2778 33760
rect 2842 33696 2858 33760
rect 2922 33696 2930 33760
rect 2610 33695 2930 33696
rect 5944 33760 6264 33761
rect 5944 33696 5952 33760
rect 6016 33696 6032 33760
rect 6096 33696 6112 33760
rect 6176 33696 6192 33760
rect 6256 33696 6264 33760
rect 5944 33695 6264 33696
rect 4277 33216 4597 33217
rect 4277 33152 4285 33216
rect 4349 33152 4365 33216
rect 4429 33152 4445 33216
rect 4509 33152 4525 33216
rect 4589 33152 4597 33216
rect 4277 33151 4597 33152
rect 7610 33216 7930 33217
rect 7610 33152 7618 33216
rect 7682 33152 7698 33216
rect 7762 33152 7778 33216
rect 7842 33152 7858 33216
rect 7922 33152 7930 33216
rect 7610 33151 7930 33152
rect 2610 32672 2930 32673
rect 2610 32608 2618 32672
rect 2682 32608 2698 32672
rect 2762 32608 2778 32672
rect 2842 32608 2858 32672
rect 2922 32608 2930 32672
rect 2610 32607 2930 32608
rect 5944 32672 6264 32673
rect 5944 32608 5952 32672
rect 6016 32608 6032 32672
rect 6096 32608 6112 32672
rect 6176 32608 6192 32672
rect 6256 32608 6264 32672
rect 5944 32607 6264 32608
rect 4277 32128 4597 32129
rect 4277 32064 4285 32128
rect 4349 32064 4365 32128
rect 4429 32064 4445 32128
rect 4509 32064 4525 32128
rect 4589 32064 4597 32128
rect 4277 32063 4597 32064
rect 7610 32128 7930 32129
rect 7610 32064 7618 32128
rect 7682 32064 7698 32128
rect 7762 32064 7778 32128
rect 7842 32064 7858 32128
rect 7922 32064 7930 32128
rect 7610 32063 7930 32064
rect 2610 31584 2930 31585
rect 2610 31520 2618 31584
rect 2682 31520 2698 31584
rect 2762 31520 2778 31584
rect 2842 31520 2858 31584
rect 2922 31520 2930 31584
rect 2610 31519 2930 31520
rect 5944 31584 6264 31585
rect 5944 31520 5952 31584
rect 6016 31520 6032 31584
rect 6096 31520 6112 31584
rect 6176 31520 6192 31584
rect 6256 31520 6264 31584
rect 5944 31519 6264 31520
rect 4277 31040 4597 31041
rect 4277 30976 4285 31040
rect 4349 30976 4365 31040
rect 4429 30976 4445 31040
rect 4509 30976 4525 31040
rect 4589 30976 4597 31040
rect 4277 30975 4597 30976
rect 7610 31040 7930 31041
rect 7610 30976 7618 31040
rect 7682 30976 7698 31040
rect 7762 30976 7778 31040
rect 7842 30976 7858 31040
rect 7922 30976 7930 31040
rect 7610 30975 7930 30976
rect 2610 30496 2930 30497
rect 2610 30432 2618 30496
rect 2682 30432 2698 30496
rect 2762 30432 2778 30496
rect 2842 30432 2858 30496
rect 2922 30432 2930 30496
rect 2610 30431 2930 30432
rect 5944 30496 6264 30497
rect 5944 30432 5952 30496
rect 6016 30432 6032 30496
rect 6096 30432 6112 30496
rect 6176 30432 6192 30496
rect 6256 30432 6264 30496
rect 5944 30431 6264 30432
rect 4277 29952 4597 29953
rect 4277 29888 4285 29952
rect 4349 29888 4365 29952
rect 4429 29888 4445 29952
rect 4509 29888 4525 29952
rect 4589 29888 4597 29952
rect 4277 29887 4597 29888
rect 7610 29952 7930 29953
rect 7610 29888 7618 29952
rect 7682 29888 7698 29952
rect 7762 29888 7778 29952
rect 7842 29888 7858 29952
rect 7922 29888 7930 29952
rect 7610 29887 7930 29888
rect 2610 29408 2930 29409
rect 2610 29344 2618 29408
rect 2682 29344 2698 29408
rect 2762 29344 2778 29408
rect 2842 29344 2858 29408
rect 2922 29344 2930 29408
rect 2610 29343 2930 29344
rect 5944 29408 6264 29409
rect 5944 29344 5952 29408
rect 6016 29344 6032 29408
rect 6096 29344 6112 29408
rect 6176 29344 6192 29408
rect 6256 29344 6264 29408
rect 5944 29343 6264 29344
rect 4277 28864 4597 28865
rect 4277 28800 4285 28864
rect 4349 28800 4365 28864
rect 4429 28800 4445 28864
rect 4509 28800 4525 28864
rect 4589 28800 4597 28864
rect 4277 28799 4597 28800
rect 7610 28864 7930 28865
rect 7610 28800 7618 28864
rect 7682 28800 7698 28864
rect 7762 28800 7778 28864
rect 7842 28800 7858 28864
rect 7922 28800 7930 28864
rect 7610 28799 7930 28800
rect 2610 28320 2930 28321
rect 2610 28256 2618 28320
rect 2682 28256 2698 28320
rect 2762 28256 2778 28320
rect 2842 28256 2858 28320
rect 2922 28256 2930 28320
rect 2610 28255 2930 28256
rect 5944 28320 6264 28321
rect 5944 28256 5952 28320
rect 6016 28256 6032 28320
rect 6096 28256 6112 28320
rect 6176 28256 6192 28320
rect 6256 28256 6264 28320
rect 5944 28255 6264 28256
rect 4277 27776 4597 27777
rect 4277 27712 4285 27776
rect 4349 27712 4365 27776
rect 4429 27712 4445 27776
rect 4509 27712 4525 27776
rect 4589 27712 4597 27776
rect 4277 27711 4597 27712
rect 7610 27776 7930 27777
rect 7610 27712 7618 27776
rect 7682 27712 7698 27776
rect 7762 27712 7778 27776
rect 7842 27712 7858 27776
rect 7922 27712 7930 27776
rect 7610 27711 7930 27712
rect 2610 27232 2930 27233
rect 2610 27168 2618 27232
rect 2682 27168 2698 27232
rect 2762 27168 2778 27232
rect 2842 27168 2858 27232
rect 2922 27168 2930 27232
rect 2610 27167 2930 27168
rect 5944 27232 6264 27233
rect 5944 27168 5952 27232
rect 6016 27168 6032 27232
rect 6096 27168 6112 27232
rect 6176 27168 6192 27232
rect 6256 27168 6264 27232
rect 5944 27167 6264 27168
rect 4277 26688 4597 26689
rect 4277 26624 4285 26688
rect 4349 26624 4365 26688
rect 4429 26624 4445 26688
rect 4509 26624 4525 26688
rect 4589 26624 4597 26688
rect 4277 26623 4597 26624
rect 7610 26688 7930 26689
rect 7610 26624 7618 26688
rect 7682 26624 7698 26688
rect 7762 26624 7778 26688
rect 7842 26624 7858 26688
rect 7922 26624 7930 26688
rect 7610 26623 7930 26624
rect 2610 26144 2930 26145
rect 2610 26080 2618 26144
rect 2682 26080 2698 26144
rect 2762 26080 2778 26144
rect 2842 26080 2858 26144
rect 2922 26080 2930 26144
rect 2610 26079 2930 26080
rect 5944 26144 6264 26145
rect 5944 26080 5952 26144
rect 6016 26080 6032 26144
rect 6096 26080 6112 26144
rect 6176 26080 6192 26144
rect 6256 26080 6264 26144
rect 5944 26079 6264 26080
rect 4277 25600 4597 25601
rect 4277 25536 4285 25600
rect 4349 25536 4365 25600
rect 4429 25536 4445 25600
rect 4509 25536 4525 25600
rect 4589 25536 4597 25600
rect 4277 25535 4597 25536
rect 7610 25600 7930 25601
rect 7610 25536 7618 25600
rect 7682 25536 7698 25600
rect 7762 25536 7778 25600
rect 7842 25536 7858 25600
rect 7922 25536 7930 25600
rect 7610 25535 7930 25536
rect 2610 25056 2930 25057
rect 2610 24992 2618 25056
rect 2682 24992 2698 25056
rect 2762 24992 2778 25056
rect 2842 24992 2858 25056
rect 2922 24992 2930 25056
rect 2610 24991 2930 24992
rect 5944 25056 6264 25057
rect 5944 24992 5952 25056
rect 6016 24992 6032 25056
rect 6096 24992 6112 25056
rect 6176 24992 6192 25056
rect 6256 24992 6264 25056
rect 5944 24991 6264 24992
rect 4277 24512 4597 24513
rect 4277 24448 4285 24512
rect 4349 24448 4365 24512
rect 4429 24448 4445 24512
rect 4509 24448 4525 24512
rect 4589 24448 4597 24512
rect 4277 24447 4597 24448
rect 7610 24512 7930 24513
rect 7610 24448 7618 24512
rect 7682 24448 7698 24512
rect 7762 24448 7778 24512
rect 7842 24448 7858 24512
rect 7922 24448 7930 24512
rect 7610 24447 7930 24448
rect 3785 24306 3851 24309
rect 62 24304 3851 24306
rect 62 24248 3790 24304
rect 3846 24248 3851 24304
rect 62 24246 3851 24248
rect 62 23792 122 24246
rect 3785 24243 3851 24246
rect 2610 23968 2930 23969
rect 2610 23904 2618 23968
rect 2682 23904 2698 23968
rect 2762 23904 2778 23968
rect 2842 23904 2858 23968
rect 2922 23904 2930 23968
rect 2610 23903 2930 23904
rect 5944 23968 6264 23969
rect 5944 23904 5952 23968
rect 6016 23904 6032 23968
rect 6096 23904 6112 23968
rect 6176 23904 6192 23968
rect 6256 23904 6264 23968
rect 5944 23903 6264 23904
rect 0 23672 480 23792
rect 4277 23424 4597 23425
rect 4277 23360 4285 23424
rect 4349 23360 4365 23424
rect 4429 23360 4445 23424
rect 4509 23360 4525 23424
rect 4589 23360 4597 23424
rect 4277 23359 4597 23360
rect 7610 23424 7930 23425
rect 7610 23360 7618 23424
rect 7682 23360 7698 23424
rect 7762 23360 7778 23424
rect 7842 23360 7858 23424
rect 7922 23360 7930 23424
rect 7610 23359 7930 23360
rect 2610 22880 2930 22881
rect 2610 22816 2618 22880
rect 2682 22816 2698 22880
rect 2762 22816 2778 22880
rect 2842 22816 2858 22880
rect 2922 22816 2930 22880
rect 2610 22815 2930 22816
rect 5944 22880 6264 22881
rect 5944 22816 5952 22880
rect 6016 22816 6032 22880
rect 6096 22816 6112 22880
rect 6176 22816 6192 22880
rect 6256 22816 6264 22880
rect 5944 22815 6264 22816
rect 4277 22336 4597 22337
rect 4277 22272 4285 22336
rect 4349 22272 4365 22336
rect 4429 22272 4445 22336
rect 4509 22272 4525 22336
rect 4589 22272 4597 22336
rect 4277 22271 4597 22272
rect 7610 22336 7930 22337
rect 7610 22272 7618 22336
rect 7682 22272 7698 22336
rect 7762 22272 7778 22336
rect 7842 22272 7858 22336
rect 7922 22272 7930 22336
rect 7610 22271 7930 22272
rect 2610 21792 2930 21793
rect 2610 21728 2618 21792
rect 2682 21728 2698 21792
rect 2762 21728 2778 21792
rect 2842 21728 2858 21792
rect 2922 21728 2930 21792
rect 2610 21727 2930 21728
rect 5944 21792 6264 21793
rect 5944 21728 5952 21792
rect 6016 21728 6032 21792
rect 6096 21728 6112 21792
rect 6176 21728 6192 21792
rect 6256 21728 6264 21792
rect 5944 21727 6264 21728
rect 4277 21248 4597 21249
rect 4277 21184 4285 21248
rect 4349 21184 4365 21248
rect 4429 21184 4445 21248
rect 4509 21184 4525 21248
rect 4589 21184 4597 21248
rect 4277 21183 4597 21184
rect 7610 21248 7930 21249
rect 7610 21184 7618 21248
rect 7682 21184 7698 21248
rect 7762 21184 7778 21248
rect 7842 21184 7858 21248
rect 7922 21184 7930 21248
rect 7610 21183 7930 21184
rect 2610 20704 2930 20705
rect 2610 20640 2618 20704
rect 2682 20640 2698 20704
rect 2762 20640 2778 20704
rect 2842 20640 2858 20704
rect 2922 20640 2930 20704
rect 2610 20639 2930 20640
rect 5944 20704 6264 20705
rect 5944 20640 5952 20704
rect 6016 20640 6032 20704
rect 6096 20640 6112 20704
rect 6176 20640 6192 20704
rect 6256 20640 6264 20704
rect 5944 20639 6264 20640
rect 4277 20160 4597 20161
rect 4277 20096 4285 20160
rect 4349 20096 4365 20160
rect 4429 20096 4445 20160
rect 4509 20096 4525 20160
rect 4589 20096 4597 20160
rect 4277 20095 4597 20096
rect 7610 20160 7930 20161
rect 7610 20096 7618 20160
rect 7682 20096 7698 20160
rect 7762 20096 7778 20160
rect 7842 20096 7858 20160
rect 7922 20096 7930 20160
rect 7610 20095 7930 20096
rect 2610 19616 2930 19617
rect 2610 19552 2618 19616
rect 2682 19552 2698 19616
rect 2762 19552 2778 19616
rect 2842 19552 2858 19616
rect 2922 19552 2930 19616
rect 2610 19551 2930 19552
rect 5944 19616 6264 19617
rect 5944 19552 5952 19616
rect 6016 19552 6032 19616
rect 6096 19552 6112 19616
rect 6176 19552 6192 19616
rect 6256 19552 6264 19616
rect 5944 19551 6264 19552
rect 4277 19072 4597 19073
rect 4277 19008 4285 19072
rect 4349 19008 4365 19072
rect 4429 19008 4445 19072
rect 4509 19008 4525 19072
rect 4589 19008 4597 19072
rect 4277 19007 4597 19008
rect 7610 19072 7930 19073
rect 7610 19008 7618 19072
rect 7682 19008 7698 19072
rect 7762 19008 7778 19072
rect 7842 19008 7858 19072
rect 7922 19008 7930 19072
rect 7610 19007 7930 19008
rect 2610 18528 2930 18529
rect 2610 18464 2618 18528
rect 2682 18464 2698 18528
rect 2762 18464 2778 18528
rect 2842 18464 2858 18528
rect 2922 18464 2930 18528
rect 2610 18463 2930 18464
rect 5944 18528 6264 18529
rect 5944 18464 5952 18528
rect 6016 18464 6032 18528
rect 6096 18464 6112 18528
rect 6176 18464 6192 18528
rect 6256 18464 6264 18528
rect 5944 18463 6264 18464
rect 4277 17984 4597 17985
rect 4277 17920 4285 17984
rect 4349 17920 4365 17984
rect 4429 17920 4445 17984
rect 4509 17920 4525 17984
rect 4589 17920 4597 17984
rect 4277 17919 4597 17920
rect 7610 17984 7930 17985
rect 7610 17920 7618 17984
rect 7682 17920 7698 17984
rect 7762 17920 7778 17984
rect 7842 17920 7858 17984
rect 7922 17920 7930 17984
rect 7610 17919 7930 17920
rect 2610 17440 2930 17441
rect 2610 17376 2618 17440
rect 2682 17376 2698 17440
rect 2762 17376 2778 17440
rect 2842 17376 2858 17440
rect 2922 17376 2930 17440
rect 2610 17375 2930 17376
rect 5944 17440 6264 17441
rect 5944 17376 5952 17440
rect 6016 17376 6032 17440
rect 6096 17376 6112 17440
rect 6176 17376 6192 17440
rect 6256 17376 6264 17440
rect 5944 17375 6264 17376
rect 4797 17234 4863 17237
rect 4797 17232 9690 17234
rect 4797 17176 4802 17232
rect 4858 17176 9690 17232
rect 4797 17174 9690 17176
rect 4797 17171 4863 17174
rect 4277 16896 4597 16897
rect 4277 16832 4285 16896
rect 4349 16832 4365 16896
rect 4429 16832 4445 16896
rect 4509 16832 4525 16896
rect 4589 16832 4597 16896
rect 4277 16831 4597 16832
rect 7610 16896 7930 16897
rect 7610 16832 7618 16896
rect 7682 16832 7698 16896
rect 7762 16832 7778 16896
rect 7842 16832 7858 16896
rect 7922 16832 7930 16896
rect 7610 16831 7930 16832
rect 9630 16720 9690 17174
rect 9520 16600 10000 16720
rect 2610 16352 2930 16353
rect 2610 16288 2618 16352
rect 2682 16288 2698 16352
rect 2762 16288 2778 16352
rect 2842 16288 2858 16352
rect 2922 16288 2930 16352
rect 2610 16287 2930 16288
rect 5944 16352 6264 16353
rect 5944 16288 5952 16352
rect 6016 16288 6032 16352
rect 6096 16288 6112 16352
rect 6176 16288 6192 16352
rect 6256 16288 6264 16352
rect 5944 16287 6264 16288
rect 4277 15808 4597 15809
rect 4277 15744 4285 15808
rect 4349 15744 4365 15808
rect 4429 15744 4445 15808
rect 4509 15744 4525 15808
rect 4589 15744 4597 15808
rect 4277 15743 4597 15744
rect 7610 15808 7930 15809
rect 7610 15744 7618 15808
rect 7682 15744 7698 15808
rect 7762 15744 7778 15808
rect 7842 15744 7858 15808
rect 7922 15744 7930 15808
rect 7610 15743 7930 15744
rect 2610 15264 2930 15265
rect 2610 15200 2618 15264
rect 2682 15200 2698 15264
rect 2762 15200 2778 15264
rect 2842 15200 2858 15264
rect 2922 15200 2930 15264
rect 2610 15199 2930 15200
rect 5944 15264 6264 15265
rect 5944 15200 5952 15264
rect 6016 15200 6032 15264
rect 6096 15200 6112 15264
rect 6176 15200 6192 15264
rect 6256 15200 6264 15264
rect 5944 15199 6264 15200
rect 4277 14720 4597 14721
rect 4277 14656 4285 14720
rect 4349 14656 4365 14720
rect 4429 14656 4445 14720
rect 4509 14656 4525 14720
rect 4589 14656 4597 14720
rect 4277 14655 4597 14656
rect 7610 14720 7930 14721
rect 7610 14656 7618 14720
rect 7682 14656 7698 14720
rect 7762 14656 7778 14720
rect 7842 14656 7858 14720
rect 7922 14656 7930 14720
rect 7610 14655 7930 14656
rect 2610 14176 2930 14177
rect 2610 14112 2618 14176
rect 2682 14112 2698 14176
rect 2762 14112 2778 14176
rect 2842 14112 2858 14176
rect 2922 14112 2930 14176
rect 2610 14111 2930 14112
rect 5944 14176 6264 14177
rect 5944 14112 5952 14176
rect 6016 14112 6032 14176
rect 6096 14112 6112 14176
rect 6176 14112 6192 14176
rect 6256 14112 6264 14176
rect 5944 14111 6264 14112
rect 4277 13632 4597 13633
rect 4277 13568 4285 13632
rect 4349 13568 4365 13632
rect 4429 13568 4445 13632
rect 4509 13568 4525 13632
rect 4589 13568 4597 13632
rect 4277 13567 4597 13568
rect 7610 13632 7930 13633
rect 7610 13568 7618 13632
rect 7682 13568 7698 13632
rect 7762 13568 7778 13632
rect 7842 13568 7858 13632
rect 7922 13568 7930 13632
rect 7610 13567 7930 13568
rect 2610 13088 2930 13089
rect 2610 13024 2618 13088
rect 2682 13024 2698 13088
rect 2762 13024 2778 13088
rect 2842 13024 2858 13088
rect 2922 13024 2930 13088
rect 2610 13023 2930 13024
rect 5944 13088 6264 13089
rect 5944 13024 5952 13088
rect 6016 13024 6032 13088
rect 6096 13024 6112 13088
rect 6176 13024 6192 13088
rect 6256 13024 6264 13088
rect 5944 13023 6264 13024
rect 4277 12544 4597 12545
rect 4277 12480 4285 12544
rect 4349 12480 4365 12544
rect 4429 12480 4445 12544
rect 4509 12480 4525 12544
rect 4589 12480 4597 12544
rect 4277 12479 4597 12480
rect 7610 12544 7930 12545
rect 7610 12480 7618 12544
rect 7682 12480 7698 12544
rect 7762 12480 7778 12544
rect 7842 12480 7858 12544
rect 7922 12480 7930 12544
rect 7610 12479 7930 12480
rect 2610 12000 2930 12001
rect 2610 11936 2618 12000
rect 2682 11936 2698 12000
rect 2762 11936 2778 12000
rect 2842 11936 2858 12000
rect 2922 11936 2930 12000
rect 2610 11935 2930 11936
rect 5944 12000 6264 12001
rect 5944 11936 5952 12000
rect 6016 11936 6032 12000
rect 6096 11936 6112 12000
rect 6176 11936 6192 12000
rect 6256 11936 6264 12000
rect 5944 11935 6264 11936
rect 4277 11456 4597 11457
rect 4277 11392 4285 11456
rect 4349 11392 4365 11456
rect 4429 11392 4445 11456
rect 4509 11392 4525 11456
rect 4589 11392 4597 11456
rect 4277 11391 4597 11392
rect 7610 11456 7930 11457
rect 7610 11392 7618 11456
rect 7682 11392 7698 11456
rect 7762 11392 7778 11456
rect 7842 11392 7858 11456
rect 7922 11392 7930 11456
rect 7610 11391 7930 11392
rect 2610 10912 2930 10913
rect 2610 10848 2618 10912
rect 2682 10848 2698 10912
rect 2762 10848 2778 10912
rect 2842 10848 2858 10912
rect 2922 10848 2930 10912
rect 2610 10847 2930 10848
rect 5944 10912 6264 10913
rect 5944 10848 5952 10912
rect 6016 10848 6032 10912
rect 6096 10848 6112 10912
rect 6176 10848 6192 10912
rect 6256 10848 6264 10912
rect 5944 10847 6264 10848
rect 4277 10368 4597 10369
rect 4277 10304 4285 10368
rect 4349 10304 4365 10368
rect 4429 10304 4445 10368
rect 4509 10304 4525 10368
rect 4589 10304 4597 10368
rect 4277 10303 4597 10304
rect 7610 10368 7930 10369
rect 7610 10304 7618 10368
rect 7682 10304 7698 10368
rect 7762 10304 7778 10368
rect 7842 10304 7858 10368
rect 7922 10304 7930 10368
rect 7610 10303 7930 10304
rect 2610 9824 2930 9825
rect 2610 9760 2618 9824
rect 2682 9760 2698 9824
rect 2762 9760 2778 9824
rect 2842 9760 2858 9824
rect 2922 9760 2930 9824
rect 2610 9759 2930 9760
rect 5944 9824 6264 9825
rect 5944 9760 5952 9824
rect 6016 9760 6032 9824
rect 6096 9760 6112 9824
rect 6176 9760 6192 9824
rect 6256 9760 6264 9824
rect 5944 9759 6264 9760
rect 4277 9280 4597 9281
rect 4277 9216 4285 9280
rect 4349 9216 4365 9280
rect 4429 9216 4445 9280
rect 4509 9216 4525 9280
rect 4589 9216 4597 9280
rect 4277 9215 4597 9216
rect 7610 9280 7930 9281
rect 7610 9216 7618 9280
rect 7682 9216 7698 9280
rect 7762 9216 7778 9280
rect 7842 9216 7858 9280
rect 7922 9216 7930 9280
rect 7610 9215 7930 9216
rect 2610 8736 2930 8737
rect 2610 8672 2618 8736
rect 2682 8672 2698 8736
rect 2762 8672 2778 8736
rect 2842 8672 2858 8736
rect 2922 8672 2930 8736
rect 2610 8671 2930 8672
rect 5944 8736 6264 8737
rect 5944 8672 5952 8736
rect 6016 8672 6032 8736
rect 6096 8672 6112 8736
rect 6176 8672 6192 8736
rect 6256 8672 6264 8736
rect 5944 8671 6264 8672
rect 4277 8192 4597 8193
rect 4277 8128 4285 8192
rect 4349 8128 4365 8192
rect 4429 8128 4445 8192
rect 4509 8128 4525 8192
rect 4589 8128 4597 8192
rect 4277 8127 4597 8128
rect 7610 8192 7930 8193
rect 7610 8128 7618 8192
rect 7682 8128 7698 8192
rect 7762 8128 7778 8192
rect 7842 8128 7858 8192
rect 7922 8128 7930 8192
rect 7610 8127 7930 8128
rect 2610 7648 2930 7649
rect 2610 7584 2618 7648
rect 2682 7584 2698 7648
rect 2762 7584 2778 7648
rect 2842 7584 2858 7648
rect 2922 7584 2930 7648
rect 2610 7583 2930 7584
rect 5944 7648 6264 7649
rect 5944 7584 5952 7648
rect 6016 7584 6032 7648
rect 6096 7584 6112 7648
rect 6176 7584 6192 7648
rect 6256 7584 6264 7648
rect 5944 7583 6264 7584
rect 4277 7104 4597 7105
rect 4277 7040 4285 7104
rect 4349 7040 4365 7104
rect 4429 7040 4445 7104
rect 4509 7040 4525 7104
rect 4589 7040 4597 7104
rect 4277 7039 4597 7040
rect 7610 7104 7930 7105
rect 7610 7040 7618 7104
rect 7682 7040 7698 7104
rect 7762 7040 7778 7104
rect 7842 7040 7858 7104
rect 7922 7040 7930 7104
rect 7610 7039 7930 7040
rect 2610 6560 2930 6561
rect 2610 6496 2618 6560
rect 2682 6496 2698 6560
rect 2762 6496 2778 6560
rect 2842 6496 2858 6560
rect 2922 6496 2930 6560
rect 2610 6495 2930 6496
rect 5944 6560 6264 6561
rect 5944 6496 5952 6560
rect 6016 6496 6032 6560
rect 6096 6496 6112 6560
rect 6176 6496 6192 6560
rect 6256 6496 6264 6560
rect 5944 6495 6264 6496
rect 4277 6016 4597 6017
rect 4277 5952 4285 6016
rect 4349 5952 4365 6016
rect 4429 5952 4445 6016
rect 4509 5952 4525 6016
rect 4589 5952 4597 6016
rect 4277 5951 4597 5952
rect 7610 6016 7930 6017
rect 7610 5952 7618 6016
rect 7682 5952 7698 6016
rect 7762 5952 7778 6016
rect 7842 5952 7858 6016
rect 7922 5952 7930 6016
rect 7610 5951 7930 5952
rect 2610 5472 2930 5473
rect 2610 5408 2618 5472
rect 2682 5408 2698 5472
rect 2762 5408 2778 5472
rect 2842 5408 2858 5472
rect 2922 5408 2930 5472
rect 2610 5407 2930 5408
rect 5944 5472 6264 5473
rect 5944 5408 5952 5472
rect 6016 5408 6032 5472
rect 6096 5408 6112 5472
rect 6176 5408 6192 5472
rect 6256 5408 6264 5472
rect 5944 5407 6264 5408
rect 4277 4928 4597 4929
rect 4277 4864 4285 4928
rect 4349 4864 4365 4928
rect 4429 4864 4445 4928
rect 4509 4864 4525 4928
rect 4589 4864 4597 4928
rect 4277 4863 4597 4864
rect 7610 4928 7930 4929
rect 7610 4864 7618 4928
rect 7682 4864 7698 4928
rect 7762 4864 7778 4928
rect 7842 4864 7858 4928
rect 7922 4864 7930 4928
rect 7610 4863 7930 4864
rect 2610 4384 2930 4385
rect 2610 4320 2618 4384
rect 2682 4320 2698 4384
rect 2762 4320 2778 4384
rect 2842 4320 2858 4384
rect 2922 4320 2930 4384
rect 2610 4319 2930 4320
rect 5944 4384 6264 4385
rect 5944 4320 5952 4384
rect 6016 4320 6032 4384
rect 6096 4320 6112 4384
rect 6176 4320 6192 4384
rect 6256 4320 6264 4384
rect 5944 4319 6264 4320
rect 4277 3840 4597 3841
rect 4277 3776 4285 3840
rect 4349 3776 4365 3840
rect 4429 3776 4445 3840
rect 4509 3776 4525 3840
rect 4589 3776 4597 3840
rect 4277 3775 4597 3776
rect 7610 3840 7930 3841
rect 7610 3776 7618 3840
rect 7682 3776 7698 3840
rect 7762 3776 7778 3840
rect 7842 3776 7858 3840
rect 7922 3776 7930 3840
rect 7610 3775 7930 3776
rect 2610 3296 2930 3297
rect 2610 3232 2618 3296
rect 2682 3232 2698 3296
rect 2762 3232 2778 3296
rect 2842 3232 2858 3296
rect 2922 3232 2930 3296
rect 2610 3231 2930 3232
rect 5944 3296 6264 3297
rect 5944 3232 5952 3296
rect 6016 3232 6032 3296
rect 6096 3232 6112 3296
rect 6176 3232 6192 3296
rect 6256 3232 6264 3296
rect 5944 3231 6264 3232
rect 4277 2752 4597 2753
rect 4277 2688 4285 2752
rect 4349 2688 4365 2752
rect 4429 2688 4445 2752
rect 4509 2688 4525 2752
rect 4589 2688 4597 2752
rect 4277 2687 4597 2688
rect 7610 2752 7930 2753
rect 7610 2688 7618 2752
rect 7682 2688 7698 2752
rect 7762 2688 7778 2752
rect 7842 2688 7858 2752
rect 7922 2688 7930 2752
rect 7610 2687 7930 2688
rect 2610 2208 2930 2209
rect 2610 2144 2618 2208
rect 2682 2144 2698 2208
rect 2762 2144 2778 2208
rect 2842 2144 2858 2208
rect 2922 2144 2930 2208
rect 2610 2143 2930 2144
rect 5944 2208 6264 2209
rect 5944 2144 5952 2208
rect 6016 2144 6032 2208
rect 6096 2144 6112 2208
rect 6176 2144 6192 2208
rect 6256 2144 6264 2208
rect 5944 2143 6264 2144
<< via3 >>
rect 2618 330780 2682 330784
rect 2618 330724 2622 330780
rect 2622 330724 2678 330780
rect 2678 330724 2682 330780
rect 2618 330720 2682 330724
rect 2698 330780 2762 330784
rect 2698 330724 2702 330780
rect 2702 330724 2758 330780
rect 2758 330724 2762 330780
rect 2698 330720 2762 330724
rect 2778 330780 2842 330784
rect 2778 330724 2782 330780
rect 2782 330724 2838 330780
rect 2838 330724 2842 330780
rect 2778 330720 2842 330724
rect 2858 330780 2922 330784
rect 2858 330724 2862 330780
rect 2862 330724 2918 330780
rect 2918 330724 2922 330780
rect 2858 330720 2922 330724
rect 5952 330780 6016 330784
rect 5952 330724 5956 330780
rect 5956 330724 6012 330780
rect 6012 330724 6016 330780
rect 5952 330720 6016 330724
rect 6032 330780 6096 330784
rect 6032 330724 6036 330780
rect 6036 330724 6092 330780
rect 6092 330724 6096 330780
rect 6032 330720 6096 330724
rect 6112 330780 6176 330784
rect 6112 330724 6116 330780
rect 6116 330724 6172 330780
rect 6172 330724 6176 330780
rect 6112 330720 6176 330724
rect 6192 330780 6256 330784
rect 6192 330724 6196 330780
rect 6196 330724 6252 330780
rect 6252 330724 6256 330780
rect 6192 330720 6256 330724
rect 4285 330236 4349 330240
rect 4285 330180 4289 330236
rect 4289 330180 4345 330236
rect 4345 330180 4349 330236
rect 4285 330176 4349 330180
rect 4365 330236 4429 330240
rect 4365 330180 4369 330236
rect 4369 330180 4425 330236
rect 4425 330180 4429 330236
rect 4365 330176 4429 330180
rect 4445 330236 4509 330240
rect 4445 330180 4449 330236
rect 4449 330180 4505 330236
rect 4505 330180 4509 330236
rect 4445 330176 4509 330180
rect 4525 330236 4589 330240
rect 4525 330180 4529 330236
rect 4529 330180 4585 330236
rect 4585 330180 4589 330236
rect 4525 330176 4589 330180
rect 7618 330236 7682 330240
rect 7618 330180 7622 330236
rect 7622 330180 7678 330236
rect 7678 330180 7682 330236
rect 7618 330176 7682 330180
rect 7698 330236 7762 330240
rect 7698 330180 7702 330236
rect 7702 330180 7758 330236
rect 7758 330180 7762 330236
rect 7698 330176 7762 330180
rect 7778 330236 7842 330240
rect 7778 330180 7782 330236
rect 7782 330180 7838 330236
rect 7838 330180 7842 330236
rect 7778 330176 7842 330180
rect 7858 330236 7922 330240
rect 7858 330180 7862 330236
rect 7862 330180 7918 330236
rect 7918 330180 7922 330236
rect 7858 330176 7922 330180
rect 2618 329692 2682 329696
rect 2618 329636 2622 329692
rect 2622 329636 2678 329692
rect 2678 329636 2682 329692
rect 2618 329632 2682 329636
rect 2698 329692 2762 329696
rect 2698 329636 2702 329692
rect 2702 329636 2758 329692
rect 2758 329636 2762 329692
rect 2698 329632 2762 329636
rect 2778 329692 2842 329696
rect 2778 329636 2782 329692
rect 2782 329636 2838 329692
rect 2838 329636 2842 329692
rect 2778 329632 2842 329636
rect 2858 329692 2922 329696
rect 2858 329636 2862 329692
rect 2862 329636 2918 329692
rect 2918 329636 2922 329692
rect 2858 329632 2922 329636
rect 5952 329692 6016 329696
rect 5952 329636 5956 329692
rect 5956 329636 6012 329692
rect 6012 329636 6016 329692
rect 5952 329632 6016 329636
rect 6032 329692 6096 329696
rect 6032 329636 6036 329692
rect 6036 329636 6092 329692
rect 6092 329636 6096 329692
rect 6032 329632 6096 329636
rect 6112 329692 6176 329696
rect 6112 329636 6116 329692
rect 6116 329636 6172 329692
rect 6172 329636 6176 329692
rect 6112 329632 6176 329636
rect 6192 329692 6256 329696
rect 6192 329636 6196 329692
rect 6196 329636 6252 329692
rect 6252 329636 6256 329692
rect 6192 329632 6256 329636
rect 4285 329148 4349 329152
rect 4285 329092 4289 329148
rect 4289 329092 4345 329148
rect 4345 329092 4349 329148
rect 4285 329088 4349 329092
rect 4365 329148 4429 329152
rect 4365 329092 4369 329148
rect 4369 329092 4425 329148
rect 4425 329092 4429 329148
rect 4365 329088 4429 329092
rect 4445 329148 4509 329152
rect 4445 329092 4449 329148
rect 4449 329092 4505 329148
rect 4505 329092 4509 329148
rect 4445 329088 4509 329092
rect 4525 329148 4589 329152
rect 4525 329092 4529 329148
rect 4529 329092 4585 329148
rect 4585 329092 4589 329148
rect 4525 329088 4589 329092
rect 7618 329148 7682 329152
rect 7618 329092 7622 329148
rect 7622 329092 7678 329148
rect 7678 329092 7682 329148
rect 7618 329088 7682 329092
rect 7698 329148 7762 329152
rect 7698 329092 7702 329148
rect 7702 329092 7758 329148
rect 7758 329092 7762 329148
rect 7698 329088 7762 329092
rect 7778 329148 7842 329152
rect 7778 329092 7782 329148
rect 7782 329092 7838 329148
rect 7838 329092 7842 329148
rect 7778 329088 7842 329092
rect 7858 329148 7922 329152
rect 7858 329092 7862 329148
rect 7862 329092 7918 329148
rect 7918 329092 7922 329148
rect 7858 329088 7922 329092
rect 2618 328604 2682 328608
rect 2618 328548 2622 328604
rect 2622 328548 2678 328604
rect 2678 328548 2682 328604
rect 2618 328544 2682 328548
rect 2698 328604 2762 328608
rect 2698 328548 2702 328604
rect 2702 328548 2758 328604
rect 2758 328548 2762 328604
rect 2698 328544 2762 328548
rect 2778 328604 2842 328608
rect 2778 328548 2782 328604
rect 2782 328548 2838 328604
rect 2838 328548 2842 328604
rect 2778 328544 2842 328548
rect 2858 328604 2922 328608
rect 2858 328548 2862 328604
rect 2862 328548 2918 328604
rect 2918 328548 2922 328604
rect 2858 328544 2922 328548
rect 5952 328604 6016 328608
rect 5952 328548 5956 328604
rect 5956 328548 6012 328604
rect 6012 328548 6016 328604
rect 5952 328544 6016 328548
rect 6032 328604 6096 328608
rect 6032 328548 6036 328604
rect 6036 328548 6092 328604
rect 6092 328548 6096 328604
rect 6032 328544 6096 328548
rect 6112 328604 6176 328608
rect 6112 328548 6116 328604
rect 6116 328548 6172 328604
rect 6172 328548 6176 328604
rect 6112 328544 6176 328548
rect 6192 328604 6256 328608
rect 6192 328548 6196 328604
rect 6196 328548 6252 328604
rect 6252 328548 6256 328604
rect 6192 328544 6256 328548
rect 4285 328060 4349 328064
rect 4285 328004 4289 328060
rect 4289 328004 4345 328060
rect 4345 328004 4349 328060
rect 4285 328000 4349 328004
rect 4365 328060 4429 328064
rect 4365 328004 4369 328060
rect 4369 328004 4425 328060
rect 4425 328004 4429 328060
rect 4365 328000 4429 328004
rect 4445 328060 4509 328064
rect 4445 328004 4449 328060
rect 4449 328004 4505 328060
rect 4505 328004 4509 328060
rect 4445 328000 4509 328004
rect 4525 328060 4589 328064
rect 4525 328004 4529 328060
rect 4529 328004 4585 328060
rect 4585 328004 4589 328060
rect 4525 328000 4589 328004
rect 7618 328060 7682 328064
rect 7618 328004 7622 328060
rect 7622 328004 7678 328060
rect 7678 328004 7682 328060
rect 7618 328000 7682 328004
rect 7698 328060 7762 328064
rect 7698 328004 7702 328060
rect 7702 328004 7758 328060
rect 7758 328004 7762 328060
rect 7698 328000 7762 328004
rect 7778 328060 7842 328064
rect 7778 328004 7782 328060
rect 7782 328004 7838 328060
rect 7838 328004 7842 328060
rect 7778 328000 7842 328004
rect 7858 328060 7922 328064
rect 7858 328004 7862 328060
rect 7862 328004 7918 328060
rect 7918 328004 7922 328060
rect 7858 328000 7922 328004
rect 2618 327516 2682 327520
rect 2618 327460 2622 327516
rect 2622 327460 2678 327516
rect 2678 327460 2682 327516
rect 2618 327456 2682 327460
rect 2698 327516 2762 327520
rect 2698 327460 2702 327516
rect 2702 327460 2758 327516
rect 2758 327460 2762 327516
rect 2698 327456 2762 327460
rect 2778 327516 2842 327520
rect 2778 327460 2782 327516
rect 2782 327460 2838 327516
rect 2838 327460 2842 327516
rect 2778 327456 2842 327460
rect 2858 327516 2922 327520
rect 2858 327460 2862 327516
rect 2862 327460 2918 327516
rect 2918 327460 2922 327516
rect 2858 327456 2922 327460
rect 5952 327516 6016 327520
rect 5952 327460 5956 327516
rect 5956 327460 6012 327516
rect 6012 327460 6016 327516
rect 5952 327456 6016 327460
rect 6032 327516 6096 327520
rect 6032 327460 6036 327516
rect 6036 327460 6092 327516
rect 6092 327460 6096 327516
rect 6032 327456 6096 327460
rect 6112 327516 6176 327520
rect 6112 327460 6116 327516
rect 6116 327460 6172 327516
rect 6172 327460 6176 327516
rect 6112 327456 6176 327460
rect 6192 327516 6256 327520
rect 6192 327460 6196 327516
rect 6196 327460 6252 327516
rect 6252 327460 6256 327516
rect 6192 327456 6256 327460
rect 4285 326972 4349 326976
rect 4285 326916 4289 326972
rect 4289 326916 4345 326972
rect 4345 326916 4349 326972
rect 4285 326912 4349 326916
rect 4365 326972 4429 326976
rect 4365 326916 4369 326972
rect 4369 326916 4425 326972
rect 4425 326916 4429 326972
rect 4365 326912 4429 326916
rect 4445 326972 4509 326976
rect 4445 326916 4449 326972
rect 4449 326916 4505 326972
rect 4505 326916 4509 326972
rect 4445 326912 4509 326916
rect 4525 326972 4589 326976
rect 4525 326916 4529 326972
rect 4529 326916 4585 326972
rect 4585 326916 4589 326972
rect 4525 326912 4589 326916
rect 7618 326972 7682 326976
rect 7618 326916 7622 326972
rect 7622 326916 7678 326972
rect 7678 326916 7682 326972
rect 7618 326912 7682 326916
rect 7698 326972 7762 326976
rect 7698 326916 7702 326972
rect 7702 326916 7758 326972
rect 7758 326916 7762 326972
rect 7698 326912 7762 326916
rect 7778 326972 7842 326976
rect 7778 326916 7782 326972
rect 7782 326916 7838 326972
rect 7838 326916 7842 326972
rect 7778 326912 7842 326916
rect 7858 326972 7922 326976
rect 7858 326916 7862 326972
rect 7862 326916 7918 326972
rect 7918 326916 7922 326972
rect 7858 326912 7922 326916
rect 2618 326428 2682 326432
rect 2618 326372 2622 326428
rect 2622 326372 2678 326428
rect 2678 326372 2682 326428
rect 2618 326368 2682 326372
rect 2698 326428 2762 326432
rect 2698 326372 2702 326428
rect 2702 326372 2758 326428
rect 2758 326372 2762 326428
rect 2698 326368 2762 326372
rect 2778 326428 2842 326432
rect 2778 326372 2782 326428
rect 2782 326372 2838 326428
rect 2838 326372 2842 326428
rect 2778 326368 2842 326372
rect 2858 326428 2922 326432
rect 2858 326372 2862 326428
rect 2862 326372 2918 326428
rect 2918 326372 2922 326428
rect 2858 326368 2922 326372
rect 5952 326428 6016 326432
rect 5952 326372 5956 326428
rect 5956 326372 6012 326428
rect 6012 326372 6016 326428
rect 5952 326368 6016 326372
rect 6032 326428 6096 326432
rect 6032 326372 6036 326428
rect 6036 326372 6092 326428
rect 6092 326372 6096 326428
rect 6032 326368 6096 326372
rect 6112 326428 6176 326432
rect 6112 326372 6116 326428
rect 6116 326372 6172 326428
rect 6172 326372 6176 326428
rect 6112 326368 6176 326372
rect 6192 326428 6256 326432
rect 6192 326372 6196 326428
rect 6196 326372 6252 326428
rect 6252 326372 6256 326428
rect 6192 326368 6256 326372
rect 4285 325884 4349 325888
rect 4285 325828 4289 325884
rect 4289 325828 4345 325884
rect 4345 325828 4349 325884
rect 4285 325824 4349 325828
rect 4365 325884 4429 325888
rect 4365 325828 4369 325884
rect 4369 325828 4425 325884
rect 4425 325828 4429 325884
rect 4365 325824 4429 325828
rect 4445 325884 4509 325888
rect 4445 325828 4449 325884
rect 4449 325828 4505 325884
rect 4505 325828 4509 325884
rect 4445 325824 4509 325828
rect 4525 325884 4589 325888
rect 4525 325828 4529 325884
rect 4529 325828 4585 325884
rect 4585 325828 4589 325884
rect 4525 325824 4589 325828
rect 7618 325884 7682 325888
rect 7618 325828 7622 325884
rect 7622 325828 7678 325884
rect 7678 325828 7682 325884
rect 7618 325824 7682 325828
rect 7698 325884 7762 325888
rect 7698 325828 7702 325884
rect 7702 325828 7758 325884
rect 7758 325828 7762 325884
rect 7698 325824 7762 325828
rect 7778 325884 7842 325888
rect 7778 325828 7782 325884
rect 7782 325828 7838 325884
rect 7838 325828 7842 325884
rect 7778 325824 7842 325828
rect 7858 325884 7922 325888
rect 7858 325828 7862 325884
rect 7862 325828 7918 325884
rect 7918 325828 7922 325884
rect 7858 325824 7922 325828
rect 2618 325340 2682 325344
rect 2618 325284 2622 325340
rect 2622 325284 2678 325340
rect 2678 325284 2682 325340
rect 2618 325280 2682 325284
rect 2698 325340 2762 325344
rect 2698 325284 2702 325340
rect 2702 325284 2758 325340
rect 2758 325284 2762 325340
rect 2698 325280 2762 325284
rect 2778 325340 2842 325344
rect 2778 325284 2782 325340
rect 2782 325284 2838 325340
rect 2838 325284 2842 325340
rect 2778 325280 2842 325284
rect 2858 325340 2922 325344
rect 2858 325284 2862 325340
rect 2862 325284 2918 325340
rect 2918 325284 2922 325340
rect 2858 325280 2922 325284
rect 5952 325340 6016 325344
rect 5952 325284 5956 325340
rect 5956 325284 6012 325340
rect 6012 325284 6016 325340
rect 5952 325280 6016 325284
rect 6032 325340 6096 325344
rect 6032 325284 6036 325340
rect 6036 325284 6092 325340
rect 6092 325284 6096 325340
rect 6032 325280 6096 325284
rect 6112 325340 6176 325344
rect 6112 325284 6116 325340
rect 6116 325284 6172 325340
rect 6172 325284 6176 325340
rect 6112 325280 6176 325284
rect 6192 325340 6256 325344
rect 6192 325284 6196 325340
rect 6196 325284 6252 325340
rect 6252 325284 6256 325340
rect 6192 325280 6256 325284
rect 4285 324796 4349 324800
rect 4285 324740 4289 324796
rect 4289 324740 4345 324796
rect 4345 324740 4349 324796
rect 4285 324736 4349 324740
rect 4365 324796 4429 324800
rect 4365 324740 4369 324796
rect 4369 324740 4425 324796
rect 4425 324740 4429 324796
rect 4365 324736 4429 324740
rect 4445 324796 4509 324800
rect 4445 324740 4449 324796
rect 4449 324740 4505 324796
rect 4505 324740 4509 324796
rect 4445 324736 4509 324740
rect 4525 324796 4589 324800
rect 4525 324740 4529 324796
rect 4529 324740 4585 324796
rect 4585 324740 4589 324796
rect 4525 324736 4589 324740
rect 7618 324796 7682 324800
rect 7618 324740 7622 324796
rect 7622 324740 7678 324796
rect 7678 324740 7682 324796
rect 7618 324736 7682 324740
rect 7698 324796 7762 324800
rect 7698 324740 7702 324796
rect 7702 324740 7758 324796
rect 7758 324740 7762 324796
rect 7698 324736 7762 324740
rect 7778 324796 7842 324800
rect 7778 324740 7782 324796
rect 7782 324740 7838 324796
rect 7838 324740 7842 324796
rect 7778 324736 7842 324740
rect 7858 324796 7922 324800
rect 7858 324740 7862 324796
rect 7862 324740 7918 324796
rect 7918 324740 7922 324796
rect 7858 324736 7922 324740
rect 2618 324252 2682 324256
rect 2618 324196 2622 324252
rect 2622 324196 2678 324252
rect 2678 324196 2682 324252
rect 2618 324192 2682 324196
rect 2698 324252 2762 324256
rect 2698 324196 2702 324252
rect 2702 324196 2758 324252
rect 2758 324196 2762 324252
rect 2698 324192 2762 324196
rect 2778 324252 2842 324256
rect 2778 324196 2782 324252
rect 2782 324196 2838 324252
rect 2838 324196 2842 324252
rect 2778 324192 2842 324196
rect 2858 324252 2922 324256
rect 2858 324196 2862 324252
rect 2862 324196 2918 324252
rect 2918 324196 2922 324252
rect 2858 324192 2922 324196
rect 5952 324252 6016 324256
rect 5952 324196 5956 324252
rect 5956 324196 6012 324252
rect 6012 324196 6016 324252
rect 5952 324192 6016 324196
rect 6032 324252 6096 324256
rect 6032 324196 6036 324252
rect 6036 324196 6092 324252
rect 6092 324196 6096 324252
rect 6032 324192 6096 324196
rect 6112 324252 6176 324256
rect 6112 324196 6116 324252
rect 6116 324196 6172 324252
rect 6172 324196 6176 324252
rect 6112 324192 6176 324196
rect 6192 324252 6256 324256
rect 6192 324196 6196 324252
rect 6196 324196 6252 324252
rect 6252 324196 6256 324252
rect 6192 324192 6256 324196
rect 4285 323708 4349 323712
rect 4285 323652 4289 323708
rect 4289 323652 4345 323708
rect 4345 323652 4349 323708
rect 4285 323648 4349 323652
rect 4365 323708 4429 323712
rect 4365 323652 4369 323708
rect 4369 323652 4425 323708
rect 4425 323652 4429 323708
rect 4365 323648 4429 323652
rect 4445 323708 4509 323712
rect 4445 323652 4449 323708
rect 4449 323652 4505 323708
rect 4505 323652 4509 323708
rect 4445 323648 4509 323652
rect 4525 323708 4589 323712
rect 4525 323652 4529 323708
rect 4529 323652 4585 323708
rect 4585 323652 4589 323708
rect 4525 323648 4589 323652
rect 7618 323708 7682 323712
rect 7618 323652 7622 323708
rect 7622 323652 7678 323708
rect 7678 323652 7682 323708
rect 7618 323648 7682 323652
rect 7698 323708 7762 323712
rect 7698 323652 7702 323708
rect 7702 323652 7758 323708
rect 7758 323652 7762 323708
rect 7698 323648 7762 323652
rect 7778 323708 7842 323712
rect 7778 323652 7782 323708
rect 7782 323652 7838 323708
rect 7838 323652 7842 323708
rect 7778 323648 7842 323652
rect 7858 323708 7922 323712
rect 7858 323652 7862 323708
rect 7862 323652 7918 323708
rect 7918 323652 7922 323708
rect 7858 323648 7922 323652
rect 2618 323164 2682 323168
rect 2618 323108 2622 323164
rect 2622 323108 2678 323164
rect 2678 323108 2682 323164
rect 2618 323104 2682 323108
rect 2698 323164 2762 323168
rect 2698 323108 2702 323164
rect 2702 323108 2758 323164
rect 2758 323108 2762 323164
rect 2698 323104 2762 323108
rect 2778 323164 2842 323168
rect 2778 323108 2782 323164
rect 2782 323108 2838 323164
rect 2838 323108 2842 323164
rect 2778 323104 2842 323108
rect 2858 323164 2922 323168
rect 2858 323108 2862 323164
rect 2862 323108 2918 323164
rect 2918 323108 2922 323164
rect 2858 323104 2922 323108
rect 5952 323164 6016 323168
rect 5952 323108 5956 323164
rect 5956 323108 6012 323164
rect 6012 323108 6016 323164
rect 5952 323104 6016 323108
rect 6032 323164 6096 323168
rect 6032 323108 6036 323164
rect 6036 323108 6092 323164
rect 6092 323108 6096 323164
rect 6032 323104 6096 323108
rect 6112 323164 6176 323168
rect 6112 323108 6116 323164
rect 6116 323108 6172 323164
rect 6172 323108 6176 323164
rect 6112 323104 6176 323108
rect 6192 323164 6256 323168
rect 6192 323108 6196 323164
rect 6196 323108 6252 323164
rect 6252 323108 6256 323164
rect 6192 323104 6256 323108
rect 4285 322620 4349 322624
rect 4285 322564 4289 322620
rect 4289 322564 4345 322620
rect 4345 322564 4349 322620
rect 4285 322560 4349 322564
rect 4365 322620 4429 322624
rect 4365 322564 4369 322620
rect 4369 322564 4425 322620
rect 4425 322564 4429 322620
rect 4365 322560 4429 322564
rect 4445 322620 4509 322624
rect 4445 322564 4449 322620
rect 4449 322564 4505 322620
rect 4505 322564 4509 322620
rect 4445 322560 4509 322564
rect 4525 322620 4589 322624
rect 4525 322564 4529 322620
rect 4529 322564 4585 322620
rect 4585 322564 4589 322620
rect 4525 322560 4589 322564
rect 7618 322620 7682 322624
rect 7618 322564 7622 322620
rect 7622 322564 7678 322620
rect 7678 322564 7682 322620
rect 7618 322560 7682 322564
rect 7698 322620 7762 322624
rect 7698 322564 7702 322620
rect 7702 322564 7758 322620
rect 7758 322564 7762 322620
rect 7698 322560 7762 322564
rect 7778 322620 7842 322624
rect 7778 322564 7782 322620
rect 7782 322564 7838 322620
rect 7838 322564 7842 322620
rect 7778 322560 7842 322564
rect 7858 322620 7922 322624
rect 7858 322564 7862 322620
rect 7862 322564 7918 322620
rect 7918 322564 7922 322620
rect 7858 322560 7922 322564
rect 2618 322076 2682 322080
rect 2618 322020 2622 322076
rect 2622 322020 2678 322076
rect 2678 322020 2682 322076
rect 2618 322016 2682 322020
rect 2698 322076 2762 322080
rect 2698 322020 2702 322076
rect 2702 322020 2758 322076
rect 2758 322020 2762 322076
rect 2698 322016 2762 322020
rect 2778 322076 2842 322080
rect 2778 322020 2782 322076
rect 2782 322020 2838 322076
rect 2838 322020 2842 322076
rect 2778 322016 2842 322020
rect 2858 322076 2922 322080
rect 2858 322020 2862 322076
rect 2862 322020 2918 322076
rect 2918 322020 2922 322076
rect 2858 322016 2922 322020
rect 5952 322076 6016 322080
rect 5952 322020 5956 322076
rect 5956 322020 6012 322076
rect 6012 322020 6016 322076
rect 5952 322016 6016 322020
rect 6032 322076 6096 322080
rect 6032 322020 6036 322076
rect 6036 322020 6092 322076
rect 6092 322020 6096 322076
rect 6032 322016 6096 322020
rect 6112 322076 6176 322080
rect 6112 322020 6116 322076
rect 6116 322020 6172 322076
rect 6172 322020 6176 322076
rect 6112 322016 6176 322020
rect 6192 322076 6256 322080
rect 6192 322020 6196 322076
rect 6196 322020 6252 322076
rect 6252 322020 6256 322076
rect 6192 322016 6256 322020
rect 4285 321532 4349 321536
rect 4285 321476 4289 321532
rect 4289 321476 4345 321532
rect 4345 321476 4349 321532
rect 4285 321472 4349 321476
rect 4365 321532 4429 321536
rect 4365 321476 4369 321532
rect 4369 321476 4425 321532
rect 4425 321476 4429 321532
rect 4365 321472 4429 321476
rect 4445 321532 4509 321536
rect 4445 321476 4449 321532
rect 4449 321476 4505 321532
rect 4505 321476 4509 321532
rect 4445 321472 4509 321476
rect 4525 321532 4589 321536
rect 4525 321476 4529 321532
rect 4529 321476 4585 321532
rect 4585 321476 4589 321532
rect 4525 321472 4589 321476
rect 7618 321532 7682 321536
rect 7618 321476 7622 321532
rect 7622 321476 7678 321532
rect 7678 321476 7682 321532
rect 7618 321472 7682 321476
rect 7698 321532 7762 321536
rect 7698 321476 7702 321532
rect 7702 321476 7758 321532
rect 7758 321476 7762 321532
rect 7698 321472 7762 321476
rect 7778 321532 7842 321536
rect 7778 321476 7782 321532
rect 7782 321476 7838 321532
rect 7838 321476 7842 321532
rect 7778 321472 7842 321476
rect 7858 321532 7922 321536
rect 7858 321476 7862 321532
rect 7862 321476 7918 321532
rect 7918 321476 7922 321532
rect 7858 321472 7922 321476
rect 2618 320988 2682 320992
rect 2618 320932 2622 320988
rect 2622 320932 2678 320988
rect 2678 320932 2682 320988
rect 2618 320928 2682 320932
rect 2698 320988 2762 320992
rect 2698 320932 2702 320988
rect 2702 320932 2758 320988
rect 2758 320932 2762 320988
rect 2698 320928 2762 320932
rect 2778 320988 2842 320992
rect 2778 320932 2782 320988
rect 2782 320932 2838 320988
rect 2838 320932 2842 320988
rect 2778 320928 2842 320932
rect 2858 320988 2922 320992
rect 2858 320932 2862 320988
rect 2862 320932 2918 320988
rect 2918 320932 2922 320988
rect 2858 320928 2922 320932
rect 5952 320988 6016 320992
rect 5952 320932 5956 320988
rect 5956 320932 6012 320988
rect 6012 320932 6016 320988
rect 5952 320928 6016 320932
rect 6032 320988 6096 320992
rect 6032 320932 6036 320988
rect 6036 320932 6092 320988
rect 6092 320932 6096 320988
rect 6032 320928 6096 320932
rect 6112 320988 6176 320992
rect 6112 320932 6116 320988
rect 6116 320932 6172 320988
rect 6172 320932 6176 320988
rect 6112 320928 6176 320932
rect 6192 320988 6256 320992
rect 6192 320932 6196 320988
rect 6196 320932 6252 320988
rect 6252 320932 6256 320988
rect 6192 320928 6256 320932
rect 4285 320444 4349 320448
rect 4285 320388 4289 320444
rect 4289 320388 4345 320444
rect 4345 320388 4349 320444
rect 4285 320384 4349 320388
rect 4365 320444 4429 320448
rect 4365 320388 4369 320444
rect 4369 320388 4425 320444
rect 4425 320388 4429 320444
rect 4365 320384 4429 320388
rect 4445 320444 4509 320448
rect 4445 320388 4449 320444
rect 4449 320388 4505 320444
rect 4505 320388 4509 320444
rect 4445 320384 4509 320388
rect 4525 320444 4589 320448
rect 4525 320388 4529 320444
rect 4529 320388 4585 320444
rect 4585 320388 4589 320444
rect 4525 320384 4589 320388
rect 7618 320444 7682 320448
rect 7618 320388 7622 320444
rect 7622 320388 7678 320444
rect 7678 320388 7682 320444
rect 7618 320384 7682 320388
rect 7698 320444 7762 320448
rect 7698 320388 7702 320444
rect 7702 320388 7758 320444
rect 7758 320388 7762 320444
rect 7698 320384 7762 320388
rect 7778 320444 7842 320448
rect 7778 320388 7782 320444
rect 7782 320388 7838 320444
rect 7838 320388 7842 320444
rect 7778 320384 7842 320388
rect 7858 320444 7922 320448
rect 7858 320388 7862 320444
rect 7862 320388 7918 320444
rect 7918 320388 7922 320444
rect 7858 320384 7922 320388
rect 2618 319900 2682 319904
rect 2618 319844 2622 319900
rect 2622 319844 2678 319900
rect 2678 319844 2682 319900
rect 2618 319840 2682 319844
rect 2698 319900 2762 319904
rect 2698 319844 2702 319900
rect 2702 319844 2758 319900
rect 2758 319844 2762 319900
rect 2698 319840 2762 319844
rect 2778 319900 2842 319904
rect 2778 319844 2782 319900
rect 2782 319844 2838 319900
rect 2838 319844 2842 319900
rect 2778 319840 2842 319844
rect 2858 319900 2922 319904
rect 2858 319844 2862 319900
rect 2862 319844 2918 319900
rect 2918 319844 2922 319900
rect 2858 319840 2922 319844
rect 5952 319900 6016 319904
rect 5952 319844 5956 319900
rect 5956 319844 6012 319900
rect 6012 319844 6016 319900
rect 5952 319840 6016 319844
rect 6032 319900 6096 319904
rect 6032 319844 6036 319900
rect 6036 319844 6092 319900
rect 6092 319844 6096 319900
rect 6032 319840 6096 319844
rect 6112 319900 6176 319904
rect 6112 319844 6116 319900
rect 6116 319844 6172 319900
rect 6172 319844 6176 319900
rect 6112 319840 6176 319844
rect 6192 319900 6256 319904
rect 6192 319844 6196 319900
rect 6196 319844 6252 319900
rect 6252 319844 6256 319900
rect 6192 319840 6256 319844
rect 4285 319356 4349 319360
rect 4285 319300 4289 319356
rect 4289 319300 4345 319356
rect 4345 319300 4349 319356
rect 4285 319296 4349 319300
rect 4365 319356 4429 319360
rect 4365 319300 4369 319356
rect 4369 319300 4425 319356
rect 4425 319300 4429 319356
rect 4365 319296 4429 319300
rect 4445 319356 4509 319360
rect 4445 319300 4449 319356
rect 4449 319300 4505 319356
rect 4505 319300 4509 319356
rect 4445 319296 4509 319300
rect 4525 319356 4589 319360
rect 4525 319300 4529 319356
rect 4529 319300 4585 319356
rect 4585 319300 4589 319356
rect 4525 319296 4589 319300
rect 7618 319356 7682 319360
rect 7618 319300 7622 319356
rect 7622 319300 7678 319356
rect 7678 319300 7682 319356
rect 7618 319296 7682 319300
rect 7698 319356 7762 319360
rect 7698 319300 7702 319356
rect 7702 319300 7758 319356
rect 7758 319300 7762 319356
rect 7698 319296 7762 319300
rect 7778 319356 7842 319360
rect 7778 319300 7782 319356
rect 7782 319300 7838 319356
rect 7838 319300 7842 319356
rect 7778 319296 7842 319300
rect 7858 319356 7922 319360
rect 7858 319300 7862 319356
rect 7862 319300 7918 319356
rect 7918 319300 7922 319356
rect 7858 319296 7922 319300
rect 2618 318812 2682 318816
rect 2618 318756 2622 318812
rect 2622 318756 2678 318812
rect 2678 318756 2682 318812
rect 2618 318752 2682 318756
rect 2698 318812 2762 318816
rect 2698 318756 2702 318812
rect 2702 318756 2758 318812
rect 2758 318756 2762 318812
rect 2698 318752 2762 318756
rect 2778 318812 2842 318816
rect 2778 318756 2782 318812
rect 2782 318756 2838 318812
rect 2838 318756 2842 318812
rect 2778 318752 2842 318756
rect 2858 318812 2922 318816
rect 2858 318756 2862 318812
rect 2862 318756 2918 318812
rect 2918 318756 2922 318812
rect 2858 318752 2922 318756
rect 5952 318812 6016 318816
rect 5952 318756 5956 318812
rect 5956 318756 6012 318812
rect 6012 318756 6016 318812
rect 5952 318752 6016 318756
rect 6032 318812 6096 318816
rect 6032 318756 6036 318812
rect 6036 318756 6092 318812
rect 6092 318756 6096 318812
rect 6032 318752 6096 318756
rect 6112 318812 6176 318816
rect 6112 318756 6116 318812
rect 6116 318756 6172 318812
rect 6172 318756 6176 318812
rect 6112 318752 6176 318756
rect 6192 318812 6256 318816
rect 6192 318756 6196 318812
rect 6196 318756 6252 318812
rect 6252 318756 6256 318812
rect 6192 318752 6256 318756
rect 4285 318268 4349 318272
rect 4285 318212 4289 318268
rect 4289 318212 4345 318268
rect 4345 318212 4349 318268
rect 4285 318208 4349 318212
rect 4365 318268 4429 318272
rect 4365 318212 4369 318268
rect 4369 318212 4425 318268
rect 4425 318212 4429 318268
rect 4365 318208 4429 318212
rect 4445 318268 4509 318272
rect 4445 318212 4449 318268
rect 4449 318212 4505 318268
rect 4505 318212 4509 318268
rect 4445 318208 4509 318212
rect 4525 318268 4589 318272
rect 4525 318212 4529 318268
rect 4529 318212 4585 318268
rect 4585 318212 4589 318268
rect 4525 318208 4589 318212
rect 7618 318268 7682 318272
rect 7618 318212 7622 318268
rect 7622 318212 7678 318268
rect 7678 318212 7682 318268
rect 7618 318208 7682 318212
rect 7698 318268 7762 318272
rect 7698 318212 7702 318268
rect 7702 318212 7758 318268
rect 7758 318212 7762 318268
rect 7698 318208 7762 318212
rect 7778 318268 7842 318272
rect 7778 318212 7782 318268
rect 7782 318212 7838 318268
rect 7838 318212 7842 318268
rect 7778 318208 7842 318212
rect 7858 318268 7922 318272
rect 7858 318212 7862 318268
rect 7862 318212 7918 318268
rect 7918 318212 7922 318268
rect 7858 318208 7922 318212
rect 2618 317724 2682 317728
rect 2618 317668 2622 317724
rect 2622 317668 2678 317724
rect 2678 317668 2682 317724
rect 2618 317664 2682 317668
rect 2698 317724 2762 317728
rect 2698 317668 2702 317724
rect 2702 317668 2758 317724
rect 2758 317668 2762 317724
rect 2698 317664 2762 317668
rect 2778 317724 2842 317728
rect 2778 317668 2782 317724
rect 2782 317668 2838 317724
rect 2838 317668 2842 317724
rect 2778 317664 2842 317668
rect 2858 317724 2922 317728
rect 2858 317668 2862 317724
rect 2862 317668 2918 317724
rect 2918 317668 2922 317724
rect 2858 317664 2922 317668
rect 5952 317724 6016 317728
rect 5952 317668 5956 317724
rect 5956 317668 6012 317724
rect 6012 317668 6016 317724
rect 5952 317664 6016 317668
rect 6032 317724 6096 317728
rect 6032 317668 6036 317724
rect 6036 317668 6092 317724
rect 6092 317668 6096 317724
rect 6032 317664 6096 317668
rect 6112 317724 6176 317728
rect 6112 317668 6116 317724
rect 6116 317668 6172 317724
rect 6172 317668 6176 317724
rect 6112 317664 6176 317668
rect 6192 317724 6256 317728
rect 6192 317668 6196 317724
rect 6196 317668 6252 317724
rect 6252 317668 6256 317724
rect 6192 317664 6256 317668
rect 4285 317180 4349 317184
rect 4285 317124 4289 317180
rect 4289 317124 4345 317180
rect 4345 317124 4349 317180
rect 4285 317120 4349 317124
rect 4365 317180 4429 317184
rect 4365 317124 4369 317180
rect 4369 317124 4425 317180
rect 4425 317124 4429 317180
rect 4365 317120 4429 317124
rect 4445 317180 4509 317184
rect 4445 317124 4449 317180
rect 4449 317124 4505 317180
rect 4505 317124 4509 317180
rect 4445 317120 4509 317124
rect 4525 317180 4589 317184
rect 4525 317124 4529 317180
rect 4529 317124 4585 317180
rect 4585 317124 4589 317180
rect 4525 317120 4589 317124
rect 7618 317180 7682 317184
rect 7618 317124 7622 317180
rect 7622 317124 7678 317180
rect 7678 317124 7682 317180
rect 7618 317120 7682 317124
rect 7698 317180 7762 317184
rect 7698 317124 7702 317180
rect 7702 317124 7758 317180
rect 7758 317124 7762 317180
rect 7698 317120 7762 317124
rect 7778 317180 7842 317184
rect 7778 317124 7782 317180
rect 7782 317124 7838 317180
rect 7838 317124 7842 317180
rect 7778 317120 7842 317124
rect 7858 317180 7922 317184
rect 7858 317124 7862 317180
rect 7862 317124 7918 317180
rect 7918 317124 7922 317180
rect 7858 317120 7922 317124
rect 2618 316636 2682 316640
rect 2618 316580 2622 316636
rect 2622 316580 2678 316636
rect 2678 316580 2682 316636
rect 2618 316576 2682 316580
rect 2698 316636 2762 316640
rect 2698 316580 2702 316636
rect 2702 316580 2758 316636
rect 2758 316580 2762 316636
rect 2698 316576 2762 316580
rect 2778 316636 2842 316640
rect 2778 316580 2782 316636
rect 2782 316580 2838 316636
rect 2838 316580 2842 316636
rect 2778 316576 2842 316580
rect 2858 316636 2922 316640
rect 2858 316580 2862 316636
rect 2862 316580 2918 316636
rect 2918 316580 2922 316636
rect 2858 316576 2922 316580
rect 5952 316636 6016 316640
rect 5952 316580 5956 316636
rect 5956 316580 6012 316636
rect 6012 316580 6016 316636
rect 5952 316576 6016 316580
rect 6032 316636 6096 316640
rect 6032 316580 6036 316636
rect 6036 316580 6092 316636
rect 6092 316580 6096 316636
rect 6032 316576 6096 316580
rect 6112 316636 6176 316640
rect 6112 316580 6116 316636
rect 6116 316580 6172 316636
rect 6172 316580 6176 316636
rect 6112 316576 6176 316580
rect 6192 316636 6256 316640
rect 6192 316580 6196 316636
rect 6196 316580 6252 316636
rect 6252 316580 6256 316636
rect 6192 316576 6256 316580
rect 4285 316092 4349 316096
rect 4285 316036 4289 316092
rect 4289 316036 4345 316092
rect 4345 316036 4349 316092
rect 4285 316032 4349 316036
rect 4365 316092 4429 316096
rect 4365 316036 4369 316092
rect 4369 316036 4425 316092
rect 4425 316036 4429 316092
rect 4365 316032 4429 316036
rect 4445 316092 4509 316096
rect 4445 316036 4449 316092
rect 4449 316036 4505 316092
rect 4505 316036 4509 316092
rect 4445 316032 4509 316036
rect 4525 316092 4589 316096
rect 4525 316036 4529 316092
rect 4529 316036 4585 316092
rect 4585 316036 4589 316092
rect 4525 316032 4589 316036
rect 7618 316092 7682 316096
rect 7618 316036 7622 316092
rect 7622 316036 7678 316092
rect 7678 316036 7682 316092
rect 7618 316032 7682 316036
rect 7698 316092 7762 316096
rect 7698 316036 7702 316092
rect 7702 316036 7758 316092
rect 7758 316036 7762 316092
rect 7698 316032 7762 316036
rect 7778 316092 7842 316096
rect 7778 316036 7782 316092
rect 7782 316036 7838 316092
rect 7838 316036 7842 316092
rect 7778 316032 7842 316036
rect 7858 316092 7922 316096
rect 7858 316036 7862 316092
rect 7862 316036 7918 316092
rect 7918 316036 7922 316092
rect 7858 316032 7922 316036
rect 2618 315548 2682 315552
rect 2618 315492 2622 315548
rect 2622 315492 2678 315548
rect 2678 315492 2682 315548
rect 2618 315488 2682 315492
rect 2698 315548 2762 315552
rect 2698 315492 2702 315548
rect 2702 315492 2758 315548
rect 2758 315492 2762 315548
rect 2698 315488 2762 315492
rect 2778 315548 2842 315552
rect 2778 315492 2782 315548
rect 2782 315492 2838 315548
rect 2838 315492 2842 315548
rect 2778 315488 2842 315492
rect 2858 315548 2922 315552
rect 2858 315492 2862 315548
rect 2862 315492 2918 315548
rect 2918 315492 2922 315548
rect 2858 315488 2922 315492
rect 5952 315548 6016 315552
rect 5952 315492 5956 315548
rect 5956 315492 6012 315548
rect 6012 315492 6016 315548
rect 5952 315488 6016 315492
rect 6032 315548 6096 315552
rect 6032 315492 6036 315548
rect 6036 315492 6092 315548
rect 6092 315492 6096 315548
rect 6032 315488 6096 315492
rect 6112 315548 6176 315552
rect 6112 315492 6116 315548
rect 6116 315492 6172 315548
rect 6172 315492 6176 315548
rect 6112 315488 6176 315492
rect 6192 315548 6256 315552
rect 6192 315492 6196 315548
rect 6196 315492 6252 315548
rect 6252 315492 6256 315548
rect 6192 315488 6256 315492
rect 4285 315004 4349 315008
rect 4285 314948 4289 315004
rect 4289 314948 4345 315004
rect 4345 314948 4349 315004
rect 4285 314944 4349 314948
rect 4365 315004 4429 315008
rect 4365 314948 4369 315004
rect 4369 314948 4425 315004
rect 4425 314948 4429 315004
rect 4365 314944 4429 314948
rect 4445 315004 4509 315008
rect 4445 314948 4449 315004
rect 4449 314948 4505 315004
rect 4505 314948 4509 315004
rect 4445 314944 4509 314948
rect 4525 315004 4589 315008
rect 4525 314948 4529 315004
rect 4529 314948 4585 315004
rect 4585 314948 4589 315004
rect 4525 314944 4589 314948
rect 7618 315004 7682 315008
rect 7618 314948 7622 315004
rect 7622 314948 7678 315004
rect 7678 314948 7682 315004
rect 7618 314944 7682 314948
rect 7698 315004 7762 315008
rect 7698 314948 7702 315004
rect 7702 314948 7758 315004
rect 7758 314948 7762 315004
rect 7698 314944 7762 314948
rect 7778 315004 7842 315008
rect 7778 314948 7782 315004
rect 7782 314948 7838 315004
rect 7838 314948 7842 315004
rect 7778 314944 7842 314948
rect 7858 315004 7922 315008
rect 7858 314948 7862 315004
rect 7862 314948 7918 315004
rect 7918 314948 7922 315004
rect 7858 314944 7922 314948
rect 2618 314460 2682 314464
rect 2618 314404 2622 314460
rect 2622 314404 2678 314460
rect 2678 314404 2682 314460
rect 2618 314400 2682 314404
rect 2698 314460 2762 314464
rect 2698 314404 2702 314460
rect 2702 314404 2758 314460
rect 2758 314404 2762 314460
rect 2698 314400 2762 314404
rect 2778 314460 2842 314464
rect 2778 314404 2782 314460
rect 2782 314404 2838 314460
rect 2838 314404 2842 314460
rect 2778 314400 2842 314404
rect 2858 314460 2922 314464
rect 2858 314404 2862 314460
rect 2862 314404 2918 314460
rect 2918 314404 2922 314460
rect 2858 314400 2922 314404
rect 5952 314460 6016 314464
rect 5952 314404 5956 314460
rect 5956 314404 6012 314460
rect 6012 314404 6016 314460
rect 5952 314400 6016 314404
rect 6032 314460 6096 314464
rect 6032 314404 6036 314460
rect 6036 314404 6092 314460
rect 6092 314404 6096 314460
rect 6032 314400 6096 314404
rect 6112 314460 6176 314464
rect 6112 314404 6116 314460
rect 6116 314404 6172 314460
rect 6172 314404 6176 314460
rect 6112 314400 6176 314404
rect 6192 314460 6256 314464
rect 6192 314404 6196 314460
rect 6196 314404 6252 314460
rect 6252 314404 6256 314460
rect 6192 314400 6256 314404
rect 4285 313916 4349 313920
rect 4285 313860 4289 313916
rect 4289 313860 4345 313916
rect 4345 313860 4349 313916
rect 4285 313856 4349 313860
rect 4365 313916 4429 313920
rect 4365 313860 4369 313916
rect 4369 313860 4425 313916
rect 4425 313860 4429 313916
rect 4365 313856 4429 313860
rect 4445 313916 4509 313920
rect 4445 313860 4449 313916
rect 4449 313860 4505 313916
rect 4505 313860 4509 313916
rect 4445 313856 4509 313860
rect 4525 313916 4589 313920
rect 4525 313860 4529 313916
rect 4529 313860 4585 313916
rect 4585 313860 4589 313916
rect 4525 313856 4589 313860
rect 7618 313916 7682 313920
rect 7618 313860 7622 313916
rect 7622 313860 7678 313916
rect 7678 313860 7682 313916
rect 7618 313856 7682 313860
rect 7698 313916 7762 313920
rect 7698 313860 7702 313916
rect 7702 313860 7758 313916
rect 7758 313860 7762 313916
rect 7698 313856 7762 313860
rect 7778 313916 7842 313920
rect 7778 313860 7782 313916
rect 7782 313860 7838 313916
rect 7838 313860 7842 313916
rect 7778 313856 7842 313860
rect 7858 313916 7922 313920
rect 7858 313860 7862 313916
rect 7862 313860 7918 313916
rect 7918 313860 7922 313916
rect 7858 313856 7922 313860
rect 2618 313372 2682 313376
rect 2618 313316 2622 313372
rect 2622 313316 2678 313372
rect 2678 313316 2682 313372
rect 2618 313312 2682 313316
rect 2698 313372 2762 313376
rect 2698 313316 2702 313372
rect 2702 313316 2758 313372
rect 2758 313316 2762 313372
rect 2698 313312 2762 313316
rect 2778 313372 2842 313376
rect 2778 313316 2782 313372
rect 2782 313316 2838 313372
rect 2838 313316 2842 313372
rect 2778 313312 2842 313316
rect 2858 313372 2922 313376
rect 2858 313316 2862 313372
rect 2862 313316 2918 313372
rect 2918 313316 2922 313372
rect 2858 313312 2922 313316
rect 5952 313372 6016 313376
rect 5952 313316 5956 313372
rect 5956 313316 6012 313372
rect 6012 313316 6016 313372
rect 5952 313312 6016 313316
rect 6032 313372 6096 313376
rect 6032 313316 6036 313372
rect 6036 313316 6092 313372
rect 6092 313316 6096 313372
rect 6032 313312 6096 313316
rect 6112 313372 6176 313376
rect 6112 313316 6116 313372
rect 6116 313316 6172 313372
rect 6172 313316 6176 313372
rect 6112 313312 6176 313316
rect 6192 313372 6256 313376
rect 6192 313316 6196 313372
rect 6196 313316 6252 313372
rect 6252 313316 6256 313372
rect 6192 313312 6256 313316
rect 4285 312828 4349 312832
rect 4285 312772 4289 312828
rect 4289 312772 4345 312828
rect 4345 312772 4349 312828
rect 4285 312768 4349 312772
rect 4365 312828 4429 312832
rect 4365 312772 4369 312828
rect 4369 312772 4425 312828
rect 4425 312772 4429 312828
rect 4365 312768 4429 312772
rect 4445 312828 4509 312832
rect 4445 312772 4449 312828
rect 4449 312772 4505 312828
rect 4505 312772 4509 312828
rect 4445 312768 4509 312772
rect 4525 312828 4589 312832
rect 4525 312772 4529 312828
rect 4529 312772 4585 312828
rect 4585 312772 4589 312828
rect 4525 312768 4589 312772
rect 7618 312828 7682 312832
rect 7618 312772 7622 312828
rect 7622 312772 7678 312828
rect 7678 312772 7682 312828
rect 7618 312768 7682 312772
rect 7698 312828 7762 312832
rect 7698 312772 7702 312828
rect 7702 312772 7758 312828
rect 7758 312772 7762 312828
rect 7698 312768 7762 312772
rect 7778 312828 7842 312832
rect 7778 312772 7782 312828
rect 7782 312772 7838 312828
rect 7838 312772 7842 312828
rect 7778 312768 7842 312772
rect 7858 312828 7922 312832
rect 7858 312772 7862 312828
rect 7862 312772 7918 312828
rect 7918 312772 7922 312828
rect 7858 312768 7922 312772
rect 2618 312284 2682 312288
rect 2618 312228 2622 312284
rect 2622 312228 2678 312284
rect 2678 312228 2682 312284
rect 2618 312224 2682 312228
rect 2698 312284 2762 312288
rect 2698 312228 2702 312284
rect 2702 312228 2758 312284
rect 2758 312228 2762 312284
rect 2698 312224 2762 312228
rect 2778 312284 2842 312288
rect 2778 312228 2782 312284
rect 2782 312228 2838 312284
rect 2838 312228 2842 312284
rect 2778 312224 2842 312228
rect 2858 312284 2922 312288
rect 2858 312228 2862 312284
rect 2862 312228 2918 312284
rect 2918 312228 2922 312284
rect 2858 312224 2922 312228
rect 5952 312284 6016 312288
rect 5952 312228 5956 312284
rect 5956 312228 6012 312284
rect 6012 312228 6016 312284
rect 5952 312224 6016 312228
rect 6032 312284 6096 312288
rect 6032 312228 6036 312284
rect 6036 312228 6092 312284
rect 6092 312228 6096 312284
rect 6032 312224 6096 312228
rect 6112 312284 6176 312288
rect 6112 312228 6116 312284
rect 6116 312228 6172 312284
rect 6172 312228 6176 312284
rect 6112 312224 6176 312228
rect 6192 312284 6256 312288
rect 6192 312228 6196 312284
rect 6196 312228 6252 312284
rect 6252 312228 6256 312284
rect 6192 312224 6256 312228
rect 4285 311740 4349 311744
rect 4285 311684 4289 311740
rect 4289 311684 4345 311740
rect 4345 311684 4349 311740
rect 4285 311680 4349 311684
rect 4365 311740 4429 311744
rect 4365 311684 4369 311740
rect 4369 311684 4425 311740
rect 4425 311684 4429 311740
rect 4365 311680 4429 311684
rect 4445 311740 4509 311744
rect 4445 311684 4449 311740
rect 4449 311684 4505 311740
rect 4505 311684 4509 311740
rect 4445 311680 4509 311684
rect 4525 311740 4589 311744
rect 4525 311684 4529 311740
rect 4529 311684 4585 311740
rect 4585 311684 4589 311740
rect 4525 311680 4589 311684
rect 7618 311740 7682 311744
rect 7618 311684 7622 311740
rect 7622 311684 7678 311740
rect 7678 311684 7682 311740
rect 7618 311680 7682 311684
rect 7698 311740 7762 311744
rect 7698 311684 7702 311740
rect 7702 311684 7758 311740
rect 7758 311684 7762 311740
rect 7698 311680 7762 311684
rect 7778 311740 7842 311744
rect 7778 311684 7782 311740
rect 7782 311684 7838 311740
rect 7838 311684 7842 311740
rect 7778 311680 7842 311684
rect 7858 311740 7922 311744
rect 7858 311684 7862 311740
rect 7862 311684 7918 311740
rect 7918 311684 7922 311740
rect 7858 311680 7922 311684
rect 2618 311196 2682 311200
rect 2618 311140 2622 311196
rect 2622 311140 2678 311196
rect 2678 311140 2682 311196
rect 2618 311136 2682 311140
rect 2698 311196 2762 311200
rect 2698 311140 2702 311196
rect 2702 311140 2758 311196
rect 2758 311140 2762 311196
rect 2698 311136 2762 311140
rect 2778 311196 2842 311200
rect 2778 311140 2782 311196
rect 2782 311140 2838 311196
rect 2838 311140 2842 311196
rect 2778 311136 2842 311140
rect 2858 311196 2922 311200
rect 2858 311140 2862 311196
rect 2862 311140 2918 311196
rect 2918 311140 2922 311196
rect 2858 311136 2922 311140
rect 5952 311196 6016 311200
rect 5952 311140 5956 311196
rect 5956 311140 6012 311196
rect 6012 311140 6016 311196
rect 5952 311136 6016 311140
rect 6032 311196 6096 311200
rect 6032 311140 6036 311196
rect 6036 311140 6092 311196
rect 6092 311140 6096 311196
rect 6032 311136 6096 311140
rect 6112 311196 6176 311200
rect 6112 311140 6116 311196
rect 6116 311140 6172 311196
rect 6172 311140 6176 311196
rect 6112 311136 6176 311140
rect 6192 311196 6256 311200
rect 6192 311140 6196 311196
rect 6196 311140 6252 311196
rect 6252 311140 6256 311196
rect 6192 311136 6256 311140
rect 4285 310652 4349 310656
rect 4285 310596 4289 310652
rect 4289 310596 4345 310652
rect 4345 310596 4349 310652
rect 4285 310592 4349 310596
rect 4365 310652 4429 310656
rect 4365 310596 4369 310652
rect 4369 310596 4425 310652
rect 4425 310596 4429 310652
rect 4365 310592 4429 310596
rect 4445 310652 4509 310656
rect 4445 310596 4449 310652
rect 4449 310596 4505 310652
rect 4505 310596 4509 310652
rect 4445 310592 4509 310596
rect 4525 310652 4589 310656
rect 4525 310596 4529 310652
rect 4529 310596 4585 310652
rect 4585 310596 4589 310652
rect 4525 310592 4589 310596
rect 7618 310652 7682 310656
rect 7618 310596 7622 310652
rect 7622 310596 7678 310652
rect 7678 310596 7682 310652
rect 7618 310592 7682 310596
rect 7698 310652 7762 310656
rect 7698 310596 7702 310652
rect 7702 310596 7758 310652
rect 7758 310596 7762 310652
rect 7698 310592 7762 310596
rect 7778 310652 7842 310656
rect 7778 310596 7782 310652
rect 7782 310596 7838 310652
rect 7838 310596 7842 310652
rect 7778 310592 7842 310596
rect 7858 310652 7922 310656
rect 7858 310596 7862 310652
rect 7862 310596 7918 310652
rect 7918 310596 7922 310652
rect 7858 310592 7922 310596
rect 2618 310108 2682 310112
rect 2618 310052 2622 310108
rect 2622 310052 2678 310108
rect 2678 310052 2682 310108
rect 2618 310048 2682 310052
rect 2698 310108 2762 310112
rect 2698 310052 2702 310108
rect 2702 310052 2758 310108
rect 2758 310052 2762 310108
rect 2698 310048 2762 310052
rect 2778 310108 2842 310112
rect 2778 310052 2782 310108
rect 2782 310052 2838 310108
rect 2838 310052 2842 310108
rect 2778 310048 2842 310052
rect 2858 310108 2922 310112
rect 2858 310052 2862 310108
rect 2862 310052 2918 310108
rect 2918 310052 2922 310108
rect 2858 310048 2922 310052
rect 5952 310108 6016 310112
rect 5952 310052 5956 310108
rect 5956 310052 6012 310108
rect 6012 310052 6016 310108
rect 5952 310048 6016 310052
rect 6032 310108 6096 310112
rect 6032 310052 6036 310108
rect 6036 310052 6092 310108
rect 6092 310052 6096 310108
rect 6032 310048 6096 310052
rect 6112 310108 6176 310112
rect 6112 310052 6116 310108
rect 6116 310052 6172 310108
rect 6172 310052 6176 310108
rect 6112 310048 6176 310052
rect 6192 310108 6256 310112
rect 6192 310052 6196 310108
rect 6196 310052 6252 310108
rect 6252 310052 6256 310108
rect 6192 310048 6256 310052
rect 4285 309564 4349 309568
rect 4285 309508 4289 309564
rect 4289 309508 4345 309564
rect 4345 309508 4349 309564
rect 4285 309504 4349 309508
rect 4365 309564 4429 309568
rect 4365 309508 4369 309564
rect 4369 309508 4425 309564
rect 4425 309508 4429 309564
rect 4365 309504 4429 309508
rect 4445 309564 4509 309568
rect 4445 309508 4449 309564
rect 4449 309508 4505 309564
rect 4505 309508 4509 309564
rect 4445 309504 4509 309508
rect 4525 309564 4589 309568
rect 4525 309508 4529 309564
rect 4529 309508 4585 309564
rect 4585 309508 4589 309564
rect 4525 309504 4589 309508
rect 7618 309564 7682 309568
rect 7618 309508 7622 309564
rect 7622 309508 7678 309564
rect 7678 309508 7682 309564
rect 7618 309504 7682 309508
rect 7698 309564 7762 309568
rect 7698 309508 7702 309564
rect 7702 309508 7758 309564
rect 7758 309508 7762 309564
rect 7698 309504 7762 309508
rect 7778 309564 7842 309568
rect 7778 309508 7782 309564
rect 7782 309508 7838 309564
rect 7838 309508 7842 309564
rect 7778 309504 7842 309508
rect 7858 309564 7922 309568
rect 7858 309508 7862 309564
rect 7862 309508 7918 309564
rect 7918 309508 7922 309564
rect 7858 309504 7922 309508
rect 2618 309020 2682 309024
rect 2618 308964 2622 309020
rect 2622 308964 2678 309020
rect 2678 308964 2682 309020
rect 2618 308960 2682 308964
rect 2698 309020 2762 309024
rect 2698 308964 2702 309020
rect 2702 308964 2758 309020
rect 2758 308964 2762 309020
rect 2698 308960 2762 308964
rect 2778 309020 2842 309024
rect 2778 308964 2782 309020
rect 2782 308964 2838 309020
rect 2838 308964 2842 309020
rect 2778 308960 2842 308964
rect 2858 309020 2922 309024
rect 2858 308964 2862 309020
rect 2862 308964 2918 309020
rect 2918 308964 2922 309020
rect 2858 308960 2922 308964
rect 5952 309020 6016 309024
rect 5952 308964 5956 309020
rect 5956 308964 6012 309020
rect 6012 308964 6016 309020
rect 5952 308960 6016 308964
rect 6032 309020 6096 309024
rect 6032 308964 6036 309020
rect 6036 308964 6092 309020
rect 6092 308964 6096 309020
rect 6032 308960 6096 308964
rect 6112 309020 6176 309024
rect 6112 308964 6116 309020
rect 6116 308964 6172 309020
rect 6172 308964 6176 309020
rect 6112 308960 6176 308964
rect 6192 309020 6256 309024
rect 6192 308964 6196 309020
rect 6196 308964 6252 309020
rect 6252 308964 6256 309020
rect 6192 308960 6256 308964
rect 4285 308476 4349 308480
rect 4285 308420 4289 308476
rect 4289 308420 4345 308476
rect 4345 308420 4349 308476
rect 4285 308416 4349 308420
rect 4365 308476 4429 308480
rect 4365 308420 4369 308476
rect 4369 308420 4425 308476
rect 4425 308420 4429 308476
rect 4365 308416 4429 308420
rect 4445 308476 4509 308480
rect 4445 308420 4449 308476
rect 4449 308420 4505 308476
rect 4505 308420 4509 308476
rect 4445 308416 4509 308420
rect 4525 308476 4589 308480
rect 4525 308420 4529 308476
rect 4529 308420 4585 308476
rect 4585 308420 4589 308476
rect 4525 308416 4589 308420
rect 7618 308476 7682 308480
rect 7618 308420 7622 308476
rect 7622 308420 7678 308476
rect 7678 308420 7682 308476
rect 7618 308416 7682 308420
rect 7698 308476 7762 308480
rect 7698 308420 7702 308476
rect 7702 308420 7758 308476
rect 7758 308420 7762 308476
rect 7698 308416 7762 308420
rect 7778 308476 7842 308480
rect 7778 308420 7782 308476
rect 7782 308420 7838 308476
rect 7838 308420 7842 308476
rect 7778 308416 7842 308420
rect 7858 308476 7922 308480
rect 7858 308420 7862 308476
rect 7862 308420 7918 308476
rect 7918 308420 7922 308476
rect 7858 308416 7922 308420
rect 2618 307932 2682 307936
rect 2618 307876 2622 307932
rect 2622 307876 2678 307932
rect 2678 307876 2682 307932
rect 2618 307872 2682 307876
rect 2698 307932 2762 307936
rect 2698 307876 2702 307932
rect 2702 307876 2758 307932
rect 2758 307876 2762 307932
rect 2698 307872 2762 307876
rect 2778 307932 2842 307936
rect 2778 307876 2782 307932
rect 2782 307876 2838 307932
rect 2838 307876 2842 307932
rect 2778 307872 2842 307876
rect 2858 307932 2922 307936
rect 2858 307876 2862 307932
rect 2862 307876 2918 307932
rect 2918 307876 2922 307932
rect 2858 307872 2922 307876
rect 5952 307932 6016 307936
rect 5952 307876 5956 307932
rect 5956 307876 6012 307932
rect 6012 307876 6016 307932
rect 5952 307872 6016 307876
rect 6032 307932 6096 307936
rect 6032 307876 6036 307932
rect 6036 307876 6092 307932
rect 6092 307876 6096 307932
rect 6032 307872 6096 307876
rect 6112 307932 6176 307936
rect 6112 307876 6116 307932
rect 6116 307876 6172 307932
rect 6172 307876 6176 307932
rect 6112 307872 6176 307876
rect 6192 307932 6256 307936
rect 6192 307876 6196 307932
rect 6196 307876 6252 307932
rect 6252 307876 6256 307932
rect 6192 307872 6256 307876
rect 4285 307388 4349 307392
rect 4285 307332 4289 307388
rect 4289 307332 4345 307388
rect 4345 307332 4349 307388
rect 4285 307328 4349 307332
rect 4365 307388 4429 307392
rect 4365 307332 4369 307388
rect 4369 307332 4425 307388
rect 4425 307332 4429 307388
rect 4365 307328 4429 307332
rect 4445 307388 4509 307392
rect 4445 307332 4449 307388
rect 4449 307332 4505 307388
rect 4505 307332 4509 307388
rect 4445 307328 4509 307332
rect 4525 307388 4589 307392
rect 4525 307332 4529 307388
rect 4529 307332 4585 307388
rect 4585 307332 4589 307388
rect 4525 307328 4589 307332
rect 7618 307388 7682 307392
rect 7618 307332 7622 307388
rect 7622 307332 7678 307388
rect 7678 307332 7682 307388
rect 7618 307328 7682 307332
rect 7698 307388 7762 307392
rect 7698 307332 7702 307388
rect 7702 307332 7758 307388
rect 7758 307332 7762 307388
rect 7698 307328 7762 307332
rect 7778 307388 7842 307392
rect 7778 307332 7782 307388
rect 7782 307332 7838 307388
rect 7838 307332 7842 307388
rect 7778 307328 7842 307332
rect 7858 307388 7922 307392
rect 7858 307332 7862 307388
rect 7862 307332 7918 307388
rect 7918 307332 7922 307388
rect 7858 307328 7922 307332
rect 2618 306844 2682 306848
rect 2618 306788 2622 306844
rect 2622 306788 2678 306844
rect 2678 306788 2682 306844
rect 2618 306784 2682 306788
rect 2698 306844 2762 306848
rect 2698 306788 2702 306844
rect 2702 306788 2758 306844
rect 2758 306788 2762 306844
rect 2698 306784 2762 306788
rect 2778 306844 2842 306848
rect 2778 306788 2782 306844
rect 2782 306788 2838 306844
rect 2838 306788 2842 306844
rect 2778 306784 2842 306788
rect 2858 306844 2922 306848
rect 2858 306788 2862 306844
rect 2862 306788 2918 306844
rect 2918 306788 2922 306844
rect 2858 306784 2922 306788
rect 5952 306844 6016 306848
rect 5952 306788 5956 306844
rect 5956 306788 6012 306844
rect 6012 306788 6016 306844
rect 5952 306784 6016 306788
rect 6032 306844 6096 306848
rect 6032 306788 6036 306844
rect 6036 306788 6092 306844
rect 6092 306788 6096 306844
rect 6032 306784 6096 306788
rect 6112 306844 6176 306848
rect 6112 306788 6116 306844
rect 6116 306788 6172 306844
rect 6172 306788 6176 306844
rect 6112 306784 6176 306788
rect 6192 306844 6256 306848
rect 6192 306788 6196 306844
rect 6196 306788 6252 306844
rect 6252 306788 6256 306844
rect 6192 306784 6256 306788
rect 4285 306300 4349 306304
rect 4285 306244 4289 306300
rect 4289 306244 4345 306300
rect 4345 306244 4349 306300
rect 4285 306240 4349 306244
rect 4365 306300 4429 306304
rect 4365 306244 4369 306300
rect 4369 306244 4425 306300
rect 4425 306244 4429 306300
rect 4365 306240 4429 306244
rect 4445 306300 4509 306304
rect 4445 306244 4449 306300
rect 4449 306244 4505 306300
rect 4505 306244 4509 306300
rect 4445 306240 4509 306244
rect 4525 306300 4589 306304
rect 4525 306244 4529 306300
rect 4529 306244 4585 306300
rect 4585 306244 4589 306300
rect 4525 306240 4589 306244
rect 7618 306300 7682 306304
rect 7618 306244 7622 306300
rect 7622 306244 7678 306300
rect 7678 306244 7682 306300
rect 7618 306240 7682 306244
rect 7698 306300 7762 306304
rect 7698 306244 7702 306300
rect 7702 306244 7758 306300
rect 7758 306244 7762 306300
rect 7698 306240 7762 306244
rect 7778 306300 7842 306304
rect 7778 306244 7782 306300
rect 7782 306244 7838 306300
rect 7838 306244 7842 306300
rect 7778 306240 7842 306244
rect 7858 306300 7922 306304
rect 7858 306244 7862 306300
rect 7862 306244 7918 306300
rect 7918 306244 7922 306300
rect 7858 306240 7922 306244
rect 2618 305756 2682 305760
rect 2618 305700 2622 305756
rect 2622 305700 2678 305756
rect 2678 305700 2682 305756
rect 2618 305696 2682 305700
rect 2698 305756 2762 305760
rect 2698 305700 2702 305756
rect 2702 305700 2758 305756
rect 2758 305700 2762 305756
rect 2698 305696 2762 305700
rect 2778 305756 2842 305760
rect 2778 305700 2782 305756
rect 2782 305700 2838 305756
rect 2838 305700 2842 305756
rect 2778 305696 2842 305700
rect 2858 305756 2922 305760
rect 2858 305700 2862 305756
rect 2862 305700 2918 305756
rect 2918 305700 2922 305756
rect 2858 305696 2922 305700
rect 5952 305756 6016 305760
rect 5952 305700 5956 305756
rect 5956 305700 6012 305756
rect 6012 305700 6016 305756
rect 5952 305696 6016 305700
rect 6032 305756 6096 305760
rect 6032 305700 6036 305756
rect 6036 305700 6092 305756
rect 6092 305700 6096 305756
rect 6032 305696 6096 305700
rect 6112 305756 6176 305760
rect 6112 305700 6116 305756
rect 6116 305700 6172 305756
rect 6172 305700 6176 305756
rect 6112 305696 6176 305700
rect 6192 305756 6256 305760
rect 6192 305700 6196 305756
rect 6196 305700 6252 305756
rect 6252 305700 6256 305756
rect 6192 305696 6256 305700
rect 4285 305212 4349 305216
rect 4285 305156 4289 305212
rect 4289 305156 4345 305212
rect 4345 305156 4349 305212
rect 4285 305152 4349 305156
rect 4365 305212 4429 305216
rect 4365 305156 4369 305212
rect 4369 305156 4425 305212
rect 4425 305156 4429 305212
rect 4365 305152 4429 305156
rect 4445 305212 4509 305216
rect 4445 305156 4449 305212
rect 4449 305156 4505 305212
rect 4505 305156 4509 305212
rect 4445 305152 4509 305156
rect 4525 305212 4589 305216
rect 4525 305156 4529 305212
rect 4529 305156 4585 305212
rect 4585 305156 4589 305212
rect 4525 305152 4589 305156
rect 7618 305212 7682 305216
rect 7618 305156 7622 305212
rect 7622 305156 7678 305212
rect 7678 305156 7682 305212
rect 7618 305152 7682 305156
rect 7698 305212 7762 305216
rect 7698 305156 7702 305212
rect 7702 305156 7758 305212
rect 7758 305156 7762 305212
rect 7698 305152 7762 305156
rect 7778 305212 7842 305216
rect 7778 305156 7782 305212
rect 7782 305156 7838 305212
rect 7838 305156 7842 305212
rect 7778 305152 7842 305156
rect 7858 305212 7922 305216
rect 7858 305156 7862 305212
rect 7862 305156 7918 305212
rect 7918 305156 7922 305212
rect 7858 305152 7922 305156
rect 2618 304668 2682 304672
rect 2618 304612 2622 304668
rect 2622 304612 2678 304668
rect 2678 304612 2682 304668
rect 2618 304608 2682 304612
rect 2698 304668 2762 304672
rect 2698 304612 2702 304668
rect 2702 304612 2758 304668
rect 2758 304612 2762 304668
rect 2698 304608 2762 304612
rect 2778 304668 2842 304672
rect 2778 304612 2782 304668
rect 2782 304612 2838 304668
rect 2838 304612 2842 304668
rect 2778 304608 2842 304612
rect 2858 304668 2922 304672
rect 2858 304612 2862 304668
rect 2862 304612 2918 304668
rect 2918 304612 2922 304668
rect 2858 304608 2922 304612
rect 5952 304668 6016 304672
rect 5952 304612 5956 304668
rect 5956 304612 6012 304668
rect 6012 304612 6016 304668
rect 5952 304608 6016 304612
rect 6032 304668 6096 304672
rect 6032 304612 6036 304668
rect 6036 304612 6092 304668
rect 6092 304612 6096 304668
rect 6032 304608 6096 304612
rect 6112 304668 6176 304672
rect 6112 304612 6116 304668
rect 6116 304612 6172 304668
rect 6172 304612 6176 304668
rect 6112 304608 6176 304612
rect 6192 304668 6256 304672
rect 6192 304612 6196 304668
rect 6196 304612 6252 304668
rect 6252 304612 6256 304668
rect 6192 304608 6256 304612
rect 4285 304124 4349 304128
rect 4285 304068 4289 304124
rect 4289 304068 4345 304124
rect 4345 304068 4349 304124
rect 4285 304064 4349 304068
rect 4365 304124 4429 304128
rect 4365 304068 4369 304124
rect 4369 304068 4425 304124
rect 4425 304068 4429 304124
rect 4365 304064 4429 304068
rect 4445 304124 4509 304128
rect 4445 304068 4449 304124
rect 4449 304068 4505 304124
rect 4505 304068 4509 304124
rect 4445 304064 4509 304068
rect 4525 304124 4589 304128
rect 4525 304068 4529 304124
rect 4529 304068 4585 304124
rect 4585 304068 4589 304124
rect 4525 304064 4589 304068
rect 7618 304124 7682 304128
rect 7618 304068 7622 304124
rect 7622 304068 7678 304124
rect 7678 304068 7682 304124
rect 7618 304064 7682 304068
rect 7698 304124 7762 304128
rect 7698 304068 7702 304124
rect 7702 304068 7758 304124
rect 7758 304068 7762 304124
rect 7698 304064 7762 304068
rect 7778 304124 7842 304128
rect 7778 304068 7782 304124
rect 7782 304068 7838 304124
rect 7838 304068 7842 304124
rect 7778 304064 7842 304068
rect 7858 304124 7922 304128
rect 7858 304068 7862 304124
rect 7862 304068 7918 304124
rect 7918 304068 7922 304124
rect 7858 304064 7922 304068
rect 2618 303580 2682 303584
rect 2618 303524 2622 303580
rect 2622 303524 2678 303580
rect 2678 303524 2682 303580
rect 2618 303520 2682 303524
rect 2698 303580 2762 303584
rect 2698 303524 2702 303580
rect 2702 303524 2758 303580
rect 2758 303524 2762 303580
rect 2698 303520 2762 303524
rect 2778 303580 2842 303584
rect 2778 303524 2782 303580
rect 2782 303524 2838 303580
rect 2838 303524 2842 303580
rect 2778 303520 2842 303524
rect 2858 303580 2922 303584
rect 2858 303524 2862 303580
rect 2862 303524 2918 303580
rect 2918 303524 2922 303580
rect 2858 303520 2922 303524
rect 5952 303580 6016 303584
rect 5952 303524 5956 303580
rect 5956 303524 6012 303580
rect 6012 303524 6016 303580
rect 5952 303520 6016 303524
rect 6032 303580 6096 303584
rect 6032 303524 6036 303580
rect 6036 303524 6092 303580
rect 6092 303524 6096 303580
rect 6032 303520 6096 303524
rect 6112 303580 6176 303584
rect 6112 303524 6116 303580
rect 6116 303524 6172 303580
rect 6172 303524 6176 303580
rect 6112 303520 6176 303524
rect 6192 303580 6256 303584
rect 6192 303524 6196 303580
rect 6196 303524 6252 303580
rect 6252 303524 6256 303580
rect 6192 303520 6256 303524
rect 4285 303036 4349 303040
rect 4285 302980 4289 303036
rect 4289 302980 4345 303036
rect 4345 302980 4349 303036
rect 4285 302976 4349 302980
rect 4365 303036 4429 303040
rect 4365 302980 4369 303036
rect 4369 302980 4425 303036
rect 4425 302980 4429 303036
rect 4365 302976 4429 302980
rect 4445 303036 4509 303040
rect 4445 302980 4449 303036
rect 4449 302980 4505 303036
rect 4505 302980 4509 303036
rect 4445 302976 4509 302980
rect 4525 303036 4589 303040
rect 4525 302980 4529 303036
rect 4529 302980 4585 303036
rect 4585 302980 4589 303036
rect 4525 302976 4589 302980
rect 7618 303036 7682 303040
rect 7618 302980 7622 303036
rect 7622 302980 7678 303036
rect 7678 302980 7682 303036
rect 7618 302976 7682 302980
rect 7698 303036 7762 303040
rect 7698 302980 7702 303036
rect 7702 302980 7758 303036
rect 7758 302980 7762 303036
rect 7698 302976 7762 302980
rect 7778 303036 7842 303040
rect 7778 302980 7782 303036
rect 7782 302980 7838 303036
rect 7838 302980 7842 303036
rect 7778 302976 7842 302980
rect 7858 303036 7922 303040
rect 7858 302980 7862 303036
rect 7862 302980 7918 303036
rect 7918 302980 7922 303036
rect 7858 302976 7922 302980
rect 2618 302492 2682 302496
rect 2618 302436 2622 302492
rect 2622 302436 2678 302492
rect 2678 302436 2682 302492
rect 2618 302432 2682 302436
rect 2698 302492 2762 302496
rect 2698 302436 2702 302492
rect 2702 302436 2758 302492
rect 2758 302436 2762 302492
rect 2698 302432 2762 302436
rect 2778 302492 2842 302496
rect 2778 302436 2782 302492
rect 2782 302436 2838 302492
rect 2838 302436 2842 302492
rect 2778 302432 2842 302436
rect 2858 302492 2922 302496
rect 2858 302436 2862 302492
rect 2862 302436 2918 302492
rect 2918 302436 2922 302492
rect 2858 302432 2922 302436
rect 5952 302492 6016 302496
rect 5952 302436 5956 302492
rect 5956 302436 6012 302492
rect 6012 302436 6016 302492
rect 5952 302432 6016 302436
rect 6032 302492 6096 302496
rect 6032 302436 6036 302492
rect 6036 302436 6092 302492
rect 6092 302436 6096 302492
rect 6032 302432 6096 302436
rect 6112 302492 6176 302496
rect 6112 302436 6116 302492
rect 6116 302436 6172 302492
rect 6172 302436 6176 302492
rect 6112 302432 6176 302436
rect 6192 302492 6256 302496
rect 6192 302436 6196 302492
rect 6196 302436 6252 302492
rect 6252 302436 6256 302492
rect 6192 302432 6256 302436
rect 4285 301948 4349 301952
rect 4285 301892 4289 301948
rect 4289 301892 4345 301948
rect 4345 301892 4349 301948
rect 4285 301888 4349 301892
rect 4365 301948 4429 301952
rect 4365 301892 4369 301948
rect 4369 301892 4425 301948
rect 4425 301892 4429 301948
rect 4365 301888 4429 301892
rect 4445 301948 4509 301952
rect 4445 301892 4449 301948
rect 4449 301892 4505 301948
rect 4505 301892 4509 301948
rect 4445 301888 4509 301892
rect 4525 301948 4589 301952
rect 4525 301892 4529 301948
rect 4529 301892 4585 301948
rect 4585 301892 4589 301948
rect 4525 301888 4589 301892
rect 7618 301948 7682 301952
rect 7618 301892 7622 301948
rect 7622 301892 7678 301948
rect 7678 301892 7682 301948
rect 7618 301888 7682 301892
rect 7698 301948 7762 301952
rect 7698 301892 7702 301948
rect 7702 301892 7758 301948
rect 7758 301892 7762 301948
rect 7698 301888 7762 301892
rect 7778 301948 7842 301952
rect 7778 301892 7782 301948
rect 7782 301892 7838 301948
rect 7838 301892 7842 301948
rect 7778 301888 7842 301892
rect 7858 301948 7922 301952
rect 7858 301892 7862 301948
rect 7862 301892 7918 301948
rect 7918 301892 7922 301948
rect 7858 301888 7922 301892
rect 2618 301404 2682 301408
rect 2618 301348 2622 301404
rect 2622 301348 2678 301404
rect 2678 301348 2682 301404
rect 2618 301344 2682 301348
rect 2698 301404 2762 301408
rect 2698 301348 2702 301404
rect 2702 301348 2758 301404
rect 2758 301348 2762 301404
rect 2698 301344 2762 301348
rect 2778 301404 2842 301408
rect 2778 301348 2782 301404
rect 2782 301348 2838 301404
rect 2838 301348 2842 301404
rect 2778 301344 2842 301348
rect 2858 301404 2922 301408
rect 2858 301348 2862 301404
rect 2862 301348 2918 301404
rect 2918 301348 2922 301404
rect 2858 301344 2922 301348
rect 5952 301404 6016 301408
rect 5952 301348 5956 301404
rect 5956 301348 6012 301404
rect 6012 301348 6016 301404
rect 5952 301344 6016 301348
rect 6032 301404 6096 301408
rect 6032 301348 6036 301404
rect 6036 301348 6092 301404
rect 6092 301348 6096 301404
rect 6032 301344 6096 301348
rect 6112 301404 6176 301408
rect 6112 301348 6116 301404
rect 6116 301348 6172 301404
rect 6172 301348 6176 301404
rect 6112 301344 6176 301348
rect 6192 301404 6256 301408
rect 6192 301348 6196 301404
rect 6196 301348 6252 301404
rect 6252 301348 6256 301404
rect 6192 301344 6256 301348
rect 4285 300860 4349 300864
rect 4285 300804 4289 300860
rect 4289 300804 4345 300860
rect 4345 300804 4349 300860
rect 4285 300800 4349 300804
rect 4365 300860 4429 300864
rect 4365 300804 4369 300860
rect 4369 300804 4425 300860
rect 4425 300804 4429 300860
rect 4365 300800 4429 300804
rect 4445 300860 4509 300864
rect 4445 300804 4449 300860
rect 4449 300804 4505 300860
rect 4505 300804 4509 300860
rect 4445 300800 4509 300804
rect 4525 300860 4589 300864
rect 4525 300804 4529 300860
rect 4529 300804 4585 300860
rect 4585 300804 4589 300860
rect 4525 300800 4589 300804
rect 7618 300860 7682 300864
rect 7618 300804 7622 300860
rect 7622 300804 7678 300860
rect 7678 300804 7682 300860
rect 7618 300800 7682 300804
rect 7698 300860 7762 300864
rect 7698 300804 7702 300860
rect 7702 300804 7758 300860
rect 7758 300804 7762 300860
rect 7698 300800 7762 300804
rect 7778 300860 7842 300864
rect 7778 300804 7782 300860
rect 7782 300804 7838 300860
rect 7838 300804 7842 300860
rect 7778 300800 7842 300804
rect 7858 300860 7922 300864
rect 7858 300804 7862 300860
rect 7862 300804 7918 300860
rect 7918 300804 7922 300860
rect 7858 300800 7922 300804
rect 2618 300316 2682 300320
rect 2618 300260 2622 300316
rect 2622 300260 2678 300316
rect 2678 300260 2682 300316
rect 2618 300256 2682 300260
rect 2698 300316 2762 300320
rect 2698 300260 2702 300316
rect 2702 300260 2758 300316
rect 2758 300260 2762 300316
rect 2698 300256 2762 300260
rect 2778 300316 2842 300320
rect 2778 300260 2782 300316
rect 2782 300260 2838 300316
rect 2838 300260 2842 300316
rect 2778 300256 2842 300260
rect 2858 300316 2922 300320
rect 2858 300260 2862 300316
rect 2862 300260 2918 300316
rect 2918 300260 2922 300316
rect 2858 300256 2922 300260
rect 5952 300316 6016 300320
rect 5952 300260 5956 300316
rect 5956 300260 6012 300316
rect 6012 300260 6016 300316
rect 5952 300256 6016 300260
rect 6032 300316 6096 300320
rect 6032 300260 6036 300316
rect 6036 300260 6092 300316
rect 6092 300260 6096 300316
rect 6032 300256 6096 300260
rect 6112 300316 6176 300320
rect 6112 300260 6116 300316
rect 6116 300260 6172 300316
rect 6172 300260 6176 300316
rect 6112 300256 6176 300260
rect 6192 300316 6256 300320
rect 6192 300260 6196 300316
rect 6196 300260 6252 300316
rect 6252 300260 6256 300316
rect 6192 300256 6256 300260
rect 4285 299772 4349 299776
rect 4285 299716 4289 299772
rect 4289 299716 4345 299772
rect 4345 299716 4349 299772
rect 4285 299712 4349 299716
rect 4365 299772 4429 299776
rect 4365 299716 4369 299772
rect 4369 299716 4425 299772
rect 4425 299716 4429 299772
rect 4365 299712 4429 299716
rect 4445 299772 4509 299776
rect 4445 299716 4449 299772
rect 4449 299716 4505 299772
rect 4505 299716 4509 299772
rect 4445 299712 4509 299716
rect 4525 299772 4589 299776
rect 4525 299716 4529 299772
rect 4529 299716 4585 299772
rect 4585 299716 4589 299772
rect 4525 299712 4589 299716
rect 7618 299772 7682 299776
rect 7618 299716 7622 299772
rect 7622 299716 7678 299772
rect 7678 299716 7682 299772
rect 7618 299712 7682 299716
rect 7698 299772 7762 299776
rect 7698 299716 7702 299772
rect 7702 299716 7758 299772
rect 7758 299716 7762 299772
rect 7698 299712 7762 299716
rect 7778 299772 7842 299776
rect 7778 299716 7782 299772
rect 7782 299716 7838 299772
rect 7838 299716 7842 299772
rect 7778 299712 7842 299716
rect 7858 299772 7922 299776
rect 7858 299716 7862 299772
rect 7862 299716 7918 299772
rect 7918 299716 7922 299772
rect 7858 299712 7922 299716
rect 2618 299228 2682 299232
rect 2618 299172 2622 299228
rect 2622 299172 2678 299228
rect 2678 299172 2682 299228
rect 2618 299168 2682 299172
rect 2698 299228 2762 299232
rect 2698 299172 2702 299228
rect 2702 299172 2758 299228
rect 2758 299172 2762 299228
rect 2698 299168 2762 299172
rect 2778 299228 2842 299232
rect 2778 299172 2782 299228
rect 2782 299172 2838 299228
rect 2838 299172 2842 299228
rect 2778 299168 2842 299172
rect 2858 299228 2922 299232
rect 2858 299172 2862 299228
rect 2862 299172 2918 299228
rect 2918 299172 2922 299228
rect 2858 299168 2922 299172
rect 5952 299228 6016 299232
rect 5952 299172 5956 299228
rect 5956 299172 6012 299228
rect 6012 299172 6016 299228
rect 5952 299168 6016 299172
rect 6032 299228 6096 299232
rect 6032 299172 6036 299228
rect 6036 299172 6092 299228
rect 6092 299172 6096 299228
rect 6032 299168 6096 299172
rect 6112 299228 6176 299232
rect 6112 299172 6116 299228
rect 6116 299172 6172 299228
rect 6172 299172 6176 299228
rect 6112 299168 6176 299172
rect 6192 299228 6256 299232
rect 6192 299172 6196 299228
rect 6196 299172 6252 299228
rect 6252 299172 6256 299228
rect 6192 299168 6256 299172
rect 4285 298684 4349 298688
rect 4285 298628 4289 298684
rect 4289 298628 4345 298684
rect 4345 298628 4349 298684
rect 4285 298624 4349 298628
rect 4365 298684 4429 298688
rect 4365 298628 4369 298684
rect 4369 298628 4425 298684
rect 4425 298628 4429 298684
rect 4365 298624 4429 298628
rect 4445 298684 4509 298688
rect 4445 298628 4449 298684
rect 4449 298628 4505 298684
rect 4505 298628 4509 298684
rect 4445 298624 4509 298628
rect 4525 298684 4589 298688
rect 4525 298628 4529 298684
rect 4529 298628 4585 298684
rect 4585 298628 4589 298684
rect 4525 298624 4589 298628
rect 7618 298684 7682 298688
rect 7618 298628 7622 298684
rect 7622 298628 7678 298684
rect 7678 298628 7682 298684
rect 7618 298624 7682 298628
rect 7698 298684 7762 298688
rect 7698 298628 7702 298684
rect 7702 298628 7758 298684
rect 7758 298628 7762 298684
rect 7698 298624 7762 298628
rect 7778 298684 7842 298688
rect 7778 298628 7782 298684
rect 7782 298628 7838 298684
rect 7838 298628 7842 298684
rect 7778 298624 7842 298628
rect 7858 298684 7922 298688
rect 7858 298628 7862 298684
rect 7862 298628 7918 298684
rect 7918 298628 7922 298684
rect 7858 298624 7922 298628
rect 2618 298140 2682 298144
rect 2618 298084 2622 298140
rect 2622 298084 2678 298140
rect 2678 298084 2682 298140
rect 2618 298080 2682 298084
rect 2698 298140 2762 298144
rect 2698 298084 2702 298140
rect 2702 298084 2758 298140
rect 2758 298084 2762 298140
rect 2698 298080 2762 298084
rect 2778 298140 2842 298144
rect 2778 298084 2782 298140
rect 2782 298084 2838 298140
rect 2838 298084 2842 298140
rect 2778 298080 2842 298084
rect 2858 298140 2922 298144
rect 2858 298084 2862 298140
rect 2862 298084 2918 298140
rect 2918 298084 2922 298140
rect 2858 298080 2922 298084
rect 5952 298140 6016 298144
rect 5952 298084 5956 298140
rect 5956 298084 6012 298140
rect 6012 298084 6016 298140
rect 5952 298080 6016 298084
rect 6032 298140 6096 298144
rect 6032 298084 6036 298140
rect 6036 298084 6092 298140
rect 6092 298084 6096 298140
rect 6032 298080 6096 298084
rect 6112 298140 6176 298144
rect 6112 298084 6116 298140
rect 6116 298084 6172 298140
rect 6172 298084 6176 298140
rect 6112 298080 6176 298084
rect 6192 298140 6256 298144
rect 6192 298084 6196 298140
rect 6196 298084 6252 298140
rect 6252 298084 6256 298140
rect 6192 298080 6256 298084
rect 4285 297596 4349 297600
rect 4285 297540 4289 297596
rect 4289 297540 4345 297596
rect 4345 297540 4349 297596
rect 4285 297536 4349 297540
rect 4365 297596 4429 297600
rect 4365 297540 4369 297596
rect 4369 297540 4425 297596
rect 4425 297540 4429 297596
rect 4365 297536 4429 297540
rect 4445 297596 4509 297600
rect 4445 297540 4449 297596
rect 4449 297540 4505 297596
rect 4505 297540 4509 297596
rect 4445 297536 4509 297540
rect 4525 297596 4589 297600
rect 4525 297540 4529 297596
rect 4529 297540 4585 297596
rect 4585 297540 4589 297596
rect 4525 297536 4589 297540
rect 7618 297596 7682 297600
rect 7618 297540 7622 297596
rect 7622 297540 7678 297596
rect 7678 297540 7682 297596
rect 7618 297536 7682 297540
rect 7698 297596 7762 297600
rect 7698 297540 7702 297596
rect 7702 297540 7758 297596
rect 7758 297540 7762 297596
rect 7698 297536 7762 297540
rect 7778 297596 7842 297600
rect 7778 297540 7782 297596
rect 7782 297540 7838 297596
rect 7838 297540 7842 297596
rect 7778 297536 7842 297540
rect 7858 297596 7922 297600
rect 7858 297540 7862 297596
rect 7862 297540 7918 297596
rect 7918 297540 7922 297596
rect 7858 297536 7922 297540
rect 2618 297052 2682 297056
rect 2618 296996 2622 297052
rect 2622 296996 2678 297052
rect 2678 296996 2682 297052
rect 2618 296992 2682 296996
rect 2698 297052 2762 297056
rect 2698 296996 2702 297052
rect 2702 296996 2758 297052
rect 2758 296996 2762 297052
rect 2698 296992 2762 296996
rect 2778 297052 2842 297056
rect 2778 296996 2782 297052
rect 2782 296996 2838 297052
rect 2838 296996 2842 297052
rect 2778 296992 2842 296996
rect 2858 297052 2922 297056
rect 2858 296996 2862 297052
rect 2862 296996 2918 297052
rect 2918 296996 2922 297052
rect 2858 296992 2922 296996
rect 5952 297052 6016 297056
rect 5952 296996 5956 297052
rect 5956 296996 6012 297052
rect 6012 296996 6016 297052
rect 5952 296992 6016 296996
rect 6032 297052 6096 297056
rect 6032 296996 6036 297052
rect 6036 296996 6092 297052
rect 6092 296996 6096 297052
rect 6032 296992 6096 296996
rect 6112 297052 6176 297056
rect 6112 296996 6116 297052
rect 6116 296996 6172 297052
rect 6172 296996 6176 297052
rect 6112 296992 6176 296996
rect 6192 297052 6256 297056
rect 6192 296996 6196 297052
rect 6196 296996 6252 297052
rect 6252 296996 6256 297052
rect 6192 296992 6256 296996
rect 4285 296508 4349 296512
rect 4285 296452 4289 296508
rect 4289 296452 4345 296508
rect 4345 296452 4349 296508
rect 4285 296448 4349 296452
rect 4365 296508 4429 296512
rect 4365 296452 4369 296508
rect 4369 296452 4425 296508
rect 4425 296452 4429 296508
rect 4365 296448 4429 296452
rect 4445 296508 4509 296512
rect 4445 296452 4449 296508
rect 4449 296452 4505 296508
rect 4505 296452 4509 296508
rect 4445 296448 4509 296452
rect 4525 296508 4589 296512
rect 4525 296452 4529 296508
rect 4529 296452 4585 296508
rect 4585 296452 4589 296508
rect 4525 296448 4589 296452
rect 7618 296508 7682 296512
rect 7618 296452 7622 296508
rect 7622 296452 7678 296508
rect 7678 296452 7682 296508
rect 7618 296448 7682 296452
rect 7698 296508 7762 296512
rect 7698 296452 7702 296508
rect 7702 296452 7758 296508
rect 7758 296452 7762 296508
rect 7698 296448 7762 296452
rect 7778 296508 7842 296512
rect 7778 296452 7782 296508
rect 7782 296452 7838 296508
rect 7838 296452 7842 296508
rect 7778 296448 7842 296452
rect 7858 296508 7922 296512
rect 7858 296452 7862 296508
rect 7862 296452 7918 296508
rect 7918 296452 7922 296508
rect 7858 296448 7922 296452
rect 2618 295964 2682 295968
rect 2618 295908 2622 295964
rect 2622 295908 2678 295964
rect 2678 295908 2682 295964
rect 2618 295904 2682 295908
rect 2698 295964 2762 295968
rect 2698 295908 2702 295964
rect 2702 295908 2758 295964
rect 2758 295908 2762 295964
rect 2698 295904 2762 295908
rect 2778 295964 2842 295968
rect 2778 295908 2782 295964
rect 2782 295908 2838 295964
rect 2838 295908 2842 295964
rect 2778 295904 2842 295908
rect 2858 295964 2922 295968
rect 2858 295908 2862 295964
rect 2862 295908 2918 295964
rect 2918 295908 2922 295964
rect 2858 295904 2922 295908
rect 5952 295964 6016 295968
rect 5952 295908 5956 295964
rect 5956 295908 6012 295964
rect 6012 295908 6016 295964
rect 5952 295904 6016 295908
rect 6032 295964 6096 295968
rect 6032 295908 6036 295964
rect 6036 295908 6092 295964
rect 6092 295908 6096 295964
rect 6032 295904 6096 295908
rect 6112 295964 6176 295968
rect 6112 295908 6116 295964
rect 6116 295908 6172 295964
rect 6172 295908 6176 295964
rect 6112 295904 6176 295908
rect 6192 295964 6256 295968
rect 6192 295908 6196 295964
rect 6196 295908 6252 295964
rect 6252 295908 6256 295964
rect 6192 295904 6256 295908
rect 4285 295420 4349 295424
rect 4285 295364 4289 295420
rect 4289 295364 4345 295420
rect 4345 295364 4349 295420
rect 4285 295360 4349 295364
rect 4365 295420 4429 295424
rect 4365 295364 4369 295420
rect 4369 295364 4425 295420
rect 4425 295364 4429 295420
rect 4365 295360 4429 295364
rect 4445 295420 4509 295424
rect 4445 295364 4449 295420
rect 4449 295364 4505 295420
rect 4505 295364 4509 295420
rect 4445 295360 4509 295364
rect 4525 295420 4589 295424
rect 4525 295364 4529 295420
rect 4529 295364 4585 295420
rect 4585 295364 4589 295420
rect 4525 295360 4589 295364
rect 7618 295420 7682 295424
rect 7618 295364 7622 295420
rect 7622 295364 7678 295420
rect 7678 295364 7682 295420
rect 7618 295360 7682 295364
rect 7698 295420 7762 295424
rect 7698 295364 7702 295420
rect 7702 295364 7758 295420
rect 7758 295364 7762 295420
rect 7698 295360 7762 295364
rect 7778 295420 7842 295424
rect 7778 295364 7782 295420
rect 7782 295364 7838 295420
rect 7838 295364 7842 295420
rect 7778 295360 7842 295364
rect 7858 295420 7922 295424
rect 7858 295364 7862 295420
rect 7862 295364 7918 295420
rect 7918 295364 7922 295420
rect 7858 295360 7922 295364
rect 2618 294876 2682 294880
rect 2618 294820 2622 294876
rect 2622 294820 2678 294876
rect 2678 294820 2682 294876
rect 2618 294816 2682 294820
rect 2698 294876 2762 294880
rect 2698 294820 2702 294876
rect 2702 294820 2758 294876
rect 2758 294820 2762 294876
rect 2698 294816 2762 294820
rect 2778 294876 2842 294880
rect 2778 294820 2782 294876
rect 2782 294820 2838 294876
rect 2838 294820 2842 294876
rect 2778 294816 2842 294820
rect 2858 294876 2922 294880
rect 2858 294820 2862 294876
rect 2862 294820 2918 294876
rect 2918 294820 2922 294876
rect 2858 294816 2922 294820
rect 5952 294876 6016 294880
rect 5952 294820 5956 294876
rect 5956 294820 6012 294876
rect 6012 294820 6016 294876
rect 5952 294816 6016 294820
rect 6032 294876 6096 294880
rect 6032 294820 6036 294876
rect 6036 294820 6092 294876
rect 6092 294820 6096 294876
rect 6032 294816 6096 294820
rect 6112 294876 6176 294880
rect 6112 294820 6116 294876
rect 6116 294820 6172 294876
rect 6172 294820 6176 294876
rect 6112 294816 6176 294820
rect 6192 294876 6256 294880
rect 6192 294820 6196 294876
rect 6196 294820 6252 294876
rect 6252 294820 6256 294876
rect 6192 294816 6256 294820
rect 4285 294332 4349 294336
rect 4285 294276 4289 294332
rect 4289 294276 4345 294332
rect 4345 294276 4349 294332
rect 4285 294272 4349 294276
rect 4365 294332 4429 294336
rect 4365 294276 4369 294332
rect 4369 294276 4425 294332
rect 4425 294276 4429 294332
rect 4365 294272 4429 294276
rect 4445 294332 4509 294336
rect 4445 294276 4449 294332
rect 4449 294276 4505 294332
rect 4505 294276 4509 294332
rect 4445 294272 4509 294276
rect 4525 294332 4589 294336
rect 4525 294276 4529 294332
rect 4529 294276 4585 294332
rect 4585 294276 4589 294332
rect 4525 294272 4589 294276
rect 7618 294332 7682 294336
rect 7618 294276 7622 294332
rect 7622 294276 7678 294332
rect 7678 294276 7682 294332
rect 7618 294272 7682 294276
rect 7698 294332 7762 294336
rect 7698 294276 7702 294332
rect 7702 294276 7758 294332
rect 7758 294276 7762 294332
rect 7698 294272 7762 294276
rect 7778 294332 7842 294336
rect 7778 294276 7782 294332
rect 7782 294276 7838 294332
rect 7838 294276 7842 294332
rect 7778 294272 7842 294276
rect 7858 294332 7922 294336
rect 7858 294276 7862 294332
rect 7862 294276 7918 294332
rect 7918 294276 7922 294332
rect 7858 294272 7922 294276
rect 2618 293788 2682 293792
rect 2618 293732 2622 293788
rect 2622 293732 2678 293788
rect 2678 293732 2682 293788
rect 2618 293728 2682 293732
rect 2698 293788 2762 293792
rect 2698 293732 2702 293788
rect 2702 293732 2758 293788
rect 2758 293732 2762 293788
rect 2698 293728 2762 293732
rect 2778 293788 2842 293792
rect 2778 293732 2782 293788
rect 2782 293732 2838 293788
rect 2838 293732 2842 293788
rect 2778 293728 2842 293732
rect 2858 293788 2922 293792
rect 2858 293732 2862 293788
rect 2862 293732 2918 293788
rect 2918 293732 2922 293788
rect 2858 293728 2922 293732
rect 5952 293788 6016 293792
rect 5952 293732 5956 293788
rect 5956 293732 6012 293788
rect 6012 293732 6016 293788
rect 5952 293728 6016 293732
rect 6032 293788 6096 293792
rect 6032 293732 6036 293788
rect 6036 293732 6092 293788
rect 6092 293732 6096 293788
rect 6032 293728 6096 293732
rect 6112 293788 6176 293792
rect 6112 293732 6116 293788
rect 6116 293732 6172 293788
rect 6172 293732 6176 293788
rect 6112 293728 6176 293732
rect 6192 293788 6256 293792
rect 6192 293732 6196 293788
rect 6196 293732 6252 293788
rect 6252 293732 6256 293788
rect 6192 293728 6256 293732
rect 4285 293244 4349 293248
rect 4285 293188 4289 293244
rect 4289 293188 4345 293244
rect 4345 293188 4349 293244
rect 4285 293184 4349 293188
rect 4365 293244 4429 293248
rect 4365 293188 4369 293244
rect 4369 293188 4425 293244
rect 4425 293188 4429 293244
rect 4365 293184 4429 293188
rect 4445 293244 4509 293248
rect 4445 293188 4449 293244
rect 4449 293188 4505 293244
rect 4505 293188 4509 293244
rect 4445 293184 4509 293188
rect 4525 293244 4589 293248
rect 4525 293188 4529 293244
rect 4529 293188 4585 293244
rect 4585 293188 4589 293244
rect 4525 293184 4589 293188
rect 7618 293244 7682 293248
rect 7618 293188 7622 293244
rect 7622 293188 7678 293244
rect 7678 293188 7682 293244
rect 7618 293184 7682 293188
rect 7698 293244 7762 293248
rect 7698 293188 7702 293244
rect 7702 293188 7758 293244
rect 7758 293188 7762 293244
rect 7698 293184 7762 293188
rect 7778 293244 7842 293248
rect 7778 293188 7782 293244
rect 7782 293188 7838 293244
rect 7838 293188 7842 293244
rect 7778 293184 7842 293188
rect 7858 293244 7922 293248
rect 7858 293188 7862 293244
rect 7862 293188 7918 293244
rect 7918 293188 7922 293244
rect 7858 293184 7922 293188
rect 2618 292700 2682 292704
rect 2618 292644 2622 292700
rect 2622 292644 2678 292700
rect 2678 292644 2682 292700
rect 2618 292640 2682 292644
rect 2698 292700 2762 292704
rect 2698 292644 2702 292700
rect 2702 292644 2758 292700
rect 2758 292644 2762 292700
rect 2698 292640 2762 292644
rect 2778 292700 2842 292704
rect 2778 292644 2782 292700
rect 2782 292644 2838 292700
rect 2838 292644 2842 292700
rect 2778 292640 2842 292644
rect 2858 292700 2922 292704
rect 2858 292644 2862 292700
rect 2862 292644 2918 292700
rect 2918 292644 2922 292700
rect 2858 292640 2922 292644
rect 5952 292700 6016 292704
rect 5952 292644 5956 292700
rect 5956 292644 6012 292700
rect 6012 292644 6016 292700
rect 5952 292640 6016 292644
rect 6032 292700 6096 292704
rect 6032 292644 6036 292700
rect 6036 292644 6092 292700
rect 6092 292644 6096 292700
rect 6032 292640 6096 292644
rect 6112 292700 6176 292704
rect 6112 292644 6116 292700
rect 6116 292644 6172 292700
rect 6172 292644 6176 292700
rect 6112 292640 6176 292644
rect 6192 292700 6256 292704
rect 6192 292644 6196 292700
rect 6196 292644 6252 292700
rect 6252 292644 6256 292700
rect 6192 292640 6256 292644
rect 4285 292156 4349 292160
rect 4285 292100 4289 292156
rect 4289 292100 4345 292156
rect 4345 292100 4349 292156
rect 4285 292096 4349 292100
rect 4365 292156 4429 292160
rect 4365 292100 4369 292156
rect 4369 292100 4425 292156
rect 4425 292100 4429 292156
rect 4365 292096 4429 292100
rect 4445 292156 4509 292160
rect 4445 292100 4449 292156
rect 4449 292100 4505 292156
rect 4505 292100 4509 292156
rect 4445 292096 4509 292100
rect 4525 292156 4589 292160
rect 4525 292100 4529 292156
rect 4529 292100 4585 292156
rect 4585 292100 4589 292156
rect 4525 292096 4589 292100
rect 7618 292156 7682 292160
rect 7618 292100 7622 292156
rect 7622 292100 7678 292156
rect 7678 292100 7682 292156
rect 7618 292096 7682 292100
rect 7698 292156 7762 292160
rect 7698 292100 7702 292156
rect 7702 292100 7758 292156
rect 7758 292100 7762 292156
rect 7698 292096 7762 292100
rect 7778 292156 7842 292160
rect 7778 292100 7782 292156
rect 7782 292100 7838 292156
rect 7838 292100 7842 292156
rect 7778 292096 7842 292100
rect 7858 292156 7922 292160
rect 7858 292100 7862 292156
rect 7862 292100 7918 292156
rect 7918 292100 7922 292156
rect 7858 292096 7922 292100
rect 2618 291612 2682 291616
rect 2618 291556 2622 291612
rect 2622 291556 2678 291612
rect 2678 291556 2682 291612
rect 2618 291552 2682 291556
rect 2698 291612 2762 291616
rect 2698 291556 2702 291612
rect 2702 291556 2758 291612
rect 2758 291556 2762 291612
rect 2698 291552 2762 291556
rect 2778 291612 2842 291616
rect 2778 291556 2782 291612
rect 2782 291556 2838 291612
rect 2838 291556 2842 291612
rect 2778 291552 2842 291556
rect 2858 291612 2922 291616
rect 2858 291556 2862 291612
rect 2862 291556 2918 291612
rect 2918 291556 2922 291612
rect 2858 291552 2922 291556
rect 5952 291612 6016 291616
rect 5952 291556 5956 291612
rect 5956 291556 6012 291612
rect 6012 291556 6016 291612
rect 5952 291552 6016 291556
rect 6032 291612 6096 291616
rect 6032 291556 6036 291612
rect 6036 291556 6092 291612
rect 6092 291556 6096 291612
rect 6032 291552 6096 291556
rect 6112 291612 6176 291616
rect 6112 291556 6116 291612
rect 6116 291556 6172 291612
rect 6172 291556 6176 291612
rect 6112 291552 6176 291556
rect 6192 291612 6256 291616
rect 6192 291556 6196 291612
rect 6196 291556 6252 291612
rect 6252 291556 6256 291612
rect 6192 291552 6256 291556
rect 4285 291068 4349 291072
rect 4285 291012 4289 291068
rect 4289 291012 4345 291068
rect 4345 291012 4349 291068
rect 4285 291008 4349 291012
rect 4365 291068 4429 291072
rect 4365 291012 4369 291068
rect 4369 291012 4425 291068
rect 4425 291012 4429 291068
rect 4365 291008 4429 291012
rect 4445 291068 4509 291072
rect 4445 291012 4449 291068
rect 4449 291012 4505 291068
rect 4505 291012 4509 291068
rect 4445 291008 4509 291012
rect 4525 291068 4589 291072
rect 4525 291012 4529 291068
rect 4529 291012 4585 291068
rect 4585 291012 4589 291068
rect 4525 291008 4589 291012
rect 7618 291068 7682 291072
rect 7618 291012 7622 291068
rect 7622 291012 7678 291068
rect 7678 291012 7682 291068
rect 7618 291008 7682 291012
rect 7698 291068 7762 291072
rect 7698 291012 7702 291068
rect 7702 291012 7758 291068
rect 7758 291012 7762 291068
rect 7698 291008 7762 291012
rect 7778 291068 7842 291072
rect 7778 291012 7782 291068
rect 7782 291012 7838 291068
rect 7838 291012 7842 291068
rect 7778 291008 7842 291012
rect 7858 291068 7922 291072
rect 7858 291012 7862 291068
rect 7862 291012 7918 291068
rect 7918 291012 7922 291068
rect 7858 291008 7922 291012
rect 2618 290524 2682 290528
rect 2618 290468 2622 290524
rect 2622 290468 2678 290524
rect 2678 290468 2682 290524
rect 2618 290464 2682 290468
rect 2698 290524 2762 290528
rect 2698 290468 2702 290524
rect 2702 290468 2758 290524
rect 2758 290468 2762 290524
rect 2698 290464 2762 290468
rect 2778 290524 2842 290528
rect 2778 290468 2782 290524
rect 2782 290468 2838 290524
rect 2838 290468 2842 290524
rect 2778 290464 2842 290468
rect 2858 290524 2922 290528
rect 2858 290468 2862 290524
rect 2862 290468 2918 290524
rect 2918 290468 2922 290524
rect 2858 290464 2922 290468
rect 5952 290524 6016 290528
rect 5952 290468 5956 290524
rect 5956 290468 6012 290524
rect 6012 290468 6016 290524
rect 5952 290464 6016 290468
rect 6032 290524 6096 290528
rect 6032 290468 6036 290524
rect 6036 290468 6092 290524
rect 6092 290468 6096 290524
rect 6032 290464 6096 290468
rect 6112 290524 6176 290528
rect 6112 290468 6116 290524
rect 6116 290468 6172 290524
rect 6172 290468 6176 290524
rect 6112 290464 6176 290468
rect 6192 290524 6256 290528
rect 6192 290468 6196 290524
rect 6196 290468 6252 290524
rect 6252 290468 6256 290524
rect 6192 290464 6256 290468
rect 4285 289980 4349 289984
rect 4285 289924 4289 289980
rect 4289 289924 4345 289980
rect 4345 289924 4349 289980
rect 4285 289920 4349 289924
rect 4365 289980 4429 289984
rect 4365 289924 4369 289980
rect 4369 289924 4425 289980
rect 4425 289924 4429 289980
rect 4365 289920 4429 289924
rect 4445 289980 4509 289984
rect 4445 289924 4449 289980
rect 4449 289924 4505 289980
rect 4505 289924 4509 289980
rect 4445 289920 4509 289924
rect 4525 289980 4589 289984
rect 4525 289924 4529 289980
rect 4529 289924 4585 289980
rect 4585 289924 4589 289980
rect 4525 289920 4589 289924
rect 7618 289980 7682 289984
rect 7618 289924 7622 289980
rect 7622 289924 7678 289980
rect 7678 289924 7682 289980
rect 7618 289920 7682 289924
rect 7698 289980 7762 289984
rect 7698 289924 7702 289980
rect 7702 289924 7758 289980
rect 7758 289924 7762 289980
rect 7698 289920 7762 289924
rect 7778 289980 7842 289984
rect 7778 289924 7782 289980
rect 7782 289924 7838 289980
rect 7838 289924 7842 289980
rect 7778 289920 7842 289924
rect 7858 289980 7922 289984
rect 7858 289924 7862 289980
rect 7862 289924 7918 289980
rect 7918 289924 7922 289980
rect 7858 289920 7922 289924
rect 2618 289436 2682 289440
rect 2618 289380 2622 289436
rect 2622 289380 2678 289436
rect 2678 289380 2682 289436
rect 2618 289376 2682 289380
rect 2698 289436 2762 289440
rect 2698 289380 2702 289436
rect 2702 289380 2758 289436
rect 2758 289380 2762 289436
rect 2698 289376 2762 289380
rect 2778 289436 2842 289440
rect 2778 289380 2782 289436
rect 2782 289380 2838 289436
rect 2838 289380 2842 289436
rect 2778 289376 2842 289380
rect 2858 289436 2922 289440
rect 2858 289380 2862 289436
rect 2862 289380 2918 289436
rect 2918 289380 2922 289436
rect 2858 289376 2922 289380
rect 5952 289436 6016 289440
rect 5952 289380 5956 289436
rect 5956 289380 6012 289436
rect 6012 289380 6016 289436
rect 5952 289376 6016 289380
rect 6032 289436 6096 289440
rect 6032 289380 6036 289436
rect 6036 289380 6092 289436
rect 6092 289380 6096 289436
rect 6032 289376 6096 289380
rect 6112 289436 6176 289440
rect 6112 289380 6116 289436
rect 6116 289380 6172 289436
rect 6172 289380 6176 289436
rect 6112 289376 6176 289380
rect 6192 289436 6256 289440
rect 6192 289380 6196 289436
rect 6196 289380 6252 289436
rect 6252 289380 6256 289436
rect 6192 289376 6256 289380
rect 4285 288892 4349 288896
rect 4285 288836 4289 288892
rect 4289 288836 4345 288892
rect 4345 288836 4349 288892
rect 4285 288832 4349 288836
rect 4365 288892 4429 288896
rect 4365 288836 4369 288892
rect 4369 288836 4425 288892
rect 4425 288836 4429 288892
rect 4365 288832 4429 288836
rect 4445 288892 4509 288896
rect 4445 288836 4449 288892
rect 4449 288836 4505 288892
rect 4505 288836 4509 288892
rect 4445 288832 4509 288836
rect 4525 288892 4589 288896
rect 4525 288836 4529 288892
rect 4529 288836 4585 288892
rect 4585 288836 4589 288892
rect 4525 288832 4589 288836
rect 7618 288892 7682 288896
rect 7618 288836 7622 288892
rect 7622 288836 7678 288892
rect 7678 288836 7682 288892
rect 7618 288832 7682 288836
rect 7698 288892 7762 288896
rect 7698 288836 7702 288892
rect 7702 288836 7758 288892
rect 7758 288836 7762 288892
rect 7698 288832 7762 288836
rect 7778 288892 7842 288896
rect 7778 288836 7782 288892
rect 7782 288836 7838 288892
rect 7838 288836 7842 288892
rect 7778 288832 7842 288836
rect 7858 288892 7922 288896
rect 7858 288836 7862 288892
rect 7862 288836 7918 288892
rect 7918 288836 7922 288892
rect 7858 288832 7922 288836
rect 2618 288348 2682 288352
rect 2618 288292 2622 288348
rect 2622 288292 2678 288348
rect 2678 288292 2682 288348
rect 2618 288288 2682 288292
rect 2698 288348 2762 288352
rect 2698 288292 2702 288348
rect 2702 288292 2758 288348
rect 2758 288292 2762 288348
rect 2698 288288 2762 288292
rect 2778 288348 2842 288352
rect 2778 288292 2782 288348
rect 2782 288292 2838 288348
rect 2838 288292 2842 288348
rect 2778 288288 2842 288292
rect 2858 288348 2922 288352
rect 2858 288292 2862 288348
rect 2862 288292 2918 288348
rect 2918 288292 2922 288348
rect 2858 288288 2922 288292
rect 5952 288348 6016 288352
rect 5952 288292 5956 288348
rect 5956 288292 6012 288348
rect 6012 288292 6016 288348
rect 5952 288288 6016 288292
rect 6032 288348 6096 288352
rect 6032 288292 6036 288348
rect 6036 288292 6092 288348
rect 6092 288292 6096 288348
rect 6032 288288 6096 288292
rect 6112 288348 6176 288352
rect 6112 288292 6116 288348
rect 6116 288292 6172 288348
rect 6172 288292 6176 288348
rect 6112 288288 6176 288292
rect 6192 288348 6256 288352
rect 6192 288292 6196 288348
rect 6196 288292 6252 288348
rect 6252 288292 6256 288348
rect 6192 288288 6256 288292
rect 4285 287804 4349 287808
rect 4285 287748 4289 287804
rect 4289 287748 4345 287804
rect 4345 287748 4349 287804
rect 4285 287744 4349 287748
rect 4365 287804 4429 287808
rect 4365 287748 4369 287804
rect 4369 287748 4425 287804
rect 4425 287748 4429 287804
rect 4365 287744 4429 287748
rect 4445 287804 4509 287808
rect 4445 287748 4449 287804
rect 4449 287748 4505 287804
rect 4505 287748 4509 287804
rect 4445 287744 4509 287748
rect 4525 287804 4589 287808
rect 4525 287748 4529 287804
rect 4529 287748 4585 287804
rect 4585 287748 4589 287804
rect 4525 287744 4589 287748
rect 7618 287804 7682 287808
rect 7618 287748 7622 287804
rect 7622 287748 7678 287804
rect 7678 287748 7682 287804
rect 7618 287744 7682 287748
rect 7698 287804 7762 287808
rect 7698 287748 7702 287804
rect 7702 287748 7758 287804
rect 7758 287748 7762 287804
rect 7698 287744 7762 287748
rect 7778 287804 7842 287808
rect 7778 287748 7782 287804
rect 7782 287748 7838 287804
rect 7838 287748 7842 287804
rect 7778 287744 7842 287748
rect 7858 287804 7922 287808
rect 7858 287748 7862 287804
rect 7862 287748 7918 287804
rect 7918 287748 7922 287804
rect 7858 287744 7922 287748
rect 2618 287260 2682 287264
rect 2618 287204 2622 287260
rect 2622 287204 2678 287260
rect 2678 287204 2682 287260
rect 2618 287200 2682 287204
rect 2698 287260 2762 287264
rect 2698 287204 2702 287260
rect 2702 287204 2758 287260
rect 2758 287204 2762 287260
rect 2698 287200 2762 287204
rect 2778 287260 2842 287264
rect 2778 287204 2782 287260
rect 2782 287204 2838 287260
rect 2838 287204 2842 287260
rect 2778 287200 2842 287204
rect 2858 287260 2922 287264
rect 2858 287204 2862 287260
rect 2862 287204 2918 287260
rect 2918 287204 2922 287260
rect 2858 287200 2922 287204
rect 5952 287260 6016 287264
rect 5952 287204 5956 287260
rect 5956 287204 6012 287260
rect 6012 287204 6016 287260
rect 5952 287200 6016 287204
rect 6032 287260 6096 287264
rect 6032 287204 6036 287260
rect 6036 287204 6092 287260
rect 6092 287204 6096 287260
rect 6032 287200 6096 287204
rect 6112 287260 6176 287264
rect 6112 287204 6116 287260
rect 6116 287204 6172 287260
rect 6172 287204 6176 287260
rect 6112 287200 6176 287204
rect 6192 287260 6256 287264
rect 6192 287204 6196 287260
rect 6196 287204 6252 287260
rect 6252 287204 6256 287260
rect 6192 287200 6256 287204
rect 4285 286716 4349 286720
rect 4285 286660 4289 286716
rect 4289 286660 4345 286716
rect 4345 286660 4349 286716
rect 4285 286656 4349 286660
rect 4365 286716 4429 286720
rect 4365 286660 4369 286716
rect 4369 286660 4425 286716
rect 4425 286660 4429 286716
rect 4365 286656 4429 286660
rect 4445 286716 4509 286720
rect 4445 286660 4449 286716
rect 4449 286660 4505 286716
rect 4505 286660 4509 286716
rect 4445 286656 4509 286660
rect 4525 286716 4589 286720
rect 4525 286660 4529 286716
rect 4529 286660 4585 286716
rect 4585 286660 4589 286716
rect 4525 286656 4589 286660
rect 7618 286716 7682 286720
rect 7618 286660 7622 286716
rect 7622 286660 7678 286716
rect 7678 286660 7682 286716
rect 7618 286656 7682 286660
rect 7698 286716 7762 286720
rect 7698 286660 7702 286716
rect 7702 286660 7758 286716
rect 7758 286660 7762 286716
rect 7698 286656 7762 286660
rect 7778 286716 7842 286720
rect 7778 286660 7782 286716
rect 7782 286660 7838 286716
rect 7838 286660 7842 286716
rect 7778 286656 7842 286660
rect 7858 286716 7922 286720
rect 7858 286660 7862 286716
rect 7862 286660 7918 286716
rect 7918 286660 7922 286716
rect 7858 286656 7922 286660
rect 2618 286172 2682 286176
rect 2618 286116 2622 286172
rect 2622 286116 2678 286172
rect 2678 286116 2682 286172
rect 2618 286112 2682 286116
rect 2698 286172 2762 286176
rect 2698 286116 2702 286172
rect 2702 286116 2758 286172
rect 2758 286116 2762 286172
rect 2698 286112 2762 286116
rect 2778 286172 2842 286176
rect 2778 286116 2782 286172
rect 2782 286116 2838 286172
rect 2838 286116 2842 286172
rect 2778 286112 2842 286116
rect 2858 286172 2922 286176
rect 2858 286116 2862 286172
rect 2862 286116 2918 286172
rect 2918 286116 2922 286172
rect 2858 286112 2922 286116
rect 5952 286172 6016 286176
rect 5952 286116 5956 286172
rect 5956 286116 6012 286172
rect 6012 286116 6016 286172
rect 5952 286112 6016 286116
rect 6032 286172 6096 286176
rect 6032 286116 6036 286172
rect 6036 286116 6092 286172
rect 6092 286116 6096 286172
rect 6032 286112 6096 286116
rect 6112 286172 6176 286176
rect 6112 286116 6116 286172
rect 6116 286116 6172 286172
rect 6172 286116 6176 286172
rect 6112 286112 6176 286116
rect 6192 286172 6256 286176
rect 6192 286116 6196 286172
rect 6196 286116 6252 286172
rect 6252 286116 6256 286172
rect 6192 286112 6256 286116
rect 4285 285628 4349 285632
rect 4285 285572 4289 285628
rect 4289 285572 4345 285628
rect 4345 285572 4349 285628
rect 4285 285568 4349 285572
rect 4365 285628 4429 285632
rect 4365 285572 4369 285628
rect 4369 285572 4425 285628
rect 4425 285572 4429 285628
rect 4365 285568 4429 285572
rect 4445 285628 4509 285632
rect 4445 285572 4449 285628
rect 4449 285572 4505 285628
rect 4505 285572 4509 285628
rect 4445 285568 4509 285572
rect 4525 285628 4589 285632
rect 4525 285572 4529 285628
rect 4529 285572 4585 285628
rect 4585 285572 4589 285628
rect 4525 285568 4589 285572
rect 7618 285628 7682 285632
rect 7618 285572 7622 285628
rect 7622 285572 7678 285628
rect 7678 285572 7682 285628
rect 7618 285568 7682 285572
rect 7698 285628 7762 285632
rect 7698 285572 7702 285628
rect 7702 285572 7758 285628
rect 7758 285572 7762 285628
rect 7698 285568 7762 285572
rect 7778 285628 7842 285632
rect 7778 285572 7782 285628
rect 7782 285572 7838 285628
rect 7838 285572 7842 285628
rect 7778 285568 7842 285572
rect 7858 285628 7922 285632
rect 7858 285572 7862 285628
rect 7862 285572 7918 285628
rect 7918 285572 7922 285628
rect 7858 285568 7922 285572
rect 2618 285084 2682 285088
rect 2618 285028 2622 285084
rect 2622 285028 2678 285084
rect 2678 285028 2682 285084
rect 2618 285024 2682 285028
rect 2698 285084 2762 285088
rect 2698 285028 2702 285084
rect 2702 285028 2758 285084
rect 2758 285028 2762 285084
rect 2698 285024 2762 285028
rect 2778 285084 2842 285088
rect 2778 285028 2782 285084
rect 2782 285028 2838 285084
rect 2838 285028 2842 285084
rect 2778 285024 2842 285028
rect 2858 285084 2922 285088
rect 2858 285028 2862 285084
rect 2862 285028 2918 285084
rect 2918 285028 2922 285084
rect 2858 285024 2922 285028
rect 5952 285084 6016 285088
rect 5952 285028 5956 285084
rect 5956 285028 6012 285084
rect 6012 285028 6016 285084
rect 5952 285024 6016 285028
rect 6032 285084 6096 285088
rect 6032 285028 6036 285084
rect 6036 285028 6092 285084
rect 6092 285028 6096 285084
rect 6032 285024 6096 285028
rect 6112 285084 6176 285088
rect 6112 285028 6116 285084
rect 6116 285028 6172 285084
rect 6172 285028 6176 285084
rect 6112 285024 6176 285028
rect 6192 285084 6256 285088
rect 6192 285028 6196 285084
rect 6196 285028 6252 285084
rect 6252 285028 6256 285084
rect 6192 285024 6256 285028
rect 4285 284540 4349 284544
rect 4285 284484 4289 284540
rect 4289 284484 4345 284540
rect 4345 284484 4349 284540
rect 4285 284480 4349 284484
rect 4365 284540 4429 284544
rect 4365 284484 4369 284540
rect 4369 284484 4425 284540
rect 4425 284484 4429 284540
rect 4365 284480 4429 284484
rect 4445 284540 4509 284544
rect 4445 284484 4449 284540
rect 4449 284484 4505 284540
rect 4505 284484 4509 284540
rect 4445 284480 4509 284484
rect 4525 284540 4589 284544
rect 4525 284484 4529 284540
rect 4529 284484 4585 284540
rect 4585 284484 4589 284540
rect 4525 284480 4589 284484
rect 7618 284540 7682 284544
rect 7618 284484 7622 284540
rect 7622 284484 7678 284540
rect 7678 284484 7682 284540
rect 7618 284480 7682 284484
rect 7698 284540 7762 284544
rect 7698 284484 7702 284540
rect 7702 284484 7758 284540
rect 7758 284484 7762 284540
rect 7698 284480 7762 284484
rect 7778 284540 7842 284544
rect 7778 284484 7782 284540
rect 7782 284484 7838 284540
rect 7838 284484 7842 284540
rect 7778 284480 7842 284484
rect 7858 284540 7922 284544
rect 7858 284484 7862 284540
rect 7862 284484 7918 284540
rect 7918 284484 7922 284540
rect 7858 284480 7922 284484
rect 2618 283996 2682 284000
rect 2618 283940 2622 283996
rect 2622 283940 2678 283996
rect 2678 283940 2682 283996
rect 2618 283936 2682 283940
rect 2698 283996 2762 284000
rect 2698 283940 2702 283996
rect 2702 283940 2758 283996
rect 2758 283940 2762 283996
rect 2698 283936 2762 283940
rect 2778 283996 2842 284000
rect 2778 283940 2782 283996
rect 2782 283940 2838 283996
rect 2838 283940 2842 283996
rect 2778 283936 2842 283940
rect 2858 283996 2922 284000
rect 2858 283940 2862 283996
rect 2862 283940 2918 283996
rect 2918 283940 2922 283996
rect 2858 283936 2922 283940
rect 5952 283996 6016 284000
rect 5952 283940 5956 283996
rect 5956 283940 6012 283996
rect 6012 283940 6016 283996
rect 5952 283936 6016 283940
rect 6032 283996 6096 284000
rect 6032 283940 6036 283996
rect 6036 283940 6092 283996
rect 6092 283940 6096 283996
rect 6032 283936 6096 283940
rect 6112 283996 6176 284000
rect 6112 283940 6116 283996
rect 6116 283940 6172 283996
rect 6172 283940 6176 283996
rect 6112 283936 6176 283940
rect 6192 283996 6256 284000
rect 6192 283940 6196 283996
rect 6196 283940 6252 283996
rect 6252 283940 6256 283996
rect 6192 283936 6256 283940
rect 4285 283452 4349 283456
rect 4285 283396 4289 283452
rect 4289 283396 4345 283452
rect 4345 283396 4349 283452
rect 4285 283392 4349 283396
rect 4365 283452 4429 283456
rect 4365 283396 4369 283452
rect 4369 283396 4425 283452
rect 4425 283396 4429 283452
rect 4365 283392 4429 283396
rect 4445 283452 4509 283456
rect 4445 283396 4449 283452
rect 4449 283396 4505 283452
rect 4505 283396 4509 283452
rect 4445 283392 4509 283396
rect 4525 283452 4589 283456
rect 4525 283396 4529 283452
rect 4529 283396 4585 283452
rect 4585 283396 4589 283452
rect 4525 283392 4589 283396
rect 7618 283452 7682 283456
rect 7618 283396 7622 283452
rect 7622 283396 7678 283452
rect 7678 283396 7682 283452
rect 7618 283392 7682 283396
rect 7698 283452 7762 283456
rect 7698 283396 7702 283452
rect 7702 283396 7758 283452
rect 7758 283396 7762 283452
rect 7698 283392 7762 283396
rect 7778 283452 7842 283456
rect 7778 283396 7782 283452
rect 7782 283396 7838 283452
rect 7838 283396 7842 283452
rect 7778 283392 7842 283396
rect 7858 283452 7922 283456
rect 7858 283396 7862 283452
rect 7862 283396 7918 283452
rect 7918 283396 7922 283452
rect 7858 283392 7922 283396
rect 2618 282908 2682 282912
rect 2618 282852 2622 282908
rect 2622 282852 2678 282908
rect 2678 282852 2682 282908
rect 2618 282848 2682 282852
rect 2698 282908 2762 282912
rect 2698 282852 2702 282908
rect 2702 282852 2758 282908
rect 2758 282852 2762 282908
rect 2698 282848 2762 282852
rect 2778 282908 2842 282912
rect 2778 282852 2782 282908
rect 2782 282852 2838 282908
rect 2838 282852 2842 282908
rect 2778 282848 2842 282852
rect 2858 282908 2922 282912
rect 2858 282852 2862 282908
rect 2862 282852 2918 282908
rect 2918 282852 2922 282908
rect 2858 282848 2922 282852
rect 5952 282908 6016 282912
rect 5952 282852 5956 282908
rect 5956 282852 6012 282908
rect 6012 282852 6016 282908
rect 5952 282848 6016 282852
rect 6032 282908 6096 282912
rect 6032 282852 6036 282908
rect 6036 282852 6092 282908
rect 6092 282852 6096 282908
rect 6032 282848 6096 282852
rect 6112 282908 6176 282912
rect 6112 282852 6116 282908
rect 6116 282852 6172 282908
rect 6172 282852 6176 282908
rect 6112 282848 6176 282852
rect 6192 282908 6256 282912
rect 6192 282852 6196 282908
rect 6196 282852 6252 282908
rect 6252 282852 6256 282908
rect 6192 282848 6256 282852
rect 4285 282364 4349 282368
rect 4285 282308 4289 282364
rect 4289 282308 4345 282364
rect 4345 282308 4349 282364
rect 4285 282304 4349 282308
rect 4365 282364 4429 282368
rect 4365 282308 4369 282364
rect 4369 282308 4425 282364
rect 4425 282308 4429 282364
rect 4365 282304 4429 282308
rect 4445 282364 4509 282368
rect 4445 282308 4449 282364
rect 4449 282308 4505 282364
rect 4505 282308 4509 282364
rect 4445 282304 4509 282308
rect 4525 282364 4589 282368
rect 4525 282308 4529 282364
rect 4529 282308 4585 282364
rect 4585 282308 4589 282364
rect 4525 282304 4589 282308
rect 7618 282364 7682 282368
rect 7618 282308 7622 282364
rect 7622 282308 7678 282364
rect 7678 282308 7682 282364
rect 7618 282304 7682 282308
rect 7698 282364 7762 282368
rect 7698 282308 7702 282364
rect 7702 282308 7758 282364
rect 7758 282308 7762 282364
rect 7698 282304 7762 282308
rect 7778 282364 7842 282368
rect 7778 282308 7782 282364
rect 7782 282308 7838 282364
rect 7838 282308 7842 282364
rect 7778 282304 7842 282308
rect 7858 282364 7922 282368
rect 7858 282308 7862 282364
rect 7862 282308 7918 282364
rect 7918 282308 7922 282364
rect 7858 282304 7922 282308
rect 2618 281820 2682 281824
rect 2618 281764 2622 281820
rect 2622 281764 2678 281820
rect 2678 281764 2682 281820
rect 2618 281760 2682 281764
rect 2698 281820 2762 281824
rect 2698 281764 2702 281820
rect 2702 281764 2758 281820
rect 2758 281764 2762 281820
rect 2698 281760 2762 281764
rect 2778 281820 2842 281824
rect 2778 281764 2782 281820
rect 2782 281764 2838 281820
rect 2838 281764 2842 281820
rect 2778 281760 2842 281764
rect 2858 281820 2922 281824
rect 2858 281764 2862 281820
rect 2862 281764 2918 281820
rect 2918 281764 2922 281820
rect 2858 281760 2922 281764
rect 5952 281820 6016 281824
rect 5952 281764 5956 281820
rect 5956 281764 6012 281820
rect 6012 281764 6016 281820
rect 5952 281760 6016 281764
rect 6032 281820 6096 281824
rect 6032 281764 6036 281820
rect 6036 281764 6092 281820
rect 6092 281764 6096 281820
rect 6032 281760 6096 281764
rect 6112 281820 6176 281824
rect 6112 281764 6116 281820
rect 6116 281764 6172 281820
rect 6172 281764 6176 281820
rect 6112 281760 6176 281764
rect 6192 281820 6256 281824
rect 6192 281764 6196 281820
rect 6196 281764 6252 281820
rect 6252 281764 6256 281820
rect 6192 281760 6256 281764
rect 4285 281276 4349 281280
rect 4285 281220 4289 281276
rect 4289 281220 4345 281276
rect 4345 281220 4349 281276
rect 4285 281216 4349 281220
rect 4365 281276 4429 281280
rect 4365 281220 4369 281276
rect 4369 281220 4425 281276
rect 4425 281220 4429 281276
rect 4365 281216 4429 281220
rect 4445 281276 4509 281280
rect 4445 281220 4449 281276
rect 4449 281220 4505 281276
rect 4505 281220 4509 281276
rect 4445 281216 4509 281220
rect 4525 281276 4589 281280
rect 4525 281220 4529 281276
rect 4529 281220 4585 281276
rect 4585 281220 4589 281276
rect 4525 281216 4589 281220
rect 7618 281276 7682 281280
rect 7618 281220 7622 281276
rect 7622 281220 7678 281276
rect 7678 281220 7682 281276
rect 7618 281216 7682 281220
rect 7698 281276 7762 281280
rect 7698 281220 7702 281276
rect 7702 281220 7758 281276
rect 7758 281220 7762 281276
rect 7698 281216 7762 281220
rect 7778 281276 7842 281280
rect 7778 281220 7782 281276
rect 7782 281220 7838 281276
rect 7838 281220 7842 281276
rect 7778 281216 7842 281220
rect 7858 281276 7922 281280
rect 7858 281220 7862 281276
rect 7862 281220 7918 281276
rect 7918 281220 7922 281276
rect 7858 281216 7922 281220
rect 2618 280732 2682 280736
rect 2618 280676 2622 280732
rect 2622 280676 2678 280732
rect 2678 280676 2682 280732
rect 2618 280672 2682 280676
rect 2698 280732 2762 280736
rect 2698 280676 2702 280732
rect 2702 280676 2758 280732
rect 2758 280676 2762 280732
rect 2698 280672 2762 280676
rect 2778 280732 2842 280736
rect 2778 280676 2782 280732
rect 2782 280676 2838 280732
rect 2838 280676 2842 280732
rect 2778 280672 2842 280676
rect 2858 280732 2922 280736
rect 2858 280676 2862 280732
rect 2862 280676 2918 280732
rect 2918 280676 2922 280732
rect 2858 280672 2922 280676
rect 5952 280732 6016 280736
rect 5952 280676 5956 280732
rect 5956 280676 6012 280732
rect 6012 280676 6016 280732
rect 5952 280672 6016 280676
rect 6032 280732 6096 280736
rect 6032 280676 6036 280732
rect 6036 280676 6092 280732
rect 6092 280676 6096 280732
rect 6032 280672 6096 280676
rect 6112 280732 6176 280736
rect 6112 280676 6116 280732
rect 6116 280676 6172 280732
rect 6172 280676 6176 280732
rect 6112 280672 6176 280676
rect 6192 280732 6256 280736
rect 6192 280676 6196 280732
rect 6196 280676 6252 280732
rect 6252 280676 6256 280732
rect 6192 280672 6256 280676
rect 4285 280188 4349 280192
rect 4285 280132 4289 280188
rect 4289 280132 4345 280188
rect 4345 280132 4349 280188
rect 4285 280128 4349 280132
rect 4365 280188 4429 280192
rect 4365 280132 4369 280188
rect 4369 280132 4425 280188
rect 4425 280132 4429 280188
rect 4365 280128 4429 280132
rect 4445 280188 4509 280192
rect 4445 280132 4449 280188
rect 4449 280132 4505 280188
rect 4505 280132 4509 280188
rect 4445 280128 4509 280132
rect 4525 280188 4589 280192
rect 4525 280132 4529 280188
rect 4529 280132 4585 280188
rect 4585 280132 4589 280188
rect 4525 280128 4589 280132
rect 7618 280188 7682 280192
rect 7618 280132 7622 280188
rect 7622 280132 7678 280188
rect 7678 280132 7682 280188
rect 7618 280128 7682 280132
rect 7698 280188 7762 280192
rect 7698 280132 7702 280188
rect 7702 280132 7758 280188
rect 7758 280132 7762 280188
rect 7698 280128 7762 280132
rect 7778 280188 7842 280192
rect 7778 280132 7782 280188
rect 7782 280132 7838 280188
rect 7838 280132 7842 280188
rect 7778 280128 7842 280132
rect 7858 280188 7922 280192
rect 7858 280132 7862 280188
rect 7862 280132 7918 280188
rect 7918 280132 7922 280188
rect 7858 280128 7922 280132
rect 2618 279644 2682 279648
rect 2618 279588 2622 279644
rect 2622 279588 2678 279644
rect 2678 279588 2682 279644
rect 2618 279584 2682 279588
rect 2698 279644 2762 279648
rect 2698 279588 2702 279644
rect 2702 279588 2758 279644
rect 2758 279588 2762 279644
rect 2698 279584 2762 279588
rect 2778 279644 2842 279648
rect 2778 279588 2782 279644
rect 2782 279588 2838 279644
rect 2838 279588 2842 279644
rect 2778 279584 2842 279588
rect 2858 279644 2922 279648
rect 2858 279588 2862 279644
rect 2862 279588 2918 279644
rect 2918 279588 2922 279644
rect 2858 279584 2922 279588
rect 5952 279644 6016 279648
rect 5952 279588 5956 279644
rect 5956 279588 6012 279644
rect 6012 279588 6016 279644
rect 5952 279584 6016 279588
rect 6032 279644 6096 279648
rect 6032 279588 6036 279644
rect 6036 279588 6092 279644
rect 6092 279588 6096 279644
rect 6032 279584 6096 279588
rect 6112 279644 6176 279648
rect 6112 279588 6116 279644
rect 6116 279588 6172 279644
rect 6172 279588 6176 279644
rect 6112 279584 6176 279588
rect 6192 279644 6256 279648
rect 6192 279588 6196 279644
rect 6196 279588 6252 279644
rect 6252 279588 6256 279644
rect 6192 279584 6256 279588
rect 4285 279100 4349 279104
rect 4285 279044 4289 279100
rect 4289 279044 4345 279100
rect 4345 279044 4349 279100
rect 4285 279040 4349 279044
rect 4365 279100 4429 279104
rect 4365 279044 4369 279100
rect 4369 279044 4425 279100
rect 4425 279044 4429 279100
rect 4365 279040 4429 279044
rect 4445 279100 4509 279104
rect 4445 279044 4449 279100
rect 4449 279044 4505 279100
rect 4505 279044 4509 279100
rect 4445 279040 4509 279044
rect 4525 279100 4589 279104
rect 4525 279044 4529 279100
rect 4529 279044 4585 279100
rect 4585 279044 4589 279100
rect 4525 279040 4589 279044
rect 7618 279100 7682 279104
rect 7618 279044 7622 279100
rect 7622 279044 7678 279100
rect 7678 279044 7682 279100
rect 7618 279040 7682 279044
rect 7698 279100 7762 279104
rect 7698 279044 7702 279100
rect 7702 279044 7758 279100
rect 7758 279044 7762 279100
rect 7698 279040 7762 279044
rect 7778 279100 7842 279104
rect 7778 279044 7782 279100
rect 7782 279044 7838 279100
rect 7838 279044 7842 279100
rect 7778 279040 7842 279044
rect 7858 279100 7922 279104
rect 7858 279044 7862 279100
rect 7862 279044 7918 279100
rect 7918 279044 7922 279100
rect 7858 279040 7922 279044
rect 2618 278556 2682 278560
rect 2618 278500 2622 278556
rect 2622 278500 2678 278556
rect 2678 278500 2682 278556
rect 2618 278496 2682 278500
rect 2698 278556 2762 278560
rect 2698 278500 2702 278556
rect 2702 278500 2758 278556
rect 2758 278500 2762 278556
rect 2698 278496 2762 278500
rect 2778 278556 2842 278560
rect 2778 278500 2782 278556
rect 2782 278500 2838 278556
rect 2838 278500 2842 278556
rect 2778 278496 2842 278500
rect 2858 278556 2922 278560
rect 2858 278500 2862 278556
rect 2862 278500 2918 278556
rect 2918 278500 2922 278556
rect 2858 278496 2922 278500
rect 5952 278556 6016 278560
rect 5952 278500 5956 278556
rect 5956 278500 6012 278556
rect 6012 278500 6016 278556
rect 5952 278496 6016 278500
rect 6032 278556 6096 278560
rect 6032 278500 6036 278556
rect 6036 278500 6092 278556
rect 6092 278500 6096 278556
rect 6032 278496 6096 278500
rect 6112 278556 6176 278560
rect 6112 278500 6116 278556
rect 6116 278500 6172 278556
rect 6172 278500 6176 278556
rect 6112 278496 6176 278500
rect 6192 278556 6256 278560
rect 6192 278500 6196 278556
rect 6196 278500 6252 278556
rect 6252 278500 6256 278556
rect 6192 278496 6256 278500
rect 4285 278012 4349 278016
rect 4285 277956 4289 278012
rect 4289 277956 4345 278012
rect 4345 277956 4349 278012
rect 4285 277952 4349 277956
rect 4365 278012 4429 278016
rect 4365 277956 4369 278012
rect 4369 277956 4425 278012
rect 4425 277956 4429 278012
rect 4365 277952 4429 277956
rect 4445 278012 4509 278016
rect 4445 277956 4449 278012
rect 4449 277956 4505 278012
rect 4505 277956 4509 278012
rect 4445 277952 4509 277956
rect 4525 278012 4589 278016
rect 4525 277956 4529 278012
rect 4529 277956 4585 278012
rect 4585 277956 4589 278012
rect 4525 277952 4589 277956
rect 7618 278012 7682 278016
rect 7618 277956 7622 278012
rect 7622 277956 7678 278012
rect 7678 277956 7682 278012
rect 7618 277952 7682 277956
rect 7698 278012 7762 278016
rect 7698 277956 7702 278012
rect 7702 277956 7758 278012
rect 7758 277956 7762 278012
rect 7698 277952 7762 277956
rect 7778 278012 7842 278016
rect 7778 277956 7782 278012
rect 7782 277956 7838 278012
rect 7838 277956 7842 278012
rect 7778 277952 7842 277956
rect 7858 278012 7922 278016
rect 7858 277956 7862 278012
rect 7862 277956 7918 278012
rect 7918 277956 7922 278012
rect 7858 277952 7922 277956
rect 2618 277468 2682 277472
rect 2618 277412 2622 277468
rect 2622 277412 2678 277468
rect 2678 277412 2682 277468
rect 2618 277408 2682 277412
rect 2698 277468 2762 277472
rect 2698 277412 2702 277468
rect 2702 277412 2758 277468
rect 2758 277412 2762 277468
rect 2698 277408 2762 277412
rect 2778 277468 2842 277472
rect 2778 277412 2782 277468
rect 2782 277412 2838 277468
rect 2838 277412 2842 277468
rect 2778 277408 2842 277412
rect 2858 277468 2922 277472
rect 2858 277412 2862 277468
rect 2862 277412 2918 277468
rect 2918 277412 2922 277468
rect 2858 277408 2922 277412
rect 5952 277468 6016 277472
rect 5952 277412 5956 277468
rect 5956 277412 6012 277468
rect 6012 277412 6016 277468
rect 5952 277408 6016 277412
rect 6032 277468 6096 277472
rect 6032 277412 6036 277468
rect 6036 277412 6092 277468
rect 6092 277412 6096 277468
rect 6032 277408 6096 277412
rect 6112 277468 6176 277472
rect 6112 277412 6116 277468
rect 6116 277412 6172 277468
rect 6172 277412 6176 277468
rect 6112 277408 6176 277412
rect 6192 277468 6256 277472
rect 6192 277412 6196 277468
rect 6196 277412 6252 277468
rect 6252 277412 6256 277468
rect 6192 277408 6256 277412
rect 4285 276924 4349 276928
rect 4285 276868 4289 276924
rect 4289 276868 4345 276924
rect 4345 276868 4349 276924
rect 4285 276864 4349 276868
rect 4365 276924 4429 276928
rect 4365 276868 4369 276924
rect 4369 276868 4425 276924
rect 4425 276868 4429 276924
rect 4365 276864 4429 276868
rect 4445 276924 4509 276928
rect 4445 276868 4449 276924
rect 4449 276868 4505 276924
rect 4505 276868 4509 276924
rect 4445 276864 4509 276868
rect 4525 276924 4589 276928
rect 4525 276868 4529 276924
rect 4529 276868 4585 276924
rect 4585 276868 4589 276924
rect 4525 276864 4589 276868
rect 7618 276924 7682 276928
rect 7618 276868 7622 276924
rect 7622 276868 7678 276924
rect 7678 276868 7682 276924
rect 7618 276864 7682 276868
rect 7698 276924 7762 276928
rect 7698 276868 7702 276924
rect 7702 276868 7758 276924
rect 7758 276868 7762 276924
rect 7698 276864 7762 276868
rect 7778 276924 7842 276928
rect 7778 276868 7782 276924
rect 7782 276868 7838 276924
rect 7838 276868 7842 276924
rect 7778 276864 7842 276868
rect 7858 276924 7922 276928
rect 7858 276868 7862 276924
rect 7862 276868 7918 276924
rect 7918 276868 7922 276924
rect 7858 276864 7922 276868
rect 2618 276380 2682 276384
rect 2618 276324 2622 276380
rect 2622 276324 2678 276380
rect 2678 276324 2682 276380
rect 2618 276320 2682 276324
rect 2698 276380 2762 276384
rect 2698 276324 2702 276380
rect 2702 276324 2758 276380
rect 2758 276324 2762 276380
rect 2698 276320 2762 276324
rect 2778 276380 2842 276384
rect 2778 276324 2782 276380
rect 2782 276324 2838 276380
rect 2838 276324 2842 276380
rect 2778 276320 2842 276324
rect 2858 276380 2922 276384
rect 2858 276324 2862 276380
rect 2862 276324 2918 276380
rect 2918 276324 2922 276380
rect 2858 276320 2922 276324
rect 5952 276380 6016 276384
rect 5952 276324 5956 276380
rect 5956 276324 6012 276380
rect 6012 276324 6016 276380
rect 5952 276320 6016 276324
rect 6032 276380 6096 276384
rect 6032 276324 6036 276380
rect 6036 276324 6092 276380
rect 6092 276324 6096 276380
rect 6032 276320 6096 276324
rect 6112 276380 6176 276384
rect 6112 276324 6116 276380
rect 6116 276324 6172 276380
rect 6172 276324 6176 276380
rect 6112 276320 6176 276324
rect 6192 276380 6256 276384
rect 6192 276324 6196 276380
rect 6196 276324 6252 276380
rect 6252 276324 6256 276380
rect 6192 276320 6256 276324
rect 4285 275836 4349 275840
rect 4285 275780 4289 275836
rect 4289 275780 4345 275836
rect 4345 275780 4349 275836
rect 4285 275776 4349 275780
rect 4365 275836 4429 275840
rect 4365 275780 4369 275836
rect 4369 275780 4425 275836
rect 4425 275780 4429 275836
rect 4365 275776 4429 275780
rect 4445 275836 4509 275840
rect 4445 275780 4449 275836
rect 4449 275780 4505 275836
rect 4505 275780 4509 275836
rect 4445 275776 4509 275780
rect 4525 275836 4589 275840
rect 4525 275780 4529 275836
rect 4529 275780 4585 275836
rect 4585 275780 4589 275836
rect 4525 275776 4589 275780
rect 7618 275836 7682 275840
rect 7618 275780 7622 275836
rect 7622 275780 7678 275836
rect 7678 275780 7682 275836
rect 7618 275776 7682 275780
rect 7698 275836 7762 275840
rect 7698 275780 7702 275836
rect 7702 275780 7758 275836
rect 7758 275780 7762 275836
rect 7698 275776 7762 275780
rect 7778 275836 7842 275840
rect 7778 275780 7782 275836
rect 7782 275780 7838 275836
rect 7838 275780 7842 275836
rect 7778 275776 7842 275780
rect 7858 275836 7922 275840
rect 7858 275780 7862 275836
rect 7862 275780 7918 275836
rect 7918 275780 7922 275836
rect 7858 275776 7922 275780
rect 2618 275292 2682 275296
rect 2618 275236 2622 275292
rect 2622 275236 2678 275292
rect 2678 275236 2682 275292
rect 2618 275232 2682 275236
rect 2698 275292 2762 275296
rect 2698 275236 2702 275292
rect 2702 275236 2758 275292
rect 2758 275236 2762 275292
rect 2698 275232 2762 275236
rect 2778 275292 2842 275296
rect 2778 275236 2782 275292
rect 2782 275236 2838 275292
rect 2838 275236 2842 275292
rect 2778 275232 2842 275236
rect 2858 275292 2922 275296
rect 2858 275236 2862 275292
rect 2862 275236 2918 275292
rect 2918 275236 2922 275292
rect 2858 275232 2922 275236
rect 5952 275292 6016 275296
rect 5952 275236 5956 275292
rect 5956 275236 6012 275292
rect 6012 275236 6016 275292
rect 5952 275232 6016 275236
rect 6032 275292 6096 275296
rect 6032 275236 6036 275292
rect 6036 275236 6092 275292
rect 6092 275236 6096 275292
rect 6032 275232 6096 275236
rect 6112 275292 6176 275296
rect 6112 275236 6116 275292
rect 6116 275236 6172 275292
rect 6172 275236 6176 275292
rect 6112 275232 6176 275236
rect 6192 275292 6256 275296
rect 6192 275236 6196 275292
rect 6196 275236 6252 275292
rect 6252 275236 6256 275292
rect 6192 275232 6256 275236
rect 4285 274748 4349 274752
rect 4285 274692 4289 274748
rect 4289 274692 4345 274748
rect 4345 274692 4349 274748
rect 4285 274688 4349 274692
rect 4365 274748 4429 274752
rect 4365 274692 4369 274748
rect 4369 274692 4425 274748
rect 4425 274692 4429 274748
rect 4365 274688 4429 274692
rect 4445 274748 4509 274752
rect 4445 274692 4449 274748
rect 4449 274692 4505 274748
rect 4505 274692 4509 274748
rect 4445 274688 4509 274692
rect 4525 274748 4589 274752
rect 4525 274692 4529 274748
rect 4529 274692 4585 274748
rect 4585 274692 4589 274748
rect 4525 274688 4589 274692
rect 7618 274748 7682 274752
rect 7618 274692 7622 274748
rect 7622 274692 7678 274748
rect 7678 274692 7682 274748
rect 7618 274688 7682 274692
rect 7698 274748 7762 274752
rect 7698 274692 7702 274748
rect 7702 274692 7758 274748
rect 7758 274692 7762 274748
rect 7698 274688 7762 274692
rect 7778 274748 7842 274752
rect 7778 274692 7782 274748
rect 7782 274692 7838 274748
rect 7838 274692 7842 274748
rect 7778 274688 7842 274692
rect 7858 274748 7922 274752
rect 7858 274692 7862 274748
rect 7862 274692 7918 274748
rect 7918 274692 7922 274748
rect 7858 274688 7922 274692
rect 2618 274204 2682 274208
rect 2618 274148 2622 274204
rect 2622 274148 2678 274204
rect 2678 274148 2682 274204
rect 2618 274144 2682 274148
rect 2698 274204 2762 274208
rect 2698 274148 2702 274204
rect 2702 274148 2758 274204
rect 2758 274148 2762 274204
rect 2698 274144 2762 274148
rect 2778 274204 2842 274208
rect 2778 274148 2782 274204
rect 2782 274148 2838 274204
rect 2838 274148 2842 274204
rect 2778 274144 2842 274148
rect 2858 274204 2922 274208
rect 2858 274148 2862 274204
rect 2862 274148 2918 274204
rect 2918 274148 2922 274204
rect 2858 274144 2922 274148
rect 5952 274204 6016 274208
rect 5952 274148 5956 274204
rect 5956 274148 6012 274204
rect 6012 274148 6016 274204
rect 5952 274144 6016 274148
rect 6032 274204 6096 274208
rect 6032 274148 6036 274204
rect 6036 274148 6092 274204
rect 6092 274148 6096 274204
rect 6032 274144 6096 274148
rect 6112 274204 6176 274208
rect 6112 274148 6116 274204
rect 6116 274148 6172 274204
rect 6172 274148 6176 274204
rect 6112 274144 6176 274148
rect 6192 274204 6256 274208
rect 6192 274148 6196 274204
rect 6196 274148 6252 274204
rect 6252 274148 6256 274204
rect 6192 274144 6256 274148
rect 4285 273660 4349 273664
rect 4285 273604 4289 273660
rect 4289 273604 4345 273660
rect 4345 273604 4349 273660
rect 4285 273600 4349 273604
rect 4365 273660 4429 273664
rect 4365 273604 4369 273660
rect 4369 273604 4425 273660
rect 4425 273604 4429 273660
rect 4365 273600 4429 273604
rect 4445 273660 4509 273664
rect 4445 273604 4449 273660
rect 4449 273604 4505 273660
rect 4505 273604 4509 273660
rect 4445 273600 4509 273604
rect 4525 273660 4589 273664
rect 4525 273604 4529 273660
rect 4529 273604 4585 273660
rect 4585 273604 4589 273660
rect 4525 273600 4589 273604
rect 7618 273660 7682 273664
rect 7618 273604 7622 273660
rect 7622 273604 7678 273660
rect 7678 273604 7682 273660
rect 7618 273600 7682 273604
rect 7698 273660 7762 273664
rect 7698 273604 7702 273660
rect 7702 273604 7758 273660
rect 7758 273604 7762 273660
rect 7698 273600 7762 273604
rect 7778 273660 7842 273664
rect 7778 273604 7782 273660
rect 7782 273604 7838 273660
rect 7838 273604 7842 273660
rect 7778 273600 7842 273604
rect 7858 273660 7922 273664
rect 7858 273604 7862 273660
rect 7862 273604 7918 273660
rect 7918 273604 7922 273660
rect 7858 273600 7922 273604
rect 2618 273116 2682 273120
rect 2618 273060 2622 273116
rect 2622 273060 2678 273116
rect 2678 273060 2682 273116
rect 2618 273056 2682 273060
rect 2698 273116 2762 273120
rect 2698 273060 2702 273116
rect 2702 273060 2758 273116
rect 2758 273060 2762 273116
rect 2698 273056 2762 273060
rect 2778 273116 2842 273120
rect 2778 273060 2782 273116
rect 2782 273060 2838 273116
rect 2838 273060 2842 273116
rect 2778 273056 2842 273060
rect 2858 273116 2922 273120
rect 2858 273060 2862 273116
rect 2862 273060 2918 273116
rect 2918 273060 2922 273116
rect 2858 273056 2922 273060
rect 5952 273116 6016 273120
rect 5952 273060 5956 273116
rect 5956 273060 6012 273116
rect 6012 273060 6016 273116
rect 5952 273056 6016 273060
rect 6032 273116 6096 273120
rect 6032 273060 6036 273116
rect 6036 273060 6092 273116
rect 6092 273060 6096 273116
rect 6032 273056 6096 273060
rect 6112 273116 6176 273120
rect 6112 273060 6116 273116
rect 6116 273060 6172 273116
rect 6172 273060 6176 273116
rect 6112 273056 6176 273060
rect 6192 273116 6256 273120
rect 6192 273060 6196 273116
rect 6196 273060 6252 273116
rect 6252 273060 6256 273116
rect 6192 273056 6256 273060
rect 4285 272572 4349 272576
rect 4285 272516 4289 272572
rect 4289 272516 4345 272572
rect 4345 272516 4349 272572
rect 4285 272512 4349 272516
rect 4365 272572 4429 272576
rect 4365 272516 4369 272572
rect 4369 272516 4425 272572
rect 4425 272516 4429 272572
rect 4365 272512 4429 272516
rect 4445 272572 4509 272576
rect 4445 272516 4449 272572
rect 4449 272516 4505 272572
rect 4505 272516 4509 272572
rect 4445 272512 4509 272516
rect 4525 272572 4589 272576
rect 4525 272516 4529 272572
rect 4529 272516 4585 272572
rect 4585 272516 4589 272572
rect 4525 272512 4589 272516
rect 7618 272572 7682 272576
rect 7618 272516 7622 272572
rect 7622 272516 7678 272572
rect 7678 272516 7682 272572
rect 7618 272512 7682 272516
rect 7698 272572 7762 272576
rect 7698 272516 7702 272572
rect 7702 272516 7758 272572
rect 7758 272516 7762 272572
rect 7698 272512 7762 272516
rect 7778 272572 7842 272576
rect 7778 272516 7782 272572
rect 7782 272516 7838 272572
rect 7838 272516 7842 272572
rect 7778 272512 7842 272516
rect 7858 272572 7922 272576
rect 7858 272516 7862 272572
rect 7862 272516 7918 272572
rect 7918 272516 7922 272572
rect 7858 272512 7922 272516
rect 2618 272028 2682 272032
rect 2618 271972 2622 272028
rect 2622 271972 2678 272028
rect 2678 271972 2682 272028
rect 2618 271968 2682 271972
rect 2698 272028 2762 272032
rect 2698 271972 2702 272028
rect 2702 271972 2758 272028
rect 2758 271972 2762 272028
rect 2698 271968 2762 271972
rect 2778 272028 2842 272032
rect 2778 271972 2782 272028
rect 2782 271972 2838 272028
rect 2838 271972 2842 272028
rect 2778 271968 2842 271972
rect 2858 272028 2922 272032
rect 2858 271972 2862 272028
rect 2862 271972 2918 272028
rect 2918 271972 2922 272028
rect 2858 271968 2922 271972
rect 5952 272028 6016 272032
rect 5952 271972 5956 272028
rect 5956 271972 6012 272028
rect 6012 271972 6016 272028
rect 5952 271968 6016 271972
rect 6032 272028 6096 272032
rect 6032 271972 6036 272028
rect 6036 271972 6092 272028
rect 6092 271972 6096 272028
rect 6032 271968 6096 271972
rect 6112 272028 6176 272032
rect 6112 271972 6116 272028
rect 6116 271972 6172 272028
rect 6172 271972 6176 272028
rect 6112 271968 6176 271972
rect 6192 272028 6256 272032
rect 6192 271972 6196 272028
rect 6196 271972 6252 272028
rect 6252 271972 6256 272028
rect 6192 271968 6256 271972
rect 4285 271484 4349 271488
rect 4285 271428 4289 271484
rect 4289 271428 4345 271484
rect 4345 271428 4349 271484
rect 4285 271424 4349 271428
rect 4365 271484 4429 271488
rect 4365 271428 4369 271484
rect 4369 271428 4425 271484
rect 4425 271428 4429 271484
rect 4365 271424 4429 271428
rect 4445 271484 4509 271488
rect 4445 271428 4449 271484
rect 4449 271428 4505 271484
rect 4505 271428 4509 271484
rect 4445 271424 4509 271428
rect 4525 271484 4589 271488
rect 4525 271428 4529 271484
rect 4529 271428 4585 271484
rect 4585 271428 4589 271484
rect 4525 271424 4589 271428
rect 7618 271484 7682 271488
rect 7618 271428 7622 271484
rect 7622 271428 7678 271484
rect 7678 271428 7682 271484
rect 7618 271424 7682 271428
rect 7698 271484 7762 271488
rect 7698 271428 7702 271484
rect 7702 271428 7758 271484
rect 7758 271428 7762 271484
rect 7698 271424 7762 271428
rect 7778 271484 7842 271488
rect 7778 271428 7782 271484
rect 7782 271428 7838 271484
rect 7838 271428 7842 271484
rect 7778 271424 7842 271428
rect 7858 271484 7922 271488
rect 7858 271428 7862 271484
rect 7862 271428 7918 271484
rect 7918 271428 7922 271484
rect 7858 271424 7922 271428
rect 2618 270940 2682 270944
rect 2618 270884 2622 270940
rect 2622 270884 2678 270940
rect 2678 270884 2682 270940
rect 2618 270880 2682 270884
rect 2698 270940 2762 270944
rect 2698 270884 2702 270940
rect 2702 270884 2758 270940
rect 2758 270884 2762 270940
rect 2698 270880 2762 270884
rect 2778 270940 2842 270944
rect 2778 270884 2782 270940
rect 2782 270884 2838 270940
rect 2838 270884 2842 270940
rect 2778 270880 2842 270884
rect 2858 270940 2922 270944
rect 2858 270884 2862 270940
rect 2862 270884 2918 270940
rect 2918 270884 2922 270940
rect 2858 270880 2922 270884
rect 5952 270940 6016 270944
rect 5952 270884 5956 270940
rect 5956 270884 6012 270940
rect 6012 270884 6016 270940
rect 5952 270880 6016 270884
rect 6032 270940 6096 270944
rect 6032 270884 6036 270940
rect 6036 270884 6092 270940
rect 6092 270884 6096 270940
rect 6032 270880 6096 270884
rect 6112 270940 6176 270944
rect 6112 270884 6116 270940
rect 6116 270884 6172 270940
rect 6172 270884 6176 270940
rect 6112 270880 6176 270884
rect 6192 270940 6256 270944
rect 6192 270884 6196 270940
rect 6196 270884 6252 270940
rect 6252 270884 6256 270940
rect 6192 270880 6256 270884
rect 4285 270396 4349 270400
rect 4285 270340 4289 270396
rect 4289 270340 4345 270396
rect 4345 270340 4349 270396
rect 4285 270336 4349 270340
rect 4365 270396 4429 270400
rect 4365 270340 4369 270396
rect 4369 270340 4425 270396
rect 4425 270340 4429 270396
rect 4365 270336 4429 270340
rect 4445 270396 4509 270400
rect 4445 270340 4449 270396
rect 4449 270340 4505 270396
rect 4505 270340 4509 270396
rect 4445 270336 4509 270340
rect 4525 270396 4589 270400
rect 4525 270340 4529 270396
rect 4529 270340 4585 270396
rect 4585 270340 4589 270396
rect 4525 270336 4589 270340
rect 7618 270396 7682 270400
rect 7618 270340 7622 270396
rect 7622 270340 7678 270396
rect 7678 270340 7682 270396
rect 7618 270336 7682 270340
rect 7698 270396 7762 270400
rect 7698 270340 7702 270396
rect 7702 270340 7758 270396
rect 7758 270340 7762 270396
rect 7698 270336 7762 270340
rect 7778 270396 7842 270400
rect 7778 270340 7782 270396
rect 7782 270340 7838 270396
rect 7838 270340 7842 270396
rect 7778 270336 7842 270340
rect 7858 270396 7922 270400
rect 7858 270340 7862 270396
rect 7862 270340 7918 270396
rect 7918 270340 7922 270396
rect 7858 270336 7922 270340
rect 2618 269852 2682 269856
rect 2618 269796 2622 269852
rect 2622 269796 2678 269852
rect 2678 269796 2682 269852
rect 2618 269792 2682 269796
rect 2698 269852 2762 269856
rect 2698 269796 2702 269852
rect 2702 269796 2758 269852
rect 2758 269796 2762 269852
rect 2698 269792 2762 269796
rect 2778 269852 2842 269856
rect 2778 269796 2782 269852
rect 2782 269796 2838 269852
rect 2838 269796 2842 269852
rect 2778 269792 2842 269796
rect 2858 269852 2922 269856
rect 2858 269796 2862 269852
rect 2862 269796 2918 269852
rect 2918 269796 2922 269852
rect 2858 269792 2922 269796
rect 5952 269852 6016 269856
rect 5952 269796 5956 269852
rect 5956 269796 6012 269852
rect 6012 269796 6016 269852
rect 5952 269792 6016 269796
rect 6032 269852 6096 269856
rect 6032 269796 6036 269852
rect 6036 269796 6092 269852
rect 6092 269796 6096 269852
rect 6032 269792 6096 269796
rect 6112 269852 6176 269856
rect 6112 269796 6116 269852
rect 6116 269796 6172 269852
rect 6172 269796 6176 269852
rect 6112 269792 6176 269796
rect 6192 269852 6256 269856
rect 6192 269796 6196 269852
rect 6196 269796 6252 269852
rect 6252 269796 6256 269852
rect 6192 269792 6256 269796
rect 4285 269308 4349 269312
rect 4285 269252 4289 269308
rect 4289 269252 4345 269308
rect 4345 269252 4349 269308
rect 4285 269248 4349 269252
rect 4365 269308 4429 269312
rect 4365 269252 4369 269308
rect 4369 269252 4425 269308
rect 4425 269252 4429 269308
rect 4365 269248 4429 269252
rect 4445 269308 4509 269312
rect 4445 269252 4449 269308
rect 4449 269252 4505 269308
rect 4505 269252 4509 269308
rect 4445 269248 4509 269252
rect 4525 269308 4589 269312
rect 4525 269252 4529 269308
rect 4529 269252 4585 269308
rect 4585 269252 4589 269308
rect 4525 269248 4589 269252
rect 7618 269308 7682 269312
rect 7618 269252 7622 269308
rect 7622 269252 7678 269308
rect 7678 269252 7682 269308
rect 7618 269248 7682 269252
rect 7698 269308 7762 269312
rect 7698 269252 7702 269308
rect 7702 269252 7758 269308
rect 7758 269252 7762 269308
rect 7698 269248 7762 269252
rect 7778 269308 7842 269312
rect 7778 269252 7782 269308
rect 7782 269252 7838 269308
rect 7838 269252 7842 269308
rect 7778 269248 7842 269252
rect 7858 269308 7922 269312
rect 7858 269252 7862 269308
rect 7862 269252 7918 269308
rect 7918 269252 7922 269308
rect 7858 269248 7922 269252
rect 2618 268764 2682 268768
rect 2618 268708 2622 268764
rect 2622 268708 2678 268764
rect 2678 268708 2682 268764
rect 2618 268704 2682 268708
rect 2698 268764 2762 268768
rect 2698 268708 2702 268764
rect 2702 268708 2758 268764
rect 2758 268708 2762 268764
rect 2698 268704 2762 268708
rect 2778 268764 2842 268768
rect 2778 268708 2782 268764
rect 2782 268708 2838 268764
rect 2838 268708 2842 268764
rect 2778 268704 2842 268708
rect 2858 268764 2922 268768
rect 2858 268708 2862 268764
rect 2862 268708 2918 268764
rect 2918 268708 2922 268764
rect 2858 268704 2922 268708
rect 5952 268764 6016 268768
rect 5952 268708 5956 268764
rect 5956 268708 6012 268764
rect 6012 268708 6016 268764
rect 5952 268704 6016 268708
rect 6032 268764 6096 268768
rect 6032 268708 6036 268764
rect 6036 268708 6092 268764
rect 6092 268708 6096 268764
rect 6032 268704 6096 268708
rect 6112 268764 6176 268768
rect 6112 268708 6116 268764
rect 6116 268708 6172 268764
rect 6172 268708 6176 268764
rect 6112 268704 6176 268708
rect 6192 268764 6256 268768
rect 6192 268708 6196 268764
rect 6196 268708 6252 268764
rect 6252 268708 6256 268764
rect 6192 268704 6256 268708
rect 4285 268220 4349 268224
rect 4285 268164 4289 268220
rect 4289 268164 4345 268220
rect 4345 268164 4349 268220
rect 4285 268160 4349 268164
rect 4365 268220 4429 268224
rect 4365 268164 4369 268220
rect 4369 268164 4425 268220
rect 4425 268164 4429 268220
rect 4365 268160 4429 268164
rect 4445 268220 4509 268224
rect 4445 268164 4449 268220
rect 4449 268164 4505 268220
rect 4505 268164 4509 268220
rect 4445 268160 4509 268164
rect 4525 268220 4589 268224
rect 4525 268164 4529 268220
rect 4529 268164 4585 268220
rect 4585 268164 4589 268220
rect 4525 268160 4589 268164
rect 7618 268220 7682 268224
rect 7618 268164 7622 268220
rect 7622 268164 7678 268220
rect 7678 268164 7682 268220
rect 7618 268160 7682 268164
rect 7698 268220 7762 268224
rect 7698 268164 7702 268220
rect 7702 268164 7758 268220
rect 7758 268164 7762 268220
rect 7698 268160 7762 268164
rect 7778 268220 7842 268224
rect 7778 268164 7782 268220
rect 7782 268164 7838 268220
rect 7838 268164 7842 268220
rect 7778 268160 7842 268164
rect 7858 268220 7922 268224
rect 7858 268164 7862 268220
rect 7862 268164 7918 268220
rect 7918 268164 7922 268220
rect 7858 268160 7922 268164
rect 2618 267676 2682 267680
rect 2618 267620 2622 267676
rect 2622 267620 2678 267676
rect 2678 267620 2682 267676
rect 2618 267616 2682 267620
rect 2698 267676 2762 267680
rect 2698 267620 2702 267676
rect 2702 267620 2758 267676
rect 2758 267620 2762 267676
rect 2698 267616 2762 267620
rect 2778 267676 2842 267680
rect 2778 267620 2782 267676
rect 2782 267620 2838 267676
rect 2838 267620 2842 267676
rect 2778 267616 2842 267620
rect 2858 267676 2922 267680
rect 2858 267620 2862 267676
rect 2862 267620 2918 267676
rect 2918 267620 2922 267676
rect 2858 267616 2922 267620
rect 5952 267676 6016 267680
rect 5952 267620 5956 267676
rect 5956 267620 6012 267676
rect 6012 267620 6016 267676
rect 5952 267616 6016 267620
rect 6032 267676 6096 267680
rect 6032 267620 6036 267676
rect 6036 267620 6092 267676
rect 6092 267620 6096 267676
rect 6032 267616 6096 267620
rect 6112 267676 6176 267680
rect 6112 267620 6116 267676
rect 6116 267620 6172 267676
rect 6172 267620 6176 267676
rect 6112 267616 6176 267620
rect 6192 267676 6256 267680
rect 6192 267620 6196 267676
rect 6196 267620 6252 267676
rect 6252 267620 6256 267676
rect 6192 267616 6256 267620
rect 4285 267132 4349 267136
rect 4285 267076 4289 267132
rect 4289 267076 4345 267132
rect 4345 267076 4349 267132
rect 4285 267072 4349 267076
rect 4365 267132 4429 267136
rect 4365 267076 4369 267132
rect 4369 267076 4425 267132
rect 4425 267076 4429 267132
rect 4365 267072 4429 267076
rect 4445 267132 4509 267136
rect 4445 267076 4449 267132
rect 4449 267076 4505 267132
rect 4505 267076 4509 267132
rect 4445 267072 4509 267076
rect 4525 267132 4589 267136
rect 4525 267076 4529 267132
rect 4529 267076 4585 267132
rect 4585 267076 4589 267132
rect 4525 267072 4589 267076
rect 7618 267132 7682 267136
rect 7618 267076 7622 267132
rect 7622 267076 7678 267132
rect 7678 267076 7682 267132
rect 7618 267072 7682 267076
rect 7698 267132 7762 267136
rect 7698 267076 7702 267132
rect 7702 267076 7758 267132
rect 7758 267076 7762 267132
rect 7698 267072 7762 267076
rect 7778 267132 7842 267136
rect 7778 267076 7782 267132
rect 7782 267076 7838 267132
rect 7838 267076 7842 267132
rect 7778 267072 7842 267076
rect 7858 267132 7922 267136
rect 7858 267076 7862 267132
rect 7862 267076 7918 267132
rect 7918 267076 7922 267132
rect 7858 267072 7922 267076
rect 2618 266588 2682 266592
rect 2618 266532 2622 266588
rect 2622 266532 2678 266588
rect 2678 266532 2682 266588
rect 2618 266528 2682 266532
rect 2698 266588 2762 266592
rect 2698 266532 2702 266588
rect 2702 266532 2758 266588
rect 2758 266532 2762 266588
rect 2698 266528 2762 266532
rect 2778 266588 2842 266592
rect 2778 266532 2782 266588
rect 2782 266532 2838 266588
rect 2838 266532 2842 266588
rect 2778 266528 2842 266532
rect 2858 266588 2922 266592
rect 2858 266532 2862 266588
rect 2862 266532 2918 266588
rect 2918 266532 2922 266588
rect 2858 266528 2922 266532
rect 5952 266588 6016 266592
rect 5952 266532 5956 266588
rect 5956 266532 6012 266588
rect 6012 266532 6016 266588
rect 5952 266528 6016 266532
rect 6032 266588 6096 266592
rect 6032 266532 6036 266588
rect 6036 266532 6092 266588
rect 6092 266532 6096 266588
rect 6032 266528 6096 266532
rect 6112 266588 6176 266592
rect 6112 266532 6116 266588
rect 6116 266532 6172 266588
rect 6172 266532 6176 266588
rect 6112 266528 6176 266532
rect 6192 266588 6256 266592
rect 6192 266532 6196 266588
rect 6196 266532 6252 266588
rect 6252 266532 6256 266588
rect 6192 266528 6256 266532
rect 4285 266044 4349 266048
rect 4285 265988 4289 266044
rect 4289 265988 4345 266044
rect 4345 265988 4349 266044
rect 4285 265984 4349 265988
rect 4365 266044 4429 266048
rect 4365 265988 4369 266044
rect 4369 265988 4425 266044
rect 4425 265988 4429 266044
rect 4365 265984 4429 265988
rect 4445 266044 4509 266048
rect 4445 265988 4449 266044
rect 4449 265988 4505 266044
rect 4505 265988 4509 266044
rect 4445 265984 4509 265988
rect 4525 266044 4589 266048
rect 4525 265988 4529 266044
rect 4529 265988 4585 266044
rect 4585 265988 4589 266044
rect 4525 265984 4589 265988
rect 7618 266044 7682 266048
rect 7618 265988 7622 266044
rect 7622 265988 7678 266044
rect 7678 265988 7682 266044
rect 7618 265984 7682 265988
rect 7698 266044 7762 266048
rect 7698 265988 7702 266044
rect 7702 265988 7758 266044
rect 7758 265988 7762 266044
rect 7698 265984 7762 265988
rect 7778 266044 7842 266048
rect 7778 265988 7782 266044
rect 7782 265988 7838 266044
rect 7838 265988 7842 266044
rect 7778 265984 7842 265988
rect 7858 266044 7922 266048
rect 7858 265988 7862 266044
rect 7862 265988 7918 266044
rect 7918 265988 7922 266044
rect 7858 265984 7922 265988
rect 2618 265500 2682 265504
rect 2618 265444 2622 265500
rect 2622 265444 2678 265500
rect 2678 265444 2682 265500
rect 2618 265440 2682 265444
rect 2698 265500 2762 265504
rect 2698 265444 2702 265500
rect 2702 265444 2758 265500
rect 2758 265444 2762 265500
rect 2698 265440 2762 265444
rect 2778 265500 2842 265504
rect 2778 265444 2782 265500
rect 2782 265444 2838 265500
rect 2838 265444 2842 265500
rect 2778 265440 2842 265444
rect 2858 265500 2922 265504
rect 2858 265444 2862 265500
rect 2862 265444 2918 265500
rect 2918 265444 2922 265500
rect 2858 265440 2922 265444
rect 5952 265500 6016 265504
rect 5952 265444 5956 265500
rect 5956 265444 6012 265500
rect 6012 265444 6016 265500
rect 5952 265440 6016 265444
rect 6032 265500 6096 265504
rect 6032 265444 6036 265500
rect 6036 265444 6092 265500
rect 6092 265444 6096 265500
rect 6032 265440 6096 265444
rect 6112 265500 6176 265504
rect 6112 265444 6116 265500
rect 6116 265444 6172 265500
rect 6172 265444 6176 265500
rect 6112 265440 6176 265444
rect 6192 265500 6256 265504
rect 6192 265444 6196 265500
rect 6196 265444 6252 265500
rect 6252 265444 6256 265500
rect 6192 265440 6256 265444
rect 4285 264956 4349 264960
rect 4285 264900 4289 264956
rect 4289 264900 4345 264956
rect 4345 264900 4349 264956
rect 4285 264896 4349 264900
rect 4365 264956 4429 264960
rect 4365 264900 4369 264956
rect 4369 264900 4425 264956
rect 4425 264900 4429 264956
rect 4365 264896 4429 264900
rect 4445 264956 4509 264960
rect 4445 264900 4449 264956
rect 4449 264900 4505 264956
rect 4505 264900 4509 264956
rect 4445 264896 4509 264900
rect 4525 264956 4589 264960
rect 4525 264900 4529 264956
rect 4529 264900 4585 264956
rect 4585 264900 4589 264956
rect 4525 264896 4589 264900
rect 7618 264956 7682 264960
rect 7618 264900 7622 264956
rect 7622 264900 7678 264956
rect 7678 264900 7682 264956
rect 7618 264896 7682 264900
rect 7698 264956 7762 264960
rect 7698 264900 7702 264956
rect 7702 264900 7758 264956
rect 7758 264900 7762 264956
rect 7698 264896 7762 264900
rect 7778 264956 7842 264960
rect 7778 264900 7782 264956
rect 7782 264900 7838 264956
rect 7838 264900 7842 264956
rect 7778 264896 7842 264900
rect 7858 264956 7922 264960
rect 7858 264900 7862 264956
rect 7862 264900 7918 264956
rect 7918 264900 7922 264956
rect 7858 264896 7922 264900
rect 2618 264412 2682 264416
rect 2618 264356 2622 264412
rect 2622 264356 2678 264412
rect 2678 264356 2682 264412
rect 2618 264352 2682 264356
rect 2698 264412 2762 264416
rect 2698 264356 2702 264412
rect 2702 264356 2758 264412
rect 2758 264356 2762 264412
rect 2698 264352 2762 264356
rect 2778 264412 2842 264416
rect 2778 264356 2782 264412
rect 2782 264356 2838 264412
rect 2838 264356 2842 264412
rect 2778 264352 2842 264356
rect 2858 264412 2922 264416
rect 2858 264356 2862 264412
rect 2862 264356 2918 264412
rect 2918 264356 2922 264412
rect 2858 264352 2922 264356
rect 5952 264412 6016 264416
rect 5952 264356 5956 264412
rect 5956 264356 6012 264412
rect 6012 264356 6016 264412
rect 5952 264352 6016 264356
rect 6032 264412 6096 264416
rect 6032 264356 6036 264412
rect 6036 264356 6092 264412
rect 6092 264356 6096 264412
rect 6032 264352 6096 264356
rect 6112 264412 6176 264416
rect 6112 264356 6116 264412
rect 6116 264356 6172 264412
rect 6172 264356 6176 264412
rect 6112 264352 6176 264356
rect 6192 264412 6256 264416
rect 6192 264356 6196 264412
rect 6196 264356 6252 264412
rect 6252 264356 6256 264412
rect 6192 264352 6256 264356
rect 4285 263868 4349 263872
rect 4285 263812 4289 263868
rect 4289 263812 4345 263868
rect 4345 263812 4349 263868
rect 4285 263808 4349 263812
rect 4365 263868 4429 263872
rect 4365 263812 4369 263868
rect 4369 263812 4425 263868
rect 4425 263812 4429 263868
rect 4365 263808 4429 263812
rect 4445 263868 4509 263872
rect 4445 263812 4449 263868
rect 4449 263812 4505 263868
rect 4505 263812 4509 263868
rect 4445 263808 4509 263812
rect 4525 263868 4589 263872
rect 4525 263812 4529 263868
rect 4529 263812 4585 263868
rect 4585 263812 4589 263868
rect 4525 263808 4589 263812
rect 7618 263868 7682 263872
rect 7618 263812 7622 263868
rect 7622 263812 7678 263868
rect 7678 263812 7682 263868
rect 7618 263808 7682 263812
rect 7698 263868 7762 263872
rect 7698 263812 7702 263868
rect 7702 263812 7758 263868
rect 7758 263812 7762 263868
rect 7698 263808 7762 263812
rect 7778 263868 7842 263872
rect 7778 263812 7782 263868
rect 7782 263812 7838 263868
rect 7838 263812 7842 263868
rect 7778 263808 7842 263812
rect 7858 263868 7922 263872
rect 7858 263812 7862 263868
rect 7862 263812 7918 263868
rect 7918 263812 7922 263868
rect 7858 263808 7922 263812
rect 2618 263324 2682 263328
rect 2618 263268 2622 263324
rect 2622 263268 2678 263324
rect 2678 263268 2682 263324
rect 2618 263264 2682 263268
rect 2698 263324 2762 263328
rect 2698 263268 2702 263324
rect 2702 263268 2758 263324
rect 2758 263268 2762 263324
rect 2698 263264 2762 263268
rect 2778 263324 2842 263328
rect 2778 263268 2782 263324
rect 2782 263268 2838 263324
rect 2838 263268 2842 263324
rect 2778 263264 2842 263268
rect 2858 263324 2922 263328
rect 2858 263268 2862 263324
rect 2862 263268 2918 263324
rect 2918 263268 2922 263324
rect 2858 263264 2922 263268
rect 5952 263324 6016 263328
rect 5952 263268 5956 263324
rect 5956 263268 6012 263324
rect 6012 263268 6016 263324
rect 5952 263264 6016 263268
rect 6032 263324 6096 263328
rect 6032 263268 6036 263324
rect 6036 263268 6092 263324
rect 6092 263268 6096 263324
rect 6032 263264 6096 263268
rect 6112 263324 6176 263328
rect 6112 263268 6116 263324
rect 6116 263268 6172 263324
rect 6172 263268 6176 263324
rect 6112 263264 6176 263268
rect 6192 263324 6256 263328
rect 6192 263268 6196 263324
rect 6196 263268 6252 263324
rect 6252 263268 6256 263324
rect 6192 263264 6256 263268
rect 4285 262780 4349 262784
rect 4285 262724 4289 262780
rect 4289 262724 4345 262780
rect 4345 262724 4349 262780
rect 4285 262720 4349 262724
rect 4365 262780 4429 262784
rect 4365 262724 4369 262780
rect 4369 262724 4425 262780
rect 4425 262724 4429 262780
rect 4365 262720 4429 262724
rect 4445 262780 4509 262784
rect 4445 262724 4449 262780
rect 4449 262724 4505 262780
rect 4505 262724 4509 262780
rect 4445 262720 4509 262724
rect 4525 262780 4589 262784
rect 4525 262724 4529 262780
rect 4529 262724 4585 262780
rect 4585 262724 4589 262780
rect 4525 262720 4589 262724
rect 7618 262780 7682 262784
rect 7618 262724 7622 262780
rect 7622 262724 7678 262780
rect 7678 262724 7682 262780
rect 7618 262720 7682 262724
rect 7698 262780 7762 262784
rect 7698 262724 7702 262780
rect 7702 262724 7758 262780
rect 7758 262724 7762 262780
rect 7698 262720 7762 262724
rect 7778 262780 7842 262784
rect 7778 262724 7782 262780
rect 7782 262724 7838 262780
rect 7838 262724 7842 262780
rect 7778 262720 7842 262724
rect 7858 262780 7922 262784
rect 7858 262724 7862 262780
rect 7862 262724 7918 262780
rect 7918 262724 7922 262780
rect 7858 262720 7922 262724
rect 2618 262236 2682 262240
rect 2618 262180 2622 262236
rect 2622 262180 2678 262236
rect 2678 262180 2682 262236
rect 2618 262176 2682 262180
rect 2698 262236 2762 262240
rect 2698 262180 2702 262236
rect 2702 262180 2758 262236
rect 2758 262180 2762 262236
rect 2698 262176 2762 262180
rect 2778 262236 2842 262240
rect 2778 262180 2782 262236
rect 2782 262180 2838 262236
rect 2838 262180 2842 262236
rect 2778 262176 2842 262180
rect 2858 262236 2922 262240
rect 2858 262180 2862 262236
rect 2862 262180 2918 262236
rect 2918 262180 2922 262236
rect 2858 262176 2922 262180
rect 5952 262236 6016 262240
rect 5952 262180 5956 262236
rect 5956 262180 6012 262236
rect 6012 262180 6016 262236
rect 5952 262176 6016 262180
rect 6032 262236 6096 262240
rect 6032 262180 6036 262236
rect 6036 262180 6092 262236
rect 6092 262180 6096 262236
rect 6032 262176 6096 262180
rect 6112 262236 6176 262240
rect 6112 262180 6116 262236
rect 6116 262180 6172 262236
rect 6172 262180 6176 262236
rect 6112 262176 6176 262180
rect 6192 262236 6256 262240
rect 6192 262180 6196 262236
rect 6196 262180 6252 262236
rect 6252 262180 6256 262236
rect 6192 262176 6256 262180
rect 4285 261692 4349 261696
rect 4285 261636 4289 261692
rect 4289 261636 4345 261692
rect 4345 261636 4349 261692
rect 4285 261632 4349 261636
rect 4365 261692 4429 261696
rect 4365 261636 4369 261692
rect 4369 261636 4425 261692
rect 4425 261636 4429 261692
rect 4365 261632 4429 261636
rect 4445 261692 4509 261696
rect 4445 261636 4449 261692
rect 4449 261636 4505 261692
rect 4505 261636 4509 261692
rect 4445 261632 4509 261636
rect 4525 261692 4589 261696
rect 4525 261636 4529 261692
rect 4529 261636 4585 261692
rect 4585 261636 4589 261692
rect 4525 261632 4589 261636
rect 7618 261692 7682 261696
rect 7618 261636 7622 261692
rect 7622 261636 7678 261692
rect 7678 261636 7682 261692
rect 7618 261632 7682 261636
rect 7698 261692 7762 261696
rect 7698 261636 7702 261692
rect 7702 261636 7758 261692
rect 7758 261636 7762 261692
rect 7698 261632 7762 261636
rect 7778 261692 7842 261696
rect 7778 261636 7782 261692
rect 7782 261636 7838 261692
rect 7838 261636 7842 261692
rect 7778 261632 7842 261636
rect 7858 261692 7922 261696
rect 7858 261636 7862 261692
rect 7862 261636 7918 261692
rect 7918 261636 7922 261692
rect 7858 261632 7922 261636
rect 2618 261148 2682 261152
rect 2618 261092 2622 261148
rect 2622 261092 2678 261148
rect 2678 261092 2682 261148
rect 2618 261088 2682 261092
rect 2698 261148 2762 261152
rect 2698 261092 2702 261148
rect 2702 261092 2758 261148
rect 2758 261092 2762 261148
rect 2698 261088 2762 261092
rect 2778 261148 2842 261152
rect 2778 261092 2782 261148
rect 2782 261092 2838 261148
rect 2838 261092 2842 261148
rect 2778 261088 2842 261092
rect 2858 261148 2922 261152
rect 2858 261092 2862 261148
rect 2862 261092 2918 261148
rect 2918 261092 2922 261148
rect 2858 261088 2922 261092
rect 5952 261148 6016 261152
rect 5952 261092 5956 261148
rect 5956 261092 6012 261148
rect 6012 261092 6016 261148
rect 5952 261088 6016 261092
rect 6032 261148 6096 261152
rect 6032 261092 6036 261148
rect 6036 261092 6092 261148
rect 6092 261092 6096 261148
rect 6032 261088 6096 261092
rect 6112 261148 6176 261152
rect 6112 261092 6116 261148
rect 6116 261092 6172 261148
rect 6172 261092 6176 261148
rect 6112 261088 6176 261092
rect 6192 261148 6256 261152
rect 6192 261092 6196 261148
rect 6196 261092 6252 261148
rect 6252 261092 6256 261148
rect 6192 261088 6256 261092
rect 4285 260604 4349 260608
rect 4285 260548 4289 260604
rect 4289 260548 4345 260604
rect 4345 260548 4349 260604
rect 4285 260544 4349 260548
rect 4365 260604 4429 260608
rect 4365 260548 4369 260604
rect 4369 260548 4425 260604
rect 4425 260548 4429 260604
rect 4365 260544 4429 260548
rect 4445 260604 4509 260608
rect 4445 260548 4449 260604
rect 4449 260548 4505 260604
rect 4505 260548 4509 260604
rect 4445 260544 4509 260548
rect 4525 260604 4589 260608
rect 4525 260548 4529 260604
rect 4529 260548 4585 260604
rect 4585 260548 4589 260604
rect 4525 260544 4589 260548
rect 7618 260604 7682 260608
rect 7618 260548 7622 260604
rect 7622 260548 7678 260604
rect 7678 260548 7682 260604
rect 7618 260544 7682 260548
rect 7698 260604 7762 260608
rect 7698 260548 7702 260604
rect 7702 260548 7758 260604
rect 7758 260548 7762 260604
rect 7698 260544 7762 260548
rect 7778 260604 7842 260608
rect 7778 260548 7782 260604
rect 7782 260548 7838 260604
rect 7838 260548 7842 260604
rect 7778 260544 7842 260548
rect 7858 260604 7922 260608
rect 7858 260548 7862 260604
rect 7862 260548 7918 260604
rect 7918 260548 7922 260604
rect 7858 260544 7922 260548
rect 2618 260060 2682 260064
rect 2618 260004 2622 260060
rect 2622 260004 2678 260060
rect 2678 260004 2682 260060
rect 2618 260000 2682 260004
rect 2698 260060 2762 260064
rect 2698 260004 2702 260060
rect 2702 260004 2758 260060
rect 2758 260004 2762 260060
rect 2698 260000 2762 260004
rect 2778 260060 2842 260064
rect 2778 260004 2782 260060
rect 2782 260004 2838 260060
rect 2838 260004 2842 260060
rect 2778 260000 2842 260004
rect 2858 260060 2922 260064
rect 2858 260004 2862 260060
rect 2862 260004 2918 260060
rect 2918 260004 2922 260060
rect 2858 260000 2922 260004
rect 5952 260060 6016 260064
rect 5952 260004 5956 260060
rect 5956 260004 6012 260060
rect 6012 260004 6016 260060
rect 5952 260000 6016 260004
rect 6032 260060 6096 260064
rect 6032 260004 6036 260060
rect 6036 260004 6092 260060
rect 6092 260004 6096 260060
rect 6032 260000 6096 260004
rect 6112 260060 6176 260064
rect 6112 260004 6116 260060
rect 6116 260004 6172 260060
rect 6172 260004 6176 260060
rect 6112 260000 6176 260004
rect 6192 260060 6256 260064
rect 6192 260004 6196 260060
rect 6196 260004 6252 260060
rect 6252 260004 6256 260060
rect 6192 260000 6256 260004
rect 4285 259516 4349 259520
rect 4285 259460 4289 259516
rect 4289 259460 4345 259516
rect 4345 259460 4349 259516
rect 4285 259456 4349 259460
rect 4365 259516 4429 259520
rect 4365 259460 4369 259516
rect 4369 259460 4425 259516
rect 4425 259460 4429 259516
rect 4365 259456 4429 259460
rect 4445 259516 4509 259520
rect 4445 259460 4449 259516
rect 4449 259460 4505 259516
rect 4505 259460 4509 259516
rect 4445 259456 4509 259460
rect 4525 259516 4589 259520
rect 4525 259460 4529 259516
rect 4529 259460 4585 259516
rect 4585 259460 4589 259516
rect 4525 259456 4589 259460
rect 7618 259516 7682 259520
rect 7618 259460 7622 259516
rect 7622 259460 7678 259516
rect 7678 259460 7682 259516
rect 7618 259456 7682 259460
rect 7698 259516 7762 259520
rect 7698 259460 7702 259516
rect 7702 259460 7758 259516
rect 7758 259460 7762 259516
rect 7698 259456 7762 259460
rect 7778 259516 7842 259520
rect 7778 259460 7782 259516
rect 7782 259460 7838 259516
rect 7838 259460 7842 259516
rect 7778 259456 7842 259460
rect 7858 259516 7922 259520
rect 7858 259460 7862 259516
rect 7862 259460 7918 259516
rect 7918 259460 7922 259516
rect 7858 259456 7922 259460
rect 2618 258972 2682 258976
rect 2618 258916 2622 258972
rect 2622 258916 2678 258972
rect 2678 258916 2682 258972
rect 2618 258912 2682 258916
rect 2698 258972 2762 258976
rect 2698 258916 2702 258972
rect 2702 258916 2758 258972
rect 2758 258916 2762 258972
rect 2698 258912 2762 258916
rect 2778 258972 2842 258976
rect 2778 258916 2782 258972
rect 2782 258916 2838 258972
rect 2838 258916 2842 258972
rect 2778 258912 2842 258916
rect 2858 258972 2922 258976
rect 2858 258916 2862 258972
rect 2862 258916 2918 258972
rect 2918 258916 2922 258972
rect 2858 258912 2922 258916
rect 5952 258972 6016 258976
rect 5952 258916 5956 258972
rect 5956 258916 6012 258972
rect 6012 258916 6016 258972
rect 5952 258912 6016 258916
rect 6032 258972 6096 258976
rect 6032 258916 6036 258972
rect 6036 258916 6092 258972
rect 6092 258916 6096 258972
rect 6032 258912 6096 258916
rect 6112 258972 6176 258976
rect 6112 258916 6116 258972
rect 6116 258916 6172 258972
rect 6172 258916 6176 258972
rect 6112 258912 6176 258916
rect 6192 258972 6256 258976
rect 6192 258916 6196 258972
rect 6196 258916 6252 258972
rect 6252 258916 6256 258972
rect 6192 258912 6256 258916
rect 4285 258428 4349 258432
rect 4285 258372 4289 258428
rect 4289 258372 4345 258428
rect 4345 258372 4349 258428
rect 4285 258368 4349 258372
rect 4365 258428 4429 258432
rect 4365 258372 4369 258428
rect 4369 258372 4425 258428
rect 4425 258372 4429 258428
rect 4365 258368 4429 258372
rect 4445 258428 4509 258432
rect 4445 258372 4449 258428
rect 4449 258372 4505 258428
rect 4505 258372 4509 258428
rect 4445 258368 4509 258372
rect 4525 258428 4589 258432
rect 4525 258372 4529 258428
rect 4529 258372 4585 258428
rect 4585 258372 4589 258428
rect 4525 258368 4589 258372
rect 7618 258428 7682 258432
rect 7618 258372 7622 258428
rect 7622 258372 7678 258428
rect 7678 258372 7682 258428
rect 7618 258368 7682 258372
rect 7698 258428 7762 258432
rect 7698 258372 7702 258428
rect 7702 258372 7758 258428
rect 7758 258372 7762 258428
rect 7698 258368 7762 258372
rect 7778 258428 7842 258432
rect 7778 258372 7782 258428
rect 7782 258372 7838 258428
rect 7838 258372 7842 258428
rect 7778 258368 7842 258372
rect 7858 258428 7922 258432
rect 7858 258372 7862 258428
rect 7862 258372 7918 258428
rect 7918 258372 7922 258428
rect 7858 258368 7922 258372
rect 2618 257884 2682 257888
rect 2618 257828 2622 257884
rect 2622 257828 2678 257884
rect 2678 257828 2682 257884
rect 2618 257824 2682 257828
rect 2698 257884 2762 257888
rect 2698 257828 2702 257884
rect 2702 257828 2758 257884
rect 2758 257828 2762 257884
rect 2698 257824 2762 257828
rect 2778 257884 2842 257888
rect 2778 257828 2782 257884
rect 2782 257828 2838 257884
rect 2838 257828 2842 257884
rect 2778 257824 2842 257828
rect 2858 257884 2922 257888
rect 2858 257828 2862 257884
rect 2862 257828 2918 257884
rect 2918 257828 2922 257884
rect 2858 257824 2922 257828
rect 5952 257884 6016 257888
rect 5952 257828 5956 257884
rect 5956 257828 6012 257884
rect 6012 257828 6016 257884
rect 5952 257824 6016 257828
rect 6032 257884 6096 257888
rect 6032 257828 6036 257884
rect 6036 257828 6092 257884
rect 6092 257828 6096 257884
rect 6032 257824 6096 257828
rect 6112 257884 6176 257888
rect 6112 257828 6116 257884
rect 6116 257828 6172 257884
rect 6172 257828 6176 257884
rect 6112 257824 6176 257828
rect 6192 257884 6256 257888
rect 6192 257828 6196 257884
rect 6196 257828 6252 257884
rect 6252 257828 6256 257884
rect 6192 257824 6256 257828
rect 4285 257340 4349 257344
rect 4285 257284 4289 257340
rect 4289 257284 4345 257340
rect 4345 257284 4349 257340
rect 4285 257280 4349 257284
rect 4365 257340 4429 257344
rect 4365 257284 4369 257340
rect 4369 257284 4425 257340
rect 4425 257284 4429 257340
rect 4365 257280 4429 257284
rect 4445 257340 4509 257344
rect 4445 257284 4449 257340
rect 4449 257284 4505 257340
rect 4505 257284 4509 257340
rect 4445 257280 4509 257284
rect 4525 257340 4589 257344
rect 4525 257284 4529 257340
rect 4529 257284 4585 257340
rect 4585 257284 4589 257340
rect 4525 257280 4589 257284
rect 7618 257340 7682 257344
rect 7618 257284 7622 257340
rect 7622 257284 7678 257340
rect 7678 257284 7682 257340
rect 7618 257280 7682 257284
rect 7698 257340 7762 257344
rect 7698 257284 7702 257340
rect 7702 257284 7758 257340
rect 7758 257284 7762 257340
rect 7698 257280 7762 257284
rect 7778 257340 7842 257344
rect 7778 257284 7782 257340
rect 7782 257284 7838 257340
rect 7838 257284 7842 257340
rect 7778 257280 7842 257284
rect 7858 257340 7922 257344
rect 7858 257284 7862 257340
rect 7862 257284 7918 257340
rect 7918 257284 7922 257340
rect 7858 257280 7922 257284
rect 2618 256796 2682 256800
rect 2618 256740 2622 256796
rect 2622 256740 2678 256796
rect 2678 256740 2682 256796
rect 2618 256736 2682 256740
rect 2698 256796 2762 256800
rect 2698 256740 2702 256796
rect 2702 256740 2758 256796
rect 2758 256740 2762 256796
rect 2698 256736 2762 256740
rect 2778 256796 2842 256800
rect 2778 256740 2782 256796
rect 2782 256740 2838 256796
rect 2838 256740 2842 256796
rect 2778 256736 2842 256740
rect 2858 256796 2922 256800
rect 2858 256740 2862 256796
rect 2862 256740 2918 256796
rect 2918 256740 2922 256796
rect 2858 256736 2922 256740
rect 5952 256796 6016 256800
rect 5952 256740 5956 256796
rect 5956 256740 6012 256796
rect 6012 256740 6016 256796
rect 5952 256736 6016 256740
rect 6032 256796 6096 256800
rect 6032 256740 6036 256796
rect 6036 256740 6092 256796
rect 6092 256740 6096 256796
rect 6032 256736 6096 256740
rect 6112 256796 6176 256800
rect 6112 256740 6116 256796
rect 6116 256740 6172 256796
rect 6172 256740 6176 256796
rect 6112 256736 6176 256740
rect 6192 256796 6256 256800
rect 6192 256740 6196 256796
rect 6196 256740 6252 256796
rect 6252 256740 6256 256796
rect 6192 256736 6256 256740
rect 4285 256252 4349 256256
rect 4285 256196 4289 256252
rect 4289 256196 4345 256252
rect 4345 256196 4349 256252
rect 4285 256192 4349 256196
rect 4365 256252 4429 256256
rect 4365 256196 4369 256252
rect 4369 256196 4425 256252
rect 4425 256196 4429 256252
rect 4365 256192 4429 256196
rect 4445 256252 4509 256256
rect 4445 256196 4449 256252
rect 4449 256196 4505 256252
rect 4505 256196 4509 256252
rect 4445 256192 4509 256196
rect 4525 256252 4589 256256
rect 4525 256196 4529 256252
rect 4529 256196 4585 256252
rect 4585 256196 4589 256252
rect 4525 256192 4589 256196
rect 7618 256252 7682 256256
rect 7618 256196 7622 256252
rect 7622 256196 7678 256252
rect 7678 256196 7682 256252
rect 7618 256192 7682 256196
rect 7698 256252 7762 256256
rect 7698 256196 7702 256252
rect 7702 256196 7758 256252
rect 7758 256196 7762 256252
rect 7698 256192 7762 256196
rect 7778 256252 7842 256256
rect 7778 256196 7782 256252
rect 7782 256196 7838 256252
rect 7838 256196 7842 256252
rect 7778 256192 7842 256196
rect 7858 256252 7922 256256
rect 7858 256196 7862 256252
rect 7862 256196 7918 256252
rect 7918 256196 7922 256252
rect 7858 256192 7922 256196
rect 2618 255708 2682 255712
rect 2618 255652 2622 255708
rect 2622 255652 2678 255708
rect 2678 255652 2682 255708
rect 2618 255648 2682 255652
rect 2698 255708 2762 255712
rect 2698 255652 2702 255708
rect 2702 255652 2758 255708
rect 2758 255652 2762 255708
rect 2698 255648 2762 255652
rect 2778 255708 2842 255712
rect 2778 255652 2782 255708
rect 2782 255652 2838 255708
rect 2838 255652 2842 255708
rect 2778 255648 2842 255652
rect 2858 255708 2922 255712
rect 2858 255652 2862 255708
rect 2862 255652 2918 255708
rect 2918 255652 2922 255708
rect 2858 255648 2922 255652
rect 5952 255708 6016 255712
rect 5952 255652 5956 255708
rect 5956 255652 6012 255708
rect 6012 255652 6016 255708
rect 5952 255648 6016 255652
rect 6032 255708 6096 255712
rect 6032 255652 6036 255708
rect 6036 255652 6092 255708
rect 6092 255652 6096 255708
rect 6032 255648 6096 255652
rect 6112 255708 6176 255712
rect 6112 255652 6116 255708
rect 6116 255652 6172 255708
rect 6172 255652 6176 255708
rect 6112 255648 6176 255652
rect 6192 255708 6256 255712
rect 6192 255652 6196 255708
rect 6196 255652 6252 255708
rect 6252 255652 6256 255708
rect 6192 255648 6256 255652
rect 4285 255164 4349 255168
rect 4285 255108 4289 255164
rect 4289 255108 4345 255164
rect 4345 255108 4349 255164
rect 4285 255104 4349 255108
rect 4365 255164 4429 255168
rect 4365 255108 4369 255164
rect 4369 255108 4425 255164
rect 4425 255108 4429 255164
rect 4365 255104 4429 255108
rect 4445 255164 4509 255168
rect 4445 255108 4449 255164
rect 4449 255108 4505 255164
rect 4505 255108 4509 255164
rect 4445 255104 4509 255108
rect 4525 255164 4589 255168
rect 4525 255108 4529 255164
rect 4529 255108 4585 255164
rect 4585 255108 4589 255164
rect 4525 255104 4589 255108
rect 7618 255164 7682 255168
rect 7618 255108 7622 255164
rect 7622 255108 7678 255164
rect 7678 255108 7682 255164
rect 7618 255104 7682 255108
rect 7698 255164 7762 255168
rect 7698 255108 7702 255164
rect 7702 255108 7758 255164
rect 7758 255108 7762 255164
rect 7698 255104 7762 255108
rect 7778 255164 7842 255168
rect 7778 255108 7782 255164
rect 7782 255108 7838 255164
rect 7838 255108 7842 255164
rect 7778 255104 7842 255108
rect 7858 255164 7922 255168
rect 7858 255108 7862 255164
rect 7862 255108 7918 255164
rect 7918 255108 7922 255164
rect 7858 255104 7922 255108
rect 2618 254620 2682 254624
rect 2618 254564 2622 254620
rect 2622 254564 2678 254620
rect 2678 254564 2682 254620
rect 2618 254560 2682 254564
rect 2698 254620 2762 254624
rect 2698 254564 2702 254620
rect 2702 254564 2758 254620
rect 2758 254564 2762 254620
rect 2698 254560 2762 254564
rect 2778 254620 2842 254624
rect 2778 254564 2782 254620
rect 2782 254564 2838 254620
rect 2838 254564 2842 254620
rect 2778 254560 2842 254564
rect 2858 254620 2922 254624
rect 2858 254564 2862 254620
rect 2862 254564 2918 254620
rect 2918 254564 2922 254620
rect 2858 254560 2922 254564
rect 5952 254620 6016 254624
rect 5952 254564 5956 254620
rect 5956 254564 6012 254620
rect 6012 254564 6016 254620
rect 5952 254560 6016 254564
rect 6032 254620 6096 254624
rect 6032 254564 6036 254620
rect 6036 254564 6092 254620
rect 6092 254564 6096 254620
rect 6032 254560 6096 254564
rect 6112 254620 6176 254624
rect 6112 254564 6116 254620
rect 6116 254564 6172 254620
rect 6172 254564 6176 254620
rect 6112 254560 6176 254564
rect 6192 254620 6256 254624
rect 6192 254564 6196 254620
rect 6196 254564 6252 254620
rect 6252 254564 6256 254620
rect 6192 254560 6256 254564
rect 4285 254076 4349 254080
rect 4285 254020 4289 254076
rect 4289 254020 4345 254076
rect 4345 254020 4349 254076
rect 4285 254016 4349 254020
rect 4365 254076 4429 254080
rect 4365 254020 4369 254076
rect 4369 254020 4425 254076
rect 4425 254020 4429 254076
rect 4365 254016 4429 254020
rect 4445 254076 4509 254080
rect 4445 254020 4449 254076
rect 4449 254020 4505 254076
rect 4505 254020 4509 254076
rect 4445 254016 4509 254020
rect 4525 254076 4589 254080
rect 4525 254020 4529 254076
rect 4529 254020 4585 254076
rect 4585 254020 4589 254076
rect 4525 254016 4589 254020
rect 7618 254076 7682 254080
rect 7618 254020 7622 254076
rect 7622 254020 7678 254076
rect 7678 254020 7682 254076
rect 7618 254016 7682 254020
rect 7698 254076 7762 254080
rect 7698 254020 7702 254076
rect 7702 254020 7758 254076
rect 7758 254020 7762 254076
rect 7698 254016 7762 254020
rect 7778 254076 7842 254080
rect 7778 254020 7782 254076
rect 7782 254020 7838 254076
rect 7838 254020 7842 254076
rect 7778 254016 7842 254020
rect 7858 254076 7922 254080
rect 7858 254020 7862 254076
rect 7862 254020 7918 254076
rect 7918 254020 7922 254076
rect 7858 254016 7922 254020
rect 2618 253532 2682 253536
rect 2618 253476 2622 253532
rect 2622 253476 2678 253532
rect 2678 253476 2682 253532
rect 2618 253472 2682 253476
rect 2698 253532 2762 253536
rect 2698 253476 2702 253532
rect 2702 253476 2758 253532
rect 2758 253476 2762 253532
rect 2698 253472 2762 253476
rect 2778 253532 2842 253536
rect 2778 253476 2782 253532
rect 2782 253476 2838 253532
rect 2838 253476 2842 253532
rect 2778 253472 2842 253476
rect 2858 253532 2922 253536
rect 2858 253476 2862 253532
rect 2862 253476 2918 253532
rect 2918 253476 2922 253532
rect 2858 253472 2922 253476
rect 5952 253532 6016 253536
rect 5952 253476 5956 253532
rect 5956 253476 6012 253532
rect 6012 253476 6016 253532
rect 5952 253472 6016 253476
rect 6032 253532 6096 253536
rect 6032 253476 6036 253532
rect 6036 253476 6092 253532
rect 6092 253476 6096 253532
rect 6032 253472 6096 253476
rect 6112 253532 6176 253536
rect 6112 253476 6116 253532
rect 6116 253476 6172 253532
rect 6172 253476 6176 253532
rect 6112 253472 6176 253476
rect 6192 253532 6256 253536
rect 6192 253476 6196 253532
rect 6196 253476 6252 253532
rect 6252 253476 6256 253532
rect 6192 253472 6256 253476
rect 4285 252988 4349 252992
rect 4285 252932 4289 252988
rect 4289 252932 4345 252988
rect 4345 252932 4349 252988
rect 4285 252928 4349 252932
rect 4365 252988 4429 252992
rect 4365 252932 4369 252988
rect 4369 252932 4425 252988
rect 4425 252932 4429 252988
rect 4365 252928 4429 252932
rect 4445 252988 4509 252992
rect 4445 252932 4449 252988
rect 4449 252932 4505 252988
rect 4505 252932 4509 252988
rect 4445 252928 4509 252932
rect 4525 252988 4589 252992
rect 4525 252932 4529 252988
rect 4529 252932 4585 252988
rect 4585 252932 4589 252988
rect 4525 252928 4589 252932
rect 7618 252988 7682 252992
rect 7618 252932 7622 252988
rect 7622 252932 7678 252988
rect 7678 252932 7682 252988
rect 7618 252928 7682 252932
rect 7698 252988 7762 252992
rect 7698 252932 7702 252988
rect 7702 252932 7758 252988
rect 7758 252932 7762 252988
rect 7698 252928 7762 252932
rect 7778 252988 7842 252992
rect 7778 252932 7782 252988
rect 7782 252932 7838 252988
rect 7838 252932 7842 252988
rect 7778 252928 7842 252932
rect 7858 252988 7922 252992
rect 7858 252932 7862 252988
rect 7862 252932 7918 252988
rect 7918 252932 7922 252988
rect 7858 252928 7922 252932
rect 2618 252444 2682 252448
rect 2618 252388 2622 252444
rect 2622 252388 2678 252444
rect 2678 252388 2682 252444
rect 2618 252384 2682 252388
rect 2698 252444 2762 252448
rect 2698 252388 2702 252444
rect 2702 252388 2758 252444
rect 2758 252388 2762 252444
rect 2698 252384 2762 252388
rect 2778 252444 2842 252448
rect 2778 252388 2782 252444
rect 2782 252388 2838 252444
rect 2838 252388 2842 252444
rect 2778 252384 2842 252388
rect 2858 252444 2922 252448
rect 2858 252388 2862 252444
rect 2862 252388 2918 252444
rect 2918 252388 2922 252444
rect 2858 252384 2922 252388
rect 5952 252444 6016 252448
rect 5952 252388 5956 252444
rect 5956 252388 6012 252444
rect 6012 252388 6016 252444
rect 5952 252384 6016 252388
rect 6032 252444 6096 252448
rect 6032 252388 6036 252444
rect 6036 252388 6092 252444
rect 6092 252388 6096 252444
rect 6032 252384 6096 252388
rect 6112 252444 6176 252448
rect 6112 252388 6116 252444
rect 6116 252388 6172 252444
rect 6172 252388 6176 252444
rect 6112 252384 6176 252388
rect 6192 252444 6256 252448
rect 6192 252388 6196 252444
rect 6196 252388 6252 252444
rect 6252 252388 6256 252444
rect 6192 252384 6256 252388
rect 4285 251900 4349 251904
rect 4285 251844 4289 251900
rect 4289 251844 4345 251900
rect 4345 251844 4349 251900
rect 4285 251840 4349 251844
rect 4365 251900 4429 251904
rect 4365 251844 4369 251900
rect 4369 251844 4425 251900
rect 4425 251844 4429 251900
rect 4365 251840 4429 251844
rect 4445 251900 4509 251904
rect 4445 251844 4449 251900
rect 4449 251844 4505 251900
rect 4505 251844 4509 251900
rect 4445 251840 4509 251844
rect 4525 251900 4589 251904
rect 4525 251844 4529 251900
rect 4529 251844 4585 251900
rect 4585 251844 4589 251900
rect 4525 251840 4589 251844
rect 7618 251900 7682 251904
rect 7618 251844 7622 251900
rect 7622 251844 7678 251900
rect 7678 251844 7682 251900
rect 7618 251840 7682 251844
rect 7698 251900 7762 251904
rect 7698 251844 7702 251900
rect 7702 251844 7758 251900
rect 7758 251844 7762 251900
rect 7698 251840 7762 251844
rect 7778 251900 7842 251904
rect 7778 251844 7782 251900
rect 7782 251844 7838 251900
rect 7838 251844 7842 251900
rect 7778 251840 7842 251844
rect 7858 251900 7922 251904
rect 7858 251844 7862 251900
rect 7862 251844 7918 251900
rect 7918 251844 7922 251900
rect 7858 251840 7922 251844
rect 2618 251356 2682 251360
rect 2618 251300 2622 251356
rect 2622 251300 2678 251356
rect 2678 251300 2682 251356
rect 2618 251296 2682 251300
rect 2698 251356 2762 251360
rect 2698 251300 2702 251356
rect 2702 251300 2758 251356
rect 2758 251300 2762 251356
rect 2698 251296 2762 251300
rect 2778 251356 2842 251360
rect 2778 251300 2782 251356
rect 2782 251300 2838 251356
rect 2838 251300 2842 251356
rect 2778 251296 2842 251300
rect 2858 251356 2922 251360
rect 2858 251300 2862 251356
rect 2862 251300 2918 251356
rect 2918 251300 2922 251356
rect 2858 251296 2922 251300
rect 5952 251356 6016 251360
rect 5952 251300 5956 251356
rect 5956 251300 6012 251356
rect 6012 251300 6016 251356
rect 5952 251296 6016 251300
rect 6032 251356 6096 251360
rect 6032 251300 6036 251356
rect 6036 251300 6092 251356
rect 6092 251300 6096 251356
rect 6032 251296 6096 251300
rect 6112 251356 6176 251360
rect 6112 251300 6116 251356
rect 6116 251300 6172 251356
rect 6172 251300 6176 251356
rect 6112 251296 6176 251300
rect 6192 251356 6256 251360
rect 6192 251300 6196 251356
rect 6196 251300 6252 251356
rect 6252 251300 6256 251356
rect 6192 251296 6256 251300
rect 4285 250812 4349 250816
rect 4285 250756 4289 250812
rect 4289 250756 4345 250812
rect 4345 250756 4349 250812
rect 4285 250752 4349 250756
rect 4365 250812 4429 250816
rect 4365 250756 4369 250812
rect 4369 250756 4425 250812
rect 4425 250756 4429 250812
rect 4365 250752 4429 250756
rect 4445 250812 4509 250816
rect 4445 250756 4449 250812
rect 4449 250756 4505 250812
rect 4505 250756 4509 250812
rect 4445 250752 4509 250756
rect 4525 250812 4589 250816
rect 4525 250756 4529 250812
rect 4529 250756 4585 250812
rect 4585 250756 4589 250812
rect 4525 250752 4589 250756
rect 7618 250812 7682 250816
rect 7618 250756 7622 250812
rect 7622 250756 7678 250812
rect 7678 250756 7682 250812
rect 7618 250752 7682 250756
rect 7698 250812 7762 250816
rect 7698 250756 7702 250812
rect 7702 250756 7758 250812
rect 7758 250756 7762 250812
rect 7698 250752 7762 250756
rect 7778 250812 7842 250816
rect 7778 250756 7782 250812
rect 7782 250756 7838 250812
rect 7838 250756 7842 250812
rect 7778 250752 7842 250756
rect 7858 250812 7922 250816
rect 7858 250756 7862 250812
rect 7862 250756 7918 250812
rect 7918 250756 7922 250812
rect 7858 250752 7922 250756
rect 2618 250268 2682 250272
rect 2618 250212 2622 250268
rect 2622 250212 2678 250268
rect 2678 250212 2682 250268
rect 2618 250208 2682 250212
rect 2698 250268 2762 250272
rect 2698 250212 2702 250268
rect 2702 250212 2758 250268
rect 2758 250212 2762 250268
rect 2698 250208 2762 250212
rect 2778 250268 2842 250272
rect 2778 250212 2782 250268
rect 2782 250212 2838 250268
rect 2838 250212 2842 250268
rect 2778 250208 2842 250212
rect 2858 250268 2922 250272
rect 2858 250212 2862 250268
rect 2862 250212 2918 250268
rect 2918 250212 2922 250268
rect 2858 250208 2922 250212
rect 5952 250268 6016 250272
rect 5952 250212 5956 250268
rect 5956 250212 6012 250268
rect 6012 250212 6016 250268
rect 5952 250208 6016 250212
rect 6032 250268 6096 250272
rect 6032 250212 6036 250268
rect 6036 250212 6092 250268
rect 6092 250212 6096 250268
rect 6032 250208 6096 250212
rect 6112 250268 6176 250272
rect 6112 250212 6116 250268
rect 6116 250212 6172 250268
rect 6172 250212 6176 250268
rect 6112 250208 6176 250212
rect 6192 250268 6256 250272
rect 6192 250212 6196 250268
rect 6196 250212 6252 250268
rect 6252 250212 6256 250268
rect 6192 250208 6256 250212
rect 4285 249724 4349 249728
rect 4285 249668 4289 249724
rect 4289 249668 4345 249724
rect 4345 249668 4349 249724
rect 4285 249664 4349 249668
rect 4365 249724 4429 249728
rect 4365 249668 4369 249724
rect 4369 249668 4425 249724
rect 4425 249668 4429 249724
rect 4365 249664 4429 249668
rect 4445 249724 4509 249728
rect 4445 249668 4449 249724
rect 4449 249668 4505 249724
rect 4505 249668 4509 249724
rect 4445 249664 4509 249668
rect 4525 249724 4589 249728
rect 4525 249668 4529 249724
rect 4529 249668 4585 249724
rect 4585 249668 4589 249724
rect 4525 249664 4589 249668
rect 7618 249724 7682 249728
rect 7618 249668 7622 249724
rect 7622 249668 7678 249724
rect 7678 249668 7682 249724
rect 7618 249664 7682 249668
rect 7698 249724 7762 249728
rect 7698 249668 7702 249724
rect 7702 249668 7758 249724
rect 7758 249668 7762 249724
rect 7698 249664 7762 249668
rect 7778 249724 7842 249728
rect 7778 249668 7782 249724
rect 7782 249668 7838 249724
rect 7838 249668 7842 249724
rect 7778 249664 7842 249668
rect 7858 249724 7922 249728
rect 7858 249668 7862 249724
rect 7862 249668 7918 249724
rect 7918 249668 7922 249724
rect 7858 249664 7922 249668
rect 2618 249180 2682 249184
rect 2618 249124 2622 249180
rect 2622 249124 2678 249180
rect 2678 249124 2682 249180
rect 2618 249120 2682 249124
rect 2698 249180 2762 249184
rect 2698 249124 2702 249180
rect 2702 249124 2758 249180
rect 2758 249124 2762 249180
rect 2698 249120 2762 249124
rect 2778 249180 2842 249184
rect 2778 249124 2782 249180
rect 2782 249124 2838 249180
rect 2838 249124 2842 249180
rect 2778 249120 2842 249124
rect 2858 249180 2922 249184
rect 2858 249124 2862 249180
rect 2862 249124 2918 249180
rect 2918 249124 2922 249180
rect 2858 249120 2922 249124
rect 5952 249180 6016 249184
rect 5952 249124 5956 249180
rect 5956 249124 6012 249180
rect 6012 249124 6016 249180
rect 5952 249120 6016 249124
rect 6032 249180 6096 249184
rect 6032 249124 6036 249180
rect 6036 249124 6092 249180
rect 6092 249124 6096 249180
rect 6032 249120 6096 249124
rect 6112 249180 6176 249184
rect 6112 249124 6116 249180
rect 6116 249124 6172 249180
rect 6172 249124 6176 249180
rect 6112 249120 6176 249124
rect 6192 249180 6256 249184
rect 6192 249124 6196 249180
rect 6196 249124 6252 249180
rect 6252 249124 6256 249180
rect 6192 249120 6256 249124
rect 4285 248636 4349 248640
rect 4285 248580 4289 248636
rect 4289 248580 4345 248636
rect 4345 248580 4349 248636
rect 4285 248576 4349 248580
rect 4365 248636 4429 248640
rect 4365 248580 4369 248636
rect 4369 248580 4425 248636
rect 4425 248580 4429 248636
rect 4365 248576 4429 248580
rect 4445 248636 4509 248640
rect 4445 248580 4449 248636
rect 4449 248580 4505 248636
rect 4505 248580 4509 248636
rect 4445 248576 4509 248580
rect 4525 248636 4589 248640
rect 4525 248580 4529 248636
rect 4529 248580 4585 248636
rect 4585 248580 4589 248636
rect 4525 248576 4589 248580
rect 7618 248636 7682 248640
rect 7618 248580 7622 248636
rect 7622 248580 7678 248636
rect 7678 248580 7682 248636
rect 7618 248576 7682 248580
rect 7698 248636 7762 248640
rect 7698 248580 7702 248636
rect 7702 248580 7758 248636
rect 7758 248580 7762 248636
rect 7698 248576 7762 248580
rect 7778 248636 7842 248640
rect 7778 248580 7782 248636
rect 7782 248580 7838 248636
rect 7838 248580 7842 248636
rect 7778 248576 7842 248580
rect 7858 248636 7922 248640
rect 7858 248580 7862 248636
rect 7862 248580 7918 248636
rect 7918 248580 7922 248636
rect 7858 248576 7922 248580
rect 2618 248092 2682 248096
rect 2618 248036 2622 248092
rect 2622 248036 2678 248092
rect 2678 248036 2682 248092
rect 2618 248032 2682 248036
rect 2698 248092 2762 248096
rect 2698 248036 2702 248092
rect 2702 248036 2758 248092
rect 2758 248036 2762 248092
rect 2698 248032 2762 248036
rect 2778 248092 2842 248096
rect 2778 248036 2782 248092
rect 2782 248036 2838 248092
rect 2838 248036 2842 248092
rect 2778 248032 2842 248036
rect 2858 248092 2922 248096
rect 2858 248036 2862 248092
rect 2862 248036 2918 248092
rect 2918 248036 2922 248092
rect 2858 248032 2922 248036
rect 5952 248092 6016 248096
rect 5952 248036 5956 248092
rect 5956 248036 6012 248092
rect 6012 248036 6016 248092
rect 5952 248032 6016 248036
rect 6032 248092 6096 248096
rect 6032 248036 6036 248092
rect 6036 248036 6092 248092
rect 6092 248036 6096 248092
rect 6032 248032 6096 248036
rect 6112 248092 6176 248096
rect 6112 248036 6116 248092
rect 6116 248036 6172 248092
rect 6172 248036 6176 248092
rect 6112 248032 6176 248036
rect 6192 248092 6256 248096
rect 6192 248036 6196 248092
rect 6196 248036 6252 248092
rect 6252 248036 6256 248092
rect 6192 248032 6256 248036
rect 4285 247548 4349 247552
rect 4285 247492 4289 247548
rect 4289 247492 4345 247548
rect 4345 247492 4349 247548
rect 4285 247488 4349 247492
rect 4365 247548 4429 247552
rect 4365 247492 4369 247548
rect 4369 247492 4425 247548
rect 4425 247492 4429 247548
rect 4365 247488 4429 247492
rect 4445 247548 4509 247552
rect 4445 247492 4449 247548
rect 4449 247492 4505 247548
rect 4505 247492 4509 247548
rect 4445 247488 4509 247492
rect 4525 247548 4589 247552
rect 4525 247492 4529 247548
rect 4529 247492 4585 247548
rect 4585 247492 4589 247548
rect 4525 247488 4589 247492
rect 7618 247548 7682 247552
rect 7618 247492 7622 247548
rect 7622 247492 7678 247548
rect 7678 247492 7682 247548
rect 7618 247488 7682 247492
rect 7698 247548 7762 247552
rect 7698 247492 7702 247548
rect 7702 247492 7758 247548
rect 7758 247492 7762 247548
rect 7698 247488 7762 247492
rect 7778 247548 7842 247552
rect 7778 247492 7782 247548
rect 7782 247492 7838 247548
rect 7838 247492 7842 247548
rect 7778 247488 7842 247492
rect 7858 247548 7922 247552
rect 7858 247492 7862 247548
rect 7862 247492 7918 247548
rect 7918 247492 7922 247548
rect 7858 247488 7922 247492
rect 2618 247004 2682 247008
rect 2618 246948 2622 247004
rect 2622 246948 2678 247004
rect 2678 246948 2682 247004
rect 2618 246944 2682 246948
rect 2698 247004 2762 247008
rect 2698 246948 2702 247004
rect 2702 246948 2758 247004
rect 2758 246948 2762 247004
rect 2698 246944 2762 246948
rect 2778 247004 2842 247008
rect 2778 246948 2782 247004
rect 2782 246948 2838 247004
rect 2838 246948 2842 247004
rect 2778 246944 2842 246948
rect 2858 247004 2922 247008
rect 2858 246948 2862 247004
rect 2862 246948 2918 247004
rect 2918 246948 2922 247004
rect 2858 246944 2922 246948
rect 5952 247004 6016 247008
rect 5952 246948 5956 247004
rect 5956 246948 6012 247004
rect 6012 246948 6016 247004
rect 5952 246944 6016 246948
rect 6032 247004 6096 247008
rect 6032 246948 6036 247004
rect 6036 246948 6092 247004
rect 6092 246948 6096 247004
rect 6032 246944 6096 246948
rect 6112 247004 6176 247008
rect 6112 246948 6116 247004
rect 6116 246948 6172 247004
rect 6172 246948 6176 247004
rect 6112 246944 6176 246948
rect 6192 247004 6256 247008
rect 6192 246948 6196 247004
rect 6196 246948 6252 247004
rect 6252 246948 6256 247004
rect 6192 246944 6256 246948
rect 4285 246460 4349 246464
rect 4285 246404 4289 246460
rect 4289 246404 4345 246460
rect 4345 246404 4349 246460
rect 4285 246400 4349 246404
rect 4365 246460 4429 246464
rect 4365 246404 4369 246460
rect 4369 246404 4425 246460
rect 4425 246404 4429 246460
rect 4365 246400 4429 246404
rect 4445 246460 4509 246464
rect 4445 246404 4449 246460
rect 4449 246404 4505 246460
rect 4505 246404 4509 246460
rect 4445 246400 4509 246404
rect 4525 246460 4589 246464
rect 4525 246404 4529 246460
rect 4529 246404 4585 246460
rect 4585 246404 4589 246460
rect 4525 246400 4589 246404
rect 7618 246460 7682 246464
rect 7618 246404 7622 246460
rect 7622 246404 7678 246460
rect 7678 246404 7682 246460
rect 7618 246400 7682 246404
rect 7698 246460 7762 246464
rect 7698 246404 7702 246460
rect 7702 246404 7758 246460
rect 7758 246404 7762 246460
rect 7698 246400 7762 246404
rect 7778 246460 7842 246464
rect 7778 246404 7782 246460
rect 7782 246404 7838 246460
rect 7838 246404 7842 246460
rect 7778 246400 7842 246404
rect 7858 246460 7922 246464
rect 7858 246404 7862 246460
rect 7862 246404 7918 246460
rect 7918 246404 7922 246460
rect 7858 246400 7922 246404
rect 2618 245916 2682 245920
rect 2618 245860 2622 245916
rect 2622 245860 2678 245916
rect 2678 245860 2682 245916
rect 2618 245856 2682 245860
rect 2698 245916 2762 245920
rect 2698 245860 2702 245916
rect 2702 245860 2758 245916
rect 2758 245860 2762 245916
rect 2698 245856 2762 245860
rect 2778 245916 2842 245920
rect 2778 245860 2782 245916
rect 2782 245860 2838 245916
rect 2838 245860 2842 245916
rect 2778 245856 2842 245860
rect 2858 245916 2922 245920
rect 2858 245860 2862 245916
rect 2862 245860 2918 245916
rect 2918 245860 2922 245916
rect 2858 245856 2922 245860
rect 5952 245916 6016 245920
rect 5952 245860 5956 245916
rect 5956 245860 6012 245916
rect 6012 245860 6016 245916
rect 5952 245856 6016 245860
rect 6032 245916 6096 245920
rect 6032 245860 6036 245916
rect 6036 245860 6092 245916
rect 6092 245860 6096 245916
rect 6032 245856 6096 245860
rect 6112 245916 6176 245920
rect 6112 245860 6116 245916
rect 6116 245860 6172 245916
rect 6172 245860 6176 245916
rect 6112 245856 6176 245860
rect 6192 245916 6256 245920
rect 6192 245860 6196 245916
rect 6196 245860 6252 245916
rect 6252 245860 6256 245916
rect 6192 245856 6256 245860
rect 4285 245372 4349 245376
rect 4285 245316 4289 245372
rect 4289 245316 4345 245372
rect 4345 245316 4349 245372
rect 4285 245312 4349 245316
rect 4365 245372 4429 245376
rect 4365 245316 4369 245372
rect 4369 245316 4425 245372
rect 4425 245316 4429 245372
rect 4365 245312 4429 245316
rect 4445 245372 4509 245376
rect 4445 245316 4449 245372
rect 4449 245316 4505 245372
rect 4505 245316 4509 245372
rect 4445 245312 4509 245316
rect 4525 245372 4589 245376
rect 4525 245316 4529 245372
rect 4529 245316 4585 245372
rect 4585 245316 4589 245372
rect 4525 245312 4589 245316
rect 7618 245372 7682 245376
rect 7618 245316 7622 245372
rect 7622 245316 7678 245372
rect 7678 245316 7682 245372
rect 7618 245312 7682 245316
rect 7698 245372 7762 245376
rect 7698 245316 7702 245372
rect 7702 245316 7758 245372
rect 7758 245316 7762 245372
rect 7698 245312 7762 245316
rect 7778 245372 7842 245376
rect 7778 245316 7782 245372
rect 7782 245316 7838 245372
rect 7838 245316 7842 245372
rect 7778 245312 7842 245316
rect 7858 245372 7922 245376
rect 7858 245316 7862 245372
rect 7862 245316 7918 245372
rect 7918 245316 7922 245372
rect 7858 245312 7922 245316
rect 2618 244828 2682 244832
rect 2618 244772 2622 244828
rect 2622 244772 2678 244828
rect 2678 244772 2682 244828
rect 2618 244768 2682 244772
rect 2698 244828 2762 244832
rect 2698 244772 2702 244828
rect 2702 244772 2758 244828
rect 2758 244772 2762 244828
rect 2698 244768 2762 244772
rect 2778 244828 2842 244832
rect 2778 244772 2782 244828
rect 2782 244772 2838 244828
rect 2838 244772 2842 244828
rect 2778 244768 2842 244772
rect 2858 244828 2922 244832
rect 2858 244772 2862 244828
rect 2862 244772 2918 244828
rect 2918 244772 2922 244828
rect 2858 244768 2922 244772
rect 5952 244828 6016 244832
rect 5952 244772 5956 244828
rect 5956 244772 6012 244828
rect 6012 244772 6016 244828
rect 5952 244768 6016 244772
rect 6032 244828 6096 244832
rect 6032 244772 6036 244828
rect 6036 244772 6092 244828
rect 6092 244772 6096 244828
rect 6032 244768 6096 244772
rect 6112 244828 6176 244832
rect 6112 244772 6116 244828
rect 6116 244772 6172 244828
rect 6172 244772 6176 244828
rect 6112 244768 6176 244772
rect 6192 244828 6256 244832
rect 6192 244772 6196 244828
rect 6196 244772 6252 244828
rect 6252 244772 6256 244828
rect 6192 244768 6256 244772
rect 4285 244284 4349 244288
rect 4285 244228 4289 244284
rect 4289 244228 4345 244284
rect 4345 244228 4349 244284
rect 4285 244224 4349 244228
rect 4365 244284 4429 244288
rect 4365 244228 4369 244284
rect 4369 244228 4425 244284
rect 4425 244228 4429 244284
rect 4365 244224 4429 244228
rect 4445 244284 4509 244288
rect 4445 244228 4449 244284
rect 4449 244228 4505 244284
rect 4505 244228 4509 244284
rect 4445 244224 4509 244228
rect 4525 244284 4589 244288
rect 4525 244228 4529 244284
rect 4529 244228 4585 244284
rect 4585 244228 4589 244284
rect 4525 244224 4589 244228
rect 7618 244284 7682 244288
rect 7618 244228 7622 244284
rect 7622 244228 7678 244284
rect 7678 244228 7682 244284
rect 7618 244224 7682 244228
rect 7698 244284 7762 244288
rect 7698 244228 7702 244284
rect 7702 244228 7758 244284
rect 7758 244228 7762 244284
rect 7698 244224 7762 244228
rect 7778 244284 7842 244288
rect 7778 244228 7782 244284
rect 7782 244228 7838 244284
rect 7838 244228 7842 244284
rect 7778 244224 7842 244228
rect 7858 244284 7922 244288
rect 7858 244228 7862 244284
rect 7862 244228 7918 244284
rect 7918 244228 7922 244284
rect 7858 244224 7922 244228
rect 2618 243740 2682 243744
rect 2618 243684 2622 243740
rect 2622 243684 2678 243740
rect 2678 243684 2682 243740
rect 2618 243680 2682 243684
rect 2698 243740 2762 243744
rect 2698 243684 2702 243740
rect 2702 243684 2758 243740
rect 2758 243684 2762 243740
rect 2698 243680 2762 243684
rect 2778 243740 2842 243744
rect 2778 243684 2782 243740
rect 2782 243684 2838 243740
rect 2838 243684 2842 243740
rect 2778 243680 2842 243684
rect 2858 243740 2922 243744
rect 2858 243684 2862 243740
rect 2862 243684 2918 243740
rect 2918 243684 2922 243740
rect 2858 243680 2922 243684
rect 5952 243740 6016 243744
rect 5952 243684 5956 243740
rect 5956 243684 6012 243740
rect 6012 243684 6016 243740
rect 5952 243680 6016 243684
rect 6032 243740 6096 243744
rect 6032 243684 6036 243740
rect 6036 243684 6092 243740
rect 6092 243684 6096 243740
rect 6032 243680 6096 243684
rect 6112 243740 6176 243744
rect 6112 243684 6116 243740
rect 6116 243684 6172 243740
rect 6172 243684 6176 243740
rect 6112 243680 6176 243684
rect 6192 243740 6256 243744
rect 6192 243684 6196 243740
rect 6196 243684 6252 243740
rect 6252 243684 6256 243740
rect 6192 243680 6256 243684
rect 4285 243196 4349 243200
rect 4285 243140 4289 243196
rect 4289 243140 4345 243196
rect 4345 243140 4349 243196
rect 4285 243136 4349 243140
rect 4365 243196 4429 243200
rect 4365 243140 4369 243196
rect 4369 243140 4425 243196
rect 4425 243140 4429 243196
rect 4365 243136 4429 243140
rect 4445 243196 4509 243200
rect 4445 243140 4449 243196
rect 4449 243140 4505 243196
rect 4505 243140 4509 243196
rect 4445 243136 4509 243140
rect 4525 243196 4589 243200
rect 4525 243140 4529 243196
rect 4529 243140 4585 243196
rect 4585 243140 4589 243196
rect 4525 243136 4589 243140
rect 7618 243196 7682 243200
rect 7618 243140 7622 243196
rect 7622 243140 7678 243196
rect 7678 243140 7682 243196
rect 7618 243136 7682 243140
rect 7698 243196 7762 243200
rect 7698 243140 7702 243196
rect 7702 243140 7758 243196
rect 7758 243140 7762 243196
rect 7698 243136 7762 243140
rect 7778 243196 7842 243200
rect 7778 243140 7782 243196
rect 7782 243140 7838 243196
rect 7838 243140 7842 243196
rect 7778 243136 7842 243140
rect 7858 243196 7922 243200
rect 7858 243140 7862 243196
rect 7862 243140 7918 243196
rect 7918 243140 7922 243196
rect 7858 243136 7922 243140
rect 2618 242652 2682 242656
rect 2618 242596 2622 242652
rect 2622 242596 2678 242652
rect 2678 242596 2682 242652
rect 2618 242592 2682 242596
rect 2698 242652 2762 242656
rect 2698 242596 2702 242652
rect 2702 242596 2758 242652
rect 2758 242596 2762 242652
rect 2698 242592 2762 242596
rect 2778 242652 2842 242656
rect 2778 242596 2782 242652
rect 2782 242596 2838 242652
rect 2838 242596 2842 242652
rect 2778 242592 2842 242596
rect 2858 242652 2922 242656
rect 2858 242596 2862 242652
rect 2862 242596 2918 242652
rect 2918 242596 2922 242652
rect 2858 242592 2922 242596
rect 5952 242652 6016 242656
rect 5952 242596 5956 242652
rect 5956 242596 6012 242652
rect 6012 242596 6016 242652
rect 5952 242592 6016 242596
rect 6032 242652 6096 242656
rect 6032 242596 6036 242652
rect 6036 242596 6092 242652
rect 6092 242596 6096 242652
rect 6032 242592 6096 242596
rect 6112 242652 6176 242656
rect 6112 242596 6116 242652
rect 6116 242596 6172 242652
rect 6172 242596 6176 242652
rect 6112 242592 6176 242596
rect 6192 242652 6256 242656
rect 6192 242596 6196 242652
rect 6196 242596 6252 242652
rect 6252 242596 6256 242652
rect 6192 242592 6256 242596
rect 4285 242108 4349 242112
rect 4285 242052 4289 242108
rect 4289 242052 4345 242108
rect 4345 242052 4349 242108
rect 4285 242048 4349 242052
rect 4365 242108 4429 242112
rect 4365 242052 4369 242108
rect 4369 242052 4425 242108
rect 4425 242052 4429 242108
rect 4365 242048 4429 242052
rect 4445 242108 4509 242112
rect 4445 242052 4449 242108
rect 4449 242052 4505 242108
rect 4505 242052 4509 242108
rect 4445 242048 4509 242052
rect 4525 242108 4589 242112
rect 4525 242052 4529 242108
rect 4529 242052 4585 242108
rect 4585 242052 4589 242108
rect 4525 242048 4589 242052
rect 7618 242108 7682 242112
rect 7618 242052 7622 242108
rect 7622 242052 7678 242108
rect 7678 242052 7682 242108
rect 7618 242048 7682 242052
rect 7698 242108 7762 242112
rect 7698 242052 7702 242108
rect 7702 242052 7758 242108
rect 7758 242052 7762 242108
rect 7698 242048 7762 242052
rect 7778 242108 7842 242112
rect 7778 242052 7782 242108
rect 7782 242052 7838 242108
rect 7838 242052 7842 242108
rect 7778 242048 7842 242052
rect 7858 242108 7922 242112
rect 7858 242052 7862 242108
rect 7862 242052 7918 242108
rect 7918 242052 7922 242108
rect 7858 242048 7922 242052
rect 2618 241564 2682 241568
rect 2618 241508 2622 241564
rect 2622 241508 2678 241564
rect 2678 241508 2682 241564
rect 2618 241504 2682 241508
rect 2698 241564 2762 241568
rect 2698 241508 2702 241564
rect 2702 241508 2758 241564
rect 2758 241508 2762 241564
rect 2698 241504 2762 241508
rect 2778 241564 2842 241568
rect 2778 241508 2782 241564
rect 2782 241508 2838 241564
rect 2838 241508 2842 241564
rect 2778 241504 2842 241508
rect 2858 241564 2922 241568
rect 2858 241508 2862 241564
rect 2862 241508 2918 241564
rect 2918 241508 2922 241564
rect 2858 241504 2922 241508
rect 5952 241564 6016 241568
rect 5952 241508 5956 241564
rect 5956 241508 6012 241564
rect 6012 241508 6016 241564
rect 5952 241504 6016 241508
rect 6032 241564 6096 241568
rect 6032 241508 6036 241564
rect 6036 241508 6092 241564
rect 6092 241508 6096 241564
rect 6032 241504 6096 241508
rect 6112 241564 6176 241568
rect 6112 241508 6116 241564
rect 6116 241508 6172 241564
rect 6172 241508 6176 241564
rect 6112 241504 6176 241508
rect 6192 241564 6256 241568
rect 6192 241508 6196 241564
rect 6196 241508 6252 241564
rect 6252 241508 6256 241564
rect 6192 241504 6256 241508
rect 4285 241020 4349 241024
rect 4285 240964 4289 241020
rect 4289 240964 4345 241020
rect 4345 240964 4349 241020
rect 4285 240960 4349 240964
rect 4365 241020 4429 241024
rect 4365 240964 4369 241020
rect 4369 240964 4425 241020
rect 4425 240964 4429 241020
rect 4365 240960 4429 240964
rect 4445 241020 4509 241024
rect 4445 240964 4449 241020
rect 4449 240964 4505 241020
rect 4505 240964 4509 241020
rect 4445 240960 4509 240964
rect 4525 241020 4589 241024
rect 4525 240964 4529 241020
rect 4529 240964 4585 241020
rect 4585 240964 4589 241020
rect 4525 240960 4589 240964
rect 7618 241020 7682 241024
rect 7618 240964 7622 241020
rect 7622 240964 7678 241020
rect 7678 240964 7682 241020
rect 7618 240960 7682 240964
rect 7698 241020 7762 241024
rect 7698 240964 7702 241020
rect 7702 240964 7758 241020
rect 7758 240964 7762 241020
rect 7698 240960 7762 240964
rect 7778 241020 7842 241024
rect 7778 240964 7782 241020
rect 7782 240964 7838 241020
rect 7838 240964 7842 241020
rect 7778 240960 7842 240964
rect 7858 241020 7922 241024
rect 7858 240964 7862 241020
rect 7862 240964 7918 241020
rect 7918 240964 7922 241020
rect 7858 240960 7922 240964
rect 2618 240476 2682 240480
rect 2618 240420 2622 240476
rect 2622 240420 2678 240476
rect 2678 240420 2682 240476
rect 2618 240416 2682 240420
rect 2698 240476 2762 240480
rect 2698 240420 2702 240476
rect 2702 240420 2758 240476
rect 2758 240420 2762 240476
rect 2698 240416 2762 240420
rect 2778 240476 2842 240480
rect 2778 240420 2782 240476
rect 2782 240420 2838 240476
rect 2838 240420 2842 240476
rect 2778 240416 2842 240420
rect 2858 240476 2922 240480
rect 2858 240420 2862 240476
rect 2862 240420 2918 240476
rect 2918 240420 2922 240476
rect 2858 240416 2922 240420
rect 5952 240476 6016 240480
rect 5952 240420 5956 240476
rect 5956 240420 6012 240476
rect 6012 240420 6016 240476
rect 5952 240416 6016 240420
rect 6032 240476 6096 240480
rect 6032 240420 6036 240476
rect 6036 240420 6092 240476
rect 6092 240420 6096 240476
rect 6032 240416 6096 240420
rect 6112 240476 6176 240480
rect 6112 240420 6116 240476
rect 6116 240420 6172 240476
rect 6172 240420 6176 240476
rect 6112 240416 6176 240420
rect 6192 240476 6256 240480
rect 6192 240420 6196 240476
rect 6196 240420 6252 240476
rect 6252 240420 6256 240476
rect 6192 240416 6256 240420
rect 4285 239932 4349 239936
rect 4285 239876 4289 239932
rect 4289 239876 4345 239932
rect 4345 239876 4349 239932
rect 4285 239872 4349 239876
rect 4365 239932 4429 239936
rect 4365 239876 4369 239932
rect 4369 239876 4425 239932
rect 4425 239876 4429 239932
rect 4365 239872 4429 239876
rect 4445 239932 4509 239936
rect 4445 239876 4449 239932
rect 4449 239876 4505 239932
rect 4505 239876 4509 239932
rect 4445 239872 4509 239876
rect 4525 239932 4589 239936
rect 4525 239876 4529 239932
rect 4529 239876 4585 239932
rect 4585 239876 4589 239932
rect 4525 239872 4589 239876
rect 7618 239932 7682 239936
rect 7618 239876 7622 239932
rect 7622 239876 7678 239932
rect 7678 239876 7682 239932
rect 7618 239872 7682 239876
rect 7698 239932 7762 239936
rect 7698 239876 7702 239932
rect 7702 239876 7758 239932
rect 7758 239876 7762 239932
rect 7698 239872 7762 239876
rect 7778 239932 7842 239936
rect 7778 239876 7782 239932
rect 7782 239876 7838 239932
rect 7838 239876 7842 239932
rect 7778 239872 7842 239876
rect 7858 239932 7922 239936
rect 7858 239876 7862 239932
rect 7862 239876 7918 239932
rect 7918 239876 7922 239932
rect 7858 239872 7922 239876
rect 2618 239388 2682 239392
rect 2618 239332 2622 239388
rect 2622 239332 2678 239388
rect 2678 239332 2682 239388
rect 2618 239328 2682 239332
rect 2698 239388 2762 239392
rect 2698 239332 2702 239388
rect 2702 239332 2758 239388
rect 2758 239332 2762 239388
rect 2698 239328 2762 239332
rect 2778 239388 2842 239392
rect 2778 239332 2782 239388
rect 2782 239332 2838 239388
rect 2838 239332 2842 239388
rect 2778 239328 2842 239332
rect 2858 239388 2922 239392
rect 2858 239332 2862 239388
rect 2862 239332 2918 239388
rect 2918 239332 2922 239388
rect 2858 239328 2922 239332
rect 5952 239388 6016 239392
rect 5952 239332 5956 239388
rect 5956 239332 6012 239388
rect 6012 239332 6016 239388
rect 5952 239328 6016 239332
rect 6032 239388 6096 239392
rect 6032 239332 6036 239388
rect 6036 239332 6092 239388
rect 6092 239332 6096 239388
rect 6032 239328 6096 239332
rect 6112 239388 6176 239392
rect 6112 239332 6116 239388
rect 6116 239332 6172 239388
rect 6172 239332 6176 239388
rect 6112 239328 6176 239332
rect 6192 239388 6256 239392
rect 6192 239332 6196 239388
rect 6196 239332 6252 239388
rect 6252 239332 6256 239388
rect 6192 239328 6256 239332
rect 4285 238844 4349 238848
rect 4285 238788 4289 238844
rect 4289 238788 4345 238844
rect 4345 238788 4349 238844
rect 4285 238784 4349 238788
rect 4365 238844 4429 238848
rect 4365 238788 4369 238844
rect 4369 238788 4425 238844
rect 4425 238788 4429 238844
rect 4365 238784 4429 238788
rect 4445 238844 4509 238848
rect 4445 238788 4449 238844
rect 4449 238788 4505 238844
rect 4505 238788 4509 238844
rect 4445 238784 4509 238788
rect 4525 238844 4589 238848
rect 4525 238788 4529 238844
rect 4529 238788 4585 238844
rect 4585 238788 4589 238844
rect 4525 238784 4589 238788
rect 7618 238844 7682 238848
rect 7618 238788 7622 238844
rect 7622 238788 7678 238844
rect 7678 238788 7682 238844
rect 7618 238784 7682 238788
rect 7698 238844 7762 238848
rect 7698 238788 7702 238844
rect 7702 238788 7758 238844
rect 7758 238788 7762 238844
rect 7698 238784 7762 238788
rect 7778 238844 7842 238848
rect 7778 238788 7782 238844
rect 7782 238788 7838 238844
rect 7838 238788 7842 238844
rect 7778 238784 7842 238788
rect 7858 238844 7922 238848
rect 7858 238788 7862 238844
rect 7862 238788 7918 238844
rect 7918 238788 7922 238844
rect 7858 238784 7922 238788
rect 2618 238300 2682 238304
rect 2618 238244 2622 238300
rect 2622 238244 2678 238300
rect 2678 238244 2682 238300
rect 2618 238240 2682 238244
rect 2698 238300 2762 238304
rect 2698 238244 2702 238300
rect 2702 238244 2758 238300
rect 2758 238244 2762 238300
rect 2698 238240 2762 238244
rect 2778 238300 2842 238304
rect 2778 238244 2782 238300
rect 2782 238244 2838 238300
rect 2838 238244 2842 238300
rect 2778 238240 2842 238244
rect 2858 238300 2922 238304
rect 2858 238244 2862 238300
rect 2862 238244 2918 238300
rect 2918 238244 2922 238300
rect 2858 238240 2922 238244
rect 5952 238300 6016 238304
rect 5952 238244 5956 238300
rect 5956 238244 6012 238300
rect 6012 238244 6016 238300
rect 5952 238240 6016 238244
rect 6032 238300 6096 238304
rect 6032 238244 6036 238300
rect 6036 238244 6092 238300
rect 6092 238244 6096 238300
rect 6032 238240 6096 238244
rect 6112 238300 6176 238304
rect 6112 238244 6116 238300
rect 6116 238244 6172 238300
rect 6172 238244 6176 238300
rect 6112 238240 6176 238244
rect 6192 238300 6256 238304
rect 6192 238244 6196 238300
rect 6196 238244 6252 238300
rect 6252 238244 6256 238300
rect 6192 238240 6256 238244
rect 4285 237756 4349 237760
rect 4285 237700 4289 237756
rect 4289 237700 4345 237756
rect 4345 237700 4349 237756
rect 4285 237696 4349 237700
rect 4365 237756 4429 237760
rect 4365 237700 4369 237756
rect 4369 237700 4425 237756
rect 4425 237700 4429 237756
rect 4365 237696 4429 237700
rect 4445 237756 4509 237760
rect 4445 237700 4449 237756
rect 4449 237700 4505 237756
rect 4505 237700 4509 237756
rect 4445 237696 4509 237700
rect 4525 237756 4589 237760
rect 4525 237700 4529 237756
rect 4529 237700 4585 237756
rect 4585 237700 4589 237756
rect 4525 237696 4589 237700
rect 7618 237756 7682 237760
rect 7618 237700 7622 237756
rect 7622 237700 7678 237756
rect 7678 237700 7682 237756
rect 7618 237696 7682 237700
rect 7698 237756 7762 237760
rect 7698 237700 7702 237756
rect 7702 237700 7758 237756
rect 7758 237700 7762 237756
rect 7698 237696 7762 237700
rect 7778 237756 7842 237760
rect 7778 237700 7782 237756
rect 7782 237700 7838 237756
rect 7838 237700 7842 237756
rect 7778 237696 7842 237700
rect 7858 237756 7922 237760
rect 7858 237700 7862 237756
rect 7862 237700 7918 237756
rect 7918 237700 7922 237756
rect 7858 237696 7922 237700
rect 2618 237212 2682 237216
rect 2618 237156 2622 237212
rect 2622 237156 2678 237212
rect 2678 237156 2682 237212
rect 2618 237152 2682 237156
rect 2698 237212 2762 237216
rect 2698 237156 2702 237212
rect 2702 237156 2758 237212
rect 2758 237156 2762 237212
rect 2698 237152 2762 237156
rect 2778 237212 2842 237216
rect 2778 237156 2782 237212
rect 2782 237156 2838 237212
rect 2838 237156 2842 237212
rect 2778 237152 2842 237156
rect 2858 237212 2922 237216
rect 2858 237156 2862 237212
rect 2862 237156 2918 237212
rect 2918 237156 2922 237212
rect 2858 237152 2922 237156
rect 5952 237212 6016 237216
rect 5952 237156 5956 237212
rect 5956 237156 6012 237212
rect 6012 237156 6016 237212
rect 5952 237152 6016 237156
rect 6032 237212 6096 237216
rect 6032 237156 6036 237212
rect 6036 237156 6092 237212
rect 6092 237156 6096 237212
rect 6032 237152 6096 237156
rect 6112 237212 6176 237216
rect 6112 237156 6116 237212
rect 6116 237156 6172 237212
rect 6172 237156 6176 237212
rect 6112 237152 6176 237156
rect 6192 237212 6256 237216
rect 6192 237156 6196 237212
rect 6196 237156 6252 237212
rect 6252 237156 6256 237212
rect 6192 237152 6256 237156
rect 4285 236668 4349 236672
rect 4285 236612 4289 236668
rect 4289 236612 4345 236668
rect 4345 236612 4349 236668
rect 4285 236608 4349 236612
rect 4365 236668 4429 236672
rect 4365 236612 4369 236668
rect 4369 236612 4425 236668
rect 4425 236612 4429 236668
rect 4365 236608 4429 236612
rect 4445 236668 4509 236672
rect 4445 236612 4449 236668
rect 4449 236612 4505 236668
rect 4505 236612 4509 236668
rect 4445 236608 4509 236612
rect 4525 236668 4589 236672
rect 4525 236612 4529 236668
rect 4529 236612 4585 236668
rect 4585 236612 4589 236668
rect 4525 236608 4589 236612
rect 7618 236668 7682 236672
rect 7618 236612 7622 236668
rect 7622 236612 7678 236668
rect 7678 236612 7682 236668
rect 7618 236608 7682 236612
rect 7698 236668 7762 236672
rect 7698 236612 7702 236668
rect 7702 236612 7758 236668
rect 7758 236612 7762 236668
rect 7698 236608 7762 236612
rect 7778 236668 7842 236672
rect 7778 236612 7782 236668
rect 7782 236612 7838 236668
rect 7838 236612 7842 236668
rect 7778 236608 7842 236612
rect 7858 236668 7922 236672
rect 7858 236612 7862 236668
rect 7862 236612 7918 236668
rect 7918 236612 7922 236668
rect 7858 236608 7922 236612
rect 2618 236124 2682 236128
rect 2618 236068 2622 236124
rect 2622 236068 2678 236124
rect 2678 236068 2682 236124
rect 2618 236064 2682 236068
rect 2698 236124 2762 236128
rect 2698 236068 2702 236124
rect 2702 236068 2758 236124
rect 2758 236068 2762 236124
rect 2698 236064 2762 236068
rect 2778 236124 2842 236128
rect 2778 236068 2782 236124
rect 2782 236068 2838 236124
rect 2838 236068 2842 236124
rect 2778 236064 2842 236068
rect 2858 236124 2922 236128
rect 2858 236068 2862 236124
rect 2862 236068 2918 236124
rect 2918 236068 2922 236124
rect 2858 236064 2922 236068
rect 5952 236124 6016 236128
rect 5952 236068 5956 236124
rect 5956 236068 6012 236124
rect 6012 236068 6016 236124
rect 5952 236064 6016 236068
rect 6032 236124 6096 236128
rect 6032 236068 6036 236124
rect 6036 236068 6092 236124
rect 6092 236068 6096 236124
rect 6032 236064 6096 236068
rect 6112 236124 6176 236128
rect 6112 236068 6116 236124
rect 6116 236068 6172 236124
rect 6172 236068 6176 236124
rect 6112 236064 6176 236068
rect 6192 236124 6256 236128
rect 6192 236068 6196 236124
rect 6196 236068 6252 236124
rect 6252 236068 6256 236124
rect 6192 236064 6256 236068
rect 4285 235580 4349 235584
rect 4285 235524 4289 235580
rect 4289 235524 4345 235580
rect 4345 235524 4349 235580
rect 4285 235520 4349 235524
rect 4365 235580 4429 235584
rect 4365 235524 4369 235580
rect 4369 235524 4425 235580
rect 4425 235524 4429 235580
rect 4365 235520 4429 235524
rect 4445 235580 4509 235584
rect 4445 235524 4449 235580
rect 4449 235524 4505 235580
rect 4505 235524 4509 235580
rect 4445 235520 4509 235524
rect 4525 235580 4589 235584
rect 4525 235524 4529 235580
rect 4529 235524 4585 235580
rect 4585 235524 4589 235580
rect 4525 235520 4589 235524
rect 7618 235580 7682 235584
rect 7618 235524 7622 235580
rect 7622 235524 7678 235580
rect 7678 235524 7682 235580
rect 7618 235520 7682 235524
rect 7698 235580 7762 235584
rect 7698 235524 7702 235580
rect 7702 235524 7758 235580
rect 7758 235524 7762 235580
rect 7698 235520 7762 235524
rect 7778 235580 7842 235584
rect 7778 235524 7782 235580
rect 7782 235524 7838 235580
rect 7838 235524 7842 235580
rect 7778 235520 7842 235524
rect 7858 235580 7922 235584
rect 7858 235524 7862 235580
rect 7862 235524 7918 235580
rect 7918 235524 7922 235580
rect 7858 235520 7922 235524
rect 2618 235036 2682 235040
rect 2618 234980 2622 235036
rect 2622 234980 2678 235036
rect 2678 234980 2682 235036
rect 2618 234976 2682 234980
rect 2698 235036 2762 235040
rect 2698 234980 2702 235036
rect 2702 234980 2758 235036
rect 2758 234980 2762 235036
rect 2698 234976 2762 234980
rect 2778 235036 2842 235040
rect 2778 234980 2782 235036
rect 2782 234980 2838 235036
rect 2838 234980 2842 235036
rect 2778 234976 2842 234980
rect 2858 235036 2922 235040
rect 2858 234980 2862 235036
rect 2862 234980 2918 235036
rect 2918 234980 2922 235036
rect 2858 234976 2922 234980
rect 5952 235036 6016 235040
rect 5952 234980 5956 235036
rect 5956 234980 6012 235036
rect 6012 234980 6016 235036
rect 5952 234976 6016 234980
rect 6032 235036 6096 235040
rect 6032 234980 6036 235036
rect 6036 234980 6092 235036
rect 6092 234980 6096 235036
rect 6032 234976 6096 234980
rect 6112 235036 6176 235040
rect 6112 234980 6116 235036
rect 6116 234980 6172 235036
rect 6172 234980 6176 235036
rect 6112 234976 6176 234980
rect 6192 235036 6256 235040
rect 6192 234980 6196 235036
rect 6196 234980 6252 235036
rect 6252 234980 6256 235036
rect 6192 234976 6256 234980
rect 4285 234492 4349 234496
rect 4285 234436 4289 234492
rect 4289 234436 4345 234492
rect 4345 234436 4349 234492
rect 4285 234432 4349 234436
rect 4365 234492 4429 234496
rect 4365 234436 4369 234492
rect 4369 234436 4425 234492
rect 4425 234436 4429 234492
rect 4365 234432 4429 234436
rect 4445 234492 4509 234496
rect 4445 234436 4449 234492
rect 4449 234436 4505 234492
rect 4505 234436 4509 234492
rect 4445 234432 4509 234436
rect 4525 234492 4589 234496
rect 4525 234436 4529 234492
rect 4529 234436 4585 234492
rect 4585 234436 4589 234492
rect 4525 234432 4589 234436
rect 7618 234492 7682 234496
rect 7618 234436 7622 234492
rect 7622 234436 7678 234492
rect 7678 234436 7682 234492
rect 7618 234432 7682 234436
rect 7698 234492 7762 234496
rect 7698 234436 7702 234492
rect 7702 234436 7758 234492
rect 7758 234436 7762 234492
rect 7698 234432 7762 234436
rect 7778 234492 7842 234496
rect 7778 234436 7782 234492
rect 7782 234436 7838 234492
rect 7838 234436 7842 234492
rect 7778 234432 7842 234436
rect 7858 234492 7922 234496
rect 7858 234436 7862 234492
rect 7862 234436 7918 234492
rect 7918 234436 7922 234492
rect 7858 234432 7922 234436
rect 2618 233948 2682 233952
rect 2618 233892 2622 233948
rect 2622 233892 2678 233948
rect 2678 233892 2682 233948
rect 2618 233888 2682 233892
rect 2698 233948 2762 233952
rect 2698 233892 2702 233948
rect 2702 233892 2758 233948
rect 2758 233892 2762 233948
rect 2698 233888 2762 233892
rect 2778 233948 2842 233952
rect 2778 233892 2782 233948
rect 2782 233892 2838 233948
rect 2838 233892 2842 233948
rect 2778 233888 2842 233892
rect 2858 233948 2922 233952
rect 2858 233892 2862 233948
rect 2862 233892 2918 233948
rect 2918 233892 2922 233948
rect 2858 233888 2922 233892
rect 5952 233948 6016 233952
rect 5952 233892 5956 233948
rect 5956 233892 6012 233948
rect 6012 233892 6016 233948
rect 5952 233888 6016 233892
rect 6032 233948 6096 233952
rect 6032 233892 6036 233948
rect 6036 233892 6092 233948
rect 6092 233892 6096 233948
rect 6032 233888 6096 233892
rect 6112 233948 6176 233952
rect 6112 233892 6116 233948
rect 6116 233892 6172 233948
rect 6172 233892 6176 233948
rect 6112 233888 6176 233892
rect 6192 233948 6256 233952
rect 6192 233892 6196 233948
rect 6196 233892 6252 233948
rect 6252 233892 6256 233948
rect 6192 233888 6256 233892
rect 4285 233404 4349 233408
rect 4285 233348 4289 233404
rect 4289 233348 4345 233404
rect 4345 233348 4349 233404
rect 4285 233344 4349 233348
rect 4365 233404 4429 233408
rect 4365 233348 4369 233404
rect 4369 233348 4425 233404
rect 4425 233348 4429 233404
rect 4365 233344 4429 233348
rect 4445 233404 4509 233408
rect 4445 233348 4449 233404
rect 4449 233348 4505 233404
rect 4505 233348 4509 233404
rect 4445 233344 4509 233348
rect 4525 233404 4589 233408
rect 4525 233348 4529 233404
rect 4529 233348 4585 233404
rect 4585 233348 4589 233404
rect 4525 233344 4589 233348
rect 7618 233404 7682 233408
rect 7618 233348 7622 233404
rect 7622 233348 7678 233404
rect 7678 233348 7682 233404
rect 7618 233344 7682 233348
rect 7698 233404 7762 233408
rect 7698 233348 7702 233404
rect 7702 233348 7758 233404
rect 7758 233348 7762 233404
rect 7698 233344 7762 233348
rect 7778 233404 7842 233408
rect 7778 233348 7782 233404
rect 7782 233348 7838 233404
rect 7838 233348 7842 233404
rect 7778 233344 7842 233348
rect 7858 233404 7922 233408
rect 7858 233348 7862 233404
rect 7862 233348 7918 233404
rect 7918 233348 7922 233404
rect 7858 233344 7922 233348
rect 2618 232860 2682 232864
rect 2618 232804 2622 232860
rect 2622 232804 2678 232860
rect 2678 232804 2682 232860
rect 2618 232800 2682 232804
rect 2698 232860 2762 232864
rect 2698 232804 2702 232860
rect 2702 232804 2758 232860
rect 2758 232804 2762 232860
rect 2698 232800 2762 232804
rect 2778 232860 2842 232864
rect 2778 232804 2782 232860
rect 2782 232804 2838 232860
rect 2838 232804 2842 232860
rect 2778 232800 2842 232804
rect 2858 232860 2922 232864
rect 2858 232804 2862 232860
rect 2862 232804 2918 232860
rect 2918 232804 2922 232860
rect 2858 232800 2922 232804
rect 5952 232860 6016 232864
rect 5952 232804 5956 232860
rect 5956 232804 6012 232860
rect 6012 232804 6016 232860
rect 5952 232800 6016 232804
rect 6032 232860 6096 232864
rect 6032 232804 6036 232860
rect 6036 232804 6092 232860
rect 6092 232804 6096 232860
rect 6032 232800 6096 232804
rect 6112 232860 6176 232864
rect 6112 232804 6116 232860
rect 6116 232804 6172 232860
rect 6172 232804 6176 232860
rect 6112 232800 6176 232804
rect 6192 232860 6256 232864
rect 6192 232804 6196 232860
rect 6196 232804 6252 232860
rect 6252 232804 6256 232860
rect 6192 232800 6256 232804
rect 4285 232316 4349 232320
rect 4285 232260 4289 232316
rect 4289 232260 4345 232316
rect 4345 232260 4349 232316
rect 4285 232256 4349 232260
rect 4365 232316 4429 232320
rect 4365 232260 4369 232316
rect 4369 232260 4425 232316
rect 4425 232260 4429 232316
rect 4365 232256 4429 232260
rect 4445 232316 4509 232320
rect 4445 232260 4449 232316
rect 4449 232260 4505 232316
rect 4505 232260 4509 232316
rect 4445 232256 4509 232260
rect 4525 232316 4589 232320
rect 4525 232260 4529 232316
rect 4529 232260 4585 232316
rect 4585 232260 4589 232316
rect 4525 232256 4589 232260
rect 7618 232316 7682 232320
rect 7618 232260 7622 232316
rect 7622 232260 7678 232316
rect 7678 232260 7682 232316
rect 7618 232256 7682 232260
rect 7698 232316 7762 232320
rect 7698 232260 7702 232316
rect 7702 232260 7758 232316
rect 7758 232260 7762 232316
rect 7698 232256 7762 232260
rect 7778 232316 7842 232320
rect 7778 232260 7782 232316
rect 7782 232260 7838 232316
rect 7838 232260 7842 232316
rect 7778 232256 7842 232260
rect 7858 232316 7922 232320
rect 7858 232260 7862 232316
rect 7862 232260 7918 232316
rect 7918 232260 7922 232316
rect 7858 232256 7922 232260
rect 2618 231772 2682 231776
rect 2618 231716 2622 231772
rect 2622 231716 2678 231772
rect 2678 231716 2682 231772
rect 2618 231712 2682 231716
rect 2698 231772 2762 231776
rect 2698 231716 2702 231772
rect 2702 231716 2758 231772
rect 2758 231716 2762 231772
rect 2698 231712 2762 231716
rect 2778 231772 2842 231776
rect 2778 231716 2782 231772
rect 2782 231716 2838 231772
rect 2838 231716 2842 231772
rect 2778 231712 2842 231716
rect 2858 231772 2922 231776
rect 2858 231716 2862 231772
rect 2862 231716 2918 231772
rect 2918 231716 2922 231772
rect 2858 231712 2922 231716
rect 5952 231772 6016 231776
rect 5952 231716 5956 231772
rect 5956 231716 6012 231772
rect 6012 231716 6016 231772
rect 5952 231712 6016 231716
rect 6032 231772 6096 231776
rect 6032 231716 6036 231772
rect 6036 231716 6092 231772
rect 6092 231716 6096 231772
rect 6032 231712 6096 231716
rect 6112 231772 6176 231776
rect 6112 231716 6116 231772
rect 6116 231716 6172 231772
rect 6172 231716 6176 231772
rect 6112 231712 6176 231716
rect 6192 231772 6256 231776
rect 6192 231716 6196 231772
rect 6196 231716 6252 231772
rect 6252 231716 6256 231772
rect 6192 231712 6256 231716
rect 4285 231228 4349 231232
rect 4285 231172 4289 231228
rect 4289 231172 4345 231228
rect 4345 231172 4349 231228
rect 4285 231168 4349 231172
rect 4365 231228 4429 231232
rect 4365 231172 4369 231228
rect 4369 231172 4425 231228
rect 4425 231172 4429 231228
rect 4365 231168 4429 231172
rect 4445 231228 4509 231232
rect 4445 231172 4449 231228
rect 4449 231172 4505 231228
rect 4505 231172 4509 231228
rect 4445 231168 4509 231172
rect 4525 231228 4589 231232
rect 4525 231172 4529 231228
rect 4529 231172 4585 231228
rect 4585 231172 4589 231228
rect 4525 231168 4589 231172
rect 7618 231228 7682 231232
rect 7618 231172 7622 231228
rect 7622 231172 7678 231228
rect 7678 231172 7682 231228
rect 7618 231168 7682 231172
rect 7698 231228 7762 231232
rect 7698 231172 7702 231228
rect 7702 231172 7758 231228
rect 7758 231172 7762 231228
rect 7698 231168 7762 231172
rect 7778 231228 7842 231232
rect 7778 231172 7782 231228
rect 7782 231172 7838 231228
rect 7838 231172 7842 231228
rect 7778 231168 7842 231172
rect 7858 231228 7922 231232
rect 7858 231172 7862 231228
rect 7862 231172 7918 231228
rect 7918 231172 7922 231228
rect 7858 231168 7922 231172
rect 2618 230684 2682 230688
rect 2618 230628 2622 230684
rect 2622 230628 2678 230684
rect 2678 230628 2682 230684
rect 2618 230624 2682 230628
rect 2698 230684 2762 230688
rect 2698 230628 2702 230684
rect 2702 230628 2758 230684
rect 2758 230628 2762 230684
rect 2698 230624 2762 230628
rect 2778 230684 2842 230688
rect 2778 230628 2782 230684
rect 2782 230628 2838 230684
rect 2838 230628 2842 230684
rect 2778 230624 2842 230628
rect 2858 230684 2922 230688
rect 2858 230628 2862 230684
rect 2862 230628 2918 230684
rect 2918 230628 2922 230684
rect 2858 230624 2922 230628
rect 5952 230684 6016 230688
rect 5952 230628 5956 230684
rect 5956 230628 6012 230684
rect 6012 230628 6016 230684
rect 5952 230624 6016 230628
rect 6032 230684 6096 230688
rect 6032 230628 6036 230684
rect 6036 230628 6092 230684
rect 6092 230628 6096 230684
rect 6032 230624 6096 230628
rect 6112 230684 6176 230688
rect 6112 230628 6116 230684
rect 6116 230628 6172 230684
rect 6172 230628 6176 230684
rect 6112 230624 6176 230628
rect 6192 230684 6256 230688
rect 6192 230628 6196 230684
rect 6196 230628 6252 230684
rect 6252 230628 6256 230684
rect 6192 230624 6256 230628
rect 4285 230140 4349 230144
rect 4285 230084 4289 230140
rect 4289 230084 4345 230140
rect 4345 230084 4349 230140
rect 4285 230080 4349 230084
rect 4365 230140 4429 230144
rect 4365 230084 4369 230140
rect 4369 230084 4425 230140
rect 4425 230084 4429 230140
rect 4365 230080 4429 230084
rect 4445 230140 4509 230144
rect 4445 230084 4449 230140
rect 4449 230084 4505 230140
rect 4505 230084 4509 230140
rect 4445 230080 4509 230084
rect 4525 230140 4589 230144
rect 4525 230084 4529 230140
rect 4529 230084 4585 230140
rect 4585 230084 4589 230140
rect 4525 230080 4589 230084
rect 7618 230140 7682 230144
rect 7618 230084 7622 230140
rect 7622 230084 7678 230140
rect 7678 230084 7682 230140
rect 7618 230080 7682 230084
rect 7698 230140 7762 230144
rect 7698 230084 7702 230140
rect 7702 230084 7758 230140
rect 7758 230084 7762 230140
rect 7698 230080 7762 230084
rect 7778 230140 7842 230144
rect 7778 230084 7782 230140
rect 7782 230084 7838 230140
rect 7838 230084 7842 230140
rect 7778 230080 7842 230084
rect 7858 230140 7922 230144
rect 7858 230084 7862 230140
rect 7862 230084 7918 230140
rect 7918 230084 7922 230140
rect 7858 230080 7922 230084
rect 2618 229596 2682 229600
rect 2618 229540 2622 229596
rect 2622 229540 2678 229596
rect 2678 229540 2682 229596
rect 2618 229536 2682 229540
rect 2698 229596 2762 229600
rect 2698 229540 2702 229596
rect 2702 229540 2758 229596
rect 2758 229540 2762 229596
rect 2698 229536 2762 229540
rect 2778 229596 2842 229600
rect 2778 229540 2782 229596
rect 2782 229540 2838 229596
rect 2838 229540 2842 229596
rect 2778 229536 2842 229540
rect 2858 229596 2922 229600
rect 2858 229540 2862 229596
rect 2862 229540 2918 229596
rect 2918 229540 2922 229596
rect 2858 229536 2922 229540
rect 5952 229596 6016 229600
rect 5952 229540 5956 229596
rect 5956 229540 6012 229596
rect 6012 229540 6016 229596
rect 5952 229536 6016 229540
rect 6032 229596 6096 229600
rect 6032 229540 6036 229596
rect 6036 229540 6092 229596
rect 6092 229540 6096 229596
rect 6032 229536 6096 229540
rect 6112 229596 6176 229600
rect 6112 229540 6116 229596
rect 6116 229540 6172 229596
rect 6172 229540 6176 229596
rect 6112 229536 6176 229540
rect 6192 229596 6256 229600
rect 6192 229540 6196 229596
rect 6196 229540 6252 229596
rect 6252 229540 6256 229596
rect 6192 229536 6256 229540
rect 4285 229052 4349 229056
rect 4285 228996 4289 229052
rect 4289 228996 4345 229052
rect 4345 228996 4349 229052
rect 4285 228992 4349 228996
rect 4365 229052 4429 229056
rect 4365 228996 4369 229052
rect 4369 228996 4425 229052
rect 4425 228996 4429 229052
rect 4365 228992 4429 228996
rect 4445 229052 4509 229056
rect 4445 228996 4449 229052
rect 4449 228996 4505 229052
rect 4505 228996 4509 229052
rect 4445 228992 4509 228996
rect 4525 229052 4589 229056
rect 4525 228996 4529 229052
rect 4529 228996 4585 229052
rect 4585 228996 4589 229052
rect 4525 228992 4589 228996
rect 7618 229052 7682 229056
rect 7618 228996 7622 229052
rect 7622 228996 7678 229052
rect 7678 228996 7682 229052
rect 7618 228992 7682 228996
rect 7698 229052 7762 229056
rect 7698 228996 7702 229052
rect 7702 228996 7758 229052
rect 7758 228996 7762 229052
rect 7698 228992 7762 228996
rect 7778 229052 7842 229056
rect 7778 228996 7782 229052
rect 7782 228996 7838 229052
rect 7838 228996 7842 229052
rect 7778 228992 7842 228996
rect 7858 229052 7922 229056
rect 7858 228996 7862 229052
rect 7862 228996 7918 229052
rect 7918 228996 7922 229052
rect 7858 228992 7922 228996
rect 2618 228508 2682 228512
rect 2618 228452 2622 228508
rect 2622 228452 2678 228508
rect 2678 228452 2682 228508
rect 2618 228448 2682 228452
rect 2698 228508 2762 228512
rect 2698 228452 2702 228508
rect 2702 228452 2758 228508
rect 2758 228452 2762 228508
rect 2698 228448 2762 228452
rect 2778 228508 2842 228512
rect 2778 228452 2782 228508
rect 2782 228452 2838 228508
rect 2838 228452 2842 228508
rect 2778 228448 2842 228452
rect 2858 228508 2922 228512
rect 2858 228452 2862 228508
rect 2862 228452 2918 228508
rect 2918 228452 2922 228508
rect 2858 228448 2922 228452
rect 5952 228508 6016 228512
rect 5952 228452 5956 228508
rect 5956 228452 6012 228508
rect 6012 228452 6016 228508
rect 5952 228448 6016 228452
rect 6032 228508 6096 228512
rect 6032 228452 6036 228508
rect 6036 228452 6092 228508
rect 6092 228452 6096 228508
rect 6032 228448 6096 228452
rect 6112 228508 6176 228512
rect 6112 228452 6116 228508
rect 6116 228452 6172 228508
rect 6172 228452 6176 228508
rect 6112 228448 6176 228452
rect 6192 228508 6256 228512
rect 6192 228452 6196 228508
rect 6196 228452 6252 228508
rect 6252 228452 6256 228508
rect 6192 228448 6256 228452
rect 4285 227964 4349 227968
rect 4285 227908 4289 227964
rect 4289 227908 4345 227964
rect 4345 227908 4349 227964
rect 4285 227904 4349 227908
rect 4365 227964 4429 227968
rect 4365 227908 4369 227964
rect 4369 227908 4425 227964
rect 4425 227908 4429 227964
rect 4365 227904 4429 227908
rect 4445 227964 4509 227968
rect 4445 227908 4449 227964
rect 4449 227908 4505 227964
rect 4505 227908 4509 227964
rect 4445 227904 4509 227908
rect 4525 227964 4589 227968
rect 4525 227908 4529 227964
rect 4529 227908 4585 227964
rect 4585 227908 4589 227964
rect 4525 227904 4589 227908
rect 7618 227964 7682 227968
rect 7618 227908 7622 227964
rect 7622 227908 7678 227964
rect 7678 227908 7682 227964
rect 7618 227904 7682 227908
rect 7698 227964 7762 227968
rect 7698 227908 7702 227964
rect 7702 227908 7758 227964
rect 7758 227908 7762 227964
rect 7698 227904 7762 227908
rect 7778 227964 7842 227968
rect 7778 227908 7782 227964
rect 7782 227908 7838 227964
rect 7838 227908 7842 227964
rect 7778 227904 7842 227908
rect 7858 227964 7922 227968
rect 7858 227908 7862 227964
rect 7862 227908 7918 227964
rect 7918 227908 7922 227964
rect 7858 227904 7922 227908
rect 2618 227420 2682 227424
rect 2618 227364 2622 227420
rect 2622 227364 2678 227420
rect 2678 227364 2682 227420
rect 2618 227360 2682 227364
rect 2698 227420 2762 227424
rect 2698 227364 2702 227420
rect 2702 227364 2758 227420
rect 2758 227364 2762 227420
rect 2698 227360 2762 227364
rect 2778 227420 2842 227424
rect 2778 227364 2782 227420
rect 2782 227364 2838 227420
rect 2838 227364 2842 227420
rect 2778 227360 2842 227364
rect 2858 227420 2922 227424
rect 2858 227364 2862 227420
rect 2862 227364 2918 227420
rect 2918 227364 2922 227420
rect 2858 227360 2922 227364
rect 5952 227420 6016 227424
rect 5952 227364 5956 227420
rect 5956 227364 6012 227420
rect 6012 227364 6016 227420
rect 5952 227360 6016 227364
rect 6032 227420 6096 227424
rect 6032 227364 6036 227420
rect 6036 227364 6092 227420
rect 6092 227364 6096 227420
rect 6032 227360 6096 227364
rect 6112 227420 6176 227424
rect 6112 227364 6116 227420
rect 6116 227364 6172 227420
rect 6172 227364 6176 227420
rect 6112 227360 6176 227364
rect 6192 227420 6256 227424
rect 6192 227364 6196 227420
rect 6196 227364 6252 227420
rect 6252 227364 6256 227420
rect 6192 227360 6256 227364
rect 4285 226876 4349 226880
rect 4285 226820 4289 226876
rect 4289 226820 4345 226876
rect 4345 226820 4349 226876
rect 4285 226816 4349 226820
rect 4365 226876 4429 226880
rect 4365 226820 4369 226876
rect 4369 226820 4425 226876
rect 4425 226820 4429 226876
rect 4365 226816 4429 226820
rect 4445 226876 4509 226880
rect 4445 226820 4449 226876
rect 4449 226820 4505 226876
rect 4505 226820 4509 226876
rect 4445 226816 4509 226820
rect 4525 226876 4589 226880
rect 4525 226820 4529 226876
rect 4529 226820 4585 226876
rect 4585 226820 4589 226876
rect 4525 226816 4589 226820
rect 7618 226876 7682 226880
rect 7618 226820 7622 226876
rect 7622 226820 7678 226876
rect 7678 226820 7682 226876
rect 7618 226816 7682 226820
rect 7698 226876 7762 226880
rect 7698 226820 7702 226876
rect 7702 226820 7758 226876
rect 7758 226820 7762 226876
rect 7698 226816 7762 226820
rect 7778 226876 7842 226880
rect 7778 226820 7782 226876
rect 7782 226820 7838 226876
rect 7838 226820 7842 226876
rect 7778 226816 7842 226820
rect 7858 226876 7922 226880
rect 7858 226820 7862 226876
rect 7862 226820 7918 226876
rect 7918 226820 7922 226876
rect 7858 226816 7922 226820
rect 2618 226332 2682 226336
rect 2618 226276 2622 226332
rect 2622 226276 2678 226332
rect 2678 226276 2682 226332
rect 2618 226272 2682 226276
rect 2698 226332 2762 226336
rect 2698 226276 2702 226332
rect 2702 226276 2758 226332
rect 2758 226276 2762 226332
rect 2698 226272 2762 226276
rect 2778 226332 2842 226336
rect 2778 226276 2782 226332
rect 2782 226276 2838 226332
rect 2838 226276 2842 226332
rect 2778 226272 2842 226276
rect 2858 226332 2922 226336
rect 2858 226276 2862 226332
rect 2862 226276 2918 226332
rect 2918 226276 2922 226332
rect 2858 226272 2922 226276
rect 5952 226332 6016 226336
rect 5952 226276 5956 226332
rect 5956 226276 6012 226332
rect 6012 226276 6016 226332
rect 5952 226272 6016 226276
rect 6032 226332 6096 226336
rect 6032 226276 6036 226332
rect 6036 226276 6092 226332
rect 6092 226276 6096 226332
rect 6032 226272 6096 226276
rect 6112 226332 6176 226336
rect 6112 226276 6116 226332
rect 6116 226276 6172 226332
rect 6172 226276 6176 226332
rect 6112 226272 6176 226276
rect 6192 226332 6256 226336
rect 6192 226276 6196 226332
rect 6196 226276 6252 226332
rect 6252 226276 6256 226332
rect 6192 226272 6256 226276
rect 4285 225788 4349 225792
rect 4285 225732 4289 225788
rect 4289 225732 4345 225788
rect 4345 225732 4349 225788
rect 4285 225728 4349 225732
rect 4365 225788 4429 225792
rect 4365 225732 4369 225788
rect 4369 225732 4425 225788
rect 4425 225732 4429 225788
rect 4365 225728 4429 225732
rect 4445 225788 4509 225792
rect 4445 225732 4449 225788
rect 4449 225732 4505 225788
rect 4505 225732 4509 225788
rect 4445 225728 4509 225732
rect 4525 225788 4589 225792
rect 4525 225732 4529 225788
rect 4529 225732 4585 225788
rect 4585 225732 4589 225788
rect 4525 225728 4589 225732
rect 7618 225788 7682 225792
rect 7618 225732 7622 225788
rect 7622 225732 7678 225788
rect 7678 225732 7682 225788
rect 7618 225728 7682 225732
rect 7698 225788 7762 225792
rect 7698 225732 7702 225788
rect 7702 225732 7758 225788
rect 7758 225732 7762 225788
rect 7698 225728 7762 225732
rect 7778 225788 7842 225792
rect 7778 225732 7782 225788
rect 7782 225732 7838 225788
rect 7838 225732 7842 225788
rect 7778 225728 7842 225732
rect 7858 225788 7922 225792
rect 7858 225732 7862 225788
rect 7862 225732 7918 225788
rect 7918 225732 7922 225788
rect 7858 225728 7922 225732
rect 2618 225244 2682 225248
rect 2618 225188 2622 225244
rect 2622 225188 2678 225244
rect 2678 225188 2682 225244
rect 2618 225184 2682 225188
rect 2698 225244 2762 225248
rect 2698 225188 2702 225244
rect 2702 225188 2758 225244
rect 2758 225188 2762 225244
rect 2698 225184 2762 225188
rect 2778 225244 2842 225248
rect 2778 225188 2782 225244
rect 2782 225188 2838 225244
rect 2838 225188 2842 225244
rect 2778 225184 2842 225188
rect 2858 225244 2922 225248
rect 2858 225188 2862 225244
rect 2862 225188 2918 225244
rect 2918 225188 2922 225244
rect 2858 225184 2922 225188
rect 5952 225244 6016 225248
rect 5952 225188 5956 225244
rect 5956 225188 6012 225244
rect 6012 225188 6016 225244
rect 5952 225184 6016 225188
rect 6032 225244 6096 225248
rect 6032 225188 6036 225244
rect 6036 225188 6092 225244
rect 6092 225188 6096 225244
rect 6032 225184 6096 225188
rect 6112 225244 6176 225248
rect 6112 225188 6116 225244
rect 6116 225188 6172 225244
rect 6172 225188 6176 225244
rect 6112 225184 6176 225188
rect 6192 225244 6256 225248
rect 6192 225188 6196 225244
rect 6196 225188 6252 225244
rect 6252 225188 6256 225244
rect 6192 225184 6256 225188
rect 4285 224700 4349 224704
rect 4285 224644 4289 224700
rect 4289 224644 4345 224700
rect 4345 224644 4349 224700
rect 4285 224640 4349 224644
rect 4365 224700 4429 224704
rect 4365 224644 4369 224700
rect 4369 224644 4425 224700
rect 4425 224644 4429 224700
rect 4365 224640 4429 224644
rect 4445 224700 4509 224704
rect 4445 224644 4449 224700
rect 4449 224644 4505 224700
rect 4505 224644 4509 224700
rect 4445 224640 4509 224644
rect 4525 224700 4589 224704
rect 4525 224644 4529 224700
rect 4529 224644 4585 224700
rect 4585 224644 4589 224700
rect 4525 224640 4589 224644
rect 7618 224700 7682 224704
rect 7618 224644 7622 224700
rect 7622 224644 7678 224700
rect 7678 224644 7682 224700
rect 7618 224640 7682 224644
rect 7698 224700 7762 224704
rect 7698 224644 7702 224700
rect 7702 224644 7758 224700
rect 7758 224644 7762 224700
rect 7698 224640 7762 224644
rect 7778 224700 7842 224704
rect 7778 224644 7782 224700
rect 7782 224644 7838 224700
rect 7838 224644 7842 224700
rect 7778 224640 7842 224644
rect 7858 224700 7922 224704
rect 7858 224644 7862 224700
rect 7862 224644 7918 224700
rect 7918 224644 7922 224700
rect 7858 224640 7922 224644
rect 2618 224156 2682 224160
rect 2618 224100 2622 224156
rect 2622 224100 2678 224156
rect 2678 224100 2682 224156
rect 2618 224096 2682 224100
rect 2698 224156 2762 224160
rect 2698 224100 2702 224156
rect 2702 224100 2758 224156
rect 2758 224100 2762 224156
rect 2698 224096 2762 224100
rect 2778 224156 2842 224160
rect 2778 224100 2782 224156
rect 2782 224100 2838 224156
rect 2838 224100 2842 224156
rect 2778 224096 2842 224100
rect 2858 224156 2922 224160
rect 2858 224100 2862 224156
rect 2862 224100 2918 224156
rect 2918 224100 2922 224156
rect 2858 224096 2922 224100
rect 5952 224156 6016 224160
rect 5952 224100 5956 224156
rect 5956 224100 6012 224156
rect 6012 224100 6016 224156
rect 5952 224096 6016 224100
rect 6032 224156 6096 224160
rect 6032 224100 6036 224156
rect 6036 224100 6092 224156
rect 6092 224100 6096 224156
rect 6032 224096 6096 224100
rect 6112 224156 6176 224160
rect 6112 224100 6116 224156
rect 6116 224100 6172 224156
rect 6172 224100 6176 224156
rect 6112 224096 6176 224100
rect 6192 224156 6256 224160
rect 6192 224100 6196 224156
rect 6196 224100 6252 224156
rect 6252 224100 6256 224156
rect 6192 224096 6256 224100
rect 4285 223612 4349 223616
rect 4285 223556 4289 223612
rect 4289 223556 4345 223612
rect 4345 223556 4349 223612
rect 4285 223552 4349 223556
rect 4365 223612 4429 223616
rect 4365 223556 4369 223612
rect 4369 223556 4425 223612
rect 4425 223556 4429 223612
rect 4365 223552 4429 223556
rect 4445 223612 4509 223616
rect 4445 223556 4449 223612
rect 4449 223556 4505 223612
rect 4505 223556 4509 223612
rect 4445 223552 4509 223556
rect 4525 223612 4589 223616
rect 4525 223556 4529 223612
rect 4529 223556 4585 223612
rect 4585 223556 4589 223612
rect 4525 223552 4589 223556
rect 7618 223612 7682 223616
rect 7618 223556 7622 223612
rect 7622 223556 7678 223612
rect 7678 223556 7682 223612
rect 7618 223552 7682 223556
rect 7698 223612 7762 223616
rect 7698 223556 7702 223612
rect 7702 223556 7758 223612
rect 7758 223556 7762 223612
rect 7698 223552 7762 223556
rect 7778 223612 7842 223616
rect 7778 223556 7782 223612
rect 7782 223556 7838 223612
rect 7838 223556 7842 223612
rect 7778 223552 7842 223556
rect 7858 223612 7922 223616
rect 7858 223556 7862 223612
rect 7862 223556 7918 223612
rect 7918 223556 7922 223612
rect 7858 223552 7922 223556
rect 2618 223068 2682 223072
rect 2618 223012 2622 223068
rect 2622 223012 2678 223068
rect 2678 223012 2682 223068
rect 2618 223008 2682 223012
rect 2698 223068 2762 223072
rect 2698 223012 2702 223068
rect 2702 223012 2758 223068
rect 2758 223012 2762 223068
rect 2698 223008 2762 223012
rect 2778 223068 2842 223072
rect 2778 223012 2782 223068
rect 2782 223012 2838 223068
rect 2838 223012 2842 223068
rect 2778 223008 2842 223012
rect 2858 223068 2922 223072
rect 2858 223012 2862 223068
rect 2862 223012 2918 223068
rect 2918 223012 2922 223068
rect 2858 223008 2922 223012
rect 5952 223068 6016 223072
rect 5952 223012 5956 223068
rect 5956 223012 6012 223068
rect 6012 223012 6016 223068
rect 5952 223008 6016 223012
rect 6032 223068 6096 223072
rect 6032 223012 6036 223068
rect 6036 223012 6092 223068
rect 6092 223012 6096 223068
rect 6032 223008 6096 223012
rect 6112 223068 6176 223072
rect 6112 223012 6116 223068
rect 6116 223012 6172 223068
rect 6172 223012 6176 223068
rect 6112 223008 6176 223012
rect 6192 223068 6256 223072
rect 6192 223012 6196 223068
rect 6196 223012 6252 223068
rect 6252 223012 6256 223068
rect 6192 223008 6256 223012
rect 4285 222524 4349 222528
rect 4285 222468 4289 222524
rect 4289 222468 4345 222524
rect 4345 222468 4349 222524
rect 4285 222464 4349 222468
rect 4365 222524 4429 222528
rect 4365 222468 4369 222524
rect 4369 222468 4425 222524
rect 4425 222468 4429 222524
rect 4365 222464 4429 222468
rect 4445 222524 4509 222528
rect 4445 222468 4449 222524
rect 4449 222468 4505 222524
rect 4505 222468 4509 222524
rect 4445 222464 4509 222468
rect 4525 222524 4589 222528
rect 4525 222468 4529 222524
rect 4529 222468 4585 222524
rect 4585 222468 4589 222524
rect 4525 222464 4589 222468
rect 7618 222524 7682 222528
rect 7618 222468 7622 222524
rect 7622 222468 7678 222524
rect 7678 222468 7682 222524
rect 7618 222464 7682 222468
rect 7698 222524 7762 222528
rect 7698 222468 7702 222524
rect 7702 222468 7758 222524
rect 7758 222468 7762 222524
rect 7698 222464 7762 222468
rect 7778 222524 7842 222528
rect 7778 222468 7782 222524
rect 7782 222468 7838 222524
rect 7838 222468 7842 222524
rect 7778 222464 7842 222468
rect 7858 222524 7922 222528
rect 7858 222468 7862 222524
rect 7862 222468 7918 222524
rect 7918 222468 7922 222524
rect 7858 222464 7922 222468
rect 2618 221980 2682 221984
rect 2618 221924 2622 221980
rect 2622 221924 2678 221980
rect 2678 221924 2682 221980
rect 2618 221920 2682 221924
rect 2698 221980 2762 221984
rect 2698 221924 2702 221980
rect 2702 221924 2758 221980
rect 2758 221924 2762 221980
rect 2698 221920 2762 221924
rect 2778 221980 2842 221984
rect 2778 221924 2782 221980
rect 2782 221924 2838 221980
rect 2838 221924 2842 221980
rect 2778 221920 2842 221924
rect 2858 221980 2922 221984
rect 2858 221924 2862 221980
rect 2862 221924 2918 221980
rect 2918 221924 2922 221980
rect 2858 221920 2922 221924
rect 5952 221980 6016 221984
rect 5952 221924 5956 221980
rect 5956 221924 6012 221980
rect 6012 221924 6016 221980
rect 5952 221920 6016 221924
rect 6032 221980 6096 221984
rect 6032 221924 6036 221980
rect 6036 221924 6092 221980
rect 6092 221924 6096 221980
rect 6032 221920 6096 221924
rect 6112 221980 6176 221984
rect 6112 221924 6116 221980
rect 6116 221924 6172 221980
rect 6172 221924 6176 221980
rect 6112 221920 6176 221924
rect 6192 221980 6256 221984
rect 6192 221924 6196 221980
rect 6196 221924 6252 221980
rect 6252 221924 6256 221980
rect 6192 221920 6256 221924
rect 4285 221436 4349 221440
rect 4285 221380 4289 221436
rect 4289 221380 4345 221436
rect 4345 221380 4349 221436
rect 4285 221376 4349 221380
rect 4365 221436 4429 221440
rect 4365 221380 4369 221436
rect 4369 221380 4425 221436
rect 4425 221380 4429 221436
rect 4365 221376 4429 221380
rect 4445 221436 4509 221440
rect 4445 221380 4449 221436
rect 4449 221380 4505 221436
rect 4505 221380 4509 221436
rect 4445 221376 4509 221380
rect 4525 221436 4589 221440
rect 4525 221380 4529 221436
rect 4529 221380 4585 221436
rect 4585 221380 4589 221436
rect 4525 221376 4589 221380
rect 7618 221436 7682 221440
rect 7618 221380 7622 221436
rect 7622 221380 7678 221436
rect 7678 221380 7682 221436
rect 7618 221376 7682 221380
rect 7698 221436 7762 221440
rect 7698 221380 7702 221436
rect 7702 221380 7758 221436
rect 7758 221380 7762 221436
rect 7698 221376 7762 221380
rect 7778 221436 7842 221440
rect 7778 221380 7782 221436
rect 7782 221380 7838 221436
rect 7838 221380 7842 221436
rect 7778 221376 7842 221380
rect 7858 221436 7922 221440
rect 7858 221380 7862 221436
rect 7862 221380 7918 221436
rect 7918 221380 7922 221436
rect 7858 221376 7922 221380
rect 2618 220892 2682 220896
rect 2618 220836 2622 220892
rect 2622 220836 2678 220892
rect 2678 220836 2682 220892
rect 2618 220832 2682 220836
rect 2698 220892 2762 220896
rect 2698 220836 2702 220892
rect 2702 220836 2758 220892
rect 2758 220836 2762 220892
rect 2698 220832 2762 220836
rect 2778 220892 2842 220896
rect 2778 220836 2782 220892
rect 2782 220836 2838 220892
rect 2838 220836 2842 220892
rect 2778 220832 2842 220836
rect 2858 220892 2922 220896
rect 2858 220836 2862 220892
rect 2862 220836 2918 220892
rect 2918 220836 2922 220892
rect 2858 220832 2922 220836
rect 5952 220892 6016 220896
rect 5952 220836 5956 220892
rect 5956 220836 6012 220892
rect 6012 220836 6016 220892
rect 5952 220832 6016 220836
rect 6032 220892 6096 220896
rect 6032 220836 6036 220892
rect 6036 220836 6092 220892
rect 6092 220836 6096 220892
rect 6032 220832 6096 220836
rect 6112 220892 6176 220896
rect 6112 220836 6116 220892
rect 6116 220836 6172 220892
rect 6172 220836 6176 220892
rect 6112 220832 6176 220836
rect 6192 220892 6256 220896
rect 6192 220836 6196 220892
rect 6196 220836 6252 220892
rect 6252 220836 6256 220892
rect 6192 220832 6256 220836
rect 4285 220348 4349 220352
rect 4285 220292 4289 220348
rect 4289 220292 4345 220348
rect 4345 220292 4349 220348
rect 4285 220288 4349 220292
rect 4365 220348 4429 220352
rect 4365 220292 4369 220348
rect 4369 220292 4425 220348
rect 4425 220292 4429 220348
rect 4365 220288 4429 220292
rect 4445 220348 4509 220352
rect 4445 220292 4449 220348
rect 4449 220292 4505 220348
rect 4505 220292 4509 220348
rect 4445 220288 4509 220292
rect 4525 220348 4589 220352
rect 4525 220292 4529 220348
rect 4529 220292 4585 220348
rect 4585 220292 4589 220348
rect 4525 220288 4589 220292
rect 7618 220348 7682 220352
rect 7618 220292 7622 220348
rect 7622 220292 7678 220348
rect 7678 220292 7682 220348
rect 7618 220288 7682 220292
rect 7698 220348 7762 220352
rect 7698 220292 7702 220348
rect 7702 220292 7758 220348
rect 7758 220292 7762 220348
rect 7698 220288 7762 220292
rect 7778 220348 7842 220352
rect 7778 220292 7782 220348
rect 7782 220292 7838 220348
rect 7838 220292 7842 220348
rect 7778 220288 7842 220292
rect 7858 220348 7922 220352
rect 7858 220292 7862 220348
rect 7862 220292 7918 220348
rect 7918 220292 7922 220348
rect 7858 220288 7922 220292
rect 2618 219804 2682 219808
rect 2618 219748 2622 219804
rect 2622 219748 2678 219804
rect 2678 219748 2682 219804
rect 2618 219744 2682 219748
rect 2698 219804 2762 219808
rect 2698 219748 2702 219804
rect 2702 219748 2758 219804
rect 2758 219748 2762 219804
rect 2698 219744 2762 219748
rect 2778 219804 2842 219808
rect 2778 219748 2782 219804
rect 2782 219748 2838 219804
rect 2838 219748 2842 219804
rect 2778 219744 2842 219748
rect 2858 219804 2922 219808
rect 2858 219748 2862 219804
rect 2862 219748 2918 219804
rect 2918 219748 2922 219804
rect 2858 219744 2922 219748
rect 5952 219804 6016 219808
rect 5952 219748 5956 219804
rect 5956 219748 6012 219804
rect 6012 219748 6016 219804
rect 5952 219744 6016 219748
rect 6032 219804 6096 219808
rect 6032 219748 6036 219804
rect 6036 219748 6092 219804
rect 6092 219748 6096 219804
rect 6032 219744 6096 219748
rect 6112 219804 6176 219808
rect 6112 219748 6116 219804
rect 6116 219748 6172 219804
rect 6172 219748 6176 219804
rect 6112 219744 6176 219748
rect 6192 219804 6256 219808
rect 6192 219748 6196 219804
rect 6196 219748 6252 219804
rect 6252 219748 6256 219804
rect 6192 219744 6256 219748
rect 4285 219260 4349 219264
rect 4285 219204 4289 219260
rect 4289 219204 4345 219260
rect 4345 219204 4349 219260
rect 4285 219200 4349 219204
rect 4365 219260 4429 219264
rect 4365 219204 4369 219260
rect 4369 219204 4425 219260
rect 4425 219204 4429 219260
rect 4365 219200 4429 219204
rect 4445 219260 4509 219264
rect 4445 219204 4449 219260
rect 4449 219204 4505 219260
rect 4505 219204 4509 219260
rect 4445 219200 4509 219204
rect 4525 219260 4589 219264
rect 4525 219204 4529 219260
rect 4529 219204 4585 219260
rect 4585 219204 4589 219260
rect 4525 219200 4589 219204
rect 7618 219260 7682 219264
rect 7618 219204 7622 219260
rect 7622 219204 7678 219260
rect 7678 219204 7682 219260
rect 7618 219200 7682 219204
rect 7698 219260 7762 219264
rect 7698 219204 7702 219260
rect 7702 219204 7758 219260
rect 7758 219204 7762 219260
rect 7698 219200 7762 219204
rect 7778 219260 7842 219264
rect 7778 219204 7782 219260
rect 7782 219204 7838 219260
rect 7838 219204 7842 219260
rect 7778 219200 7842 219204
rect 7858 219260 7922 219264
rect 7858 219204 7862 219260
rect 7862 219204 7918 219260
rect 7918 219204 7922 219260
rect 7858 219200 7922 219204
rect 2618 218716 2682 218720
rect 2618 218660 2622 218716
rect 2622 218660 2678 218716
rect 2678 218660 2682 218716
rect 2618 218656 2682 218660
rect 2698 218716 2762 218720
rect 2698 218660 2702 218716
rect 2702 218660 2758 218716
rect 2758 218660 2762 218716
rect 2698 218656 2762 218660
rect 2778 218716 2842 218720
rect 2778 218660 2782 218716
rect 2782 218660 2838 218716
rect 2838 218660 2842 218716
rect 2778 218656 2842 218660
rect 2858 218716 2922 218720
rect 2858 218660 2862 218716
rect 2862 218660 2918 218716
rect 2918 218660 2922 218716
rect 2858 218656 2922 218660
rect 5952 218716 6016 218720
rect 5952 218660 5956 218716
rect 5956 218660 6012 218716
rect 6012 218660 6016 218716
rect 5952 218656 6016 218660
rect 6032 218716 6096 218720
rect 6032 218660 6036 218716
rect 6036 218660 6092 218716
rect 6092 218660 6096 218716
rect 6032 218656 6096 218660
rect 6112 218716 6176 218720
rect 6112 218660 6116 218716
rect 6116 218660 6172 218716
rect 6172 218660 6176 218716
rect 6112 218656 6176 218660
rect 6192 218716 6256 218720
rect 6192 218660 6196 218716
rect 6196 218660 6252 218716
rect 6252 218660 6256 218716
rect 6192 218656 6256 218660
rect 4285 218172 4349 218176
rect 4285 218116 4289 218172
rect 4289 218116 4345 218172
rect 4345 218116 4349 218172
rect 4285 218112 4349 218116
rect 4365 218172 4429 218176
rect 4365 218116 4369 218172
rect 4369 218116 4425 218172
rect 4425 218116 4429 218172
rect 4365 218112 4429 218116
rect 4445 218172 4509 218176
rect 4445 218116 4449 218172
rect 4449 218116 4505 218172
rect 4505 218116 4509 218172
rect 4445 218112 4509 218116
rect 4525 218172 4589 218176
rect 4525 218116 4529 218172
rect 4529 218116 4585 218172
rect 4585 218116 4589 218172
rect 4525 218112 4589 218116
rect 7618 218172 7682 218176
rect 7618 218116 7622 218172
rect 7622 218116 7678 218172
rect 7678 218116 7682 218172
rect 7618 218112 7682 218116
rect 7698 218172 7762 218176
rect 7698 218116 7702 218172
rect 7702 218116 7758 218172
rect 7758 218116 7762 218172
rect 7698 218112 7762 218116
rect 7778 218172 7842 218176
rect 7778 218116 7782 218172
rect 7782 218116 7838 218172
rect 7838 218116 7842 218172
rect 7778 218112 7842 218116
rect 7858 218172 7922 218176
rect 7858 218116 7862 218172
rect 7862 218116 7918 218172
rect 7918 218116 7922 218172
rect 7858 218112 7922 218116
rect 2618 217628 2682 217632
rect 2618 217572 2622 217628
rect 2622 217572 2678 217628
rect 2678 217572 2682 217628
rect 2618 217568 2682 217572
rect 2698 217628 2762 217632
rect 2698 217572 2702 217628
rect 2702 217572 2758 217628
rect 2758 217572 2762 217628
rect 2698 217568 2762 217572
rect 2778 217628 2842 217632
rect 2778 217572 2782 217628
rect 2782 217572 2838 217628
rect 2838 217572 2842 217628
rect 2778 217568 2842 217572
rect 2858 217628 2922 217632
rect 2858 217572 2862 217628
rect 2862 217572 2918 217628
rect 2918 217572 2922 217628
rect 2858 217568 2922 217572
rect 5952 217628 6016 217632
rect 5952 217572 5956 217628
rect 5956 217572 6012 217628
rect 6012 217572 6016 217628
rect 5952 217568 6016 217572
rect 6032 217628 6096 217632
rect 6032 217572 6036 217628
rect 6036 217572 6092 217628
rect 6092 217572 6096 217628
rect 6032 217568 6096 217572
rect 6112 217628 6176 217632
rect 6112 217572 6116 217628
rect 6116 217572 6172 217628
rect 6172 217572 6176 217628
rect 6112 217568 6176 217572
rect 6192 217628 6256 217632
rect 6192 217572 6196 217628
rect 6196 217572 6252 217628
rect 6252 217572 6256 217628
rect 6192 217568 6256 217572
rect 4285 217084 4349 217088
rect 4285 217028 4289 217084
rect 4289 217028 4345 217084
rect 4345 217028 4349 217084
rect 4285 217024 4349 217028
rect 4365 217084 4429 217088
rect 4365 217028 4369 217084
rect 4369 217028 4425 217084
rect 4425 217028 4429 217084
rect 4365 217024 4429 217028
rect 4445 217084 4509 217088
rect 4445 217028 4449 217084
rect 4449 217028 4505 217084
rect 4505 217028 4509 217084
rect 4445 217024 4509 217028
rect 4525 217084 4589 217088
rect 4525 217028 4529 217084
rect 4529 217028 4585 217084
rect 4585 217028 4589 217084
rect 4525 217024 4589 217028
rect 7618 217084 7682 217088
rect 7618 217028 7622 217084
rect 7622 217028 7678 217084
rect 7678 217028 7682 217084
rect 7618 217024 7682 217028
rect 7698 217084 7762 217088
rect 7698 217028 7702 217084
rect 7702 217028 7758 217084
rect 7758 217028 7762 217084
rect 7698 217024 7762 217028
rect 7778 217084 7842 217088
rect 7778 217028 7782 217084
rect 7782 217028 7838 217084
rect 7838 217028 7842 217084
rect 7778 217024 7842 217028
rect 7858 217084 7922 217088
rect 7858 217028 7862 217084
rect 7862 217028 7918 217084
rect 7918 217028 7922 217084
rect 7858 217024 7922 217028
rect 2618 216540 2682 216544
rect 2618 216484 2622 216540
rect 2622 216484 2678 216540
rect 2678 216484 2682 216540
rect 2618 216480 2682 216484
rect 2698 216540 2762 216544
rect 2698 216484 2702 216540
rect 2702 216484 2758 216540
rect 2758 216484 2762 216540
rect 2698 216480 2762 216484
rect 2778 216540 2842 216544
rect 2778 216484 2782 216540
rect 2782 216484 2838 216540
rect 2838 216484 2842 216540
rect 2778 216480 2842 216484
rect 2858 216540 2922 216544
rect 2858 216484 2862 216540
rect 2862 216484 2918 216540
rect 2918 216484 2922 216540
rect 2858 216480 2922 216484
rect 5952 216540 6016 216544
rect 5952 216484 5956 216540
rect 5956 216484 6012 216540
rect 6012 216484 6016 216540
rect 5952 216480 6016 216484
rect 6032 216540 6096 216544
rect 6032 216484 6036 216540
rect 6036 216484 6092 216540
rect 6092 216484 6096 216540
rect 6032 216480 6096 216484
rect 6112 216540 6176 216544
rect 6112 216484 6116 216540
rect 6116 216484 6172 216540
rect 6172 216484 6176 216540
rect 6112 216480 6176 216484
rect 6192 216540 6256 216544
rect 6192 216484 6196 216540
rect 6196 216484 6252 216540
rect 6252 216484 6256 216540
rect 6192 216480 6256 216484
rect 4285 215996 4349 216000
rect 4285 215940 4289 215996
rect 4289 215940 4345 215996
rect 4345 215940 4349 215996
rect 4285 215936 4349 215940
rect 4365 215996 4429 216000
rect 4365 215940 4369 215996
rect 4369 215940 4425 215996
rect 4425 215940 4429 215996
rect 4365 215936 4429 215940
rect 4445 215996 4509 216000
rect 4445 215940 4449 215996
rect 4449 215940 4505 215996
rect 4505 215940 4509 215996
rect 4445 215936 4509 215940
rect 4525 215996 4589 216000
rect 4525 215940 4529 215996
rect 4529 215940 4585 215996
rect 4585 215940 4589 215996
rect 4525 215936 4589 215940
rect 7618 215996 7682 216000
rect 7618 215940 7622 215996
rect 7622 215940 7678 215996
rect 7678 215940 7682 215996
rect 7618 215936 7682 215940
rect 7698 215996 7762 216000
rect 7698 215940 7702 215996
rect 7702 215940 7758 215996
rect 7758 215940 7762 215996
rect 7698 215936 7762 215940
rect 7778 215996 7842 216000
rect 7778 215940 7782 215996
rect 7782 215940 7838 215996
rect 7838 215940 7842 215996
rect 7778 215936 7842 215940
rect 7858 215996 7922 216000
rect 7858 215940 7862 215996
rect 7862 215940 7918 215996
rect 7918 215940 7922 215996
rect 7858 215936 7922 215940
rect 2618 215452 2682 215456
rect 2618 215396 2622 215452
rect 2622 215396 2678 215452
rect 2678 215396 2682 215452
rect 2618 215392 2682 215396
rect 2698 215452 2762 215456
rect 2698 215396 2702 215452
rect 2702 215396 2758 215452
rect 2758 215396 2762 215452
rect 2698 215392 2762 215396
rect 2778 215452 2842 215456
rect 2778 215396 2782 215452
rect 2782 215396 2838 215452
rect 2838 215396 2842 215452
rect 2778 215392 2842 215396
rect 2858 215452 2922 215456
rect 2858 215396 2862 215452
rect 2862 215396 2918 215452
rect 2918 215396 2922 215452
rect 2858 215392 2922 215396
rect 5952 215452 6016 215456
rect 5952 215396 5956 215452
rect 5956 215396 6012 215452
rect 6012 215396 6016 215452
rect 5952 215392 6016 215396
rect 6032 215452 6096 215456
rect 6032 215396 6036 215452
rect 6036 215396 6092 215452
rect 6092 215396 6096 215452
rect 6032 215392 6096 215396
rect 6112 215452 6176 215456
rect 6112 215396 6116 215452
rect 6116 215396 6172 215452
rect 6172 215396 6176 215452
rect 6112 215392 6176 215396
rect 6192 215452 6256 215456
rect 6192 215396 6196 215452
rect 6196 215396 6252 215452
rect 6252 215396 6256 215452
rect 6192 215392 6256 215396
rect 4285 214908 4349 214912
rect 4285 214852 4289 214908
rect 4289 214852 4345 214908
rect 4345 214852 4349 214908
rect 4285 214848 4349 214852
rect 4365 214908 4429 214912
rect 4365 214852 4369 214908
rect 4369 214852 4425 214908
rect 4425 214852 4429 214908
rect 4365 214848 4429 214852
rect 4445 214908 4509 214912
rect 4445 214852 4449 214908
rect 4449 214852 4505 214908
rect 4505 214852 4509 214908
rect 4445 214848 4509 214852
rect 4525 214908 4589 214912
rect 4525 214852 4529 214908
rect 4529 214852 4585 214908
rect 4585 214852 4589 214908
rect 4525 214848 4589 214852
rect 7618 214908 7682 214912
rect 7618 214852 7622 214908
rect 7622 214852 7678 214908
rect 7678 214852 7682 214908
rect 7618 214848 7682 214852
rect 7698 214908 7762 214912
rect 7698 214852 7702 214908
rect 7702 214852 7758 214908
rect 7758 214852 7762 214908
rect 7698 214848 7762 214852
rect 7778 214908 7842 214912
rect 7778 214852 7782 214908
rect 7782 214852 7838 214908
rect 7838 214852 7842 214908
rect 7778 214848 7842 214852
rect 7858 214908 7922 214912
rect 7858 214852 7862 214908
rect 7862 214852 7918 214908
rect 7918 214852 7922 214908
rect 7858 214848 7922 214852
rect 2618 214364 2682 214368
rect 2618 214308 2622 214364
rect 2622 214308 2678 214364
rect 2678 214308 2682 214364
rect 2618 214304 2682 214308
rect 2698 214364 2762 214368
rect 2698 214308 2702 214364
rect 2702 214308 2758 214364
rect 2758 214308 2762 214364
rect 2698 214304 2762 214308
rect 2778 214364 2842 214368
rect 2778 214308 2782 214364
rect 2782 214308 2838 214364
rect 2838 214308 2842 214364
rect 2778 214304 2842 214308
rect 2858 214364 2922 214368
rect 2858 214308 2862 214364
rect 2862 214308 2918 214364
rect 2918 214308 2922 214364
rect 2858 214304 2922 214308
rect 5952 214364 6016 214368
rect 5952 214308 5956 214364
rect 5956 214308 6012 214364
rect 6012 214308 6016 214364
rect 5952 214304 6016 214308
rect 6032 214364 6096 214368
rect 6032 214308 6036 214364
rect 6036 214308 6092 214364
rect 6092 214308 6096 214364
rect 6032 214304 6096 214308
rect 6112 214364 6176 214368
rect 6112 214308 6116 214364
rect 6116 214308 6172 214364
rect 6172 214308 6176 214364
rect 6112 214304 6176 214308
rect 6192 214364 6256 214368
rect 6192 214308 6196 214364
rect 6196 214308 6252 214364
rect 6252 214308 6256 214364
rect 6192 214304 6256 214308
rect 4285 213820 4349 213824
rect 4285 213764 4289 213820
rect 4289 213764 4345 213820
rect 4345 213764 4349 213820
rect 4285 213760 4349 213764
rect 4365 213820 4429 213824
rect 4365 213764 4369 213820
rect 4369 213764 4425 213820
rect 4425 213764 4429 213820
rect 4365 213760 4429 213764
rect 4445 213820 4509 213824
rect 4445 213764 4449 213820
rect 4449 213764 4505 213820
rect 4505 213764 4509 213820
rect 4445 213760 4509 213764
rect 4525 213820 4589 213824
rect 4525 213764 4529 213820
rect 4529 213764 4585 213820
rect 4585 213764 4589 213820
rect 4525 213760 4589 213764
rect 7618 213820 7682 213824
rect 7618 213764 7622 213820
rect 7622 213764 7678 213820
rect 7678 213764 7682 213820
rect 7618 213760 7682 213764
rect 7698 213820 7762 213824
rect 7698 213764 7702 213820
rect 7702 213764 7758 213820
rect 7758 213764 7762 213820
rect 7698 213760 7762 213764
rect 7778 213820 7842 213824
rect 7778 213764 7782 213820
rect 7782 213764 7838 213820
rect 7838 213764 7842 213820
rect 7778 213760 7842 213764
rect 7858 213820 7922 213824
rect 7858 213764 7862 213820
rect 7862 213764 7918 213820
rect 7918 213764 7922 213820
rect 7858 213760 7922 213764
rect 2618 213276 2682 213280
rect 2618 213220 2622 213276
rect 2622 213220 2678 213276
rect 2678 213220 2682 213276
rect 2618 213216 2682 213220
rect 2698 213276 2762 213280
rect 2698 213220 2702 213276
rect 2702 213220 2758 213276
rect 2758 213220 2762 213276
rect 2698 213216 2762 213220
rect 2778 213276 2842 213280
rect 2778 213220 2782 213276
rect 2782 213220 2838 213276
rect 2838 213220 2842 213276
rect 2778 213216 2842 213220
rect 2858 213276 2922 213280
rect 2858 213220 2862 213276
rect 2862 213220 2918 213276
rect 2918 213220 2922 213276
rect 2858 213216 2922 213220
rect 5952 213276 6016 213280
rect 5952 213220 5956 213276
rect 5956 213220 6012 213276
rect 6012 213220 6016 213276
rect 5952 213216 6016 213220
rect 6032 213276 6096 213280
rect 6032 213220 6036 213276
rect 6036 213220 6092 213276
rect 6092 213220 6096 213276
rect 6032 213216 6096 213220
rect 6112 213276 6176 213280
rect 6112 213220 6116 213276
rect 6116 213220 6172 213276
rect 6172 213220 6176 213276
rect 6112 213216 6176 213220
rect 6192 213276 6256 213280
rect 6192 213220 6196 213276
rect 6196 213220 6252 213276
rect 6252 213220 6256 213276
rect 6192 213216 6256 213220
rect 4285 212732 4349 212736
rect 4285 212676 4289 212732
rect 4289 212676 4345 212732
rect 4345 212676 4349 212732
rect 4285 212672 4349 212676
rect 4365 212732 4429 212736
rect 4365 212676 4369 212732
rect 4369 212676 4425 212732
rect 4425 212676 4429 212732
rect 4365 212672 4429 212676
rect 4445 212732 4509 212736
rect 4445 212676 4449 212732
rect 4449 212676 4505 212732
rect 4505 212676 4509 212732
rect 4445 212672 4509 212676
rect 4525 212732 4589 212736
rect 4525 212676 4529 212732
rect 4529 212676 4585 212732
rect 4585 212676 4589 212732
rect 4525 212672 4589 212676
rect 7618 212732 7682 212736
rect 7618 212676 7622 212732
rect 7622 212676 7678 212732
rect 7678 212676 7682 212732
rect 7618 212672 7682 212676
rect 7698 212732 7762 212736
rect 7698 212676 7702 212732
rect 7702 212676 7758 212732
rect 7758 212676 7762 212732
rect 7698 212672 7762 212676
rect 7778 212732 7842 212736
rect 7778 212676 7782 212732
rect 7782 212676 7838 212732
rect 7838 212676 7842 212732
rect 7778 212672 7842 212676
rect 7858 212732 7922 212736
rect 7858 212676 7862 212732
rect 7862 212676 7918 212732
rect 7918 212676 7922 212732
rect 7858 212672 7922 212676
rect 2618 212188 2682 212192
rect 2618 212132 2622 212188
rect 2622 212132 2678 212188
rect 2678 212132 2682 212188
rect 2618 212128 2682 212132
rect 2698 212188 2762 212192
rect 2698 212132 2702 212188
rect 2702 212132 2758 212188
rect 2758 212132 2762 212188
rect 2698 212128 2762 212132
rect 2778 212188 2842 212192
rect 2778 212132 2782 212188
rect 2782 212132 2838 212188
rect 2838 212132 2842 212188
rect 2778 212128 2842 212132
rect 2858 212188 2922 212192
rect 2858 212132 2862 212188
rect 2862 212132 2918 212188
rect 2918 212132 2922 212188
rect 2858 212128 2922 212132
rect 5952 212188 6016 212192
rect 5952 212132 5956 212188
rect 5956 212132 6012 212188
rect 6012 212132 6016 212188
rect 5952 212128 6016 212132
rect 6032 212188 6096 212192
rect 6032 212132 6036 212188
rect 6036 212132 6092 212188
rect 6092 212132 6096 212188
rect 6032 212128 6096 212132
rect 6112 212188 6176 212192
rect 6112 212132 6116 212188
rect 6116 212132 6172 212188
rect 6172 212132 6176 212188
rect 6112 212128 6176 212132
rect 6192 212188 6256 212192
rect 6192 212132 6196 212188
rect 6196 212132 6252 212188
rect 6252 212132 6256 212188
rect 6192 212128 6256 212132
rect 4285 211644 4349 211648
rect 4285 211588 4289 211644
rect 4289 211588 4345 211644
rect 4345 211588 4349 211644
rect 4285 211584 4349 211588
rect 4365 211644 4429 211648
rect 4365 211588 4369 211644
rect 4369 211588 4425 211644
rect 4425 211588 4429 211644
rect 4365 211584 4429 211588
rect 4445 211644 4509 211648
rect 4445 211588 4449 211644
rect 4449 211588 4505 211644
rect 4505 211588 4509 211644
rect 4445 211584 4509 211588
rect 4525 211644 4589 211648
rect 4525 211588 4529 211644
rect 4529 211588 4585 211644
rect 4585 211588 4589 211644
rect 4525 211584 4589 211588
rect 7618 211644 7682 211648
rect 7618 211588 7622 211644
rect 7622 211588 7678 211644
rect 7678 211588 7682 211644
rect 7618 211584 7682 211588
rect 7698 211644 7762 211648
rect 7698 211588 7702 211644
rect 7702 211588 7758 211644
rect 7758 211588 7762 211644
rect 7698 211584 7762 211588
rect 7778 211644 7842 211648
rect 7778 211588 7782 211644
rect 7782 211588 7838 211644
rect 7838 211588 7842 211644
rect 7778 211584 7842 211588
rect 7858 211644 7922 211648
rect 7858 211588 7862 211644
rect 7862 211588 7918 211644
rect 7918 211588 7922 211644
rect 7858 211584 7922 211588
rect 2618 211100 2682 211104
rect 2618 211044 2622 211100
rect 2622 211044 2678 211100
rect 2678 211044 2682 211100
rect 2618 211040 2682 211044
rect 2698 211100 2762 211104
rect 2698 211044 2702 211100
rect 2702 211044 2758 211100
rect 2758 211044 2762 211100
rect 2698 211040 2762 211044
rect 2778 211100 2842 211104
rect 2778 211044 2782 211100
rect 2782 211044 2838 211100
rect 2838 211044 2842 211100
rect 2778 211040 2842 211044
rect 2858 211100 2922 211104
rect 2858 211044 2862 211100
rect 2862 211044 2918 211100
rect 2918 211044 2922 211100
rect 2858 211040 2922 211044
rect 5952 211100 6016 211104
rect 5952 211044 5956 211100
rect 5956 211044 6012 211100
rect 6012 211044 6016 211100
rect 5952 211040 6016 211044
rect 6032 211100 6096 211104
rect 6032 211044 6036 211100
rect 6036 211044 6092 211100
rect 6092 211044 6096 211100
rect 6032 211040 6096 211044
rect 6112 211100 6176 211104
rect 6112 211044 6116 211100
rect 6116 211044 6172 211100
rect 6172 211044 6176 211100
rect 6112 211040 6176 211044
rect 6192 211100 6256 211104
rect 6192 211044 6196 211100
rect 6196 211044 6252 211100
rect 6252 211044 6256 211100
rect 6192 211040 6256 211044
rect 4285 210556 4349 210560
rect 4285 210500 4289 210556
rect 4289 210500 4345 210556
rect 4345 210500 4349 210556
rect 4285 210496 4349 210500
rect 4365 210556 4429 210560
rect 4365 210500 4369 210556
rect 4369 210500 4425 210556
rect 4425 210500 4429 210556
rect 4365 210496 4429 210500
rect 4445 210556 4509 210560
rect 4445 210500 4449 210556
rect 4449 210500 4505 210556
rect 4505 210500 4509 210556
rect 4445 210496 4509 210500
rect 4525 210556 4589 210560
rect 4525 210500 4529 210556
rect 4529 210500 4585 210556
rect 4585 210500 4589 210556
rect 4525 210496 4589 210500
rect 7618 210556 7682 210560
rect 7618 210500 7622 210556
rect 7622 210500 7678 210556
rect 7678 210500 7682 210556
rect 7618 210496 7682 210500
rect 7698 210556 7762 210560
rect 7698 210500 7702 210556
rect 7702 210500 7758 210556
rect 7758 210500 7762 210556
rect 7698 210496 7762 210500
rect 7778 210556 7842 210560
rect 7778 210500 7782 210556
rect 7782 210500 7838 210556
rect 7838 210500 7842 210556
rect 7778 210496 7842 210500
rect 7858 210556 7922 210560
rect 7858 210500 7862 210556
rect 7862 210500 7918 210556
rect 7918 210500 7922 210556
rect 7858 210496 7922 210500
rect 2618 210012 2682 210016
rect 2618 209956 2622 210012
rect 2622 209956 2678 210012
rect 2678 209956 2682 210012
rect 2618 209952 2682 209956
rect 2698 210012 2762 210016
rect 2698 209956 2702 210012
rect 2702 209956 2758 210012
rect 2758 209956 2762 210012
rect 2698 209952 2762 209956
rect 2778 210012 2842 210016
rect 2778 209956 2782 210012
rect 2782 209956 2838 210012
rect 2838 209956 2842 210012
rect 2778 209952 2842 209956
rect 2858 210012 2922 210016
rect 2858 209956 2862 210012
rect 2862 209956 2918 210012
rect 2918 209956 2922 210012
rect 2858 209952 2922 209956
rect 5952 210012 6016 210016
rect 5952 209956 5956 210012
rect 5956 209956 6012 210012
rect 6012 209956 6016 210012
rect 5952 209952 6016 209956
rect 6032 210012 6096 210016
rect 6032 209956 6036 210012
rect 6036 209956 6092 210012
rect 6092 209956 6096 210012
rect 6032 209952 6096 209956
rect 6112 210012 6176 210016
rect 6112 209956 6116 210012
rect 6116 209956 6172 210012
rect 6172 209956 6176 210012
rect 6112 209952 6176 209956
rect 6192 210012 6256 210016
rect 6192 209956 6196 210012
rect 6196 209956 6252 210012
rect 6252 209956 6256 210012
rect 6192 209952 6256 209956
rect 4285 209468 4349 209472
rect 4285 209412 4289 209468
rect 4289 209412 4345 209468
rect 4345 209412 4349 209468
rect 4285 209408 4349 209412
rect 4365 209468 4429 209472
rect 4365 209412 4369 209468
rect 4369 209412 4425 209468
rect 4425 209412 4429 209468
rect 4365 209408 4429 209412
rect 4445 209468 4509 209472
rect 4445 209412 4449 209468
rect 4449 209412 4505 209468
rect 4505 209412 4509 209468
rect 4445 209408 4509 209412
rect 4525 209468 4589 209472
rect 4525 209412 4529 209468
rect 4529 209412 4585 209468
rect 4585 209412 4589 209468
rect 4525 209408 4589 209412
rect 7618 209468 7682 209472
rect 7618 209412 7622 209468
rect 7622 209412 7678 209468
rect 7678 209412 7682 209468
rect 7618 209408 7682 209412
rect 7698 209468 7762 209472
rect 7698 209412 7702 209468
rect 7702 209412 7758 209468
rect 7758 209412 7762 209468
rect 7698 209408 7762 209412
rect 7778 209468 7842 209472
rect 7778 209412 7782 209468
rect 7782 209412 7838 209468
rect 7838 209412 7842 209468
rect 7778 209408 7842 209412
rect 7858 209468 7922 209472
rect 7858 209412 7862 209468
rect 7862 209412 7918 209468
rect 7918 209412 7922 209468
rect 7858 209408 7922 209412
rect 2618 208924 2682 208928
rect 2618 208868 2622 208924
rect 2622 208868 2678 208924
rect 2678 208868 2682 208924
rect 2618 208864 2682 208868
rect 2698 208924 2762 208928
rect 2698 208868 2702 208924
rect 2702 208868 2758 208924
rect 2758 208868 2762 208924
rect 2698 208864 2762 208868
rect 2778 208924 2842 208928
rect 2778 208868 2782 208924
rect 2782 208868 2838 208924
rect 2838 208868 2842 208924
rect 2778 208864 2842 208868
rect 2858 208924 2922 208928
rect 2858 208868 2862 208924
rect 2862 208868 2918 208924
rect 2918 208868 2922 208924
rect 2858 208864 2922 208868
rect 5952 208924 6016 208928
rect 5952 208868 5956 208924
rect 5956 208868 6012 208924
rect 6012 208868 6016 208924
rect 5952 208864 6016 208868
rect 6032 208924 6096 208928
rect 6032 208868 6036 208924
rect 6036 208868 6092 208924
rect 6092 208868 6096 208924
rect 6032 208864 6096 208868
rect 6112 208924 6176 208928
rect 6112 208868 6116 208924
rect 6116 208868 6172 208924
rect 6172 208868 6176 208924
rect 6112 208864 6176 208868
rect 6192 208924 6256 208928
rect 6192 208868 6196 208924
rect 6196 208868 6252 208924
rect 6252 208868 6256 208924
rect 6192 208864 6256 208868
rect 4285 208380 4349 208384
rect 4285 208324 4289 208380
rect 4289 208324 4345 208380
rect 4345 208324 4349 208380
rect 4285 208320 4349 208324
rect 4365 208380 4429 208384
rect 4365 208324 4369 208380
rect 4369 208324 4425 208380
rect 4425 208324 4429 208380
rect 4365 208320 4429 208324
rect 4445 208380 4509 208384
rect 4445 208324 4449 208380
rect 4449 208324 4505 208380
rect 4505 208324 4509 208380
rect 4445 208320 4509 208324
rect 4525 208380 4589 208384
rect 4525 208324 4529 208380
rect 4529 208324 4585 208380
rect 4585 208324 4589 208380
rect 4525 208320 4589 208324
rect 7618 208380 7682 208384
rect 7618 208324 7622 208380
rect 7622 208324 7678 208380
rect 7678 208324 7682 208380
rect 7618 208320 7682 208324
rect 7698 208380 7762 208384
rect 7698 208324 7702 208380
rect 7702 208324 7758 208380
rect 7758 208324 7762 208380
rect 7698 208320 7762 208324
rect 7778 208380 7842 208384
rect 7778 208324 7782 208380
rect 7782 208324 7838 208380
rect 7838 208324 7842 208380
rect 7778 208320 7842 208324
rect 7858 208380 7922 208384
rect 7858 208324 7862 208380
rect 7862 208324 7918 208380
rect 7918 208324 7922 208380
rect 7858 208320 7922 208324
rect 2618 207836 2682 207840
rect 2618 207780 2622 207836
rect 2622 207780 2678 207836
rect 2678 207780 2682 207836
rect 2618 207776 2682 207780
rect 2698 207836 2762 207840
rect 2698 207780 2702 207836
rect 2702 207780 2758 207836
rect 2758 207780 2762 207836
rect 2698 207776 2762 207780
rect 2778 207836 2842 207840
rect 2778 207780 2782 207836
rect 2782 207780 2838 207836
rect 2838 207780 2842 207836
rect 2778 207776 2842 207780
rect 2858 207836 2922 207840
rect 2858 207780 2862 207836
rect 2862 207780 2918 207836
rect 2918 207780 2922 207836
rect 2858 207776 2922 207780
rect 5952 207836 6016 207840
rect 5952 207780 5956 207836
rect 5956 207780 6012 207836
rect 6012 207780 6016 207836
rect 5952 207776 6016 207780
rect 6032 207836 6096 207840
rect 6032 207780 6036 207836
rect 6036 207780 6092 207836
rect 6092 207780 6096 207836
rect 6032 207776 6096 207780
rect 6112 207836 6176 207840
rect 6112 207780 6116 207836
rect 6116 207780 6172 207836
rect 6172 207780 6176 207836
rect 6112 207776 6176 207780
rect 6192 207836 6256 207840
rect 6192 207780 6196 207836
rect 6196 207780 6252 207836
rect 6252 207780 6256 207836
rect 6192 207776 6256 207780
rect 4285 207292 4349 207296
rect 4285 207236 4289 207292
rect 4289 207236 4345 207292
rect 4345 207236 4349 207292
rect 4285 207232 4349 207236
rect 4365 207292 4429 207296
rect 4365 207236 4369 207292
rect 4369 207236 4425 207292
rect 4425 207236 4429 207292
rect 4365 207232 4429 207236
rect 4445 207292 4509 207296
rect 4445 207236 4449 207292
rect 4449 207236 4505 207292
rect 4505 207236 4509 207292
rect 4445 207232 4509 207236
rect 4525 207292 4589 207296
rect 4525 207236 4529 207292
rect 4529 207236 4585 207292
rect 4585 207236 4589 207292
rect 4525 207232 4589 207236
rect 7618 207292 7682 207296
rect 7618 207236 7622 207292
rect 7622 207236 7678 207292
rect 7678 207236 7682 207292
rect 7618 207232 7682 207236
rect 7698 207292 7762 207296
rect 7698 207236 7702 207292
rect 7702 207236 7758 207292
rect 7758 207236 7762 207292
rect 7698 207232 7762 207236
rect 7778 207292 7842 207296
rect 7778 207236 7782 207292
rect 7782 207236 7838 207292
rect 7838 207236 7842 207292
rect 7778 207232 7842 207236
rect 7858 207292 7922 207296
rect 7858 207236 7862 207292
rect 7862 207236 7918 207292
rect 7918 207236 7922 207292
rect 7858 207232 7922 207236
rect 2618 206748 2682 206752
rect 2618 206692 2622 206748
rect 2622 206692 2678 206748
rect 2678 206692 2682 206748
rect 2618 206688 2682 206692
rect 2698 206748 2762 206752
rect 2698 206692 2702 206748
rect 2702 206692 2758 206748
rect 2758 206692 2762 206748
rect 2698 206688 2762 206692
rect 2778 206748 2842 206752
rect 2778 206692 2782 206748
rect 2782 206692 2838 206748
rect 2838 206692 2842 206748
rect 2778 206688 2842 206692
rect 2858 206748 2922 206752
rect 2858 206692 2862 206748
rect 2862 206692 2918 206748
rect 2918 206692 2922 206748
rect 2858 206688 2922 206692
rect 5952 206748 6016 206752
rect 5952 206692 5956 206748
rect 5956 206692 6012 206748
rect 6012 206692 6016 206748
rect 5952 206688 6016 206692
rect 6032 206748 6096 206752
rect 6032 206692 6036 206748
rect 6036 206692 6092 206748
rect 6092 206692 6096 206748
rect 6032 206688 6096 206692
rect 6112 206748 6176 206752
rect 6112 206692 6116 206748
rect 6116 206692 6172 206748
rect 6172 206692 6176 206748
rect 6112 206688 6176 206692
rect 6192 206748 6256 206752
rect 6192 206692 6196 206748
rect 6196 206692 6252 206748
rect 6252 206692 6256 206748
rect 6192 206688 6256 206692
rect 4285 206204 4349 206208
rect 4285 206148 4289 206204
rect 4289 206148 4345 206204
rect 4345 206148 4349 206204
rect 4285 206144 4349 206148
rect 4365 206204 4429 206208
rect 4365 206148 4369 206204
rect 4369 206148 4425 206204
rect 4425 206148 4429 206204
rect 4365 206144 4429 206148
rect 4445 206204 4509 206208
rect 4445 206148 4449 206204
rect 4449 206148 4505 206204
rect 4505 206148 4509 206204
rect 4445 206144 4509 206148
rect 4525 206204 4589 206208
rect 4525 206148 4529 206204
rect 4529 206148 4585 206204
rect 4585 206148 4589 206204
rect 4525 206144 4589 206148
rect 7618 206204 7682 206208
rect 7618 206148 7622 206204
rect 7622 206148 7678 206204
rect 7678 206148 7682 206204
rect 7618 206144 7682 206148
rect 7698 206204 7762 206208
rect 7698 206148 7702 206204
rect 7702 206148 7758 206204
rect 7758 206148 7762 206204
rect 7698 206144 7762 206148
rect 7778 206204 7842 206208
rect 7778 206148 7782 206204
rect 7782 206148 7838 206204
rect 7838 206148 7842 206204
rect 7778 206144 7842 206148
rect 7858 206204 7922 206208
rect 7858 206148 7862 206204
rect 7862 206148 7918 206204
rect 7918 206148 7922 206204
rect 7858 206144 7922 206148
rect 2618 205660 2682 205664
rect 2618 205604 2622 205660
rect 2622 205604 2678 205660
rect 2678 205604 2682 205660
rect 2618 205600 2682 205604
rect 2698 205660 2762 205664
rect 2698 205604 2702 205660
rect 2702 205604 2758 205660
rect 2758 205604 2762 205660
rect 2698 205600 2762 205604
rect 2778 205660 2842 205664
rect 2778 205604 2782 205660
rect 2782 205604 2838 205660
rect 2838 205604 2842 205660
rect 2778 205600 2842 205604
rect 2858 205660 2922 205664
rect 2858 205604 2862 205660
rect 2862 205604 2918 205660
rect 2918 205604 2922 205660
rect 2858 205600 2922 205604
rect 5952 205660 6016 205664
rect 5952 205604 5956 205660
rect 5956 205604 6012 205660
rect 6012 205604 6016 205660
rect 5952 205600 6016 205604
rect 6032 205660 6096 205664
rect 6032 205604 6036 205660
rect 6036 205604 6092 205660
rect 6092 205604 6096 205660
rect 6032 205600 6096 205604
rect 6112 205660 6176 205664
rect 6112 205604 6116 205660
rect 6116 205604 6172 205660
rect 6172 205604 6176 205660
rect 6112 205600 6176 205604
rect 6192 205660 6256 205664
rect 6192 205604 6196 205660
rect 6196 205604 6252 205660
rect 6252 205604 6256 205660
rect 6192 205600 6256 205604
rect 4285 205116 4349 205120
rect 4285 205060 4289 205116
rect 4289 205060 4345 205116
rect 4345 205060 4349 205116
rect 4285 205056 4349 205060
rect 4365 205116 4429 205120
rect 4365 205060 4369 205116
rect 4369 205060 4425 205116
rect 4425 205060 4429 205116
rect 4365 205056 4429 205060
rect 4445 205116 4509 205120
rect 4445 205060 4449 205116
rect 4449 205060 4505 205116
rect 4505 205060 4509 205116
rect 4445 205056 4509 205060
rect 4525 205116 4589 205120
rect 4525 205060 4529 205116
rect 4529 205060 4585 205116
rect 4585 205060 4589 205116
rect 4525 205056 4589 205060
rect 7618 205116 7682 205120
rect 7618 205060 7622 205116
rect 7622 205060 7678 205116
rect 7678 205060 7682 205116
rect 7618 205056 7682 205060
rect 7698 205116 7762 205120
rect 7698 205060 7702 205116
rect 7702 205060 7758 205116
rect 7758 205060 7762 205116
rect 7698 205056 7762 205060
rect 7778 205116 7842 205120
rect 7778 205060 7782 205116
rect 7782 205060 7838 205116
rect 7838 205060 7842 205116
rect 7778 205056 7842 205060
rect 7858 205116 7922 205120
rect 7858 205060 7862 205116
rect 7862 205060 7918 205116
rect 7918 205060 7922 205116
rect 7858 205056 7922 205060
rect 2618 204572 2682 204576
rect 2618 204516 2622 204572
rect 2622 204516 2678 204572
rect 2678 204516 2682 204572
rect 2618 204512 2682 204516
rect 2698 204572 2762 204576
rect 2698 204516 2702 204572
rect 2702 204516 2758 204572
rect 2758 204516 2762 204572
rect 2698 204512 2762 204516
rect 2778 204572 2842 204576
rect 2778 204516 2782 204572
rect 2782 204516 2838 204572
rect 2838 204516 2842 204572
rect 2778 204512 2842 204516
rect 2858 204572 2922 204576
rect 2858 204516 2862 204572
rect 2862 204516 2918 204572
rect 2918 204516 2922 204572
rect 2858 204512 2922 204516
rect 5952 204572 6016 204576
rect 5952 204516 5956 204572
rect 5956 204516 6012 204572
rect 6012 204516 6016 204572
rect 5952 204512 6016 204516
rect 6032 204572 6096 204576
rect 6032 204516 6036 204572
rect 6036 204516 6092 204572
rect 6092 204516 6096 204572
rect 6032 204512 6096 204516
rect 6112 204572 6176 204576
rect 6112 204516 6116 204572
rect 6116 204516 6172 204572
rect 6172 204516 6176 204572
rect 6112 204512 6176 204516
rect 6192 204572 6256 204576
rect 6192 204516 6196 204572
rect 6196 204516 6252 204572
rect 6252 204516 6256 204572
rect 6192 204512 6256 204516
rect 4285 204028 4349 204032
rect 4285 203972 4289 204028
rect 4289 203972 4345 204028
rect 4345 203972 4349 204028
rect 4285 203968 4349 203972
rect 4365 204028 4429 204032
rect 4365 203972 4369 204028
rect 4369 203972 4425 204028
rect 4425 203972 4429 204028
rect 4365 203968 4429 203972
rect 4445 204028 4509 204032
rect 4445 203972 4449 204028
rect 4449 203972 4505 204028
rect 4505 203972 4509 204028
rect 4445 203968 4509 203972
rect 4525 204028 4589 204032
rect 4525 203972 4529 204028
rect 4529 203972 4585 204028
rect 4585 203972 4589 204028
rect 4525 203968 4589 203972
rect 7618 204028 7682 204032
rect 7618 203972 7622 204028
rect 7622 203972 7678 204028
rect 7678 203972 7682 204028
rect 7618 203968 7682 203972
rect 7698 204028 7762 204032
rect 7698 203972 7702 204028
rect 7702 203972 7758 204028
rect 7758 203972 7762 204028
rect 7698 203968 7762 203972
rect 7778 204028 7842 204032
rect 7778 203972 7782 204028
rect 7782 203972 7838 204028
rect 7838 203972 7842 204028
rect 7778 203968 7842 203972
rect 7858 204028 7922 204032
rect 7858 203972 7862 204028
rect 7862 203972 7918 204028
rect 7918 203972 7922 204028
rect 7858 203968 7922 203972
rect 2618 203484 2682 203488
rect 2618 203428 2622 203484
rect 2622 203428 2678 203484
rect 2678 203428 2682 203484
rect 2618 203424 2682 203428
rect 2698 203484 2762 203488
rect 2698 203428 2702 203484
rect 2702 203428 2758 203484
rect 2758 203428 2762 203484
rect 2698 203424 2762 203428
rect 2778 203484 2842 203488
rect 2778 203428 2782 203484
rect 2782 203428 2838 203484
rect 2838 203428 2842 203484
rect 2778 203424 2842 203428
rect 2858 203484 2922 203488
rect 2858 203428 2862 203484
rect 2862 203428 2918 203484
rect 2918 203428 2922 203484
rect 2858 203424 2922 203428
rect 5952 203484 6016 203488
rect 5952 203428 5956 203484
rect 5956 203428 6012 203484
rect 6012 203428 6016 203484
rect 5952 203424 6016 203428
rect 6032 203484 6096 203488
rect 6032 203428 6036 203484
rect 6036 203428 6092 203484
rect 6092 203428 6096 203484
rect 6032 203424 6096 203428
rect 6112 203484 6176 203488
rect 6112 203428 6116 203484
rect 6116 203428 6172 203484
rect 6172 203428 6176 203484
rect 6112 203424 6176 203428
rect 6192 203484 6256 203488
rect 6192 203428 6196 203484
rect 6196 203428 6252 203484
rect 6252 203428 6256 203484
rect 6192 203424 6256 203428
rect 4285 202940 4349 202944
rect 4285 202884 4289 202940
rect 4289 202884 4345 202940
rect 4345 202884 4349 202940
rect 4285 202880 4349 202884
rect 4365 202940 4429 202944
rect 4365 202884 4369 202940
rect 4369 202884 4425 202940
rect 4425 202884 4429 202940
rect 4365 202880 4429 202884
rect 4445 202940 4509 202944
rect 4445 202884 4449 202940
rect 4449 202884 4505 202940
rect 4505 202884 4509 202940
rect 4445 202880 4509 202884
rect 4525 202940 4589 202944
rect 4525 202884 4529 202940
rect 4529 202884 4585 202940
rect 4585 202884 4589 202940
rect 4525 202880 4589 202884
rect 7618 202940 7682 202944
rect 7618 202884 7622 202940
rect 7622 202884 7678 202940
rect 7678 202884 7682 202940
rect 7618 202880 7682 202884
rect 7698 202940 7762 202944
rect 7698 202884 7702 202940
rect 7702 202884 7758 202940
rect 7758 202884 7762 202940
rect 7698 202880 7762 202884
rect 7778 202940 7842 202944
rect 7778 202884 7782 202940
rect 7782 202884 7838 202940
rect 7838 202884 7842 202940
rect 7778 202880 7842 202884
rect 7858 202940 7922 202944
rect 7858 202884 7862 202940
rect 7862 202884 7918 202940
rect 7918 202884 7922 202940
rect 7858 202880 7922 202884
rect 2618 202396 2682 202400
rect 2618 202340 2622 202396
rect 2622 202340 2678 202396
rect 2678 202340 2682 202396
rect 2618 202336 2682 202340
rect 2698 202396 2762 202400
rect 2698 202340 2702 202396
rect 2702 202340 2758 202396
rect 2758 202340 2762 202396
rect 2698 202336 2762 202340
rect 2778 202396 2842 202400
rect 2778 202340 2782 202396
rect 2782 202340 2838 202396
rect 2838 202340 2842 202396
rect 2778 202336 2842 202340
rect 2858 202396 2922 202400
rect 2858 202340 2862 202396
rect 2862 202340 2918 202396
rect 2918 202340 2922 202396
rect 2858 202336 2922 202340
rect 5952 202396 6016 202400
rect 5952 202340 5956 202396
rect 5956 202340 6012 202396
rect 6012 202340 6016 202396
rect 5952 202336 6016 202340
rect 6032 202396 6096 202400
rect 6032 202340 6036 202396
rect 6036 202340 6092 202396
rect 6092 202340 6096 202396
rect 6032 202336 6096 202340
rect 6112 202396 6176 202400
rect 6112 202340 6116 202396
rect 6116 202340 6172 202396
rect 6172 202340 6176 202396
rect 6112 202336 6176 202340
rect 6192 202396 6256 202400
rect 6192 202340 6196 202396
rect 6196 202340 6252 202396
rect 6252 202340 6256 202396
rect 6192 202336 6256 202340
rect 4285 201852 4349 201856
rect 4285 201796 4289 201852
rect 4289 201796 4345 201852
rect 4345 201796 4349 201852
rect 4285 201792 4349 201796
rect 4365 201852 4429 201856
rect 4365 201796 4369 201852
rect 4369 201796 4425 201852
rect 4425 201796 4429 201852
rect 4365 201792 4429 201796
rect 4445 201852 4509 201856
rect 4445 201796 4449 201852
rect 4449 201796 4505 201852
rect 4505 201796 4509 201852
rect 4445 201792 4509 201796
rect 4525 201852 4589 201856
rect 4525 201796 4529 201852
rect 4529 201796 4585 201852
rect 4585 201796 4589 201852
rect 4525 201792 4589 201796
rect 7618 201852 7682 201856
rect 7618 201796 7622 201852
rect 7622 201796 7678 201852
rect 7678 201796 7682 201852
rect 7618 201792 7682 201796
rect 7698 201852 7762 201856
rect 7698 201796 7702 201852
rect 7702 201796 7758 201852
rect 7758 201796 7762 201852
rect 7698 201792 7762 201796
rect 7778 201852 7842 201856
rect 7778 201796 7782 201852
rect 7782 201796 7838 201852
rect 7838 201796 7842 201852
rect 7778 201792 7842 201796
rect 7858 201852 7922 201856
rect 7858 201796 7862 201852
rect 7862 201796 7918 201852
rect 7918 201796 7922 201852
rect 7858 201792 7922 201796
rect 2618 201308 2682 201312
rect 2618 201252 2622 201308
rect 2622 201252 2678 201308
rect 2678 201252 2682 201308
rect 2618 201248 2682 201252
rect 2698 201308 2762 201312
rect 2698 201252 2702 201308
rect 2702 201252 2758 201308
rect 2758 201252 2762 201308
rect 2698 201248 2762 201252
rect 2778 201308 2842 201312
rect 2778 201252 2782 201308
rect 2782 201252 2838 201308
rect 2838 201252 2842 201308
rect 2778 201248 2842 201252
rect 2858 201308 2922 201312
rect 2858 201252 2862 201308
rect 2862 201252 2918 201308
rect 2918 201252 2922 201308
rect 2858 201248 2922 201252
rect 5952 201308 6016 201312
rect 5952 201252 5956 201308
rect 5956 201252 6012 201308
rect 6012 201252 6016 201308
rect 5952 201248 6016 201252
rect 6032 201308 6096 201312
rect 6032 201252 6036 201308
rect 6036 201252 6092 201308
rect 6092 201252 6096 201308
rect 6032 201248 6096 201252
rect 6112 201308 6176 201312
rect 6112 201252 6116 201308
rect 6116 201252 6172 201308
rect 6172 201252 6176 201308
rect 6112 201248 6176 201252
rect 6192 201308 6256 201312
rect 6192 201252 6196 201308
rect 6196 201252 6252 201308
rect 6252 201252 6256 201308
rect 6192 201248 6256 201252
rect 4285 200764 4349 200768
rect 4285 200708 4289 200764
rect 4289 200708 4345 200764
rect 4345 200708 4349 200764
rect 4285 200704 4349 200708
rect 4365 200764 4429 200768
rect 4365 200708 4369 200764
rect 4369 200708 4425 200764
rect 4425 200708 4429 200764
rect 4365 200704 4429 200708
rect 4445 200764 4509 200768
rect 4445 200708 4449 200764
rect 4449 200708 4505 200764
rect 4505 200708 4509 200764
rect 4445 200704 4509 200708
rect 4525 200764 4589 200768
rect 4525 200708 4529 200764
rect 4529 200708 4585 200764
rect 4585 200708 4589 200764
rect 4525 200704 4589 200708
rect 7618 200764 7682 200768
rect 7618 200708 7622 200764
rect 7622 200708 7678 200764
rect 7678 200708 7682 200764
rect 7618 200704 7682 200708
rect 7698 200764 7762 200768
rect 7698 200708 7702 200764
rect 7702 200708 7758 200764
rect 7758 200708 7762 200764
rect 7698 200704 7762 200708
rect 7778 200764 7842 200768
rect 7778 200708 7782 200764
rect 7782 200708 7838 200764
rect 7838 200708 7842 200764
rect 7778 200704 7842 200708
rect 7858 200764 7922 200768
rect 7858 200708 7862 200764
rect 7862 200708 7918 200764
rect 7918 200708 7922 200764
rect 7858 200704 7922 200708
rect 2618 200220 2682 200224
rect 2618 200164 2622 200220
rect 2622 200164 2678 200220
rect 2678 200164 2682 200220
rect 2618 200160 2682 200164
rect 2698 200220 2762 200224
rect 2698 200164 2702 200220
rect 2702 200164 2758 200220
rect 2758 200164 2762 200220
rect 2698 200160 2762 200164
rect 2778 200220 2842 200224
rect 2778 200164 2782 200220
rect 2782 200164 2838 200220
rect 2838 200164 2842 200220
rect 2778 200160 2842 200164
rect 2858 200220 2922 200224
rect 2858 200164 2862 200220
rect 2862 200164 2918 200220
rect 2918 200164 2922 200220
rect 2858 200160 2922 200164
rect 5952 200220 6016 200224
rect 5952 200164 5956 200220
rect 5956 200164 6012 200220
rect 6012 200164 6016 200220
rect 5952 200160 6016 200164
rect 6032 200220 6096 200224
rect 6032 200164 6036 200220
rect 6036 200164 6092 200220
rect 6092 200164 6096 200220
rect 6032 200160 6096 200164
rect 6112 200220 6176 200224
rect 6112 200164 6116 200220
rect 6116 200164 6172 200220
rect 6172 200164 6176 200220
rect 6112 200160 6176 200164
rect 6192 200220 6256 200224
rect 6192 200164 6196 200220
rect 6196 200164 6252 200220
rect 6252 200164 6256 200220
rect 6192 200160 6256 200164
rect 4285 199676 4349 199680
rect 4285 199620 4289 199676
rect 4289 199620 4345 199676
rect 4345 199620 4349 199676
rect 4285 199616 4349 199620
rect 4365 199676 4429 199680
rect 4365 199620 4369 199676
rect 4369 199620 4425 199676
rect 4425 199620 4429 199676
rect 4365 199616 4429 199620
rect 4445 199676 4509 199680
rect 4445 199620 4449 199676
rect 4449 199620 4505 199676
rect 4505 199620 4509 199676
rect 4445 199616 4509 199620
rect 4525 199676 4589 199680
rect 4525 199620 4529 199676
rect 4529 199620 4585 199676
rect 4585 199620 4589 199676
rect 4525 199616 4589 199620
rect 7618 199676 7682 199680
rect 7618 199620 7622 199676
rect 7622 199620 7678 199676
rect 7678 199620 7682 199676
rect 7618 199616 7682 199620
rect 7698 199676 7762 199680
rect 7698 199620 7702 199676
rect 7702 199620 7758 199676
rect 7758 199620 7762 199676
rect 7698 199616 7762 199620
rect 7778 199676 7842 199680
rect 7778 199620 7782 199676
rect 7782 199620 7838 199676
rect 7838 199620 7842 199676
rect 7778 199616 7842 199620
rect 7858 199676 7922 199680
rect 7858 199620 7862 199676
rect 7862 199620 7918 199676
rect 7918 199620 7922 199676
rect 7858 199616 7922 199620
rect 2618 199132 2682 199136
rect 2618 199076 2622 199132
rect 2622 199076 2678 199132
rect 2678 199076 2682 199132
rect 2618 199072 2682 199076
rect 2698 199132 2762 199136
rect 2698 199076 2702 199132
rect 2702 199076 2758 199132
rect 2758 199076 2762 199132
rect 2698 199072 2762 199076
rect 2778 199132 2842 199136
rect 2778 199076 2782 199132
rect 2782 199076 2838 199132
rect 2838 199076 2842 199132
rect 2778 199072 2842 199076
rect 2858 199132 2922 199136
rect 2858 199076 2862 199132
rect 2862 199076 2918 199132
rect 2918 199076 2922 199132
rect 2858 199072 2922 199076
rect 5952 199132 6016 199136
rect 5952 199076 5956 199132
rect 5956 199076 6012 199132
rect 6012 199076 6016 199132
rect 5952 199072 6016 199076
rect 6032 199132 6096 199136
rect 6032 199076 6036 199132
rect 6036 199076 6092 199132
rect 6092 199076 6096 199132
rect 6032 199072 6096 199076
rect 6112 199132 6176 199136
rect 6112 199076 6116 199132
rect 6116 199076 6172 199132
rect 6172 199076 6176 199132
rect 6112 199072 6176 199076
rect 6192 199132 6256 199136
rect 6192 199076 6196 199132
rect 6196 199076 6252 199132
rect 6252 199076 6256 199132
rect 6192 199072 6256 199076
rect 4285 198588 4349 198592
rect 4285 198532 4289 198588
rect 4289 198532 4345 198588
rect 4345 198532 4349 198588
rect 4285 198528 4349 198532
rect 4365 198588 4429 198592
rect 4365 198532 4369 198588
rect 4369 198532 4425 198588
rect 4425 198532 4429 198588
rect 4365 198528 4429 198532
rect 4445 198588 4509 198592
rect 4445 198532 4449 198588
rect 4449 198532 4505 198588
rect 4505 198532 4509 198588
rect 4445 198528 4509 198532
rect 4525 198588 4589 198592
rect 4525 198532 4529 198588
rect 4529 198532 4585 198588
rect 4585 198532 4589 198588
rect 4525 198528 4589 198532
rect 7618 198588 7682 198592
rect 7618 198532 7622 198588
rect 7622 198532 7678 198588
rect 7678 198532 7682 198588
rect 7618 198528 7682 198532
rect 7698 198588 7762 198592
rect 7698 198532 7702 198588
rect 7702 198532 7758 198588
rect 7758 198532 7762 198588
rect 7698 198528 7762 198532
rect 7778 198588 7842 198592
rect 7778 198532 7782 198588
rect 7782 198532 7838 198588
rect 7838 198532 7842 198588
rect 7778 198528 7842 198532
rect 7858 198588 7922 198592
rect 7858 198532 7862 198588
rect 7862 198532 7918 198588
rect 7918 198532 7922 198588
rect 7858 198528 7922 198532
rect 2618 198044 2682 198048
rect 2618 197988 2622 198044
rect 2622 197988 2678 198044
rect 2678 197988 2682 198044
rect 2618 197984 2682 197988
rect 2698 198044 2762 198048
rect 2698 197988 2702 198044
rect 2702 197988 2758 198044
rect 2758 197988 2762 198044
rect 2698 197984 2762 197988
rect 2778 198044 2842 198048
rect 2778 197988 2782 198044
rect 2782 197988 2838 198044
rect 2838 197988 2842 198044
rect 2778 197984 2842 197988
rect 2858 198044 2922 198048
rect 2858 197988 2862 198044
rect 2862 197988 2918 198044
rect 2918 197988 2922 198044
rect 2858 197984 2922 197988
rect 5952 198044 6016 198048
rect 5952 197988 5956 198044
rect 5956 197988 6012 198044
rect 6012 197988 6016 198044
rect 5952 197984 6016 197988
rect 6032 198044 6096 198048
rect 6032 197988 6036 198044
rect 6036 197988 6092 198044
rect 6092 197988 6096 198044
rect 6032 197984 6096 197988
rect 6112 198044 6176 198048
rect 6112 197988 6116 198044
rect 6116 197988 6172 198044
rect 6172 197988 6176 198044
rect 6112 197984 6176 197988
rect 6192 198044 6256 198048
rect 6192 197988 6196 198044
rect 6196 197988 6252 198044
rect 6252 197988 6256 198044
rect 6192 197984 6256 197988
rect 4285 197500 4349 197504
rect 4285 197444 4289 197500
rect 4289 197444 4345 197500
rect 4345 197444 4349 197500
rect 4285 197440 4349 197444
rect 4365 197500 4429 197504
rect 4365 197444 4369 197500
rect 4369 197444 4425 197500
rect 4425 197444 4429 197500
rect 4365 197440 4429 197444
rect 4445 197500 4509 197504
rect 4445 197444 4449 197500
rect 4449 197444 4505 197500
rect 4505 197444 4509 197500
rect 4445 197440 4509 197444
rect 4525 197500 4589 197504
rect 4525 197444 4529 197500
rect 4529 197444 4585 197500
rect 4585 197444 4589 197500
rect 4525 197440 4589 197444
rect 7618 197500 7682 197504
rect 7618 197444 7622 197500
rect 7622 197444 7678 197500
rect 7678 197444 7682 197500
rect 7618 197440 7682 197444
rect 7698 197500 7762 197504
rect 7698 197444 7702 197500
rect 7702 197444 7758 197500
rect 7758 197444 7762 197500
rect 7698 197440 7762 197444
rect 7778 197500 7842 197504
rect 7778 197444 7782 197500
rect 7782 197444 7838 197500
rect 7838 197444 7842 197500
rect 7778 197440 7842 197444
rect 7858 197500 7922 197504
rect 7858 197444 7862 197500
rect 7862 197444 7918 197500
rect 7918 197444 7922 197500
rect 7858 197440 7922 197444
rect 2618 196956 2682 196960
rect 2618 196900 2622 196956
rect 2622 196900 2678 196956
rect 2678 196900 2682 196956
rect 2618 196896 2682 196900
rect 2698 196956 2762 196960
rect 2698 196900 2702 196956
rect 2702 196900 2758 196956
rect 2758 196900 2762 196956
rect 2698 196896 2762 196900
rect 2778 196956 2842 196960
rect 2778 196900 2782 196956
rect 2782 196900 2838 196956
rect 2838 196900 2842 196956
rect 2778 196896 2842 196900
rect 2858 196956 2922 196960
rect 2858 196900 2862 196956
rect 2862 196900 2918 196956
rect 2918 196900 2922 196956
rect 2858 196896 2922 196900
rect 5952 196956 6016 196960
rect 5952 196900 5956 196956
rect 5956 196900 6012 196956
rect 6012 196900 6016 196956
rect 5952 196896 6016 196900
rect 6032 196956 6096 196960
rect 6032 196900 6036 196956
rect 6036 196900 6092 196956
rect 6092 196900 6096 196956
rect 6032 196896 6096 196900
rect 6112 196956 6176 196960
rect 6112 196900 6116 196956
rect 6116 196900 6172 196956
rect 6172 196900 6176 196956
rect 6112 196896 6176 196900
rect 6192 196956 6256 196960
rect 6192 196900 6196 196956
rect 6196 196900 6252 196956
rect 6252 196900 6256 196956
rect 6192 196896 6256 196900
rect 4285 196412 4349 196416
rect 4285 196356 4289 196412
rect 4289 196356 4345 196412
rect 4345 196356 4349 196412
rect 4285 196352 4349 196356
rect 4365 196412 4429 196416
rect 4365 196356 4369 196412
rect 4369 196356 4425 196412
rect 4425 196356 4429 196412
rect 4365 196352 4429 196356
rect 4445 196412 4509 196416
rect 4445 196356 4449 196412
rect 4449 196356 4505 196412
rect 4505 196356 4509 196412
rect 4445 196352 4509 196356
rect 4525 196412 4589 196416
rect 4525 196356 4529 196412
rect 4529 196356 4585 196412
rect 4585 196356 4589 196412
rect 4525 196352 4589 196356
rect 7618 196412 7682 196416
rect 7618 196356 7622 196412
rect 7622 196356 7678 196412
rect 7678 196356 7682 196412
rect 7618 196352 7682 196356
rect 7698 196412 7762 196416
rect 7698 196356 7702 196412
rect 7702 196356 7758 196412
rect 7758 196356 7762 196412
rect 7698 196352 7762 196356
rect 7778 196412 7842 196416
rect 7778 196356 7782 196412
rect 7782 196356 7838 196412
rect 7838 196356 7842 196412
rect 7778 196352 7842 196356
rect 7858 196412 7922 196416
rect 7858 196356 7862 196412
rect 7862 196356 7918 196412
rect 7918 196356 7922 196412
rect 7858 196352 7922 196356
rect 2618 195868 2682 195872
rect 2618 195812 2622 195868
rect 2622 195812 2678 195868
rect 2678 195812 2682 195868
rect 2618 195808 2682 195812
rect 2698 195868 2762 195872
rect 2698 195812 2702 195868
rect 2702 195812 2758 195868
rect 2758 195812 2762 195868
rect 2698 195808 2762 195812
rect 2778 195868 2842 195872
rect 2778 195812 2782 195868
rect 2782 195812 2838 195868
rect 2838 195812 2842 195868
rect 2778 195808 2842 195812
rect 2858 195868 2922 195872
rect 2858 195812 2862 195868
rect 2862 195812 2918 195868
rect 2918 195812 2922 195868
rect 2858 195808 2922 195812
rect 5952 195868 6016 195872
rect 5952 195812 5956 195868
rect 5956 195812 6012 195868
rect 6012 195812 6016 195868
rect 5952 195808 6016 195812
rect 6032 195868 6096 195872
rect 6032 195812 6036 195868
rect 6036 195812 6092 195868
rect 6092 195812 6096 195868
rect 6032 195808 6096 195812
rect 6112 195868 6176 195872
rect 6112 195812 6116 195868
rect 6116 195812 6172 195868
rect 6172 195812 6176 195868
rect 6112 195808 6176 195812
rect 6192 195868 6256 195872
rect 6192 195812 6196 195868
rect 6196 195812 6252 195868
rect 6252 195812 6256 195868
rect 6192 195808 6256 195812
rect 4285 195324 4349 195328
rect 4285 195268 4289 195324
rect 4289 195268 4345 195324
rect 4345 195268 4349 195324
rect 4285 195264 4349 195268
rect 4365 195324 4429 195328
rect 4365 195268 4369 195324
rect 4369 195268 4425 195324
rect 4425 195268 4429 195324
rect 4365 195264 4429 195268
rect 4445 195324 4509 195328
rect 4445 195268 4449 195324
rect 4449 195268 4505 195324
rect 4505 195268 4509 195324
rect 4445 195264 4509 195268
rect 4525 195324 4589 195328
rect 4525 195268 4529 195324
rect 4529 195268 4585 195324
rect 4585 195268 4589 195324
rect 4525 195264 4589 195268
rect 7618 195324 7682 195328
rect 7618 195268 7622 195324
rect 7622 195268 7678 195324
rect 7678 195268 7682 195324
rect 7618 195264 7682 195268
rect 7698 195324 7762 195328
rect 7698 195268 7702 195324
rect 7702 195268 7758 195324
rect 7758 195268 7762 195324
rect 7698 195264 7762 195268
rect 7778 195324 7842 195328
rect 7778 195268 7782 195324
rect 7782 195268 7838 195324
rect 7838 195268 7842 195324
rect 7778 195264 7842 195268
rect 7858 195324 7922 195328
rect 7858 195268 7862 195324
rect 7862 195268 7918 195324
rect 7918 195268 7922 195324
rect 7858 195264 7922 195268
rect 2618 194780 2682 194784
rect 2618 194724 2622 194780
rect 2622 194724 2678 194780
rect 2678 194724 2682 194780
rect 2618 194720 2682 194724
rect 2698 194780 2762 194784
rect 2698 194724 2702 194780
rect 2702 194724 2758 194780
rect 2758 194724 2762 194780
rect 2698 194720 2762 194724
rect 2778 194780 2842 194784
rect 2778 194724 2782 194780
rect 2782 194724 2838 194780
rect 2838 194724 2842 194780
rect 2778 194720 2842 194724
rect 2858 194780 2922 194784
rect 2858 194724 2862 194780
rect 2862 194724 2918 194780
rect 2918 194724 2922 194780
rect 2858 194720 2922 194724
rect 5952 194780 6016 194784
rect 5952 194724 5956 194780
rect 5956 194724 6012 194780
rect 6012 194724 6016 194780
rect 5952 194720 6016 194724
rect 6032 194780 6096 194784
rect 6032 194724 6036 194780
rect 6036 194724 6092 194780
rect 6092 194724 6096 194780
rect 6032 194720 6096 194724
rect 6112 194780 6176 194784
rect 6112 194724 6116 194780
rect 6116 194724 6172 194780
rect 6172 194724 6176 194780
rect 6112 194720 6176 194724
rect 6192 194780 6256 194784
rect 6192 194724 6196 194780
rect 6196 194724 6252 194780
rect 6252 194724 6256 194780
rect 6192 194720 6256 194724
rect 4285 194236 4349 194240
rect 4285 194180 4289 194236
rect 4289 194180 4345 194236
rect 4345 194180 4349 194236
rect 4285 194176 4349 194180
rect 4365 194236 4429 194240
rect 4365 194180 4369 194236
rect 4369 194180 4425 194236
rect 4425 194180 4429 194236
rect 4365 194176 4429 194180
rect 4445 194236 4509 194240
rect 4445 194180 4449 194236
rect 4449 194180 4505 194236
rect 4505 194180 4509 194236
rect 4445 194176 4509 194180
rect 4525 194236 4589 194240
rect 4525 194180 4529 194236
rect 4529 194180 4585 194236
rect 4585 194180 4589 194236
rect 4525 194176 4589 194180
rect 7618 194236 7682 194240
rect 7618 194180 7622 194236
rect 7622 194180 7678 194236
rect 7678 194180 7682 194236
rect 7618 194176 7682 194180
rect 7698 194236 7762 194240
rect 7698 194180 7702 194236
rect 7702 194180 7758 194236
rect 7758 194180 7762 194236
rect 7698 194176 7762 194180
rect 7778 194236 7842 194240
rect 7778 194180 7782 194236
rect 7782 194180 7838 194236
rect 7838 194180 7842 194236
rect 7778 194176 7842 194180
rect 7858 194236 7922 194240
rect 7858 194180 7862 194236
rect 7862 194180 7918 194236
rect 7918 194180 7922 194236
rect 7858 194176 7922 194180
rect 2618 193692 2682 193696
rect 2618 193636 2622 193692
rect 2622 193636 2678 193692
rect 2678 193636 2682 193692
rect 2618 193632 2682 193636
rect 2698 193692 2762 193696
rect 2698 193636 2702 193692
rect 2702 193636 2758 193692
rect 2758 193636 2762 193692
rect 2698 193632 2762 193636
rect 2778 193692 2842 193696
rect 2778 193636 2782 193692
rect 2782 193636 2838 193692
rect 2838 193636 2842 193692
rect 2778 193632 2842 193636
rect 2858 193692 2922 193696
rect 2858 193636 2862 193692
rect 2862 193636 2918 193692
rect 2918 193636 2922 193692
rect 2858 193632 2922 193636
rect 5952 193692 6016 193696
rect 5952 193636 5956 193692
rect 5956 193636 6012 193692
rect 6012 193636 6016 193692
rect 5952 193632 6016 193636
rect 6032 193692 6096 193696
rect 6032 193636 6036 193692
rect 6036 193636 6092 193692
rect 6092 193636 6096 193692
rect 6032 193632 6096 193636
rect 6112 193692 6176 193696
rect 6112 193636 6116 193692
rect 6116 193636 6172 193692
rect 6172 193636 6176 193692
rect 6112 193632 6176 193636
rect 6192 193692 6256 193696
rect 6192 193636 6196 193692
rect 6196 193636 6252 193692
rect 6252 193636 6256 193692
rect 6192 193632 6256 193636
rect 4285 193148 4349 193152
rect 4285 193092 4289 193148
rect 4289 193092 4345 193148
rect 4345 193092 4349 193148
rect 4285 193088 4349 193092
rect 4365 193148 4429 193152
rect 4365 193092 4369 193148
rect 4369 193092 4425 193148
rect 4425 193092 4429 193148
rect 4365 193088 4429 193092
rect 4445 193148 4509 193152
rect 4445 193092 4449 193148
rect 4449 193092 4505 193148
rect 4505 193092 4509 193148
rect 4445 193088 4509 193092
rect 4525 193148 4589 193152
rect 4525 193092 4529 193148
rect 4529 193092 4585 193148
rect 4585 193092 4589 193148
rect 4525 193088 4589 193092
rect 7618 193148 7682 193152
rect 7618 193092 7622 193148
rect 7622 193092 7678 193148
rect 7678 193092 7682 193148
rect 7618 193088 7682 193092
rect 7698 193148 7762 193152
rect 7698 193092 7702 193148
rect 7702 193092 7758 193148
rect 7758 193092 7762 193148
rect 7698 193088 7762 193092
rect 7778 193148 7842 193152
rect 7778 193092 7782 193148
rect 7782 193092 7838 193148
rect 7838 193092 7842 193148
rect 7778 193088 7842 193092
rect 7858 193148 7922 193152
rect 7858 193092 7862 193148
rect 7862 193092 7918 193148
rect 7918 193092 7922 193148
rect 7858 193088 7922 193092
rect 2618 192604 2682 192608
rect 2618 192548 2622 192604
rect 2622 192548 2678 192604
rect 2678 192548 2682 192604
rect 2618 192544 2682 192548
rect 2698 192604 2762 192608
rect 2698 192548 2702 192604
rect 2702 192548 2758 192604
rect 2758 192548 2762 192604
rect 2698 192544 2762 192548
rect 2778 192604 2842 192608
rect 2778 192548 2782 192604
rect 2782 192548 2838 192604
rect 2838 192548 2842 192604
rect 2778 192544 2842 192548
rect 2858 192604 2922 192608
rect 2858 192548 2862 192604
rect 2862 192548 2918 192604
rect 2918 192548 2922 192604
rect 2858 192544 2922 192548
rect 5952 192604 6016 192608
rect 5952 192548 5956 192604
rect 5956 192548 6012 192604
rect 6012 192548 6016 192604
rect 5952 192544 6016 192548
rect 6032 192604 6096 192608
rect 6032 192548 6036 192604
rect 6036 192548 6092 192604
rect 6092 192548 6096 192604
rect 6032 192544 6096 192548
rect 6112 192604 6176 192608
rect 6112 192548 6116 192604
rect 6116 192548 6172 192604
rect 6172 192548 6176 192604
rect 6112 192544 6176 192548
rect 6192 192604 6256 192608
rect 6192 192548 6196 192604
rect 6196 192548 6252 192604
rect 6252 192548 6256 192604
rect 6192 192544 6256 192548
rect 4285 192060 4349 192064
rect 4285 192004 4289 192060
rect 4289 192004 4345 192060
rect 4345 192004 4349 192060
rect 4285 192000 4349 192004
rect 4365 192060 4429 192064
rect 4365 192004 4369 192060
rect 4369 192004 4425 192060
rect 4425 192004 4429 192060
rect 4365 192000 4429 192004
rect 4445 192060 4509 192064
rect 4445 192004 4449 192060
rect 4449 192004 4505 192060
rect 4505 192004 4509 192060
rect 4445 192000 4509 192004
rect 4525 192060 4589 192064
rect 4525 192004 4529 192060
rect 4529 192004 4585 192060
rect 4585 192004 4589 192060
rect 4525 192000 4589 192004
rect 7618 192060 7682 192064
rect 7618 192004 7622 192060
rect 7622 192004 7678 192060
rect 7678 192004 7682 192060
rect 7618 192000 7682 192004
rect 7698 192060 7762 192064
rect 7698 192004 7702 192060
rect 7702 192004 7758 192060
rect 7758 192004 7762 192060
rect 7698 192000 7762 192004
rect 7778 192060 7842 192064
rect 7778 192004 7782 192060
rect 7782 192004 7838 192060
rect 7838 192004 7842 192060
rect 7778 192000 7842 192004
rect 7858 192060 7922 192064
rect 7858 192004 7862 192060
rect 7862 192004 7918 192060
rect 7918 192004 7922 192060
rect 7858 192000 7922 192004
rect 2618 191516 2682 191520
rect 2618 191460 2622 191516
rect 2622 191460 2678 191516
rect 2678 191460 2682 191516
rect 2618 191456 2682 191460
rect 2698 191516 2762 191520
rect 2698 191460 2702 191516
rect 2702 191460 2758 191516
rect 2758 191460 2762 191516
rect 2698 191456 2762 191460
rect 2778 191516 2842 191520
rect 2778 191460 2782 191516
rect 2782 191460 2838 191516
rect 2838 191460 2842 191516
rect 2778 191456 2842 191460
rect 2858 191516 2922 191520
rect 2858 191460 2862 191516
rect 2862 191460 2918 191516
rect 2918 191460 2922 191516
rect 2858 191456 2922 191460
rect 5952 191516 6016 191520
rect 5952 191460 5956 191516
rect 5956 191460 6012 191516
rect 6012 191460 6016 191516
rect 5952 191456 6016 191460
rect 6032 191516 6096 191520
rect 6032 191460 6036 191516
rect 6036 191460 6092 191516
rect 6092 191460 6096 191516
rect 6032 191456 6096 191460
rect 6112 191516 6176 191520
rect 6112 191460 6116 191516
rect 6116 191460 6172 191516
rect 6172 191460 6176 191516
rect 6112 191456 6176 191460
rect 6192 191516 6256 191520
rect 6192 191460 6196 191516
rect 6196 191460 6252 191516
rect 6252 191460 6256 191516
rect 6192 191456 6256 191460
rect 4285 190972 4349 190976
rect 4285 190916 4289 190972
rect 4289 190916 4345 190972
rect 4345 190916 4349 190972
rect 4285 190912 4349 190916
rect 4365 190972 4429 190976
rect 4365 190916 4369 190972
rect 4369 190916 4425 190972
rect 4425 190916 4429 190972
rect 4365 190912 4429 190916
rect 4445 190972 4509 190976
rect 4445 190916 4449 190972
rect 4449 190916 4505 190972
rect 4505 190916 4509 190972
rect 4445 190912 4509 190916
rect 4525 190972 4589 190976
rect 4525 190916 4529 190972
rect 4529 190916 4585 190972
rect 4585 190916 4589 190972
rect 4525 190912 4589 190916
rect 7618 190972 7682 190976
rect 7618 190916 7622 190972
rect 7622 190916 7678 190972
rect 7678 190916 7682 190972
rect 7618 190912 7682 190916
rect 7698 190972 7762 190976
rect 7698 190916 7702 190972
rect 7702 190916 7758 190972
rect 7758 190916 7762 190972
rect 7698 190912 7762 190916
rect 7778 190972 7842 190976
rect 7778 190916 7782 190972
rect 7782 190916 7838 190972
rect 7838 190916 7842 190972
rect 7778 190912 7842 190916
rect 7858 190972 7922 190976
rect 7858 190916 7862 190972
rect 7862 190916 7918 190972
rect 7918 190916 7922 190972
rect 7858 190912 7922 190916
rect 2618 190428 2682 190432
rect 2618 190372 2622 190428
rect 2622 190372 2678 190428
rect 2678 190372 2682 190428
rect 2618 190368 2682 190372
rect 2698 190428 2762 190432
rect 2698 190372 2702 190428
rect 2702 190372 2758 190428
rect 2758 190372 2762 190428
rect 2698 190368 2762 190372
rect 2778 190428 2842 190432
rect 2778 190372 2782 190428
rect 2782 190372 2838 190428
rect 2838 190372 2842 190428
rect 2778 190368 2842 190372
rect 2858 190428 2922 190432
rect 2858 190372 2862 190428
rect 2862 190372 2918 190428
rect 2918 190372 2922 190428
rect 2858 190368 2922 190372
rect 5952 190428 6016 190432
rect 5952 190372 5956 190428
rect 5956 190372 6012 190428
rect 6012 190372 6016 190428
rect 5952 190368 6016 190372
rect 6032 190428 6096 190432
rect 6032 190372 6036 190428
rect 6036 190372 6092 190428
rect 6092 190372 6096 190428
rect 6032 190368 6096 190372
rect 6112 190428 6176 190432
rect 6112 190372 6116 190428
rect 6116 190372 6172 190428
rect 6172 190372 6176 190428
rect 6112 190368 6176 190372
rect 6192 190428 6256 190432
rect 6192 190372 6196 190428
rect 6196 190372 6252 190428
rect 6252 190372 6256 190428
rect 6192 190368 6256 190372
rect 4285 189884 4349 189888
rect 4285 189828 4289 189884
rect 4289 189828 4345 189884
rect 4345 189828 4349 189884
rect 4285 189824 4349 189828
rect 4365 189884 4429 189888
rect 4365 189828 4369 189884
rect 4369 189828 4425 189884
rect 4425 189828 4429 189884
rect 4365 189824 4429 189828
rect 4445 189884 4509 189888
rect 4445 189828 4449 189884
rect 4449 189828 4505 189884
rect 4505 189828 4509 189884
rect 4445 189824 4509 189828
rect 4525 189884 4589 189888
rect 4525 189828 4529 189884
rect 4529 189828 4585 189884
rect 4585 189828 4589 189884
rect 4525 189824 4589 189828
rect 7618 189884 7682 189888
rect 7618 189828 7622 189884
rect 7622 189828 7678 189884
rect 7678 189828 7682 189884
rect 7618 189824 7682 189828
rect 7698 189884 7762 189888
rect 7698 189828 7702 189884
rect 7702 189828 7758 189884
rect 7758 189828 7762 189884
rect 7698 189824 7762 189828
rect 7778 189884 7842 189888
rect 7778 189828 7782 189884
rect 7782 189828 7838 189884
rect 7838 189828 7842 189884
rect 7778 189824 7842 189828
rect 7858 189884 7922 189888
rect 7858 189828 7862 189884
rect 7862 189828 7918 189884
rect 7918 189828 7922 189884
rect 7858 189824 7922 189828
rect 2618 189340 2682 189344
rect 2618 189284 2622 189340
rect 2622 189284 2678 189340
rect 2678 189284 2682 189340
rect 2618 189280 2682 189284
rect 2698 189340 2762 189344
rect 2698 189284 2702 189340
rect 2702 189284 2758 189340
rect 2758 189284 2762 189340
rect 2698 189280 2762 189284
rect 2778 189340 2842 189344
rect 2778 189284 2782 189340
rect 2782 189284 2838 189340
rect 2838 189284 2842 189340
rect 2778 189280 2842 189284
rect 2858 189340 2922 189344
rect 2858 189284 2862 189340
rect 2862 189284 2918 189340
rect 2918 189284 2922 189340
rect 2858 189280 2922 189284
rect 5952 189340 6016 189344
rect 5952 189284 5956 189340
rect 5956 189284 6012 189340
rect 6012 189284 6016 189340
rect 5952 189280 6016 189284
rect 6032 189340 6096 189344
rect 6032 189284 6036 189340
rect 6036 189284 6092 189340
rect 6092 189284 6096 189340
rect 6032 189280 6096 189284
rect 6112 189340 6176 189344
rect 6112 189284 6116 189340
rect 6116 189284 6172 189340
rect 6172 189284 6176 189340
rect 6112 189280 6176 189284
rect 6192 189340 6256 189344
rect 6192 189284 6196 189340
rect 6196 189284 6252 189340
rect 6252 189284 6256 189340
rect 6192 189280 6256 189284
rect 4285 188796 4349 188800
rect 4285 188740 4289 188796
rect 4289 188740 4345 188796
rect 4345 188740 4349 188796
rect 4285 188736 4349 188740
rect 4365 188796 4429 188800
rect 4365 188740 4369 188796
rect 4369 188740 4425 188796
rect 4425 188740 4429 188796
rect 4365 188736 4429 188740
rect 4445 188796 4509 188800
rect 4445 188740 4449 188796
rect 4449 188740 4505 188796
rect 4505 188740 4509 188796
rect 4445 188736 4509 188740
rect 4525 188796 4589 188800
rect 4525 188740 4529 188796
rect 4529 188740 4585 188796
rect 4585 188740 4589 188796
rect 4525 188736 4589 188740
rect 7618 188796 7682 188800
rect 7618 188740 7622 188796
rect 7622 188740 7678 188796
rect 7678 188740 7682 188796
rect 7618 188736 7682 188740
rect 7698 188796 7762 188800
rect 7698 188740 7702 188796
rect 7702 188740 7758 188796
rect 7758 188740 7762 188796
rect 7698 188736 7762 188740
rect 7778 188796 7842 188800
rect 7778 188740 7782 188796
rect 7782 188740 7838 188796
rect 7838 188740 7842 188796
rect 7778 188736 7842 188740
rect 7858 188796 7922 188800
rect 7858 188740 7862 188796
rect 7862 188740 7918 188796
rect 7918 188740 7922 188796
rect 7858 188736 7922 188740
rect 2618 188252 2682 188256
rect 2618 188196 2622 188252
rect 2622 188196 2678 188252
rect 2678 188196 2682 188252
rect 2618 188192 2682 188196
rect 2698 188252 2762 188256
rect 2698 188196 2702 188252
rect 2702 188196 2758 188252
rect 2758 188196 2762 188252
rect 2698 188192 2762 188196
rect 2778 188252 2842 188256
rect 2778 188196 2782 188252
rect 2782 188196 2838 188252
rect 2838 188196 2842 188252
rect 2778 188192 2842 188196
rect 2858 188252 2922 188256
rect 2858 188196 2862 188252
rect 2862 188196 2918 188252
rect 2918 188196 2922 188252
rect 2858 188192 2922 188196
rect 5952 188252 6016 188256
rect 5952 188196 5956 188252
rect 5956 188196 6012 188252
rect 6012 188196 6016 188252
rect 5952 188192 6016 188196
rect 6032 188252 6096 188256
rect 6032 188196 6036 188252
rect 6036 188196 6092 188252
rect 6092 188196 6096 188252
rect 6032 188192 6096 188196
rect 6112 188252 6176 188256
rect 6112 188196 6116 188252
rect 6116 188196 6172 188252
rect 6172 188196 6176 188252
rect 6112 188192 6176 188196
rect 6192 188252 6256 188256
rect 6192 188196 6196 188252
rect 6196 188196 6252 188252
rect 6252 188196 6256 188252
rect 6192 188192 6256 188196
rect 4285 187708 4349 187712
rect 4285 187652 4289 187708
rect 4289 187652 4345 187708
rect 4345 187652 4349 187708
rect 4285 187648 4349 187652
rect 4365 187708 4429 187712
rect 4365 187652 4369 187708
rect 4369 187652 4425 187708
rect 4425 187652 4429 187708
rect 4365 187648 4429 187652
rect 4445 187708 4509 187712
rect 4445 187652 4449 187708
rect 4449 187652 4505 187708
rect 4505 187652 4509 187708
rect 4445 187648 4509 187652
rect 4525 187708 4589 187712
rect 4525 187652 4529 187708
rect 4529 187652 4585 187708
rect 4585 187652 4589 187708
rect 4525 187648 4589 187652
rect 7618 187708 7682 187712
rect 7618 187652 7622 187708
rect 7622 187652 7678 187708
rect 7678 187652 7682 187708
rect 7618 187648 7682 187652
rect 7698 187708 7762 187712
rect 7698 187652 7702 187708
rect 7702 187652 7758 187708
rect 7758 187652 7762 187708
rect 7698 187648 7762 187652
rect 7778 187708 7842 187712
rect 7778 187652 7782 187708
rect 7782 187652 7838 187708
rect 7838 187652 7842 187708
rect 7778 187648 7842 187652
rect 7858 187708 7922 187712
rect 7858 187652 7862 187708
rect 7862 187652 7918 187708
rect 7918 187652 7922 187708
rect 7858 187648 7922 187652
rect 2618 187164 2682 187168
rect 2618 187108 2622 187164
rect 2622 187108 2678 187164
rect 2678 187108 2682 187164
rect 2618 187104 2682 187108
rect 2698 187164 2762 187168
rect 2698 187108 2702 187164
rect 2702 187108 2758 187164
rect 2758 187108 2762 187164
rect 2698 187104 2762 187108
rect 2778 187164 2842 187168
rect 2778 187108 2782 187164
rect 2782 187108 2838 187164
rect 2838 187108 2842 187164
rect 2778 187104 2842 187108
rect 2858 187164 2922 187168
rect 2858 187108 2862 187164
rect 2862 187108 2918 187164
rect 2918 187108 2922 187164
rect 2858 187104 2922 187108
rect 5952 187164 6016 187168
rect 5952 187108 5956 187164
rect 5956 187108 6012 187164
rect 6012 187108 6016 187164
rect 5952 187104 6016 187108
rect 6032 187164 6096 187168
rect 6032 187108 6036 187164
rect 6036 187108 6092 187164
rect 6092 187108 6096 187164
rect 6032 187104 6096 187108
rect 6112 187164 6176 187168
rect 6112 187108 6116 187164
rect 6116 187108 6172 187164
rect 6172 187108 6176 187164
rect 6112 187104 6176 187108
rect 6192 187164 6256 187168
rect 6192 187108 6196 187164
rect 6196 187108 6252 187164
rect 6252 187108 6256 187164
rect 6192 187104 6256 187108
rect 4285 186620 4349 186624
rect 4285 186564 4289 186620
rect 4289 186564 4345 186620
rect 4345 186564 4349 186620
rect 4285 186560 4349 186564
rect 4365 186620 4429 186624
rect 4365 186564 4369 186620
rect 4369 186564 4425 186620
rect 4425 186564 4429 186620
rect 4365 186560 4429 186564
rect 4445 186620 4509 186624
rect 4445 186564 4449 186620
rect 4449 186564 4505 186620
rect 4505 186564 4509 186620
rect 4445 186560 4509 186564
rect 4525 186620 4589 186624
rect 4525 186564 4529 186620
rect 4529 186564 4585 186620
rect 4585 186564 4589 186620
rect 4525 186560 4589 186564
rect 7618 186620 7682 186624
rect 7618 186564 7622 186620
rect 7622 186564 7678 186620
rect 7678 186564 7682 186620
rect 7618 186560 7682 186564
rect 7698 186620 7762 186624
rect 7698 186564 7702 186620
rect 7702 186564 7758 186620
rect 7758 186564 7762 186620
rect 7698 186560 7762 186564
rect 7778 186620 7842 186624
rect 7778 186564 7782 186620
rect 7782 186564 7838 186620
rect 7838 186564 7842 186620
rect 7778 186560 7842 186564
rect 7858 186620 7922 186624
rect 7858 186564 7862 186620
rect 7862 186564 7918 186620
rect 7918 186564 7922 186620
rect 7858 186560 7922 186564
rect 2618 186076 2682 186080
rect 2618 186020 2622 186076
rect 2622 186020 2678 186076
rect 2678 186020 2682 186076
rect 2618 186016 2682 186020
rect 2698 186076 2762 186080
rect 2698 186020 2702 186076
rect 2702 186020 2758 186076
rect 2758 186020 2762 186076
rect 2698 186016 2762 186020
rect 2778 186076 2842 186080
rect 2778 186020 2782 186076
rect 2782 186020 2838 186076
rect 2838 186020 2842 186076
rect 2778 186016 2842 186020
rect 2858 186076 2922 186080
rect 2858 186020 2862 186076
rect 2862 186020 2918 186076
rect 2918 186020 2922 186076
rect 2858 186016 2922 186020
rect 5952 186076 6016 186080
rect 5952 186020 5956 186076
rect 5956 186020 6012 186076
rect 6012 186020 6016 186076
rect 5952 186016 6016 186020
rect 6032 186076 6096 186080
rect 6032 186020 6036 186076
rect 6036 186020 6092 186076
rect 6092 186020 6096 186076
rect 6032 186016 6096 186020
rect 6112 186076 6176 186080
rect 6112 186020 6116 186076
rect 6116 186020 6172 186076
rect 6172 186020 6176 186076
rect 6112 186016 6176 186020
rect 6192 186076 6256 186080
rect 6192 186020 6196 186076
rect 6196 186020 6252 186076
rect 6252 186020 6256 186076
rect 6192 186016 6256 186020
rect 4285 185532 4349 185536
rect 4285 185476 4289 185532
rect 4289 185476 4345 185532
rect 4345 185476 4349 185532
rect 4285 185472 4349 185476
rect 4365 185532 4429 185536
rect 4365 185476 4369 185532
rect 4369 185476 4425 185532
rect 4425 185476 4429 185532
rect 4365 185472 4429 185476
rect 4445 185532 4509 185536
rect 4445 185476 4449 185532
rect 4449 185476 4505 185532
rect 4505 185476 4509 185532
rect 4445 185472 4509 185476
rect 4525 185532 4589 185536
rect 4525 185476 4529 185532
rect 4529 185476 4585 185532
rect 4585 185476 4589 185532
rect 4525 185472 4589 185476
rect 7618 185532 7682 185536
rect 7618 185476 7622 185532
rect 7622 185476 7678 185532
rect 7678 185476 7682 185532
rect 7618 185472 7682 185476
rect 7698 185532 7762 185536
rect 7698 185476 7702 185532
rect 7702 185476 7758 185532
rect 7758 185476 7762 185532
rect 7698 185472 7762 185476
rect 7778 185532 7842 185536
rect 7778 185476 7782 185532
rect 7782 185476 7838 185532
rect 7838 185476 7842 185532
rect 7778 185472 7842 185476
rect 7858 185532 7922 185536
rect 7858 185476 7862 185532
rect 7862 185476 7918 185532
rect 7918 185476 7922 185532
rect 7858 185472 7922 185476
rect 2618 184988 2682 184992
rect 2618 184932 2622 184988
rect 2622 184932 2678 184988
rect 2678 184932 2682 184988
rect 2618 184928 2682 184932
rect 2698 184988 2762 184992
rect 2698 184932 2702 184988
rect 2702 184932 2758 184988
rect 2758 184932 2762 184988
rect 2698 184928 2762 184932
rect 2778 184988 2842 184992
rect 2778 184932 2782 184988
rect 2782 184932 2838 184988
rect 2838 184932 2842 184988
rect 2778 184928 2842 184932
rect 2858 184988 2922 184992
rect 2858 184932 2862 184988
rect 2862 184932 2918 184988
rect 2918 184932 2922 184988
rect 2858 184928 2922 184932
rect 5952 184988 6016 184992
rect 5952 184932 5956 184988
rect 5956 184932 6012 184988
rect 6012 184932 6016 184988
rect 5952 184928 6016 184932
rect 6032 184988 6096 184992
rect 6032 184932 6036 184988
rect 6036 184932 6092 184988
rect 6092 184932 6096 184988
rect 6032 184928 6096 184932
rect 6112 184988 6176 184992
rect 6112 184932 6116 184988
rect 6116 184932 6172 184988
rect 6172 184932 6176 184988
rect 6112 184928 6176 184932
rect 6192 184988 6256 184992
rect 6192 184932 6196 184988
rect 6196 184932 6252 184988
rect 6252 184932 6256 184988
rect 6192 184928 6256 184932
rect 4285 184444 4349 184448
rect 4285 184388 4289 184444
rect 4289 184388 4345 184444
rect 4345 184388 4349 184444
rect 4285 184384 4349 184388
rect 4365 184444 4429 184448
rect 4365 184388 4369 184444
rect 4369 184388 4425 184444
rect 4425 184388 4429 184444
rect 4365 184384 4429 184388
rect 4445 184444 4509 184448
rect 4445 184388 4449 184444
rect 4449 184388 4505 184444
rect 4505 184388 4509 184444
rect 4445 184384 4509 184388
rect 4525 184444 4589 184448
rect 4525 184388 4529 184444
rect 4529 184388 4585 184444
rect 4585 184388 4589 184444
rect 4525 184384 4589 184388
rect 7618 184444 7682 184448
rect 7618 184388 7622 184444
rect 7622 184388 7678 184444
rect 7678 184388 7682 184444
rect 7618 184384 7682 184388
rect 7698 184444 7762 184448
rect 7698 184388 7702 184444
rect 7702 184388 7758 184444
rect 7758 184388 7762 184444
rect 7698 184384 7762 184388
rect 7778 184444 7842 184448
rect 7778 184388 7782 184444
rect 7782 184388 7838 184444
rect 7838 184388 7842 184444
rect 7778 184384 7842 184388
rect 7858 184444 7922 184448
rect 7858 184388 7862 184444
rect 7862 184388 7918 184444
rect 7918 184388 7922 184444
rect 7858 184384 7922 184388
rect 2618 183900 2682 183904
rect 2618 183844 2622 183900
rect 2622 183844 2678 183900
rect 2678 183844 2682 183900
rect 2618 183840 2682 183844
rect 2698 183900 2762 183904
rect 2698 183844 2702 183900
rect 2702 183844 2758 183900
rect 2758 183844 2762 183900
rect 2698 183840 2762 183844
rect 2778 183900 2842 183904
rect 2778 183844 2782 183900
rect 2782 183844 2838 183900
rect 2838 183844 2842 183900
rect 2778 183840 2842 183844
rect 2858 183900 2922 183904
rect 2858 183844 2862 183900
rect 2862 183844 2918 183900
rect 2918 183844 2922 183900
rect 2858 183840 2922 183844
rect 5952 183900 6016 183904
rect 5952 183844 5956 183900
rect 5956 183844 6012 183900
rect 6012 183844 6016 183900
rect 5952 183840 6016 183844
rect 6032 183900 6096 183904
rect 6032 183844 6036 183900
rect 6036 183844 6092 183900
rect 6092 183844 6096 183900
rect 6032 183840 6096 183844
rect 6112 183900 6176 183904
rect 6112 183844 6116 183900
rect 6116 183844 6172 183900
rect 6172 183844 6176 183900
rect 6112 183840 6176 183844
rect 6192 183900 6256 183904
rect 6192 183844 6196 183900
rect 6196 183844 6252 183900
rect 6252 183844 6256 183900
rect 6192 183840 6256 183844
rect 4285 183356 4349 183360
rect 4285 183300 4289 183356
rect 4289 183300 4345 183356
rect 4345 183300 4349 183356
rect 4285 183296 4349 183300
rect 4365 183356 4429 183360
rect 4365 183300 4369 183356
rect 4369 183300 4425 183356
rect 4425 183300 4429 183356
rect 4365 183296 4429 183300
rect 4445 183356 4509 183360
rect 4445 183300 4449 183356
rect 4449 183300 4505 183356
rect 4505 183300 4509 183356
rect 4445 183296 4509 183300
rect 4525 183356 4589 183360
rect 4525 183300 4529 183356
rect 4529 183300 4585 183356
rect 4585 183300 4589 183356
rect 4525 183296 4589 183300
rect 7618 183356 7682 183360
rect 7618 183300 7622 183356
rect 7622 183300 7678 183356
rect 7678 183300 7682 183356
rect 7618 183296 7682 183300
rect 7698 183356 7762 183360
rect 7698 183300 7702 183356
rect 7702 183300 7758 183356
rect 7758 183300 7762 183356
rect 7698 183296 7762 183300
rect 7778 183356 7842 183360
rect 7778 183300 7782 183356
rect 7782 183300 7838 183356
rect 7838 183300 7842 183356
rect 7778 183296 7842 183300
rect 7858 183356 7922 183360
rect 7858 183300 7862 183356
rect 7862 183300 7918 183356
rect 7918 183300 7922 183356
rect 7858 183296 7922 183300
rect 2618 182812 2682 182816
rect 2618 182756 2622 182812
rect 2622 182756 2678 182812
rect 2678 182756 2682 182812
rect 2618 182752 2682 182756
rect 2698 182812 2762 182816
rect 2698 182756 2702 182812
rect 2702 182756 2758 182812
rect 2758 182756 2762 182812
rect 2698 182752 2762 182756
rect 2778 182812 2842 182816
rect 2778 182756 2782 182812
rect 2782 182756 2838 182812
rect 2838 182756 2842 182812
rect 2778 182752 2842 182756
rect 2858 182812 2922 182816
rect 2858 182756 2862 182812
rect 2862 182756 2918 182812
rect 2918 182756 2922 182812
rect 2858 182752 2922 182756
rect 5952 182812 6016 182816
rect 5952 182756 5956 182812
rect 5956 182756 6012 182812
rect 6012 182756 6016 182812
rect 5952 182752 6016 182756
rect 6032 182812 6096 182816
rect 6032 182756 6036 182812
rect 6036 182756 6092 182812
rect 6092 182756 6096 182812
rect 6032 182752 6096 182756
rect 6112 182812 6176 182816
rect 6112 182756 6116 182812
rect 6116 182756 6172 182812
rect 6172 182756 6176 182812
rect 6112 182752 6176 182756
rect 6192 182812 6256 182816
rect 6192 182756 6196 182812
rect 6196 182756 6252 182812
rect 6252 182756 6256 182812
rect 6192 182752 6256 182756
rect 4285 182268 4349 182272
rect 4285 182212 4289 182268
rect 4289 182212 4345 182268
rect 4345 182212 4349 182268
rect 4285 182208 4349 182212
rect 4365 182268 4429 182272
rect 4365 182212 4369 182268
rect 4369 182212 4425 182268
rect 4425 182212 4429 182268
rect 4365 182208 4429 182212
rect 4445 182268 4509 182272
rect 4445 182212 4449 182268
rect 4449 182212 4505 182268
rect 4505 182212 4509 182268
rect 4445 182208 4509 182212
rect 4525 182268 4589 182272
rect 4525 182212 4529 182268
rect 4529 182212 4585 182268
rect 4585 182212 4589 182268
rect 4525 182208 4589 182212
rect 7618 182268 7682 182272
rect 7618 182212 7622 182268
rect 7622 182212 7678 182268
rect 7678 182212 7682 182268
rect 7618 182208 7682 182212
rect 7698 182268 7762 182272
rect 7698 182212 7702 182268
rect 7702 182212 7758 182268
rect 7758 182212 7762 182268
rect 7698 182208 7762 182212
rect 7778 182268 7842 182272
rect 7778 182212 7782 182268
rect 7782 182212 7838 182268
rect 7838 182212 7842 182268
rect 7778 182208 7842 182212
rect 7858 182268 7922 182272
rect 7858 182212 7862 182268
rect 7862 182212 7918 182268
rect 7918 182212 7922 182268
rect 7858 182208 7922 182212
rect 2618 181724 2682 181728
rect 2618 181668 2622 181724
rect 2622 181668 2678 181724
rect 2678 181668 2682 181724
rect 2618 181664 2682 181668
rect 2698 181724 2762 181728
rect 2698 181668 2702 181724
rect 2702 181668 2758 181724
rect 2758 181668 2762 181724
rect 2698 181664 2762 181668
rect 2778 181724 2842 181728
rect 2778 181668 2782 181724
rect 2782 181668 2838 181724
rect 2838 181668 2842 181724
rect 2778 181664 2842 181668
rect 2858 181724 2922 181728
rect 2858 181668 2862 181724
rect 2862 181668 2918 181724
rect 2918 181668 2922 181724
rect 2858 181664 2922 181668
rect 5952 181724 6016 181728
rect 5952 181668 5956 181724
rect 5956 181668 6012 181724
rect 6012 181668 6016 181724
rect 5952 181664 6016 181668
rect 6032 181724 6096 181728
rect 6032 181668 6036 181724
rect 6036 181668 6092 181724
rect 6092 181668 6096 181724
rect 6032 181664 6096 181668
rect 6112 181724 6176 181728
rect 6112 181668 6116 181724
rect 6116 181668 6172 181724
rect 6172 181668 6176 181724
rect 6112 181664 6176 181668
rect 6192 181724 6256 181728
rect 6192 181668 6196 181724
rect 6196 181668 6252 181724
rect 6252 181668 6256 181724
rect 6192 181664 6256 181668
rect 4285 181180 4349 181184
rect 4285 181124 4289 181180
rect 4289 181124 4345 181180
rect 4345 181124 4349 181180
rect 4285 181120 4349 181124
rect 4365 181180 4429 181184
rect 4365 181124 4369 181180
rect 4369 181124 4425 181180
rect 4425 181124 4429 181180
rect 4365 181120 4429 181124
rect 4445 181180 4509 181184
rect 4445 181124 4449 181180
rect 4449 181124 4505 181180
rect 4505 181124 4509 181180
rect 4445 181120 4509 181124
rect 4525 181180 4589 181184
rect 4525 181124 4529 181180
rect 4529 181124 4585 181180
rect 4585 181124 4589 181180
rect 4525 181120 4589 181124
rect 7618 181180 7682 181184
rect 7618 181124 7622 181180
rect 7622 181124 7678 181180
rect 7678 181124 7682 181180
rect 7618 181120 7682 181124
rect 7698 181180 7762 181184
rect 7698 181124 7702 181180
rect 7702 181124 7758 181180
rect 7758 181124 7762 181180
rect 7698 181120 7762 181124
rect 7778 181180 7842 181184
rect 7778 181124 7782 181180
rect 7782 181124 7838 181180
rect 7838 181124 7842 181180
rect 7778 181120 7842 181124
rect 7858 181180 7922 181184
rect 7858 181124 7862 181180
rect 7862 181124 7918 181180
rect 7918 181124 7922 181180
rect 7858 181120 7922 181124
rect 2618 180636 2682 180640
rect 2618 180580 2622 180636
rect 2622 180580 2678 180636
rect 2678 180580 2682 180636
rect 2618 180576 2682 180580
rect 2698 180636 2762 180640
rect 2698 180580 2702 180636
rect 2702 180580 2758 180636
rect 2758 180580 2762 180636
rect 2698 180576 2762 180580
rect 2778 180636 2842 180640
rect 2778 180580 2782 180636
rect 2782 180580 2838 180636
rect 2838 180580 2842 180636
rect 2778 180576 2842 180580
rect 2858 180636 2922 180640
rect 2858 180580 2862 180636
rect 2862 180580 2918 180636
rect 2918 180580 2922 180636
rect 2858 180576 2922 180580
rect 5952 180636 6016 180640
rect 5952 180580 5956 180636
rect 5956 180580 6012 180636
rect 6012 180580 6016 180636
rect 5952 180576 6016 180580
rect 6032 180636 6096 180640
rect 6032 180580 6036 180636
rect 6036 180580 6092 180636
rect 6092 180580 6096 180636
rect 6032 180576 6096 180580
rect 6112 180636 6176 180640
rect 6112 180580 6116 180636
rect 6116 180580 6172 180636
rect 6172 180580 6176 180636
rect 6112 180576 6176 180580
rect 6192 180636 6256 180640
rect 6192 180580 6196 180636
rect 6196 180580 6252 180636
rect 6252 180580 6256 180636
rect 6192 180576 6256 180580
rect 4285 180092 4349 180096
rect 4285 180036 4289 180092
rect 4289 180036 4345 180092
rect 4345 180036 4349 180092
rect 4285 180032 4349 180036
rect 4365 180092 4429 180096
rect 4365 180036 4369 180092
rect 4369 180036 4425 180092
rect 4425 180036 4429 180092
rect 4365 180032 4429 180036
rect 4445 180092 4509 180096
rect 4445 180036 4449 180092
rect 4449 180036 4505 180092
rect 4505 180036 4509 180092
rect 4445 180032 4509 180036
rect 4525 180092 4589 180096
rect 4525 180036 4529 180092
rect 4529 180036 4585 180092
rect 4585 180036 4589 180092
rect 4525 180032 4589 180036
rect 7618 180092 7682 180096
rect 7618 180036 7622 180092
rect 7622 180036 7678 180092
rect 7678 180036 7682 180092
rect 7618 180032 7682 180036
rect 7698 180092 7762 180096
rect 7698 180036 7702 180092
rect 7702 180036 7758 180092
rect 7758 180036 7762 180092
rect 7698 180032 7762 180036
rect 7778 180092 7842 180096
rect 7778 180036 7782 180092
rect 7782 180036 7838 180092
rect 7838 180036 7842 180092
rect 7778 180032 7842 180036
rect 7858 180092 7922 180096
rect 7858 180036 7862 180092
rect 7862 180036 7918 180092
rect 7918 180036 7922 180092
rect 7858 180032 7922 180036
rect 2618 179548 2682 179552
rect 2618 179492 2622 179548
rect 2622 179492 2678 179548
rect 2678 179492 2682 179548
rect 2618 179488 2682 179492
rect 2698 179548 2762 179552
rect 2698 179492 2702 179548
rect 2702 179492 2758 179548
rect 2758 179492 2762 179548
rect 2698 179488 2762 179492
rect 2778 179548 2842 179552
rect 2778 179492 2782 179548
rect 2782 179492 2838 179548
rect 2838 179492 2842 179548
rect 2778 179488 2842 179492
rect 2858 179548 2922 179552
rect 2858 179492 2862 179548
rect 2862 179492 2918 179548
rect 2918 179492 2922 179548
rect 2858 179488 2922 179492
rect 5952 179548 6016 179552
rect 5952 179492 5956 179548
rect 5956 179492 6012 179548
rect 6012 179492 6016 179548
rect 5952 179488 6016 179492
rect 6032 179548 6096 179552
rect 6032 179492 6036 179548
rect 6036 179492 6092 179548
rect 6092 179492 6096 179548
rect 6032 179488 6096 179492
rect 6112 179548 6176 179552
rect 6112 179492 6116 179548
rect 6116 179492 6172 179548
rect 6172 179492 6176 179548
rect 6112 179488 6176 179492
rect 6192 179548 6256 179552
rect 6192 179492 6196 179548
rect 6196 179492 6252 179548
rect 6252 179492 6256 179548
rect 6192 179488 6256 179492
rect 4285 179004 4349 179008
rect 4285 178948 4289 179004
rect 4289 178948 4345 179004
rect 4345 178948 4349 179004
rect 4285 178944 4349 178948
rect 4365 179004 4429 179008
rect 4365 178948 4369 179004
rect 4369 178948 4425 179004
rect 4425 178948 4429 179004
rect 4365 178944 4429 178948
rect 4445 179004 4509 179008
rect 4445 178948 4449 179004
rect 4449 178948 4505 179004
rect 4505 178948 4509 179004
rect 4445 178944 4509 178948
rect 4525 179004 4589 179008
rect 4525 178948 4529 179004
rect 4529 178948 4585 179004
rect 4585 178948 4589 179004
rect 4525 178944 4589 178948
rect 7618 179004 7682 179008
rect 7618 178948 7622 179004
rect 7622 178948 7678 179004
rect 7678 178948 7682 179004
rect 7618 178944 7682 178948
rect 7698 179004 7762 179008
rect 7698 178948 7702 179004
rect 7702 178948 7758 179004
rect 7758 178948 7762 179004
rect 7698 178944 7762 178948
rect 7778 179004 7842 179008
rect 7778 178948 7782 179004
rect 7782 178948 7838 179004
rect 7838 178948 7842 179004
rect 7778 178944 7842 178948
rect 7858 179004 7922 179008
rect 7858 178948 7862 179004
rect 7862 178948 7918 179004
rect 7918 178948 7922 179004
rect 7858 178944 7922 178948
rect 2618 178460 2682 178464
rect 2618 178404 2622 178460
rect 2622 178404 2678 178460
rect 2678 178404 2682 178460
rect 2618 178400 2682 178404
rect 2698 178460 2762 178464
rect 2698 178404 2702 178460
rect 2702 178404 2758 178460
rect 2758 178404 2762 178460
rect 2698 178400 2762 178404
rect 2778 178460 2842 178464
rect 2778 178404 2782 178460
rect 2782 178404 2838 178460
rect 2838 178404 2842 178460
rect 2778 178400 2842 178404
rect 2858 178460 2922 178464
rect 2858 178404 2862 178460
rect 2862 178404 2918 178460
rect 2918 178404 2922 178460
rect 2858 178400 2922 178404
rect 5952 178460 6016 178464
rect 5952 178404 5956 178460
rect 5956 178404 6012 178460
rect 6012 178404 6016 178460
rect 5952 178400 6016 178404
rect 6032 178460 6096 178464
rect 6032 178404 6036 178460
rect 6036 178404 6092 178460
rect 6092 178404 6096 178460
rect 6032 178400 6096 178404
rect 6112 178460 6176 178464
rect 6112 178404 6116 178460
rect 6116 178404 6172 178460
rect 6172 178404 6176 178460
rect 6112 178400 6176 178404
rect 6192 178460 6256 178464
rect 6192 178404 6196 178460
rect 6196 178404 6252 178460
rect 6252 178404 6256 178460
rect 6192 178400 6256 178404
rect 4285 177916 4349 177920
rect 4285 177860 4289 177916
rect 4289 177860 4345 177916
rect 4345 177860 4349 177916
rect 4285 177856 4349 177860
rect 4365 177916 4429 177920
rect 4365 177860 4369 177916
rect 4369 177860 4425 177916
rect 4425 177860 4429 177916
rect 4365 177856 4429 177860
rect 4445 177916 4509 177920
rect 4445 177860 4449 177916
rect 4449 177860 4505 177916
rect 4505 177860 4509 177916
rect 4445 177856 4509 177860
rect 4525 177916 4589 177920
rect 4525 177860 4529 177916
rect 4529 177860 4585 177916
rect 4585 177860 4589 177916
rect 4525 177856 4589 177860
rect 7618 177916 7682 177920
rect 7618 177860 7622 177916
rect 7622 177860 7678 177916
rect 7678 177860 7682 177916
rect 7618 177856 7682 177860
rect 7698 177916 7762 177920
rect 7698 177860 7702 177916
rect 7702 177860 7758 177916
rect 7758 177860 7762 177916
rect 7698 177856 7762 177860
rect 7778 177916 7842 177920
rect 7778 177860 7782 177916
rect 7782 177860 7838 177916
rect 7838 177860 7842 177916
rect 7778 177856 7842 177860
rect 7858 177916 7922 177920
rect 7858 177860 7862 177916
rect 7862 177860 7918 177916
rect 7918 177860 7922 177916
rect 7858 177856 7922 177860
rect 2618 177372 2682 177376
rect 2618 177316 2622 177372
rect 2622 177316 2678 177372
rect 2678 177316 2682 177372
rect 2618 177312 2682 177316
rect 2698 177372 2762 177376
rect 2698 177316 2702 177372
rect 2702 177316 2758 177372
rect 2758 177316 2762 177372
rect 2698 177312 2762 177316
rect 2778 177372 2842 177376
rect 2778 177316 2782 177372
rect 2782 177316 2838 177372
rect 2838 177316 2842 177372
rect 2778 177312 2842 177316
rect 2858 177372 2922 177376
rect 2858 177316 2862 177372
rect 2862 177316 2918 177372
rect 2918 177316 2922 177372
rect 2858 177312 2922 177316
rect 5952 177372 6016 177376
rect 5952 177316 5956 177372
rect 5956 177316 6012 177372
rect 6012 177316 6016 177372
rect 5952 177312 6016 177316
rect 6032 177372 6096 177376
rect 6032 177316 6036 177372
rect 6036 177316 6092 177372
rect 6092 177316 6096 177372
rect 6032 177312 6096 177316
rect 6112 177372 6176 177376
rect 6112 177316 6116 177372
rect 6116 177316 6172 177372
rect 6172 177316 6176 177372
rect 6112 177312 6176 177316
rect 6192 177372 6256 177376
rect 6192 177316 6196 177372
rect 6196 177316 6252 177372
rect 6252 177316 6256 177372
rect 6192 177312 6256 177316
rect 4285 176828 4349 176832
rect 4285 176772 4289 176828
rect 4289 176772 4345 176828
rect 4345 176772 4349 176828
rect 4285 176768 4349 176772
rect 4365 176828 4429 176832
rect 4365 176772 4369 176828
rect 4369 176772 4425 176828
rect 4425 176772 4429 176828
rect 4365 176768 4429 176772
rect 4445 176828 4509 176832
rect 4445 176772 4449 176828
rect 4449 176772 4505 176828
rect 4505 176772 4509 176828
rect 4445 176768 4509 176772
rect 4525 176828 4589 176832
rect 4525 176772 4529 176828
rect 4529 176772 4585 176828
rect 4585 176772 4589 176828
rect 4525 176768 4589 176772
rect 7618 176828 7682 176832
rect 7618 176772 7622 176828
rect 7622 176772 7678 176828
rect 7678 176772 7682 176828
rect 7618 176768 7682 176772
rect 7698 176828 7762 176832
rect 7698 176772 7702 176828
rect 7702 176772 7758 176828
rect 7758 176772 7762 176828
rect 7698 176768 7762 176772
rect 7778 176828 7842 176832
rect 7778 176772 7782 176828
rect 7782 176772 7838 176828
rect 7838 176772 7842 176828
rect 7778 176768 7842 176772
rect 7858 176828 7922 176832
rect 7858 176772 7862 176828
rect 7862 176772 7918 176828
rect 7918 176772 7922 176828
rect 7858 176768 7922 176772
rect 2618 176284 2682 176288
rect 2618 176228 2622 176284
rect 2622 176228 2678 176284
rect 2678 176228 2682 176284
rect 2618 176224 2682 176228
rect 2698 176284 2762 176288
rect 2698 176228 2702 176284
rect 2702 176228 2758 176284
rect 2758 176228 2762 176284
rect 2698 176224 2762 176228
rect 2778 176284 2842 176288
rect 2778 176228 2782 176284
rect 2782 176228 2838 176284
rect 2838 176228 2842 176284
rect 2778 176224 2842 176228
rect 2858 176284 2922 176288
rect 2858 176228 2862 176284
rect 2862 176228 2918 176284
rect 2918 176228 2922 176284
rect 2858 176224 2922 176228
rect 5952 176284 6016 176288
rect 5952 176228 5956 176284
rect 5956 176228 6012 176284
rect 6012 176228 6016 176284
rect 5952 176224 6016 176228
rect 6032 176284 6096 176288
rect 6032 176228 6036 176284
rect 6036 176228 6092 176284
rect 6092 176228 6096 176284
rect 6032 176224 6096 176228
rect 6112 176284 6176 176288
rect 6112 176228 6116 176284
rect 6116 176228 6172 176284
rect 6172 176228 6176 176284
rect 6112 176224 6176 176228
rect 6192 176284 6256 176288
rect 6192 176228 6196 176284
rect 6196 176228 6252 176284
rect 6252 176228 6256 176284
rect 6192 176224 6256 176228
rect 4285 175740 4349 175744
rect 4285 175684 4289 175740
rect 4289 175684 4345 175740
rect 4345 175684 4349 175740
rect 4285 175680 4349 175684
rect 4365 175740 4429 175744
rect 4365 175684 4369 175740
rect 4369 175684 4425 175740
rect 4425 175684 4429 175740
rect 4365 175680 4429 175684
rect 4445 175740 4509 175744
rect 4445 175684 4449 175740
rect 4449 175684 4505 175740
rect 4505 175684 4509 175740
rect 4445 175680 4509 175684
rect 4525 175740 4589 175744
rect 4525 175684 4529 175740
rect 4529 175684 4585 175740
rect 4585 175684 4589 175740
rect 4525 175680 4589 175684
rect 7618 175740 7682 175744
rect 7618 175684 7622 175740
rect 7622 175684 7678 175740
rect 7678 175684 7682 175740
rect 7618 175680 7682 175684
rect 7698 175740 7762 175744
rect 7698 175684 7702 175740
rect 7702 175684 7758 175740
rect 7758 175684 7762 175740
rect 7698 175680 7762 175684
rect 7778 175740 7842 175744
rect 7778 175684 7782 175740
rect 7782 175684 7838 175740
rect 7838 175684 7842 175740
rect 7778 175680 7842 175684
rect 7858 175740 7922 175744
rect 7858 175684 7862 175740
rect 7862 175684 7918 175740
rect 7918 175684 7922 175740
rect 7858 175680 7922 175684
rect 2618 175196 2682 175200
rect 2618 175140 2622 175196
rect 2622 175140 2678 175196
rect 2678 175140 2682 175196
rect 2618 175136 2682 175140
rect 2698 175196 2762 175200
rect 2698 175140 2702 175196
rect 2702 175140 2758 175196
rect 2758 175140 2762 175196
rect 2698 175136 2762 175140
rect 2778 175196 2842 175200
rect 2778 175140 2782 175196
rect 2782 175140 2838 175196
rect 2838 175140 2842 175196
rect 2778 175136 2842 175140
rect 2858 175196 2922 175200
rect 2858 175140 2862 175196
rect 2862 175140 2918 175196
rect 2918 175140 2922 175196
rect 2858 175136 2922 175140
rect 5952 175196 6016 175200
rect 5952 175140 5956 175196
rect 5956 175140 6012 175196
rect 6012 175140 6016 175196
rect 5952 175136 6016 175140
rect 6032 175196 6096 175200
rect 6032 175140 6036 175196
rect 6036 175140 6092 175196
rect 6092 175140 6096 175196
rect 6032 175136 6096 175140
rect 6112 175196 6176 175200
rect 6112 175140 6116 175196
rect 6116 175140 6172 175196
rect 6172 175140 6176 175196
rect 6112 175136 6176 175140
rect 6192 175196 6256 175200
rect 6192 175140 6196 175196
rect 6196 175140 6252 175196
rect 6252 175140 6256 175196
rect 6192 175136 6256 175140
rect 4285 174652 4349 174656
rect 4285 174596 4289 174652
rect 4289 174596 4345 174652
rect 4345 174596 4349 174652
rect 4285 174592 4349 174596
rect 4365 174652 4429 174656
rect 4365 174596 4369 174652
rect 4369 174596 4425 174652
rect 4425 174596 4429 174652
rect 4365 174592 4429 174596
rect 4445 174652 4509 174656
rect 4445 174596 4449 174652
rect 4449 174596 4505 174652
rect 4505 174596 4509 174652
rect 4445 174592 4509 174596
rect 4525 174652 4589 174656
rect 4525 174596 4529 174652
rect 4529 174596 4585 174652
rect 4585 174596 4589 174652
rect 4525 174592 4589 174596
rect 7618 174652 7682 174656
rect 7618 174596 7622 174652
rect 7622 174596 7678 174652
rect 7678 174596 7682 174652
rect 7618 174592 7682 174596
rect 7698 174652 7762 174656
rect 7698 174596 7702 174652
rect 7702 174596 7758 174652
rect 7758 174596 7762 174652
rect 7698 174592 7762 174596
rect 7778 174652 7842 174656
rect 7778 174596 7782 174652
rect 7782 174596 7838 174652
rect 7838 174596 7842 174652
rect 7778 174592 7842 174596
rect 7858 174652 7922 174656
rect 7858 174596 7862 174652
rect 7862 174596 7918 174652
rect 7918 174596 7922 174652
rect 7858 174592 7922 174596
rect 2618 174108 2682 174112
rect 2618 174052 2622 174108
rect 2622 174052 2678 174108
rect 2678 174052 2682 174108
rect 2618 174048 2682 174052
rect 2698 174108 2762 174112
rect 2698 174052 2702 174108
rect 2702 174052 2758 174108
rect 2758 174052 2762 174108
rect 2698 174048 2762 174052
rect 2778 174108 2842 174112
rect 2778 174052 2782 174108
rect 2782 174052 2838 174108
rect 2838 174052 2842 174108
rect 2778 174048 2842 174052
rect 2858 174108 2922 174112
rect 2858 174052 2862 174108
rect 2862 174052 2918 174108
rect 2918 174052 2922 174108
rect 2858 174048 2922 174052
rect 5952 174108 6016 174112
rect 5952 174052 5956 174108
rect 5956 174052 6012 174108
rect 6012 174052 6016 174108
rect 5952 174048 6016 174052
rect 6032 174108 6096 174112
rect 6032 174052 6036 174108
rect 6036 174052 6092 174108
rect 6092 174052 6096 174108
rect 6032 174048 6096 174052
rect 6112 174108 6176 174112
rect 6112 174052 6116 174108
rect 6116 174052 6172 174108
rect 6172 174052 6176 174108
rect 6112 174048 6176 174052
rect 6192 174108 6256 174112
rect 6192 174052 6196 174108
rect 6196 174052 6252 174108
rect 6252 174052 6256 174108
rect 6192 174048 6256 174052
rect 4285 173564 4349 173568
rect 4285 173508 4289 173564
rect 4289 173508 4345 173564
rect 4345 173508 4349 173564
rect 4285 173504 4349 173508
rect 4365 173564 4429 173568
rect 4365 173508 4369 173564
rect 4369 173508 4425 173564
rect 4425 173508 4429 173564
rect 4365 173504 4429 173508
rect 4445 173564 4509 173568
rect 4445 173508 4449 173564
rect 4449 173508 4505 173564
rect 4505 173508 4509 173564
rect 4445 173504 4509 173508
rect 4525 173564 4589 173568
rect 4525 173508 4529 173564
rect 4529 173508 4585 173564
rect 4585 173508 4589 173564
rect 4525 173504 4589 173508
rect 7618 173564 7682 173568
rect 7618 173508 7622 173564
rect 7622 173508 7678 173564
rect 7678 173508 7682 173564
rect 7618 173504 7682 173508
rect 7698 173564 7762 173568
rect 7698 173508 7702 173564
rect 7702 173508 7758 173564
rect 7758 173508 7762 173564
rect 7698 173504 7762 173508
rect 7778 173564 7842 173568
rect 7778 173508 7782 173564
rect 7782 173508 7838 173564
rect 7838 173508 7842 173564
rect 7778 173504 7842 173508
rect 7858 173564 7922 173568
rect 7858 173508 7862 173564
rect 7862 173508 7918 173564
rect 7918 173508 7922 173564
rect 7858 173504 7922 173508
rect 2618 173020 2682 173024
rect 2618 172964 2622 173020
rect 2622 172964 2678 173020
rect 2678 172964 2682 173020
rect 2618 172960 2682 172964
rect 2698 173020 2762 173024
rect 2698 172964 2702 173020
rect 2702 172964 2758 173020
rect 2758 172964 2762 173020
rect 2698 172960 2762 172964
rect 2778 173020 2842 173024
rect 2778 172964 2782 173020
rect 2782 172964 2838 173020
rect 2838 172964 2842 173020
rect 2778 172960 2842 172964
rect 2858 173020 2922 173024
rect 2858 172964 2862 173020
rect 2862 172964 2918 173020
rect 2918 172964 2922 173020
rect 2858 172960 2922 172964
rect 5952 173020 6016 173024
rect 5952 172964 5956 173020
rect 5956 172964 6012 173020
rect 6012 172964 6016 173020
rect 5952 172960 6016 172964
rect 6032 173020 6096 173024
rect 6032 172964 6036 173020
rect 6036 172964 6092 173020
rect 6092 172964 6096 173020
rect 6032 172960 6096 172964
rect 6112 173020 6176 173024
rect 6112 172964 6116 173020
rect 6116 172964 6172 173020
rect 6172 172964 6176 173020
rect 6112 172960 6176 172964
rect 6192 173020 6256 173024
rect 6192 172964 6196 173020
rect 6196 172964 6252 173020
rect 6252 172964 6256 173020
rect 6192 172960 6256 172964
rect 4285 172476 4349 172480
rect 4285 172420 4289 172476
rect 4289 172420 4345 172476
rect 4345 172420 4349 172476
rect 4285 172416 4349 172420
rect 4365 172476 4429 172480
rect 4365 172420 4369 172476
rect 4369 172420 4425 172476
rect 4425 172420 4429 172476
rect 4365 172416 4429 172420
rect 4445 172476 4509 172480
rect 4445 172420 4449 172476
rect 4449 172420 4505 172476
rect 4505 172420 4509 172476
rect 4445 172416 4509 172420
rect 4525 172476 4589 172480
rect 4525 172420 4529 172476
rect 4529 172420 4585 172476
rect 4585 172420 4589 172476
rect 4525 172416 4589 172420
rect 7618 172476 7682 172480
rect 7618 172420 7622 172476
rect 7622 172420 7678 172476
rect 7678 172420 7682 172476
rect 7618 172416 7682 172420
rect 7698 172476 7762 172480
rect 7698 172420 7702 172476
rect 7702 172420 7758 172476
rect 7758 172420 7762 172476
rect 7698 172416 7762 172420
rect 7778 172476 7842 172480
rect 7778 172420 7782 172476
rect 7782 172420 7838 172476
rect 7838 172420 7842 172476
rect 7778 172416 7842 172420
rect 7858 172476 7922 172480
rect 7858 172420 7862 172476
rect 7862 172420 7918 172476
rect 7918 172420 7922 172476
rect 7858 172416 7922 172420
rect 2618 171932 2682 171936
rect 2618 171876 2622 171932
rect 2622 171876 2678 171932
rect 2678 171876 2682 171932
rect 2618 171872 2682 171876
rect 2698 171932 2762 171936
rect 2698 171876 2702 171932
rect 2702 171876 2758 171932
rect 2758 171876 2762 171932
rect 2698 171872 2762 171876
rect 2778 171932 2842 171936
rect 2778 171876 2782 171932
rect 2782 171876 2838 171932
rect 2838 171876 2842 171932
rect 2778 171872 2842 171876
rect 2858 171932 2922 171936
rect 2858 171876 2862 171932
rect 2862 171876 2918 171932
rect 2918 171876 2922 171932
rect 2858 171872 2922 171876
rect 5952 171932 6016 171936
rect 5952 171876 5956 171932
rect 5956 171876 6012 171932
rect 6012 171876 6016 171932
rect 5952 171872 6016 171876
rect 6032 171932 6096 171936
rect 6032 171876 6036 171932
rect 6036 171876 6092 171932
rect 6092 171876 6096 171932
rect 6032 171872 6096 171876
rect 6112 171932 6176 171936
rect 6112 171876 6116 171932
rect 6116 171876 6172 171932
rect 6172 171876 6176 171932
rect 6112 171872 6176 171876
rect 6192 171932 6256 171936
rect 6192 171876 6196 171932
rect 6196 171876 6252 171932
rect 6252 171876 6256 171932
rect 6192 171872 6256 171876
rect 4285 171388 4349 171392
rect 4285 171332 4289 171388
rect 4289 171332 4345 171388
rect 4345 171332 4349 171388
rect 4285 171328 4349 171332
rect 4365 171388 4429 171392
rect 4365 171332 4369 171388
rect 4369 171332 4425 171388
rect 4425 171332 4429 171388
rect 4365 171328 4429 171332
rect 4445 171388 4509 171392
rect 4445 171332 4449 171388
rect 4449 171332 4505 171388
rect 4505 171332 4509 171388
rect 4445 171328 4509 171332
rect 4525 171388 4589 171392
rect 4525 171332 4529 171388
rect 4529 171332 4585 171388
rect 4585 171332 4589 171388
rect 4525 171328 4589 171332
rect 7618 171388 7682 171392
rect 7618 171332 7622 171388
rect 7622 171332 7678 171388
rect 7678 171332 7682 171388
rect 7618 171328 7682 171332
rect 7698 171388 7762 171392
rect 7698 171332 7702 171388
rect 7702 171332 7758 171388
rect 7758 171332 7762 171388
rect 7698 171328 7762 171332
rect 7778 171388 7842 171392
rect 7778 171332 7782 171388
rect 7782 171332 7838 171388
rect 7838 171332 7842 171388
rect 7778 171328 7842 171332
rect 7858 171388 7922 171392
rect 7858 171332 7862 171388
rect 7862 171332 7918 171388
rect 7918 171332 7922 171388
rect 7858 171328 7922 171332
rect 2618 170844 2682 170848
rect 2618 170788 2622 170844
rect 2622 170788 2678 170844
rect 2678 170788 2682 170844
rect 2618 170784 2682 170788
rect 2698 170844 2762 170848
rect 2698 170788 2702 170844
rect 2702 170788 2758 170844
rect 2758 170788 2762 170844
rect 2698 170784 2762 170788
rect 2778 170844 2842 170848
rect 2778 170788 2782 170844
rect 2782 170788 2838 170844
rect 2838 170788 2842 170844
rect 2778 170784 2842 170788
rect 2858 170844 2922 170848
rect 2858 170788 2862 170844
rect 2862 170788 2918 170844
rect 2918 170788 2922 170844
rect 2858 170784 2922 170788
rect 5952 170844 6016 170848
rect 5952 170788 5956 170844
rect 5956 170788 6012 170844
rect 6012 170788 6016 170844
rect 5952 170784 6016 170788
rect 6032 170844 6096 170848
rect 6032 170788 6036 170844
rect 6036 170788 6092 170844
rect 6092 170788 6096 170844
rect 6032 170784 6096 170788
rect 6112 170844 6176 170848
rect 6112 170788 6116 170844
rect 6116 170788 6172 170844
rect 6172 170788 6176 170844
rect 6112 170784 6176 170788
rect 6192 170844 6256 170848
rect 6192 170788 6196 170844
rect 6196 170788 6252 170844
rect 6252 170788 6256 170844
rect 6192 170784 6256 170788
rect 4285 170300 4349 170304
rect 4285 170244 4289 170300
rect 4289 170244 4345 170300
rect 4345 170244 4349 170300
rect 4285 170240 4349 170244
rect 4365 170300 4429 170304
rect 4365 170244 4369 170300
rect 4369 170244 4425 170300
rect 4425 170244 4429 170300
rect 4365 170240 4429 170244
rect 4445 170300 4509 170304
rect 4445 170244 4449 170300
rect 4449 170244 4505 170300
rect 4505 170244 4509 170300
rect 4445 170240 4509 170244
rect 4525 170300 4589 170304
rect 4525 170244 4529 170300
rect 4529 170244 4585 170300
rect 4585 170244 4589 170300
rect 4525 170240 4589 170244
rect 7618 170300 7682 170304
rect 7618 170244 7622 170300
rect 7622 170244 7678 170300
rect 7678 170244 7682 170300
rect 7618 170240 7682 170244
rect 7698 170300 7762 170304
rect 7698 170244 7702 170300
rect 7702 170244 7758 170300
rect 7758 170244 7762 170300
rect 7698 170240 7762 170244
rect 7778 170300 7842 170304
rect 7778 170244 7782 170300
rect 7782 170244 7838 170300
rect 7838 170244 7842 170300
rect 7778 170240 7842 170244
rect 7858 170300 7922 170304
rect 7858 170244 7862 170300
rect 7862 170244 7918 170300
rect 7918 170244 7922 170300
rect 7858 170240 7922 170244
rect 2618 169756 2682 169760
rect 2618 169700 2622 169756
rect 2622 169700 2678 169756
rect 2678 169700 2682 169756
rect 2618 169696 2682 169700
rect 2698 169756 2762 169760
rect 2698 169700 2702 169756
rect 2702 169700 2758 169756
rect 2758 169700 2762 169756
rect 2698 169696 2762 169700
rect 2778 169756 2842 169760
rect 2778 169700 2782 169756
rect 2782 169700 2838 169756
rect 2838 169700 2842 169756
rect 2778 169696 2842 169700
rect 2858 169756 2922 169760
rect 2858 169700 2862 169756
rect 2862 169700 2918 169756
rect 2918 169700 2922 169756
rect 2858 169696 2922 169700
rect 5952 169756 6016 169760
rect 5952 169700 5956 169756
rect 5956 169700 6012 169756
rect 6012 169700 6016 169756
rect 5952 169696 6016 169700
rect 6032 169756 6096 169760
rect 6032 169700 6036 169756
rect 6036 169700 6092 169756
rect 6092 169700 6096 169756
rect 6032 169696 6096 169700
rect 6112 169756 6176 169760
rect 6112 169700 6116 169756
rect 6116 169700 6172 169756
rect 6172 169700 6176 169756
rect 6112 169696 6176 169700
rect 6192 169756 6256 169760
rect 6192 169700 6196 169756
rect 6196 169700 6252 169756
rect 6252 169700 6256 169756
rect 6192 169696 6256 169700
rect 4285 169212 4349 169216
rect 4285 169156 4289 169212
rect 4289 169156 4345 169212
rect 4345 169156 4349 169212
rect 4285 169152 4349 169156
rect 4365 169212 4429 169216
rect 4365 169156 4369 169212
rect 4369 169156 4425 169212
rect 4425 169156 4429 169212
rect 4365 169152 4429 169156
rect 4445 169212 4509 169216
rect 4445 169156 4449 169212
rect 4449 169156 4505 169212
rect 4505 169156 4509 169212
rect 4445 169152 4509 169156
rect 4525 169212 4589 169216
rect 4525 169156 4529 169212
rect 4529 169156 4585 169212
rect 4585 169156 4589 169212
rect 4525 169152 4589 169156
rect 7618 169212 7682 169216
rect 7618 169156 7622 169212
rect 7622 169156 7678 169212
rect 7678 169156 7682 169212
rect 7618 169152 7682 169156
rect 7698 169212 7762 169216
rect 7698 169156 7702 169212
rect 7702 169156 7758 169212
rect 7758 169156 7762 169212
rect 7698 169152 7762 169156
rect 7778 169212 7842 169216
rect 7778 169156 7782 169212
rect 7782 169156 7838 169212
rect 7838 169156 7842 169212
rect 7778 169152 7842 169156
rect 7858 169212 7922 169216
rect 7858 169156 7862 169212
rect 7862 169156 7918 169212
rect 7918 169156 7922 169212
rect 7858 169152 7922 169156
rect 2618 168668 2682 168672
rect 2618 168612 2622 168668
rect 2622 168612 2678 168668
rect 2678 168612 2682 168668
rect 2618 168608 2682 168612
rect 2698 168668 2762 168672
rect 2698 168612 2702 168668
rect 2702 168612 2758 168668
rect 2758 168612 2762 168668
rect 2698 168608 2762 168612
rect 2778 168668 2842 168672
rect 2778 168612 2782 168668
rect 2782 168612 2838 168668
rect 2838 168612 2842 168668
rect 2778 168608 2842 168612
rect 2858 168668 2922 168672
rect 2858 168612 2862 168668
rect 2862 168612 2918 168668
rect 2918 168612 2922 168668
rect 2858 168608 2922 168612
rect 5952 168668 6016 168672
rect 5952 168612 5956 168668
rect 5956 168612 6012 168668
rect 6012 168612 6016 168668
rect 5952 168608 6016 168612
rect 6032 168668 6096 168672
rect 6032 168612 6036 168668
rect 6036 168612 6092 168668
rect 6092 168612 6096 168668
rect 6032 168608 6096 168612
rect 6112 168668 6176 168672
rect 6112 168612 6116 168668
rect 6116 168612 6172 168668
rect 6172 168612 6176 168668
rect 6112 168608 6176 168612
rect 6192 168668 6256 168672
rect 6192 168612 6196 168668
rect 6196 168612 6252 168668
rect 6252 168612 6256 168668
rect 6192 168608 6256 168612
rect 4285 168124 4349 168128
rect 4285 168068 4289 168124
rect 4289 168068 4345 168124
rect 4345 168068 4349 168124
rect 4285 168064 4349 168068
rect 4365 168124 4429 168128
rect 4365 168068 4369 168124
rect 4369 168068 4425 168124
rect 4425 168068 4429 168124
rect 4365 168064 4429 168068
rect 4445 168124 4509 168128
rect 4445 168068 4449 168124
rect 4449 168068 4505 168124
rect 4505 168068 4509 168124
rect 4445 168064 4509 168068
rect 4525 168124 4589 168128
rect 4525 168068 4529 168124
rect 4529 168068 4585 168124
rect 4585 168068 4589 168124
rect 4525 168064 4589 168068
rect 7618 168124 7682 168128
rect 7618 168068 7622 168124
rect 7622 168068 7678 168124
rect 7678 168068 7682 168124
rect 7618 168064 7682 168068
rect 7698 168124 7762 168128
rect 7698 168068 7702 168124
rect 7702 168068 7758 168124
rect 7758 168068 7762 168124
rect 7698 168064 7762 168068
rect 7778 168124 7842 168128
rect 7778 168068 7782 168124
rect 7782 168068 7838 168124
rect 7838 168068 7842 168124
rect 7778 168064 7842 168068
rect 7858 168124 7922 168128
rect 7858 168068 7862 168124
rect 7862 168068 7918 168124
rect 7918 168068 7922 168124
rect 7858 168064 7922 168068
rect 2618 167580 2682 167584
rect 2618 167524 2622 167580
rect 2622 167524 2678 167580
rect 2678 167524 2682 167580
rect 2618 167520 2682 167524
rect 2698 167580 2762 167584
rect 2698 167524 2702 167580
rect 2702 167524 2758 167580
rect 2758 167524 2762 167580
rect 2698 167520 2762 167524
rect 2778 167580 2842 167584
rect 2778 167524 2782 167580
rect 2782 167524 2838 167580
rect 2838 167524 2842 167580
rect 2778 167520 2842 167524
rect 2858 167580 2922 167584
rect 2858 167524 2862 167580
rect 2862 167524 2918 167580
rect 2918 167524 2922 167580
rect 2858 167520 2922 167524
rect 5952 167580 6016 167584
rect 5952 167524 5956 167580
rect 5956 167524 6012 167580
rect 6012 167524 6016 167580
rect 5952 167520 6016 167524
rect 6032 167580 6096 167584
rect 6032 167524 6036 167580
rect 6036 167524 6092 167580
rect 6092 167524 6096 167580
rect 6032 167520 6096 167524
rect 6112 167580 6176 167584
rect 6112 167524 6116 167580
rect 6116 167524 6172 167580
rect 6172 167524 6176 167580
rect 6112 167520 6176 167524
rect 6192 167580 6256 167584
rect 6192 167524 6196 167580
rect 6196 167524 6252 167580
rect 6252 167524 6256 167580
rect 6192 167520 6256 167524
rect 4285 167036 4349 167040
rect 4285 166980 4289 167036
rect 4289 166980 4345 167036
rect 4345 166980 4349 167036
rect 4285 166976 4349 166980
rect 4365 167036 4429 167040
rect 4365 166980 4369 167036
rect 4369 166980 4425 167036
rect 4425 166980 4429 167036
rect 4365 166976 4429 166980
rect 4445 167036 4509 167040
rect 4445 166980 4449 167036
rect 4449 166980 4505 167036
rect 4505 166980 4509 167036
rect 4445 166976 4509 166980
rect 4525 167036 4589 167040
rect 4525 166980 4529 167036
rect 4529 166980 4585 167036
rect 4585 166980 4589 167036
rect 4525 166976 4589 166980
rect 7618 167036 7682 167040
rect 7618 166980 7622 167036
rect 7622 166980 7678 167036
rect 7678 166980 7682 167036
rect 7618 166976 7682 166980
rect 7698 167036 7762 167040
rect 7698 166980 7702 167036
rect 7702 166980 7758 167036
rect 7758 166980 7762 167036
rect 7698 166976 7762 166980
rect 7778 167036 7842 167040
rect 7778 166980 7782 167036
rect 7782 166980 7838 167036
rect 7838 166980 7842 167036
rect 7778 166976 7842 166980
rect 7858 167036 7922 167040
rect 7858 166980 7862 167036
rect 7862 166980 7918 167036
rect 7918 166980 7922 167036
rect 7858 166976 7922 166980
rect 2618 166492 2682 166496
rect 2618 166436 2622 166492
rect 2622 166436 2678 166492
rect 2678 166436 2682 166492
rect 2618 166432 2682 166436
rect 2698 166492 2762 166496
rect 2698 166436 2702 166492
rect 2702 166436 2758 166492
rect 2758 166436 2762 166492
rect 2698 166432 2762 166436
rect 2778 166492 2842 166496
rect 2778 166436 2782 166492
rect 2782 166436 2838 166492
rect 2838 166436 2842 166492
rect 2778 166432 2842 166436
rect 2858 166492 2922 166496
rect 2858 166436 2862 166492
rect 2862 166436 2918 166492
rect 2918 166436 2922 166492
rect 2858 166432 2922 166436
rect 5952 166492 6016 166496
rect 5952 166436 5956 166492
rect 5956 166436 6012 166492
rect 6012 166436 6016 166492
rect 5952 166432 6016 166436
rect 6032 166492 6096 166496
rect 6032 166436 6036 166492
rect 6036 166436 6092 166492
rect 6092 166436 6096 166492
rect 6032 166432 6096 166436
rect 6112 166492 6176 166496
rect 6112 166436 6116 166492
rect 6116 166436 6172 166492
rect 6172 166436 6176 166492
rect 6112 166432 6176 166436
rect 6192 166492 6256 166496
rect 6192 166436 6196 166492
rect 6196 166436 6252 166492
rect 6252 166436 6256 166492
rect 6192 166432 6256 166436
rect 4285 165948 4349 165952
rect 4285 165892 4289 165948
rect 4289 165892 4345 165948
rect 4345 165892 4349 165948
rect 4285 165888 4349 165892
rect 4365 165948 4429 165952
rect 4365 165892 4369 165948
rect 4369 165892 4425 165948
rect 4425 165892 4429 165948
rect 4365 165888 4429 165892
rect 4445 165948 4509 165952
rect 4445 165892 4449 165948
rect 4449 165892 4505 165948
rect 4505 165892 4509 165948
rect 4445 165888 4509 165892
rect 4525 165948 4589 165952
rect 4525 165892 4529 165948
rect 4529 165892 4585 165948
rect 4585 165892 4589 165948
rect 4525 165888 4589 165892
rect 7618 165948 7682 165952
rect 7618 165892 7622 165948
rect 7622 165892 7678 165948
rect 7678 165892 7682 165948
rect 7618 165888 7682 165892
rect 7698 165948 7762 165952
rect 7698 165892 7702 165948
rect 7702 165892 7758 165948
rect 7758 165892 7762 165948
rect 7698 165888 7762 165892
rect 7778 165948 7842 165952
rect 7778 165892 7782 165948
rect 7782 165892 7838 165948
rect 7838 165892 7842 165948
rect 7778 165888 7842 165892
rect 7858 165948 7922 165952
rect 7858 165892 7862 165948
rect 7862 165892 7918 165948
rect 7918 165892 7922 165948
rect 7858 165888 7922 165892
rect 2618 165404 2682 165408
rect 2618 165348 2622 165404
rect 2622 165348 2678 165404
rect 2678 165348 2682 165404
rect 2618 165344 2682 165348
rect 2698 165404 2762 165408
rect 2698 165348 2702 165404
rect 2702 165348 2758 165404
rect 2758 165348 2762 165404
rect 2698 165344 2762 165348
rect 2778 165404 2842 165408
rect 2778 165348 2782 165404
rect 2782 165348 2838 165404
rect 2838 165348 2842 165404
rect 2778 165344 2842 165348
rect 2858 165404 2922 165408
rect 2858 165348 2862 165404
rect 2862 165348 2918 165404
rect 2918 165348 2922 165404
rect 2858 165344 2922 165348
rect 5952 165404 6016 165408
rect 5952 165348 5956 165404
rect 5956 165348 6012 165404
rect 6012 165348 6016 165404
rect 5952 165344 6016 165348
rect 6032 165404 6096 165408
rect 6032 165348 6036 165404
rect 6036 165348 6092 165404
rect 6092 165348 6096 165404
rect 6032 165344 6096 165348
rect 6112 165404 6176 165408
rect 6112 165348 6116 165404
rect 6116 165348 6172 165404
rect 6172 165348 6176 165404
rect 6112 165344 6176 165348
rect 6192 165404 6256 165408
rect 6192 165348 6196 165404
rect 6196 165348 6252 165404
rect 6252 165348 6256 165404
rect 6192 165344 6256 165348
rect 4285 164860 4349 164864
rect 4285 164804 4289 164860
rect 4289 164804 4345 164860
rect 4345 164804 4349 164860
rect 4285 164800 4349 164804
rect 4365 164860 4429 164864
rect 4365 164804 4369 164860
rect 4369 164804 4425 164860
rect 4425 164804 4429 164860
rect 4365 164800 4429 164804
rect 4445 164860 4509 164864
rect 4445 164804 4449 164860
rect 4449 164804 4505 164860
rect 4505 164804 4509 164860
rect 4445 164800 4509 164804
rect 4525 164860 4589 164864
rect 4525 164804 4529 164860
rect 4529 164804 4585 164860
rect 4585 164804 4589 164860
rect 4525 164800 4589 164804
rect 7618 164860 7682 164864
rect 7618 164804 7622 164860
rect 7622 164804 7678 164860
rect 7678 164804 7682 164860
rect 7618 164800 7682 164804
rect 7698 164860 7762 164864
rect 7698 164804 7702 164860
rect 7702 164804 7758 164860
rect 7758 164804 7762 164860
rect 7698 164800 7762 164804
rect 7778 164860 7842 164864
rect 7778 164804 7782 164860
rect 7782 164804 7838 164860
rect 7838 164804 7842 164860
rect 7778 164800 7842 164804
rect 7858 164860 7922 164864
rect 7858 164804 7862 164860
rect 7862 164804 7918 164860
rect 7918 164804 7922 164860
rect 7858 164800 7922 164804
rect 2618 164316 2682 164320
rect 2618 164260 2622 164316
rect 2622 164260 2678 164316
rect 2678 164260 2682 164316
rect 2618 164256 2682 164260
rect 2698 164316 2762 164320
rect 2698 164260 2702 164316
rect 2702 164260 2758 164316
rect 2758 164260 2762 164316
rect 2698 164256 2762 164260
rect 2778 164316 2842 164320
rect 2778 164260 2782 164316
rect 2782 164260 2838 164316
rect 2838 164260 2842 164316
rect 2778 164256 2842 164260
rect 2858 164316 2922 164320
rect 2858 164260 2862 164316
rect 2862 164260 2918 164316
rect 2918 164260 2922 164316
rect 2858 164256 2922 164260
rect 5952 164316 6016 164320
rect 5952 164260 5956 164316
rect 5956 164260 6012 164316
rect 6012 164260 6016 164316
rect 5952 164256 6016 164260
rect 6032 164316 6096 164320
rect 6032 164260 6036 164316
rect 6036 164260 6092 164316
rect 6092 164260 6096 164316
rect 6032 164256 6096 164260
rect 6112 164316 6176 164320
rect 6112 164260 6116 164316
rect 6116 164260 6172 164316
rect 6172 164260 6176 164316
rect 6112 164256 6176 164260
rect 6192 164316 6256 164320
rect 6192 164260 6196 164316
rect 6196 164260 6252 164316
rect 6252 164260 6256 164316
rect 6192 164256 6256 164260
rect 4285 163772 4349 163776
rect 4285 163716 4289 163772
rect 4289 163716 4345 163772
rect 4345 163716 4349 163772
rect 4285 163712 4349 163716
rect 4365 163772 4429 163776
rect 4365 163716 4369 163772
rect 4369 163716 4425 163772
rect 4425 163716 4429 163772
rect 4365 163712 4429 163716
rect 4445 163772 4509 163776
rect 4445 163716 4449 163772
rect 4449 163716 4505 163772
rect 4505 163716 4509 163772
rect 4445 163712 4509 163716
rect 4525 163772 4589 163776
rect 4525 163716 4529 163772
rect 4529 163716 4585 163772
rect 4585 163716 4589 163772
rect 4525 163712 4589 163716
rect 7618 163772 7682 163776
rect 7618 163716 7622 163772
rect 7622 163716 7678 163772
rect 7678 163716 7682 163772
rect 7618 163712 7682 163716
rect 7698 163772 7762 163776
rect 7698 163716 7702 163772
rect 7702 163716 7758 163772
rect 7758 163716 7762 163772
rect 7698 163712 7762 163716
rect 7778 163772 7842 163776
rect 7778 163716 7782 163772
rect 7782 163716 7838 163772
rect 7838 163716 7842 163772
rect 7778 163712 7842 163716
rect 7858 163772 7922 163776
rect 7858 163716 7862 163772
rect 7862 163716 7918 163772
rect 7918 163716 7922 163772
rect 7858 163712 7922 163716
rect 2618 163228 2682 163232
rect 2618 163172 2622 163228
rect 2622 163172 2678 163228
rect 2678 163172 2682 163228
rect 2618 163168 2682 163172
rect 2698 163228 2762 163232
rect 2698 163172 2702 163228
rect 2702 163172 2758 163228
rect 2758 163172 2762 163228
rect 2698 163168 2762 163172
rect 2778 163228 2842 163232
rect 2778 163172 2782 163228
rect 2782 163172 2838 163228
rect 2838 163172 2842 163228
rect 2778 163168 2842 163172
rect 2858 163228 2922 163232
rect 2858 163172 2862 163228
rect 2862 163172 2918 163228
rect 2918 163172 2922 163228
rect 2858 163168 2922 163172
rect 5952 163228 6016 163232
rect 5952 163172 5956 163228
rect 5956 163172 6012 163228
rect 6012 163172 6016 163228
rect 5952 163168 6016 163172
rect 6032 163228 6096 163232
rect 6032 163172 6036 163228
rect 6036 163172 6092 163228
rect 6092 163172 6096 163228
rect 6032 163168 6096 163172
rect 6112 163228 6176 163232
rect 6112 163172 6116 163228
rect 6116 163172 6172 163228
rect 6172 163172 6176 163228
rect 6112 163168 6176 163172
rect 6192 163228 6256 163232
rect 6192 163172 6196 163228
rect 6196 163172 6252 163228
rect 6252 163172 6256 163228
rect 6192 163168 6256 163172
rect 4285 162684 4349 162688
rect 4285 162628 4289 162684
rect 4289 162628 4345 162684
rect 4345 162628 4349 162684
rect 4285 162624 4349 162628
rect 4365 162684 4429 162688
rect 4365 162628 4369 162684
rect 4369 162628 4425 162684
rect 4425 162628 4429 162684
rect 4365 162624 4429 162628
rect 4445 162684 4509 162688
rect 4445 162628 4449 162684
rect 4449 162628 4505 162684
rect 4505 162628 4509 162684
rect 4445 162624 4509 162628
rect 4525 162684 4589 162688
rect 4525 162628 4529 162684
rect 4529 162628 4585 162684
rect 4585 162628 4589 162684
rect 4525 162624 4589 162628
rect 7618 162684 7682 162688
rect 7618 162628 7622 162684
rect 7622 162628 7678 162684
rect 7678 162628 7682 162684
rect 7618 162624 7682 162628
rect 7698 162684 7762 162688
rect 7698 162628 7702 162684
rect 7702 162628 7758 162684
rect 7758 162628 7762 162684
rect 7698 162624 7762 162628
rect 7778 162684 7842 162688
rect 7778 162628 7782 162684
rect 7782 162628 7838 162684
rect 7838 162628 7842 162684
rect 7778 162624 7842 162628
rect 7858 162684 7922 162688
rect 7858 162628 7862 162684
rect 7862 162628 7918 162684
rect 7918 162628 7922 162684
rect 7858 162624 7922 162628
rect 2618 162140 2682 162144
rect 2618 162084 2622 162140
rect 2622 162084 2678 162140
rect 2678 162084 2682 162140
rect 2618 162080 2682 162084
rect 2698 162140 2762 162144
rect 2698 162084 2702 162140
rect 2702 162084 2758 162140
rect 2758 162084 2762 162140
rect 2698 162080 2762 162084
rect 2778 162140 2842 162144
rect 2778 162084 2782 162140
rect 2782 162084 2838 162140
rect 2838 162084 2842 162140
rect 2778 162080 2842 162084
rect 2858 162140 2922 162144
rect 2858 162084 2862 162140
rect 2862 162084 2918 162140
rect 2918 162084 2922 162140
rect 2858 162080 2922 162084
rect 5952 162140 6016 162144
rect 5952 162084 5956 162140
rect 5956 162084 6012 162140
rect 6012 162084 6016 162140
rect 5952 162080 6016 162084
rect 6032 162140 6096 162144
rect 6032 162084 6036 162140
rect 6036 162084 6092 162140
rect 6092 162084 6096 162140
rect 6032 162080 6096 162084
rect 6112 162140 6176 162144
rect 6112 162084 6116 162140
rect 6116 162084 6172 162140
rect 6172 162084 6176 162140
rect 6112 162080 6176 162084
rect 6192 162140 6256 162144
rect 6192 162084 6196 162140
rect 6196 162084 6252 162140
rect 6252 162084 6256 162140
rect 6192 162080 6256 162084
rect 4285 161596 4349 161600
rect 4285 161540 4289 161596
rect 4289 161540 4345 161596
rect 4345 161540 4349 161596
rect 4285 161536 4349 161540
rect 4365 161596 4429 161600
rect 4365 161540 4369 161596
rect 4369 161540 4425 161596
rect 4425 161540 4429 161596
rect 4365 161536 4429 161540
rect 4445 161596 4509 161600
rect 4445 161540 4449 161596
rect 4449 161540 4505 161596
rect 4505 161540 4509 161596
rect 4445 161536 4509 161540
rect 4525 161596 4589 161600
rect 4525 161540 4529 161596
rect 4529 161540 4585 161596
rect 4585 161540 4589 161596
rect 4525 161536 4589 161540
rect 7618 161596 7682 161600
rect 7618 161540 7622 161596
rect 7622 161540 7678 161596
rect 7678 161540 7682 161596
rect 7618 161536 7682 161540
rect 7698 161596 7762 161600
rect 7698 161540 7702 161596
rect 7702 161540 7758 161596
rect 7758 161540 7762 161596
rect 7698 161536 7762 161540
rect 7778 161596 7842 161600
rect 7778 161540 7782 161596
rect 7782 161540 7838 161596
rect 7838 161540 7842 161596
rect 7778 161536 7842 161540
rect 7858 161596 7922 161600
rect 7858 161540 7862 161596
rect 7862 161540 7918 161596
rect 7918 161540 7922 161596
rect 7858 161536 7922 161540
rect 2618 161052 2682 161056
rect 2618 160996 2622 161052
rect 2622 160996 2678 161052
rect 2678 160996 2682 161052
rect 2618 160992 2682 160996
rect 2698 161052 2762 161056
rect 2698 160996 2702 161052
rect 2702 160996 2758 161052
rect 2758 160996 2762 161052
rect 2698 160992 2762 160996
rect 2778 161052 2842 161056
rect 2778 160996 2782 161052
rect 2782 160996 2838 161052
rect 2838 160996 2842 161052
rect 2778 160992 2842 160996
rect 2858 161052 2922 161056
rect 2858 160996 2862 161052
rect 2862 160996 2918 161052
rect 2918 160996 2922 161052
rect 2858 160992 2922 160996
rect 5952 161052 6016 161056
rect 5952 160996 5956 161052
rect 5956 160996 6012 161052
rect 6012 160996 6016 161052
rect 5952 160992 6016 160996
rect 6032 161052 6096 161056
rect 6032 160996 6036 161052
rect 6036 160996 6092 161052
rect 6092 160996 6096 161052
rect 6032 160992 6096 160996
rect 6112 161052 6176 161056
rect 6112 160996 6116 161052
rect 6116 160996 6172 161052
rect 6172 160996 6176 161052
rect 6112 160992 6176 160996
rect 6192 161052 6256 161056
rect 6192 160996 6196 161052
rect 6196 160996 6252 161052
rect 6252 160996 6256 161052
rect 6192 160992 6256 160996
rect 4285 160508 4349 160512
rect 4285 160452 4289 160508
rect 4289 160452 4345 160508
rect 4345 160452 4349 160508
rect 4285 160448 4349 160452
rect 4365 160508 4429 160512
rect 4365 160452 4369 160508
rect 4369 160452 4425 160508
rect 4425 160452 4429 160508
rect 4365 160448 4429 160452
rect 4445 160508 4509 160512
rect 4445 160452 4449 160508
rect 4449 160452 4505 160508
rect 4505 160452 4509 160508
rect 4445 160448 4509 160452
rect 4525 160508 4589 160512
rect 4525 160452 4529 160508
rect 4529 160452 4585 160508
rect 4585 160452 4589 160508
rect 4525 160448 4589 160452
rect 7618 160508 7682 160512
rect 7618 160452 7622 160508
rect 7622 160452 7678 160508
rect 7678 160452 7682 160508
rect 7618 160448 7682 160452
rect 7698 160508 7762 160512
rect 7698 160452 7702 160508
rect 7702 160452 7758 160508
rect 7758 160452 7762 160508
rect 7698 160448 7762 160452
rect 7778 160508 7842 160512
rect 7778 160452 7782 160508
rect 7782 160452 7838 160508
rect 7838 160452 7842 160508
rect 7778 160448 7842 160452
rect 7858 160508 7922 160512
rect 7858 160452 7862 160508
rect 7862 160452 7918 160508
rect 7918 160452 7922 160508
rect 7858 160448 7922 160452
rect 2618 159964 2682 159968
rect 2618 159908 2622 159964
rect 2622 159908 2678 159964
rect 2678 159908 2682 159964
rect 2618 159904 2682 159908
rect 2698 159964 2762 159968
rect 2698 159908 2702 159964
rect 2702 159908 2758 159964
rect 2758 159908 2762 159964
rect 2698 159904 2762 159908
rect 2778 159964 2842 159968
rect 2778 159908 2782 159964
rect 2782 159908 2838 159964
rect 2838 159908 2842 159964
rect 2778 159904 2842 159908
rect 2858 159964 2922 159968
rect 2858 159908 2862 159964
rect 2862 159908 2918 159964
rect 2918 159908 2922 159964
rect 2858 159904 2922 159908
rect 5952 159964 6016 159968
rect 5952 159908 5956 159964
rect 5956 159908 6012 159964
rect 6012 159908 6016 159964
rect 5952 159904 6016 159908
rect 6032 159964 6096 159968
rect 6032 159908 6036 159964
rect 6036 159908 6092 159964
rect 6092 159908 6096 159964
rect 6032 159904 6096 159908
rect 6112 159964 6176 159968
rect 6112 159908 6116 159964
rect 6116 159908 6172 159964
rect 6172 159908 6176 159964
rect 6112 159904 6176 159908
rect 6192 159964 6256 159968
rect 6192 159908 6196 159964
rect 6196 159908 6252 159964
rect 6252 159908 6256 159964
rect 6192 159904 6256 159908
rect 4285 159420 4349 159424
rect 4285 159364 4289 159420
rect 4289 159364 4345 159420
rect 4345 159364 4349 159420
rect 4285 159360 4349 159364
rect 4365 159420 4429 159424
rect 4365 159364 4369 159420
rect 4369 159364 4425 159420
rect 4425 159364 4429 159420
rect 4365 159360 4429 159364
rect 4445 159420 4509 159424
rect 4445 159364 4449 159420
rect 4449 159364 4505 159420
rect 4505 159364 4509 159420
rect 4445 159360 4509 159364
rect 4525 159420 4589 159424
rect 4525 159364 4529 159420
rect 4529 159364 4585 159420
rect 4585 159364 4589 159420
rect 4525 159360 4589 159364
rect 7618 159420 7682 159424
rect 7618 159364 7622 159420
rect 7622 159364 7678 159420
rect 7678 159364 7682 159420
rect 7618 159360 7682 159364
rect 7698 159420 7762 159424
rect 7698 159364 7702 159420
rect 7702 159364 7758 159420
rect 7758 159364 7762 159420
rect 7698 159360 7762 159364
rect 7778 159420 7842 159424
rect 7778 159364 7782 159420
rect 7782 159364 7838 159420
rect 7838 159364 7842 159420
rect 7778 159360 7842 159364
rect 7858 159420 7922 159424
rect 7858 159364 7862 159420
rect 7862 159364 7918 159420
rect 7918 159364 7922 159420
rect 7858 159360 7922 159364
rect 2618 158876 2682 158880
rect 2618 158820 2622 158876
rect 2622 158820 2678 158876
rect 2678 158820 2682 158876
rect 2618 158816 2682 158820
rect 2698 158876 2762 158880
rect 2698 158820 2702 158876
rect 2702 158820 2758 158876
rect 2758 158820 2762 158876
rect 2698 158816 2762 158820
rect 2778 158876 2842 158880
rect 2778 158820 2782 158876
rect 2782 158820 2838 158876
rect 2838 158820 2842 158876
rect 2778 158816 2842 158820
rect 2858 158876 2922 158880
rect 2858 158820 2862 158876
rect 2862 158820 2918 158876
rect 2918 158820 2922 158876
rect 2858 158816 2922 158820
rect 5952 158876 6016 158880
rect 5952 158820 5956 158876
rect 5956 158820 6012 158876
rect 6012 158820 6016 158876
rect 5952 158816 6016 158820
rect 6032 158876 6096 158880
rect 6032 158820 6036 158876
rect 6036 158820 6092 158876
rect 6092 158820 6096 158876
rect 6032 158816 6096 158820
rect 6112 158876 6176 158880
rect 6112 158820 6116 158876
rect 6116 158820 6172 158876
rect 6172 158820 6176 158876
rect 6112 158816 6176 158820
rect 6192 158876 6256 158880
rect 6192 158820 6196 158876
rect 6196 158820 6252 158876
rect 6252 158820 6256 158876
rect 6192 158816 6256 158820
rect 4285 158332 4349 158336
rect 4285 158276 4289 158332
rect 4289 158276 4345 158332
rect 4345 158276 4349 158332
rect 4285 158272 4349 158276
rect 4365 158332 4429 158336
rect 4365 158276 4369 158332
rect 4369 158276 4425 158332
rect 4425 158276 4429 158332
rect 4365 158272 4429 158276
rect 4445 158332 4509 158336
rect 4445 158276 4449 158332
rect 4449 158276 4505 158332
rect 4505 158276 4509 158332
rect 4445 158272 4509 158276
rect 4525 158332 4589 158336
rect 4525 158276 4529 158332
rect 4529 158276 4585 158332
rect 4585 158276 4589 158332
rect 4525 158272 4589 158276
rect 7618 158332 7682 158336
rect 7618 158276 7622 158332
rect 7622 158276 7678 158332
rect 7678 158276 7682 158332
rect 7618 158272 7682 158276
rect 7698 158332 7762 158336
rect 7698 158276 7702 158332
rect 7702 158276 7758 158332
rect 7758 158276 7762 158332
rect 7698 158272 7762 158276
rect 7778 158332 7842 158336
rect 7778 158276 7782 158332
rect 7782 158276 7838 158332
rect 7838 158276 7842 158332
rect 7778 158272 7842 158276
rect 7858 158332 7922 158336
rect 7858 158276 7862 158332
rect 7862 158276 7918 158332
rect 7918 158276 7922 158332
rect 7858 158272 7922 158276
rect 2618 157788 2682 157792
rect 2618 157732 2622 157788
rect 2622 157732 2678 157788
rect 2678 157732 2682 157788
rect 2618 157728 2682 157732
rect 2698 157788 2762 157792
rect 2698 157732 2702 157788
rect 2702 157732 2758 157788
rect 2758 157732 2762 157788
rect 2698 157728 2762 157732
rect 2778 157788 2842 157792
rect 2778 157732 2782 157788
rect 2782 157732 2838 157788
rect 2838 157732 2842 157788
rect 2778 157728 2842 157732
rect 2858 157788 2922 157792
rect 2858 157732 2862 157788
rect 2862 157732 2918 157788
rect 2918 157732 2922 157788
rect 2858 157728 2922 157732
rect 5952 157788 6016 157792
rect 5952 157732 5956 157788
rect 5956 157732 6012 157788
rect 6012 157732 6016 157788
rect 5952 157728 6016 157732
rect 6032 157788 6096 157792
rect 6032 157732 6036 157788
rect 6036 157732 6092 157788
rect 6092 157732 6096 157788
rect 6032 157728 6096 157732
rect 6112 157788 6176 157792
rect 6112 157732 6116 157788
rect 6116 157732 6172 157788
rect 6172 157732 6176 157788
rect 6112 157728 6176 157732
rect 6192 157788 6256 157792
rect 6192 157732 6196 157788
rect 6196 157732 6252 157788
rect 6252 157732 6256 157788
rect 6192 157728 6256 157732
rect 4285 157244 4349 157248
rect 4285 157188 4289 157244
rect 4289 157188 4345 157244
rect 4345 157188 4349 157244
rect 4285 157184 4349 157188
rect 4365 157244 4429 157248
rect 4365 157188 4369 157244
rect 4369 157188 4425 157244
rect 4425 157188 4429 157244
rect 4365 157184 4429 157188
rect 4445 157244 4509 157248
rect 4445 157188 4449 157244
rect 4449 157188 4505 157244
rect 4505 157188 4509 157244
rect 4445 157184 4509 157188
rect 4525 157244 4589 157248
rect 4525 157188 4529 157244
rect 4529 157188 4585 157244
rect 4585 157188 4589 157244
rect 4525 157184 4589 157188
rect 7618 157244 7682 157248
rect 7618 157188 7622 157244
rect 7622 157188 7678 157244
rect 7678 157188 7682 157244
rect 7618 157184 7682 157188
rect 7698 157244 7762 157248
rect 7698 157188 7702 157244
rect 7702 157188 7758 157244
rect 7758 157188 7762 157244
rect 7698 157184 7762 157188
rect 7778 157244 7842 157248
rect 7778 157188 7782 157244
rect 7782 157188 7838 157244
rect 7838 157188 7842 157244
rect 7778 157184 7842 157188
rect 7858 157244 7922 157248
rect 7858 157188 7862 157244
rect 7862 157188 7918 157244
rect 7918 157188 7922 157244
rect 7858 157184 7922 157188
rect 2618 156700 2682 156704
rect 2618 156644 2622 156700
rect 2622 156644 2678 156700
rect 2678 156644 2682 156700
rect 2618 156640 2682 156644
rect 2698 156700 2762 156704
rect 2698 156644 2702 156700
rect 2702 156644 2758 156700
rect 2758 156644 2762 156700
rect 2698 156640 2762 156644
rect 2778 156700 2842 156704
rect 2778 156644 2782 156700
rect 2782 156644 2838 156700
rect 2838 156644 2842 156700
rect 2778 156640 2842 156644
rect 2858 156700 2922 156704
rect 2858 156644 2862 156700
rect 2862 156644 2918 156700
rect 2918 156644 2922 156700
rect 2858 156640 2922 156644
rect 5952 156700 6016 156704
rect 5952 156644 5956 156700
rect 5956 156644 6012 156700
rect 6012 156644 6016 156700
rect 5952 156640 6016 156644
rect 6032 156700 6096 156704
rect 6032 156644 6036 156700
rect 6036 156644 6092 156700
rect 6092 156644 6096 156700
rect 6032 156640 6096 156644
rect 6112 156700 6176 156704
rect 6112 156644 6116 156700
rect 6116 156644 6172 156700
rect 6172 156644 6176 156700
rect 6112 156640 6176 156644
rect 6192 156700 6256 156704
rect 6192 156644 6196 156700
rect 6196 156644 6252 156700
rect 6252 156644 6256 156700
rect 6192 156640 6256 156644
rect 4285 156156 4349 156160
rect 4285 156100 4289 156156
rect 4289 156100 4345 156156
rect 4345 156100 4349 156156
rect 4285 156096 4349 156100
rect 4365 156156 4429 156160
rect 4365 156100 4369 156156
rect 4369 156100 4425 156156
rect 4425 156100 4429 156156
rect 4365 156096 4429 156100
rect 4445 156156 4509 156160
rect 4445 156100 4449 156156
rect 4449 156100 4505 156156
rect 4505 156100 4509 156156
rect 4445 156096 4509 156100
rect 4525 156156 4589 156160
rect 4525 156100 4529 156156
rect 4529 156100 4585 156156
rect 4585 156100 4589 156156
rect 4525 156096 4589 156100
rect 7618 156156 7682 156160
rect 7618 156100 7622 156156
rect 7622 156100 7678 156156
rect 7678 156100 7682 156156
rect 7618 156096 7682 156100
rect 7698 156156 7762 156160
rect 7698 156100 7702 156156
rect 7702 156100 7758 156156
rect 7758 156100 7762 156156
rect 7698 156096 7762 156100
rect 7778 156156 7842 156160
rect 7778 156100 7782 156156
rect 7782 156100 7838 156156
rect 7838 156100 7842 156156
rect 7778 156096 7842 156100
rect 7858 156156 7922 156160
rect 7858 156100 7862 156156
rect 7862 156100 7918 156156
rect 7918 156100 7922 156156
rect 7858 156096 7922 156100
rect 2618 155612 2682 155616
rect 2618 155556 2622 155612
rect 2622 155556 2678 155612
rect 2678 155556 2682 155612
rect 2618 155552 2682 155556
rect 2698 155612 2762 155616
rect 2698 155556 2702 155612
rect 2702 155556 2758 155612
rect 2758 155556 2762 155612
rect 2698 155552 2762 155556
rect 2778 155612 2842 155616
rect 2778 155556 2782 155612
rect 2782 155556 2838 155612
rect 2838 155556 2842 155612
rect 2778 155552 2842 155556
rect 2858 155612 2922 155616
rect 2858 155556 2862 155612
rect 2862 155556 2918 155612
rect 2918 155556 2922 155612
rect 2858 155552 2922 155556
rect 5952 155612 6016 155616
rect 5952 155556 5956 155612
rect 5956 155556 6012 155612
rect 6012 155556 6016 155612
rect 5952 155552 6016 155556
rect 6032 155612 6096 155616
rect 6032 155556 6036 155612
rect 6036 155556 6092 155612
rect 6092 155556 6096 155612
rect 6032 155552 6096 155556
rect 6112 155612 6176 155616
rect 6112 155556 6116 155612
rect 6116 155556 6172 155612
rect 6172 155556 6176 155612
rect 6112 155552 6176 155556
rect 6192 155612 6256 155616
rect 6192 155556 6196 155612
rect 6196 155556 6252 155612
rect 6252 155556 6256 155612
rect 6192 155552 6256 155556
rect 4285 155068 4349 155072
rect 4285 155012 4289 155068
rect 4289 155012 4345 155068
rect 4345 155012 4349 155068
rect 4285 155008 4349 155012
rect 4365 155068 4429 155072
rect 4365 155012 4369 155068
rect 4369 155012 4425 155068
rect 4425 155012 4429 155068
rect 4365 155008 4429 155012
rect 4445 155068 4509 155072
rect 4445 155012 4449 155068
rect 4449 155012 4505 155068
rect 4505 155012 4509 155068
rect 4445 155008 4509 155012
rect 4525 155068 4589 155072
rect 4525 155012 4529 155068
rect 4529 155012 4585 155068
rect 4585 155012 4589 155068
rect 4525 155008 4589 155012
rect 7618 155068 7682 155072
rect 7618 155012 7622 155068
rect 7622 155012 7678 155068
rect 7678 155012 7682 155068
rect 7618 155008 7682 155012
rect 7698 155068 7762 155072
rect 7698 155012 7702 155068
rect 7702 155012 7758 155068
rect 7758 155012 7762 155068
rect 7698 155008 7762 155012
rect 7778 155068 7842 155072
rect 7778 155012 7782 155068
rect 7782 155012 7838 155068
rect 7838 155012 7842 155068
rect 7778 155008 7842 155012
rect 7858 155068 7922 155072
rect 7858 155012 7862 155068
rect 7862 155012 7918 155068
rect 7918 155012 7922 155068
rect 7858 155008 7922 155012
rect 2618 154524 2682 154528
rect 2618 154468 2622 154524
rect 2622 154468 2678 154524
rect 2678 154468 2682 154524
rect 2618 154464 2682 154468
rect 2698 154524 2762 154528
rect 2698 154468 2702 154524
rect 2702 154468 2758 154524
rect 2758 154468 2762 154524
rect 2698 154464 2762 154468
rect 2778 154524 2842 154528
rect 2778 154468 2782 154524
rect 2782 154468 2838 154524
rect 2838 154468 2842 154524
rect 2778 154464 2842 154468
rect 2858 154524 2922 154528
rect 2858 154468 2862 154524
rect 2862 154468 2918 154524
rect 2918 154468 2922 154524
rect 2858 154464 2922 154468
rect 5952 154524 6016 154528
rect 5952 154468 5956 154524
rect 5956 154468 6012 154524
rect 6012 154468 6016 154524
rect 5952 154464 6016 154468
rect 6032 154524 6096 154528
rect 6032 154468 6036 154524
rect 6036 154468 6092 154524
rect 6092 154468 6096 154524
rect 6032 154464 6096 154468
rect 6112 154524 6176 154528
rect 6112 154468 6116 154524
rect 6116 154468 6172 154524
rect 6172 154468 6176 154524
rect 6112 154464 6176 154468
rect 6192 154524 6256 154528
rect 6192 154468 6196 154524
rect 6196 154468 6252 154524
rect 6252 154468 6256 154524
rect 6192 154464 6256 154468
rect 4285 153980 4349 153984
rect 4285 153924 4289 153980
rect 4289 153924 4345 153980
rect 4345 153924 4349 153980
rect 4285 153920 4349 153924
rect 4365 153980 4429 153984
rect 4365 153924 4369 153980
rect 4369 153924 4425 153980
rect 4425 153924 4429 153980
rect 4365 153920 4429 153924
rect 4445 153980 4509 153984
rect 4445 153924 4449 153980
rect 4449 153924 4505 153980
rect 4505 153924 4509 153980
rect 4445 153920 4509 153924
rect 4525 153980 4589 153984
rect 4525 153924 4529 153980
rect 4529 153924 4585 153980
rect 4585 153924 4589 153980
rect 4525 153920 4589 153924
rect 7618 153980 7682 153984
rect 7618 153924 7622 153980
rect 7622 153924 7678 153980
rect 7678 153924 7682 153980
rect 7618 153920 7682 153924
rect 7698 153980 7762 153984
rect 7698 153924 7702 153980
rect 7702 153924 7758 153980
rect 7758 153924 7762 153980
rect 7698 153920 7762 153924
rect 7778 153980 7842 153984
rect 7778 153924 7782 153980
rect 7782 153924 7838 153980
rect 7838 153924 7842 153980
rect 7778 153920 7842 153924
rect 7858 153980 7922 153984
rect 7858 153924 7862 153980
rect 7862 153924 7918 153980
rect 7918 153924 7922 153980
rect 7858 153920 7922 153924
rect 2618 153436 2682 153440
rect 2618 153380 2622 153436
rect 2622 153380 2678 153436
rect 2678 153380 2682 153436
rect 2618 153376 2682 153380
rect 2698 153436 2762 153440
rect 2698 153380 2702 153436
rect 2702 153380 2758 153436
rect 2758 153380 2762 153436
rect 2698 153376 2762 153380
rect 2778 153436 2842 153440
rect 2778 153380 2782 153436
rect 2782 153380 2838 153436
rect 2838 153380 2842 153436
rect 2778 153376 2842 153380
rect 2858 153436 2922 153440
rect 2858 153380 2862 153436
rect 2862 153380 2918 153436
rect 2918 153380 2922 153436
rect 2858 153376 2922 153380
rect 5952 153436 6016 153440
rect 5952 153380 5956 153436
rect 5956 153380 6012 153436
rect 6012 153380 6016 153436
rect 5952 153376 6016 153380
rect 6032 153436 6096 153440
rect 6032 153380 6036 153436
rect 6036 153380 6092 153436
rect 6092 153380 6096 153436
rect 6032 153376 6096 153380
rect 6112 153436 6176 153440
rect 6112 153380 6116 153436
rect 6116 153380 6172 153436
rect 6172 153380 6176 153436
rect 6112 153376 6176 153380
rect 6192 153436 6256 153440
rect 6192 153380 6196 153436
rect 6196 153380 6252 153436
rect 6252 153380 6256 153436
rect 6192 153376 6256 153380
rect 4285 152892 4349 152896
rect 4285 152836 4289 152892
rect 4289 152836 4345 152892
rect 4345 152836 4349 152892
rect 4285 152832 4349 152836
rect 4365 152892 4429 152896
rect 4365 152836 4369 152892
rect 4369 152836 4425 152892
rect 4425 152836 4429 152892
rect 4365 152832 4429 152836
rect 4445 152892 4509 152896
rect 4445 152836 4449 152892
rect 4449 152836 4505 152892
rect 4505 152836 4509 152892
rect 4445 152832 4509 152836
rect 4525 152892 4589 152896
rect 4525 152836 4529 152892
rect 4529 152836 4585 152892
rect 4585 152836 4589 152892
rect 4525 152832 4589 152836
rect 7618 152892 7682 152896
rect 7618 152836 7622 152892
rect 7622 152836 7678 152892
rect 7678 152836 7682 152892
rect 7618 152832 7682 152836
rect 7698 152892 7762 152896
rect 7698 152836 7702 152892
rect 7702 152836 7758 152892
rect 7758 152836 7762 152892
rect 7698 152832 7762 152836
rect 7778 152892 7842 152896
rect 7778 152836 7782 152892
rect 7782 152836 7838 152892
rect 7838 152836 7842 152892
rect 7778 152832 7842 152836
rect 7858 152892 7922 152896
rect 7858 152836 7862 152892
rect 7862 152836 7918 152892
rect 7918 152836 7922 152892
rect 7858 152832 7922 152836
rect 2618 152348 2682 152352
rect 2618 152292 2622 152348
rect 2622 152292 2678 152348
rect 2678 152292 2682 152348
rect 2618 152288 2682 152292
rect 2698 152348 2762 152352
rect 2698 152292 2702 152348
rect 2702 152292 2758 152348
rect 2758 152292 2762 152348
rect 2698 152288 2762 152292
rect 2778 152348 2842 152352
rect 2778 152292 2782 152348
rect 2782 152292 2838 152348
rect 2838 152292 2842 152348
rect 2778 152288 2842 152292
rect 2858 152348 2922 152352
rect 2858 152292 2862 152348
rect 2862 152292 2918 152348
rect 2918 152292 2922 152348
rect 2858 152288 2922 152292
rect 5952 152348 6016 152352
rect 5952 152292 5956 152348
rect 5956 152292 6012 152348
rect 6012 152292 6016 152348
rect 5952 152288 6016 152292
rect 6032 152348 6096 152352
rect 6032 152292 6036 152348
rect 6036 152292 6092 152348
rect 6092 152292 6096 152348
rect 6032 152288 6096 152292
rect 6112 152348 6176 152352
rect 6112 152292 6116 152348
rect 6116 152292 6172 152348
rect 6172 152292 6176 152348
rect 6112 152288 6176 152292
rect 6192 152348 6256 152352
rect 6192 152292 6196 152348
rect 6196 152292 6252 152348
rect 6252 152292 6256 152348
rect 6192 152288 6256 152292
rect 4285 151804 4349 151808
rect 4285 151748 4289 151804
rect 4289 151748 4345 151804
rect 4345 151748 4349 151804
rect 4285 151744 4349 151748
rect 4365 151804 4429 151808
rect 4365 151748 4369 151804
rect 4369 151748 4425 151804
rect 4425 151748 4429 151804
rect 4365 151744 4429 151748
rect 4445 151804 4509 151808
rect 4445 151748 4449 151804
rect 4449 151748 4505 151804
rect 4505 151748 4509 151804
rect 4445 151744 4509 151748
rect 4525 151804 4589 151808
rect 4525 151748 4529 151804
rect 4529 151748 4585 151804
rect 4585 151748 4589 151804
rect 4525 151744 4589 151748
rect 7618 151804 7682 151808
rect 7618 151748 7622 151804
rect 7622 151748 7678 151804
rect 7678 151748 7682 151804
rect 7618 151744 7682 151748
rect 7698 151804 7762 151808
rect 7698 151748 7702 151804
rect 7702 151748 7758 151804
rect 7758 151748 7762 151804
rect 7698 151744 7762 151748
rect 7778 151804 7842 151808
rect 7778 151748 7782 151804
rect 7782 151748 7838 151804
rect 7838 151748 7842 151804
rect 7778 151744 7842 151748
rect 7858 151804 7922 151808
rect 7858 151748 7862 151804
rect 7862 151748 7918 151804
rect 7918 151748 7922 151804
rect 7858 151744 7922 151748
rect 2618 151260 2682 151264
rect 2618 151204 2622 151260
rect 2622 151204 2678 151260
rect 2678 151204 2682 151260
rect 2618 151200 2682 151204
rect 2698 151260 2762 151264
rect 2698 151204 2702 151260
rect 2702 151204 2758 151260
rect 2758 151204 2762 151260
rect 2698 151200 2762 151204
rect 2778 151260 2842 151264
rect 2778 151204 2782 151260
rect 2782 151204 2838 151260
rect 2838 151204 2842 151260
rect 2778 151200 2842 151204
rect 2858 151260 2922 151264
rect 2858 151204 2862 151260
rect 2862 151204 2918 151260
rect 2918 151204 2922 151260
rect 2858 151200 2922 151204
rect 5952 151260 6016 151264
rect 5952 151204 5956 151260
rect 5956 151204 6012 151260
rect 6012 151204 6016 151260
rect 5952 151200 6016 151204
rect 6032 151260 6096 151264
rect 6032 151204 6036 151260
rect 6036 151204 6092 151260
rect 6092 151204 6096 151260
rect 6032 151200 6096 151204
rect 6112 151260 6176 151264
rect 6112 151204 6116 151260
rect 6116 151204 6172 151260
rect 6172 151204 6176 151260
rect 6112 151200 6176 151204
rect 6192 151260 6256 151264
rect 6192 151204 6196 151260
rect 6196 151204 6252 151260
rect 6252 151204 6256 151260
rect 6192 151200 6256 151204
rect 4285 150716 4349 150720
rect 4285 150660 4289 150716
rect 4289 150660 4345 150716
rect 4345 150660 4349 150716
rect 4285 150656 4349 150660
rect 4365 150716 4429 150720
rect 4365 150660 4369 150716
rect 4369 150660 4425 150716
rect 4425 150660 4429 150716
rect 4365 150656 4429 150660
rect 4445 150716 4509 150720
rect 4445 150660 4449 150716
rect 4449 150660 4505 150716
rect 4505 150660 4509 150716
rect 4445 150656 4509 150660
rect 4525 150716 4589 150720
rect 4525 150660 4529 150716
rect 4529 150660 4585 150716
rect 4585 150660 4589 150716
rect 4525 150656 4589 150660
rect 7618 150716 7682 150720
rect 7618 150660 7622 150716
rect 7622 150660 7678 150716
rect 7678 150660 7682 150716
rect 7618 150656 7682 150660
rect 7698 150716 7762 150720
rect 7698 150660 7702 150716
rect 7702 150660 7758 150716
rect 7758 150660 7762 150716
rect 7698 150656 7762 150660
rect 7778 150716 7842 150720
rect 7778 150660 7782 150716
rect 7782 150660 7838 150716
rect 7838 150660 7842 150716
rect 7778 150656 7842 150660
rect 7858 150716 7922 150720
rect 7858 150660 7862 150716
rect 7862 150660 7918 150716
rect 7918 150660 7922 150716
rect 7858 150656 7922 150660
rect 2618 150172 2682 150176
rect 2618 150116 2622 150172
rect 2622 150116 2678 150172
rect 2678 150116 2682 150172
rect 2618 150112 2682 150116
rect 2698 150172 2762 150176
rect 2698 150116 2702 150172
rect 2702 150116 2758 150172
rect 2758 150116 2762 150172
rect 2698 150112 2762 150116
rect 2778 150172 2842 150176
rect 2778 150116 2782 150172
rect 2782 150116 2838 150172
rect 2838 150116 2842 150172
rect 2778 150112 2842 150116
rect 2858 150172 2922 150176
rect 2858 150116 2862 150172
rect 2862 150116 2918 150172
rect 2918 150116 2922 150172
rect 2858 150112 2922 150116
rect 5952 150172 6016 150176
rect 5952 150116 5956 150172
rect 5956 150116 6012 150172
rect 6012 150116 6016 150172
rect 5952 150112 6016 150116
rect 6032 150172 6096 150176
rect 6032 150116 6036 150172
rect 6036 150116 6092 150172
rect 6092 150116 6096 150172
rect 6032 150112 6096 150116
rect 6112 150172 6176 150176
rect 6112 150116 6116 150172
rect 6116 150116 6172 150172
rect 6172 150116 6176 150172
rect 6112 150112 6176 150116
rect 6192 150172 6256 150176
rect 6192 150116 6196 150172
rect 6196 150116 6252 150172
rect 6252 150116 6256 150172
rect 6192 150112 6256 150116
rect 4285 149628 4349 149632
rect 4285 149572 4289 149628
rect 4289 149572 4345 149628
rect 4345 149572 4349 149628
rect 4285 149568 4349 149572
rect 4365 149628 4429 149632
rect 4365 149572 4369 149628
rect 4369 149572 4425 149628
rect 4425 149572 4429 149628
rect 4365 149568 4429 149572
rect 4445 149628 4509 149632
rect 4445 149572 4449 149628
rect 4449 149572 4505 149628
rect 4505 149572 4509 149628
rect 4445 149568 4509 149572
rect 4525 149628 4589 149632
rect 4525 149572 4529 149628
rect 4529 149572 4585 149628
rect 4585 149572 4589 149628
rect 4525 149568 4589 149572
rect 7618 149628 7682 149632
rect 7618 149572 7622 149628
rect 7622 149572 7678 149628
rect 7678 149572 7682 149628
rect 7618 149568 7682 149572
rect 7698 149628 7762 149632
rect 7698 149572 7702 149628
rect 7702 149572 7758 149628
rect 7758 149572 7762 149628
rect 7698 149568 7762 149572
rect 7778 149628 7842 149632
rect 7778 149572 7782 149628
rect 7782 149572 7838 149628
rect 7838 149572 7842 149628
rect 7778 149568 7842 149572
rect 7858 149628 7922 149632
rect 7858 149572 7862 149628
rect 7862 149572 7918 149628
rect 7918 149572 7922 149628
rect 7858 149568 7922 149572
rect 2618 149084 2682 149088
rect 2618 149028 2622 149084
rect 2622 149028 2678 149084
rect 2678 149028 2682 149084
rect 2618 149024 2682 149028
rect 2698 149084 2762 149088
rect 2698 149028 2702 149084
rect 2702 149028 2758 149084
rect 2758 149028 2762 149084
rect 2698 149024 2762 149028
rect 2778 149084 2842 149088
rect 2778 149028 2782 149084
rect 2782 149028 2838 149084
rect 2838 149028 2842 149084
rect 2778 149024 2842 149028
rect 2858 149084 2922 149088
rect 2858 149028 2862 149084
rect 2862 149028 2918 149084
rect 2918 149028 2922 149084
rect 2858 149024 2922 149028
rect 5952 149084 6016 149088
rect 5952 149028 5956 149084
rect 5956 149028 6012 149084
rect 6012 149028 6016 149084
rect 5952 149024 6016 149028
rect 6032 149084 6096 149088
rect 6032 149028 6036 149084
rect 6036 149028 6092 149084
rect 6092 149028 6096 149084
rect 6032 149024 6096 149028
rect 6112 149084 6176 149088
rect 6112 149028 6116 149084
rect 6116 149028 6172 149084
rect 6172 149028 6176 149084
rect 6112 149024 6176 149028
rect 6192 149084 6256 149088
rect 6192 149028 6196 149084
rect 6196 149028 6252 149084
rect 6252 149028 6256 149084
rect 6192 149024 6256 149028
rect 4285 148540 4349 148544
rect 4285 148484 4289 148540
rect 4289 148484 4345 148540
rect 4345 148484 4349 148540
rect 4285 148480 4349 148484
rect 4365 148540 4429 148544
rect 4365 148484 4369 148540
rect 4369 148484 4425 148540
rect 4425 148484 4429 148540
rect 4365 148480 4429 148484
rect 4445 148540 4509 148544
rect 4445 148484 4449 148540
rect 4449 148484 4505 148540
rect 4505 148484 4509 148540
rect 4445 148480 4509 148484
rect 4525 148540 4589 148544
rect 4525 148484 4529 148540
rect 4529 148484 4585 148540
rect 4585 148484 4589 148540
rect 4525 148480 4589 148484
rect 7618 148540 7682 148544
rect 7618 148484 7622 148540
rect 7622 148484 7678 148540
rect 7678 148484 7682 148540
rect 7618 148480 7682 148484
rect 7698 148540 7762 148544
rect 7698 148484 7702 148540
rect 7702 148484 7758 148540
rect 7758 148484 7762 148540
rect 7698 148480 7762 148484
rect 7778 148540 7842 148544
rect 7778 148484 7782 148540
rect 7782 148484 7838 148540
rect 7838 148484 7842 148540
rect 7778 148480 7842 148484
rect 7858 148540 7922 148544
rect 7858 148484 7862 148540
rect 7862 148484 7918 148540
rect 7918 148484 7922 148540
rect 7858 148480 7922 148484
rect 2618 147996 2682 148000
rect 2618 147940 2622 147996
rect 2622 147940 2678 147996
rect 2678 147940 2682 147996
rect 2618 147936 2682 147940
rect 2698 147996 2762 148000
rect 2698 147940 2702 147996
rect 2702 147940 2758 147996
rect 2758 147940 2762 147996
rect 2698 147936 2762 147940
rect 2778 147996 2842 148000
rect 2778 147940 2782 147996
rect 2782 147940 2838 147996
rect 2838 147940 2842 147996
rect 2778 147936 2842 147940
rect 2858 147996 2922 148000
rect 2858 147940 2862 147996
rect 2862 147940 2918 147996
rect 2918 147940 2922 147996
rect 2858 147936 2922 147940
rect 5952 147996 6016 148000
rect 5952 147940 5956 147996
rect 5956 147940 6012 147996
rect 6012 147940 6016 147996
rect 5952 147936 6016 147940
rect 6032 147996 6096 148000
rect 6032 147940 6036 147996
rect 6036 147940 6092 147996
rect 6092 147940 6096 147996
rect 6032 147936 6096 147940
rect 6112 147996 6176 148000
rect 6112 147940 6116 147996
rect 6116 147940 6172 147996
rect 6172 147940 6176 147996
rect 6112 147936 6176 147940
rect 6192 147996 6256 148000
rect 6192 147940 6196 147996
rect 6196 147940 6252 147996
rect 6252 147940 6256 147996
rect 6192 147936 6256 147940
rect 4285 147452 4349 147456
rect 4285 147396 4289 147452
rect 4289 147396 4345 147452
rect 4345 147396 4349 147452
rect 4285 147392 4349 147396
rect 4365 147452 4429 147456
rect 4365 147396 4369 147452
rect 4369 147396 4425 147452
rect 4425 147396 4429 147452
rect 4365 147392 4429 147396
rect 4445 147452 4509 147456
rect 4445 147396 4449 147452
rect 4449 147396 4505 147452
rect 4505 147396 4509 147452
rect 4445 147392 4509 147396
rect 4525 147452 4589 147456
rect 4525 147396 4529 147452
rect 4529 147396 4585 147452
rect 4585 147396 4589 147452
rect 4525 147392 4589 147396
rect 7618 147452 7682 147456
rect 7618 147396 7622 147452
rect 7622 147396 7678 147452
rect 7678 147396 7682 147452
rect 7618 147392 7682 147396
rect 7698 147452 7762 147456
rect 7698 147396 7702 147452
rect 7702 147396 7758 147452
rect 7758 147396 7762 147452
rect 7698 147392 7762 147396
rect 7778 147452 7842 147456
rect 7778 147396 7782 147452
rect 7782 147396 7838 147452
rect 7838 147396 7842 147452
rect 7778 147392 7842 147396
rect 7858 147452 7922 147456
rect 7858 147396 7862 147452
rect 7862 147396 7918 147452
rect 7918 147396 7922 147452
rect 7858 147392 7922 147396
rect 2618 146908 2682 146912
rect 2618 146852 2622 146908
rect 2622 146852 2678 146908
rect 2678 146852 2682 146908
rect 2618 146848 2682 146852
rect 2698 146908 2762 146912
rect 2698 146852 2702 146908
rect 2702 146852 2758 146908
rect 2758 146852 2762 146908
rect 2698 146848 2762 146852
rect 2778 146908 2842 146912
rect 2778 146852 2782 146908
rect 2782 146852 2838 146908
rect 2838 146852 2842 146908
rect 2778 146848 2842 146852
rect 2858 146908 2922 146912
rect 2858 146852 2862 146908
rect 2862 146852 2918 146908
rect 2918 146852 2922 146908
rect 2858 146848 2922 146852
rect 5952 146908 6016 146912
rect 5952 146852 5956 146908
rect 5956 146852 6012 146908
rect 6012 146852 6016 146908
rect 5952 146848 6016 146852
rect 6032 146908 6096 146912
rect 6032 146852 6036 146908
rect 6036 146852 6092 146908
rect 6092 146852 6096 146908
rect 6032 146848 6096 146852
rect 6112 146908 6176 146912
rect 6112 146852 6116 146908
rect 6116 146852 6172 146908
rect 6172 146852 6176 146908
rect 6112 146848 6176 146852
rect 6192 146908 6256 146912
rect 6192 146852 6196 146908
rect 6196 146852 6252 146908
rect 6252 146852 6256 146908
rect 6192 146848 6256 146852
rect 4285 146364 4349 146368
rect 4285 146308 4289 146364
rect 4289 146308 4345 146364
rect 4345 146308 4349 146364
rect 4285 146304 4349 146308
rect 4365 146364 4429 146368
rect 4365 146308 4369 146364
rect 4369 146308 4425 146364
rect 4425 146308 4429 146364
rect 4365 146304 4429 146308
rect 4445 146364 4509 146368
rect 4445 146308 4449 146364
rect 4449 146308 4505 146364
rect 4505 146308 4509 146364
rect 4445 146304 4509 146308
rect 4525 146364 4589 146368
rect 4525 146308 4529 146364
rect 4529 146308 4585 146364
rect 4585 146308 4589 146364
rect 4525 146304 4589 146308
rect 7618 146364 7682 146368
rect 7618 146308 7622 146364
rect 7622 146308 7678 146364
rect 7678 146308 7682 146364
rect 7618 146304 7682 146308
rect 7698 146364 7762 146368
rect 7698 146308 7702 146364
rect 7702 146308 7758 146364
rect 7758 146308 7762 146364
rect 7698 146304 7762 146308
rect 7778 146364 7842 146368
rect 7778 146308 7782 146364
rect 7782 146308 7838 146364
rect 7838 146308 7842 146364
rect 7778 146304 7842 146308
rect 7858 146364 7922 146368
rect 7858 146308 7862 146364
rect 7862 146308 7918 146364
rect 7918 146308 7922 146364
rect 7858 146304 7922 146308
rect 2618 145820 2682 145824
rect 2618 145764 2622 145820
rect 2622 145764 2678 145820
rect 2678 145764 2682 145820
rect 2618 145760 2682 145764
rect 2698 145820 2762 145824
rect 2698 145764 2702 145820
rect 2702 145764 2758 145820
rect 2758 145764 2762 145820
rect 2698 145760 2762 145764
rect 2778 145820 2842 145824
rect 2778 145764 2782 145820
rect 2782 145764 2838 145820
rect 2838 145764 2842 145820
rect 2778 145760 2842 145764
rect 2858 145820 2922 145824
rect 2858 145764 2862 145820
rect 2862 145764 2918 145820
rect 2918 145764 2922 145820
rect 2858 145760 2922 145764
rect 5952 145820 6016 145824
rect 5952 145764 5956 145820
rect 5956 145764 6012 145820
rect 6012 145764 6016 145820
rect 5952 145760 6016 145764
rect 6032 145820 6096 145824
rect 6032 145764 6036 145820
rect 6036 145764 6092 145820
rect 6092 145764 6096 145820
rect 6032 145760 6096 145764
rect 6112 145820 6176 145824
rect 6112 145764 6116 145820
rect 6116 145764 6172 145820
rect 6172 145764 6176 145820
rect 6112 145760 6176 145764
rect 6192 145820 6256 145824
rect 6192 145764 6196 145820
rect 6196 145764 6252 145820
rect 6252 145764 6256 145820
rect 6192 145760 6256 145764
rect 4285 145276 4349 145280
rect 4285 145220 4289 145276
rect 4289 145220 4345 145276
rect 4345 145220 4349 145276
rect 4285 145216 4349 145220
rect 4365 145276 4429 145280
rect 4365 145220 4369 145276
rect 4369 145220 4425 145276
rect 4425 145220 4429 145276
rect 4365 145216 4429 145220
rect 4445 145276 4509 145280
rect 4445 145220 4449 145276
rect 4449 145220 4505 145276
rect 4505 145220 4509 145276
rect 4445 145216 4509 145220
rect 4525 145276 4589 145280
rect 4525 145220 4529 145276
rect 4529 145220 4585 145276
rect 4585 145220 4589 145276
rect 4525 145216 4589 145220
rect 7618 145276 7682 145280
rect 7618 145220 7622 145276
rect 7622 145220 7678 145276
rect 7678 145220 7682 145276
rect 7618 145216 7682 145220
rect 7698 145276 7762 145280
rect 7698 145220 7702 145276
rect 7702 145220 7758 145276
rect 7758 145220 7762 145276
rect 7698 145216 7762 145220
rect 7778 145276 7842 145280
rect 7778 145220 7782 145276
rect 7782 145220 7838 145276
rect 7838 145220 7842 145276
rect 7778 145216 7842 145220
rect 7858 145276 7922 145280
rect 7858 145220 7862 145276
rect 7862 145220 7918 145276
rect 7918 145220 7922 145276
rect 7858 145216 7922 145220
rect 2618 144732 2682 144736
rect 2618 144676 2622 144732
rect 2622 144676 2678 144732
rect 2678 144676 2682 144732
rect 2618 144672 2682 144676
rect 2698 144732 2762 144736
rect 2698 144676 2702 144732
rect 2702 144676 2758 144732
rect 2758 144676 2762 144732
rect 2698 144672 2762 144676
rect 2778 144732 2842 144736
rect 2778 144676 2782 144732
rect 2782 144676 2838 144732
rect 2838 144676 2842 144732
rect 2778 144672 2842 144676
rect 2858 144732 2922 144736
rect 2858 144676 2862 144732
rect 2862 144676 2918 144732
rect 2918 144676 2922 144732
rect 2858 144672 2922 144676
rect 5952 144732 6016 144736
rect 5952 144676 5956 144732
rect 5956 144676 6012 144732
rect 6012 144676 6016 144732
rect 5952 144672 6016 144676
rect 6032 144732 6096 144736
rect 6032 144676 6036 144732
rect 6036 144676 6092 144732
rect 6092 144676 6096 144732
rect 6032 144672 6096 144676
rect 6112 144732 6176 144736
rect 6112 144676 6116 144732
rect 6116 144676 6172 144732
rect 6172 144676 6176 144732
rect 6112 144672 6176 144676
rect 6192 144732 6256 144736
rect 6192 144676 6196 144732
rect 6196 144676 6252 144732
rect 6252 144676 6256 144732
rect 6192 144672 6256 144676
rect 4285 144188 4349 144192
rect 4285 144132 4289 144188
rect 4289 144132 4345 144188
rect 4345 144132 4349 144188
rect 4285 144128 4349 144132
rect 4365 144188 4429 144192
rect 4365 144132 4369 144188
rect 4369 144132 4425 144188
rect 4425 144132 4429 144188
rect 4365 144128 4429 144132
rect 4445 144188 4509 144192
rect 4445 144132 4449 144188
rect 4449 144132 4505 144188
rect 4505 144132 4509 144188
rect 4445 144128 4509 144132
rect 4525 144188 4589 144192
rect 4525 144132 4529 144188
rect 4529 144132 4585 144188
rect 4585 144132 4589 144188
rect 4525 144128 4589 144132
rect 7618 144188 7682 144192
rect 7618 144132 7622 144188
rect 7622 144132 7678 144188
rect 7678 144132 7682 144188
rect 7618 144128 7682 144132
rect 7698 144188 7762 144192
rect 7698 144132 7702 144188
rect 7702 144132 7758 144188
rect 7758 144132 7762 144188
rect 7698 144128 7762 144132
rect 7778 144188 7842 144192
rect 7778 144132 7782 144188
rect 7782 144132 7838 144188
rect 7838 144132 7842 144188
rect 7778 144128 7842 144132
rect 7858 144188 7922 144192
rect 7858 144132 7862 144188
rect 7862 144132 7918 144188
rect 7918 144132 7922 144188
rect 7858 144128 7922 144132
rect 2618 143644 2682 143648
rect 2618 143588 2622 143644
rect 2622 143588 2678 143644
rect 2678 143588 2682 143644
rect 2618 143584 2682 143588
rect 2698 143644 2762 143648
rect 2698 143588 2702 143644
rect 2702 143588 2758 143644
rect 2758 143588 2762 143644
rect 2698 143584 2762 143588
rect 2778 143644 2842 143648
rect 2778 143588 2782 143644
rect 2782 143588 2838 143644
rect 2838 143588 2842 143644
rect 2778 143584 2842 143588
rect 2858 143644 2922 143648
rect 2858 143588 2862 143644
rect 2862 143588 2918 143644
rect 2918 143588 2922 143644
rect 2858 143584 2922 143588
rect 5952 143644 6016 143648
rect 5952 143588 5956 143644
rect 5956 143588 6012 143644
rect 6012 143588 6016 143644
rect 5952 143584 6016 143588
rect 6032 143644 6096 143648
rect 6032 143588 6036 143644
rect 6036 143588 6092 143644
rect 6092 143588 6096 143644
rect 6032 143584 6096 143588
rect 6112 143644 6176 143648
rect 6112 143588 6116 143644
rect 6116 143588 6172 143644
rect 6172 143588 6176 143644
rect 6112 143584 6176 143588
rect 6192 143644 6256 143648
rect 6192 143588 6196 143644
rect 6196 143588 6252 143644
rect 6252 143588 6256 143644
rect 6192 143584 6256 143588
rect 4285 143100 4349 143104
rect 4285 143044 4289 143100
rect 4289 143044 4345 143100
rect 4345 143044 4349 143100
rect 4285 143040 4349 143044
rect 4365 143100 4429 143104
rect 4365 143044 4369 143100
rect 4369 143044 4425 143100
rect 4425 143044 4429 143100
rect 4365 143040 4429 143044
rect 4445 143100 4509 143104
rect 4445 143044 4449 143100
rect 4449 143044 4505 143100
rect 4505 143044 4509 143100
rect 4445 143040 4509 143044
rect 4525 143100 4589 143104
rect 4525 143044 4529 143100
rect 4529 143044 4585 143100
rect 4585 143044 4589 143100
rect 4525 143040 4589 143044
rect 7618 143100 7682 143104
rect 7618 143044 7622 143100
rect 7622 143044 7678 143100
rect 7678 143044 7682 143100
rect 7618 143040 7682 143044
rect 7698 143100 7762 143104
rect 7698 143044 7702 143100
rect 7702 143044 7758 143100
rect 7758 143044 7762 143100
rect 7698 143040 7762 143044
rect 7778 143100 7842 143104
rect 7778 143044 7782 143100
rect 7782 143044 7838 143100
rect 7838 143044 7842 143100
rect 7778 143040 7842 143044
rect 7858 143100 7922 143104
rect 7858 143044 7862 143100
rect 7862 143044 7918 143100
rect 7918 143044 7922 143100
rect 7858 143040 7922 143044
rect 2618 142556 2682 142560
rect 2618 142500 2622 142556
rect 2622 142500 2678 142556
rect 2678 142500 2682 142556
rect 2618 142496 2682 142500
rect 2698 142556 2762 142560
rect 2698 142500 2702 142556
rect 2702 142500 2758 142556
rect 2758 142500 2762 142556
rect 2698 142496 2762 142500
rect 2778 142556 2842 142560
rect 2778 142500 2782 142556
rect 2782 142500 2838 142556
rect 2838 142500 2842 142556
rect 2778 142496 2842 142500
rect 2858 142556 2922 142560
rect 2858 142500 2862 142556
rect 2862 142500 2918 142556
rect 2918 142500 2922 142556
rect 2858 142496 2922 142500
rect 5952 142556 6016 142560
rect 5952 142500 5956 142556
rect 5956 142500 6012 142556
rect 6012 142500 6016 142556
rect 5952 142496 6016 142500
rect 6032 142556 6096 142560
rect 6032 142500 6036 142556
rect 6036 142500 6092 142556
rect 6092 142500 6096 142556
rect 6032 142496 6096 142500
rect 6112 142556 6176 142560
rect 6112 142500 6116 142556
rect 6116 142500 6172 142556
rect 6172 142500 6176 142556
rect 6112 142496 6176 142500
rect 6192 142556 6256 142560
rect 6192 142500 6196 142556
rect 6196 142500 6252 142556
rect 6252 142500 6256 142556
rect 6192 142496 6256 142500
rect 4285 142012 4349 142016
rect 4285 141956 4289 142012
rect 4289 141956 4345 142012
rect 4345 141956 4349 142012
rect 4285 141952 4349 141956
rect 4365 142012 4429 142016
rect 4365 141956 4369 142012
rect 4369 141956 4425 142012
rect 4425 141956 4429 142012
rect 4365 141952 4429 141956
rect 4445 142012 4509 142016
rect 4445 141956 4449 142012
rect 4449 141956 4505 142012
rect 4505 141956 4509 142012
rect 4445 141952 4509 141956
rect 4525 142012 4589 142016
rect 4525 141956 4529 142012
rect 4529 141956 4585 142012
rect 4585 141956 4589 142012
rect 4525 141952 4589 141956
rect 7618 142012 7682 142016
rect 7618 141956 7622 142012
rect 7622 141956 7678 142012
rect 7678 141956 7682 142012
rect 7618 141952 7682 141956
rect 7698 142012 7762 142016
rect 7698 141956 7702 142012
rect 7702 141956 7758 142012
rect 7758 141956 7762 142012
rect 7698 141952 7762 141956
rect 7778 142012 7842 142016
rect 7778 141956 7782 142012
rect 7782 141956 7838 142012
rect 7838 141956 7842 142012
rect 7778 141952 7842 141956
rect 7858 142012 7922 142016
rect 7858 141956 7862 142012
rect 7862 141956 7918 142012
rect 7918 141956 7922 142012
rect 7858 141952 7922 141956
rect 2618 141468 2682 141472
rect 2618 141412 2622 141468
rect 2622 141412 2678 141468
rect 2678 141412 2682 141468
rect 2618 141408 2682 141412
rect 2698 141468 2762 141472
rect 2698 141412 2702 141468
rect 2702 141412 2758 141468
rect 2758 141412 2762 141468
rect 2698 141408 2762 141412
rect 2778 141468 2842 141472
rect 2778 141412 2782 141468
rect 2782 141412 2838 141468
rect 2838 141412 2842 141468
rect 2778 141408 2842 141412
rect 2858 141468 2922 141472
rect 2858 141412 2862 141468
rect 2862 141412 2918 141468
rect 2918 141412 2922 141468
rect 2858 141408 2922 141412
rect 5952 141468 6016 141472
rect 5952 141412 5956 141468
rect 5956 141412 6012 141468
rect 6012 141412 6016 141468
rect 5952 141408 6016 141412
rect 6032 141468 6096 141472
rect 6032 141412 6036 141468
rect 6036 141412 6092 141468
rect 6092 141412 6096 141468
rect 6032 141408 6096 141412
rect 6112 141468 6176 141472
rect 6112 141412 6116 141468
rect 6116 141412 6172 141468
rect 6172 141412 6176 141468
rect 6112 141408 6176 141412
rect 6192 141468 6256 141472
rect 6192 141412 6196 141468
rect 6196 141412 6252 141468
rect 6252 141412 6256 141468
rect 6192 141408 6256 141412
rect 4285 140924 4349 140928
rect 4285 140868 4289 140924
rect 4289 140868 4345 140924
rect 4345 140868 4349 140924
rect 4285 140864 4349 140868
rect 4365 140924 4429 140928
rect 4365 140868 4369 140924
rect 4369 140868 4425 140924
rect 4425 140868 4429 140924
rect 4365 140864 4429 140868
rect 4445 140924 4509 140928
rect 4445 140868 4449 140924
rect 4449 140868 4505 140924
rect 4505 140868 4509 140924
rect 4445 140864 4509 140868
rect 4525 140924 4589 140928
rect 4525 140868 4529 140924
rect 4529 140868 4585 140924
rect 4585 140868 4589 140924
rect 4525 140864 4589 140868
rect 7618 140924 7682 140928
rect 7618 140868 7622 140924
rect 7622 140868 7678 140924
rect 7678 140868 7682 140924
rect 7618 140864 7682 140868
rect 7698 140924 7762 140928
rect 7698 140868 7702 140924
rect 7702 140868 7758 140924
rect 7758 140868 7762 140924
rect 7698 140864 7762 140868
rect 7778 140924 7842 140928
rect 7778 140868 7782 140924
rect 7782 140868 7838 140924
rect 7838 140868 7842 140924
rect 7778 140864 7842 140868
rect 7858 140924 7922 140928
rect 7858 140868 7862 140924
rect 7862 140868 7918 140924
rect 7918 140868 7922 140924
rect 7858 140864 7922 140868
rect 2618 140380 2682 140384
rect 2618 140324 2622 140380
rect 2622 140324 2678 140380
rect 2678 140324 2682 140380
rect 2618 140320 2682 140324
rect 2698 140380 2762 140384
rect 2698 140324 2702 140380
rect 2702 140324 2758 140380
rect 2758 140324 2762 140380
rect 2698 140320 2762 140324
rect 2778 140380 2842 140384
rect 2778 140324 2782 140380
rect 2782 140324 2838 140380
rect 2838 140324 2842 140380
rect 2778 140320 2842 140324
rect 2858 140380 2922 140384
rect 2858 140324 2862 140380
rect 2862 140324 2918 140380
rect 2918 140324 2922 140380
rect 2858 140320 2922 140324
rect 5952 140380 6016 140384
rect 5952 140324 5956 140380
rect 5956 140324 6012 140380
rect 6012 140324 6016 140380
rect 5952 140320 6016 140324
rect 6032 140380 6096 140384
rect 6032 140324 6036 140380
rect 6036 140324 6092 140380
rect 6092 140324 6096 140380
rect 6032 140320 6096 140324
rect 6112 140380 6176 140384
rect 6112 140324 6116 140380
rect 6116 140324 6172 140380
rect 6172 140324 6176 140380
rect 6112 140320 6176 140324
rect 6192 140380 6256 140384
rect 6192 140324 6196 140380
rect 6196 140324 6252 140380
rect 6252 140324 6256 140380
rect 6192 140320 6256 140324
rect 4285 139836 4349 139840
rect 4285 139780 4289 139836
rect 4289 139780 4345 139836
rect 4345 139780 4349 139836
rect 4285 139776 4349 139780
rect 4365 139836 4429 139840
rect 4365 139780 4369 139836
rect 4369 139780 4425 139836
rect 4425 139780 4429 139836
rect 4365 139776 4429 139780
rect 4445 139836 4509 139840
rect 4445 139780 4449 139836
rect 4449 139780 4505 139836
rect 4505 139780 4509 139836
rect 4445 139776 4509 139780
rect 4525 139836 4589 139840
rect 4525 139780 4529 139836
rect 4529 139780 4585 139836
rect 4585 139780 4589 139836
rect 4525 139776 4589 139780
rect 7618 139836 7682 139840
rect 7618 139780 7622 139836
rect 7622 139780 7678 139836
rect 7678 139780 7682 139836
rect 7618 139776 7682 139780
rect 7698 139836 7762 139840
rect 7698 139780 7702 139836
rect 7702 139780 7758 139836
rect 7758 139780 7762 139836
rect 7698 139776 7762 139780
rect 7778 139836 7842 139840
rect 7778 139780 7782 139836
rect 7782 139780 7838 139836
rect 7838 139780 7842 139836
rect 7778 139776 7842 139780
rect 7858 139836 7922 139840
rect 7858 139780 7862 139836
rect 7862 139780 7918 139836
rect 7918 139780 7922 139836
rect 7858 139776 7922 139780
rect 2618 139292 2682 139296
rect 2618 139236 2622 139292
rect 2622 139236 2678 139292
rect 2678 139236 2682 139292
rect 2618 139232 2682 139236
rect 2698 139292 2762 139296
rect 2698 139236 2702 139292
rect 2702 139236 2758 139292
rect 2758 139236 2762 139292
rect 2698 139232 2762 139236
rect 2778 139292 2842 139296
rect 2778 139236 2782 139292
rect 2782 139236 2838 139292
rect 2838 139236 2842 139292
rect 2778 139232 2842 139236
rect 2858 139292 2922 139296
rect 2858 139236 2862 139292
rect 2862 139236 2918 139292
rect 2918 139236 2922 139292
rect 2858 139232 2922 139236
rect 5952 139292 6016 139296
rect 5952 139236 5956 139292
rect 5956 139236 6012 139292
rect 6012 139236 6016 139292
rect 5952 139232 6016 139236
rect 6032 139292 6096 139296
rect 6032 139236 6036 139292
rect 6036 139236 6092 139292
rect 6092 139236 6096 139292
rect 6032 139232 6096 139236
rect 6112 139292 6176 139296
rect 6112 139236 6116 139292
rect 6116 139236 6172 139292
rect 6172 139236 6176 139292
rect 6112 139232 6176 139236
rect 6192 139292 6256 139296
rect 6192 139236 6196 139292
rect 6196 139236 6252 139292
rect 6252 139236 6256 139292
rect 6192 139232 6256 139236
rect 4285 138748 4349 138752
rect 4285 138692 4289 138748
rect 4289 138692 4345 138748
rect 4345 138692 4349 138748
rect 4285 138688 4349 138692
rect 4365 138748 4429 138752
rect 4365 138692 4369 138748
rect 4369 138692 4425 138748
rect 4425 138692 4429 138748
rect 4365 138688 4429 138692
rect 4445 138748 4509 138752
rect 4445 138692 4449 138748
rect 4449 138692 4505 138748
rect 4505 138692 4509 138748
rect 4445 138688 4509 138692
rect 4525 138748 4589 138752
rect 4525 138692 4529 138748
rect 4529 138692 4585 138748
rect 4585 138692 4589 138748
rect 4525 138688 4589 138692
rect 7618 138748 7682 138752
rect 7618 138692 7622 138748
rect 7622 138692 7678 138748
rect 7678 138692 7682 138748
rect 7618 138688 7682 138692
rect 7698 138748 7762 138752
rect 7698 138692 7702 138748
rect 7702 138692 7758 138748
rect 7758 138692 7762 138748
rect 7698 138688 7762 138692
rect 7778 138748 7842 138752
rect 7778 138692 7782 138748
rect 7782 138692 7838 138748
rect 7838 138692 7842 138748
rect 7778 138688 7842 138692
rect 7858 138748 7922 138752
rect 7858 138692 7862 138748
rect 7862 138692 7918 138748
rect 7918 138692 7922 138748
rect 7858 138688 7922 138692
rect 2618 138204 2682 138208
rect 2618 138148 2622 138204
rect 2622 138148 2678 138204
rect 2678 138148 2682 138204
rect 2618 138144 2682 138148
rect 2698 138204 2762 138208
rect 2698 138148 2702 138204
rect 2702 138148 2758 138204
rect 2758 138148 2762 138204
rect 2698 138144 2762 138148
rect 2778 138204 2842 138208
rect 2778 138148 2782 138204
rect 2782 138148 2838 138204
rect 2838 138148 2842 138204
rect 2778 138144 2842 138148
rect 2858 138204 2922 138208
rect 2858 138148 2862 138204
rect 2862 138148 2918 138204
rect 2918 138148 2922 138204
rect 2858 138144 2922 138148
rect 5952 138204 6016 138208
rect 5952 138148 5956 138204
rect 5956 138148 6012 138204
rect 6012 138148 6016 138204
rect 5952 138144 6016 138148
rect 6032 138204 6096 138208
rect 6032 138148 6036 138204
rect 6036 138148 6092 138204
rect 6092 138148 6096 138204
rect 6032 138144 6096 138148
rect 6112 138204 6176 138208
rect 6112 138148 6116 138204
rect 6116 138148 6172 138204
rect 6172 138148 6176 138204
rect 6112 138144 6176 138148
rect 6192 138204 6256 138208
rect 6192 138148 6196 138204
rect 6196 138148 6252 138204
rect 6252 138148 6256 138204
rect 6192 138144 6256 138148
rect 4285 137660 4349 137664
rect 4285 137604 4289 137660
rect 4289 137604 4345 137660
rect 4345 137604 4349 137660
rect 4285 137600 4349 137604
rect 4365 137660 4429 137664
rect 4365 137604 4369 137660
rect 4369 137604 4425 137660
rect 4425 137604 4429 137660
rect 4365 137600 4429 137604
rect 4445 137660 4509 137664
rect 4445 137604 4449 137660
rect 4449 137604 4505 137660
rect 4505 137604 4509 137660
rect 4445 137600 4509 137604
rect 4525 137660 4589 137664
rect 4525 137604 4529 137660
rect 4529 137604 4585 137660
rect 4585 137604 4589 137660
rect 4525 137600 4589 137604
rect 7618 137660 7682 137664
rect 7618 137604 7622 137660
rect 7622 137604 7678 137660
rect 7678 137604 7682 137660
rect 7618 137600 7682 137604
rect 7698 137660 7762 137664
rect 7698 137604 7702 137660
rect 7702 137604 7758 137660
rect 7758 137604 7762 137660
rect 7698 137600 7762 137604
rect 7778 137660 7842 137664
rect 7778 137604 7782 137660
rect 7782 137604 7838 137660
rect 7838 137604 7842 137660
rect 7778 137600 7842 137604
rect 7858 137660 7922 137664
rect 7858 137604 7862 137660
rect 7862 137604 7918 137660
rect 7918 137604 7922 137660
rect 7858 137600 7922 137604
rect 2618 137116 2682 137120
rect 2618 137060 2622 137116
rect 2622 137060 2678 137116
rect 2678 137060 2682 137116
rect 2618 137056 2682 137060
rect 2698 137116 2762 137120
rect 2698 137060 2702 137116
rect 2702 137060 2758 137116
rect 2758 137060 2762 137116
rect 2698 137056 2762 137060
rect 2778 137116 2842 137120
rect 2778 137060 2782 137116
rect 2782 137060 2838 137116
rect 2838 137060 2842 137116
rect 2778 137056 2842 137060
rect 2858 137116 2922 137120
rect 2858 137060 2862 137116
rect 2862 137060 2918 137116
rect 2918 137060 2922 137116
rect 2858 137056 2922 137060
rect 5952 137116 6016 137120
rect 5952 137060 5956 137116
rect 5956 137060 6012 137116
rect 6012 137060 6016 137116
rect 5952 137056 6016 137060
rect 6032 137116 6096 137120
rect 6032 137060 6036 137116
rect 6036 137060 6092 137116
rect 6092 137060 6096 137116
rect 6032 137056 6096 137060
rect 6112 137116 6176 137120
rect 6112 137060 6116 137116
rect 6116 137060 6172 137116
rect 6172 137060 6176 137116
rect 6112 137056 6176 137060
rect 6192 137116 6256 137120
rect 6192 137060 6196 137116
rect 6196 137060 6252 137116
rect 6252 137060 6256 137116
rect 6192 137056 6256 137060
rect 4285 136572 4349 136576
rect 4285 136516 4289 136572
rect 4289 136516 4345 136572
rect 4345 136516 4349 136572
rect 4285 136512 4349 136516
rect 4365 136572 4429 136576
rect 4365 136516 4369 136572
rect 4369 136516 4425 136572
rect 4425 136516 4429 136572
rect 4365 136512 4429 136516
rect 4445 136572 4509 136576
rect 4445 136516 4449 136572
rect 4449 136516 4505 136572
rect 4505 136516 4509 136572
rect 4445 136512 4509 136516
rect 4525 136572 4589 136576
rect 4525 136516 4529 136572
rect 4529 136516 4585 136572
rect 4585 136516 4589 136572
rect 4525 136512 4589 136516
rect 7618 136572 7682 136576
rect 7618 136516 7622 136572
rect 7622 136516 7678 136572
rect 7678 136516 7682 136572
rect 7618 136512 7682 136516
rect 7698 136572 7762 136576
rect 7698 136516 7702 136572
rect 7702 136516 7758 136572
rect 7758 136516 7762 136572
rect 7698 136512 7762 136516
rect 7778 136572 7842 136576
rect 7778 136516 7782 136572
rect 7782 136516 7838 136572
rect 7838 136516 7842 136572
rect 7778 136512 7842 136516
rect 7858 136572 7922 136576
rect 7858 136516 7862 136572
rect 7862 136516 7918 136572
rect 7918 136516 7922 136572
rect 7858 136512 7922 136516
rect 2618 136028 2682 136032
rect 2618 135972 2622 136028
rect 2622 135972 2678 136028
rect 2678 135972 2682 136028
rect 2618 135968 2682 135972
rect 2698 136028 2762 136032
rect 2698 135972 2702 136028
rect 2702 135972 2758 136028
rect 2758 135972 2762 136028
rect 2698 135968 2762 135972
rect 2778 136028 2842 136032
rect 2778 135972 2782 136028
rect 2782 135972 2838 136028
rect 2838 135972 2842 136028
rect 2778 135968 2842 135972
rect 2858 136028 2922 136032
rect 2858 135972 2862 136028
rect 2862 135972 2918 136028
rect 2918 135972 2922 136028
rect 2858 135968 2922 135972
rect 5952 136028 6016 136032
rect 5952 135972 5956 136028
rect 5956 135972 6012 136028
rect 6012 135972 6016 136028
rect 5952 135968 6016 135972
rect 6032 136028 6096 136032
rect 6032 135972 6036 136028
rect 6036 135972 6092 136028
rect 6092 135972 6096 136028
rect 6032 135968 6096 135972
rect 6112 136028 6176 136032
rect 6112 135972 6116 136028
rect 6116 135972 6172 136028
rect 6172 135972 6176 136028
rect 6112 135968 6176 135972
rect 6192 136028 6256 136032
rect 6192 135972 6196 136028
rect 6196 135972 6252 136028
rect 6252 135972 6256 136028
rect 6192 135968 6256 135972
rect 4285 135484 4349 135488
rect 4285 135428 4289 135484
rect 4289 135428 4345 135484
rect 4345 135428 4349 135484
rect 4285 135424 4349 135428
rect 4365 135484 4429 135488
rect 4365 135428 4369 135484
rect 4369 135428 4425 135484
rect 4425 135428 4429 135484
rect 4365 135424 4429 135428
rect 4445 135484 4509 135488
rect 4445 135428 4449 135484
rect 4449 135428 4505 135484
rect 4505 135428 4509 135484
rect 4445 135424 4509 135428
rect 4525 135484 4589 135488
rect 4525 135428 4529 135484
rect 4529 135428 4585 135484
rect 4585 135428 4589 135484
rect 4525 135424 4589 135428
rect 7618 135484 7682 135488
rect 7618 135428 7622 135484
rect 7622 135428 7678 135484
rect 7678 135428 7682 135484
rect 7618 135424 7682 135428
rect 7698 135484 7762 135488
rect 7698 135428 7702 135484
rect 7702 135428 7758 135484
rect 7758 135428 7762 135484
rect 7698 135424 7762 135428
rect 7778 135484 7842 135488
rect 7778 135428 7782 135484
rect 7782 135428 7838 135484
rect 7838 135428 7842 135484
rect 7778 135424 7842 135428
rect 7858 135484 7922 135488
rect 7858 135428 7862 135484
rect 7862 135428 7918 135484
rect 7918 135428 7922 135484
rect 7858 135424 7922 135428
rect 2618 134940 2682 134944
rect 2618 134884 2622 134940
rect 2622 134884 2678 134940
rect 2678 134884 2682 134940
rect 2618 134880 2682 134884
rect 2698 134940 2762 134944
rect 2698 134884 2702 134940
rect 2702 134884 2758 134940
rect 2758 134884 2762 134940
rect 2698 134880 2762 134884
rect 2778 134940 2842 134944
rect 2778 134884 2782 134940
rect 2782 134884 2838 134940
rect 2838 134884 2842 134940
rect 2778 134880 2842 134884
rect 2858 134940 2922 134944
rect 2858 134884 2862 134940
rect 2862 134884 2918 134940
rect 2918 134884 2922 134940
rect 2858 134880 2922 134884
rect 5952 134940 6016 134944
rect 5952 134884 5956 134940
rect 5956 134884 6012 134940
rect 6012 134884 6016 134940
rect 5952 134880 6016 134884
rect 6032 134940 6096 134944
rect 6032 134884 6036 134940
rect 6036 134884 6092 134940
rect 6092 134884 6096 134940
rect 6032 134880 6096 134884
rect 6112 134940 6176 134944
rect 6112 134884 6116 134940
rect 6116 134884 6172 134940
rect 6172 134884 6176 134940
rect 6112 134880 6176 134884
rect 6192 134940 6256 134944
rect 6192 134884 6196 134940
rect 6196 134884 6252 134940
rect 6252 134884 6256 134940
rect 6192 134880 6256 134884
rect 4285 134396 4349 134400
rect 4285 134340 4289 134396
rect 4289 134340 4345 134396
rect 4345 134340 4349 134396
rect 4285 134336 4349 134340
rect 4365 134396 4429 134400
rect 4365 134340 4369 134396
rect 4369 134340 4425 134396
rect 4425 134340 4429 134396
rect 4365 134336 4429 134340
rect 4445 134396 4509 134400
rect 4445 134340 4449 134396
rect 4449 134340 4505 134396
rect 4505 134340 4509 134396
rect 4445 134336 4509 134340
rect 4525 134396 4589 134400
rect 4525 134340 4529 134396
rect 4529 134340 4585 134396
rect 4585 134340 4589 134396
rect 4525 134336 4589 134340
rect 7618 134396 7682 134400
rect 7618 134340 7622 134396
rect 7622 134340 7678 134396
rect 7678 134340 7682 134396
rect 7618 134336 7682 134340
rect 7698 134396 7762 134400
rect 7698 134340 7702 134396
rect 7702 134340 7758 134396
rect 7758 134340 7762 134396
rect 7698 134336 7762 134340
rect 7778 134396 7842 134400
rect 7778 134340 7782 134396
rect 7782 134340 7838 134396
rect 7838 134340 7842 134396
rect 7778 134336 7842 134340
rect 7858 134396 7922 134400
rect 7858 134340 7862 134396
rect 7862 134340 7918 134396
rect 7918 134340 7922 134396
rect 7858 134336 7922 134340
rect 2618 133852 2682 133856
rect 2618 133796 2622 133852
rect 2622 133796 2678 133852
rect 2678 133796 2682 133852
rect 2618 133792 2682 133796
rect 2698 133852 2762 133856
rect 2698 133796 2702 133852
rect 2702 133796 2758 133852
rect 2758 133796 2762 133852
rect 2698 133792 2762 133796
rect 2778 133852 2842 133856
rect 2778 133796 2782 133852
rect 2782 133796 2838 133852
rect 2838 133796 2842 133852
rect 2778 133792 2842 133796
rect 2858 133852 2922 133856
rect 2858 133796 2862 133852
rect 2862 133796 2918 133852
rect 2918 133796 2922 133852
rect 2858 133792 2922 133796
rect 5952 133852 6016 133856
rect 5952 133796 5956 133852
rect 5956 133796 6012 133852
rect 6012 133796 6016 133852
rect 5952 133792 6016 133796
rect 6032 133852 6096 133856
rect 6032 133796 6036 133852
rect 6036 133796 6092 133852
rect 6092 133796 6096 133852
rect 6032 133792 6096 133796
rect 6112 133852 6176 133856
rect 6112 133796 6116 133852
rect 6116 133796 6172 133852
rect 6172 133796 6176 133852
rect 6112 133792 6176 133796
rect 6192 133852 6256 133856
rect 6192 133796 6196 133852
rect 6196 133796 6252 133852
rect 6252 133796 6256 133852
rect 6192 133792 6256 133796
rect 4285 133308 4349 133312
rect 4285 133252 4289 133308
rect 4289 133252 4345 133308
rect 4345 133252 4349 133308
rect 4285 133248 4349 133252
rect 4365 133308 4429 133312
rect 4365 133252 4369 133308
rect 4369 133252 4425 133308
rect 4425 133252 4429 133308
rect 4365 133248 4429 133252
rect 4445 133308 4509 133312
rect 4445 133252 4449 133308
rect 4449 133252 4505 133308
rect 4505 133252 4509 133308
rect 4445 133248 4509 133252
rect 4525 133308 4589 133312
rect 4525 133252 4529 133308
rect 4529 133252 4585 133308
rect 4585 133252 4589 133308
rect 4525 133248 4589 133252
rect 7618 133308 7682 133312
rect 7618 133252 7622 133308
rect 7622 133252 7678 133308
rect 7678 133252 7682 133308
rect 7618 133248 7682 133252
rect 7698 133308 7762 133312
rect 7698 133252 7702 133308
rect 7702 133252 7758 133308
rect 7758 133252 7762 133308
rect 7698 133248 7762 133252
rect 7778 133308 7842 133312
rect 7778 133252 7782 133308
rect 7782 133252 7838 133308
rect 7838 133252 7842 133308
rect 7778 133248 7842 133252
rect 7858 133308 7922 133312
rect 7858 133252 7862 133308
rect 7862 133252 7918 133308
rect 7918 133252 7922 133308
rect 7858 133248 7922 133252
rect 2618 132764 2682 132768
rect 2618 132708 2622 132764
rect 2622 132708 2678 132764
rect 2678 132708 2682 132764
rect 2618 132704 2682 132708
rect 2698 132764 2762 132768
rect 2698 132708 2702 132764
rect 2702 132708 2758 132764
rect 2758 132708 2762 132764
rect 2698 132704 2762 132708
rect 2778 132764 2842 132768
rect 2778 132708 2782 132764
rect 2782 132708 2838 132764
rect 2838 132708 2842 132764
rect 2778 132704 2842 132708
rect 2858 132764 2922 132768
rect 2858 132708 2862 132764
rect 2862 132708 2918 132764
rect 2918 132708 2922 132764
rect 2858 132704 2922 132708
rect 5952 132764 6016 132768
rect 5952 132708 5956 132764
rect 5956 132708 6012 132764
rect 6012 132708 6016 132764
rect 5952 132704 6016 132708
rect 6032 132764 6096 132768
rect 6032 132708 6036 132764
rect 6036 132708 6092 132764
rect 6092 132708 6096 132764
rect 6032 132704 6096 132708
rect 6112 132764 6176 132768
rect 6112 132708 6116 132764
rect 6116 132708 6172 132764
rect 6172 132708 6176 132764
rect 6112 132704 6176 132708
rect 6192 132764 6256 132768
rect 6192 132708 6196 132764
rect 6196 132708 6252 132764
rect 6252 132708 6256 132764
rect 6192 132704 6256 132708
rect 4285 132220 4349 132224
rect 4285 132164 4289 132220
rect 4289 132164 4345 132220
rect 4345 132164 4349 132220
rect 4285 132160 4349 132164
rect 4365 132220 4429 132224
rect 4365 132164 4369 132220
rect 4369 132164 4425 132220
rect 4425 132164 4429 132220
rect 4365 132160 4429 132164
rect 4445 132220 4509 132224
rect 4445 132164 4449 132220
rect 4449 132164 4505 132220
rect 4505 132164 4509 132220
rect 4445 132160 4509 132164
rect 4525 132220 4589 132224
rect 4525 132164 4529 132220
rect 4529 132164 4585 132220
rect 4585 132164 4589 132220
rect 4525 132160 4589 132164
rect 7618 132220 7682 132224
rect 7618 132164 7622 132220
rect 7622 132164 7678 132220
rect 7678 132164 7682 132220
rect 7618 132160 7682 132164
rect 7698 132220 7762 132224
rect 7698 132164 7702 132220
rect 7702 132164 7758 132220
rect 7758 132164 7762 132220
rect 7698 132160 7762 132164
rect 7778 132220 7842 132224
rect 7778 132164 7782 132220
rect 7782 132164 7838 132220
rect 7838 132164 7842 132220
rect 7778 132160 7842 132164
rect 7858 132220 7922 132224
rect 7858 132164 7862 132220
rect 7862 132164 7918 132220
rect 7918 132164 7922 132220
rect 7858 132160 7922 132164
rect 2618 131676 2682 131680
rect 2618 131620 2622 131676
rect 2622 131620 2678 131676
rect 2678 131620 2682 131676
rect 2618 131616 2682 131620
rect 2698 131676 2762 131680
rect 2698 131620 2702 131676
rect 2702 131620 2758 131676
rect 2758 131620 2762 131676
rect 2698 131616 2762 131620
rect 2778 131676 2842 131680
rect 2778 131620 2782 131676
rect 2782 131620 2838 131676
rect 2838 131620 2842 131676
rect 2778 131616 2842 131620
rect 2858 131676 2922 131680
rect 2858 131620 2862 131676
rect 2862 131620 2918 131676
rect 2918 131620 2922 131676
rect 2858 131616 2922 131620
rect 5952 131676 6016 131680
rect 5952 131620 5956 131676
rect 5956 131620 6012 131676
rect 6012 131620 6016 131676
rect 5952 131616 6016 131620
rect 6032 131676 6096 131680
rect 6032 131620 6036 131676
rect 6036 131620 6092 131676
rect 6092 131620 6096 131676
rect 6032 131616 6096 131620
rect 6112 131676 6176 131680
rect 6112 131620 6116 131676
rect 6116 131620 6172 131676
rect 6172 131620 6176 131676
rect 6112 131616 6176 131620
rect 6192 131676 6256 131680
rect 6192 131620 6196 131676
rect 6196 131620 6252 131676
rect 6252 131620 6256 131676
rect 6192 131616 6256 131620
rect 4285 131132 4349 131136
rect 4285 131076 4289 131132
rect 4289 131076 4345 131132
rect 4345 131076 4349 131132
rect 4285 131072 4349 131076
rect 4365 131132 4429 131136
rect 4365 131076 4369 131132
rect 4369 131076 4425 131132
rect 4425 131076 4429 131132
rect 4365 131072 4429 131076
rect 4445 131132 4509 131136
rect 4445 131076 4449 131132
rect 4449 131076 4505 131132
rect 4505 131076 4509 131132
rect 4445 131072 4509 131076
rect 4525 131132 4589 131136
rect 4525 131076 4529 131132
rect 4529 131076 4585 131132
rect 4585 131076 4589 131132
rect 4525 131072 4589 131076
rect 7618 131132 7682 131136
rect 7618 131076 7622 131132
rect 7622 131076 7678 131132
rect 7678 131076 7682 131132
rect 7618 131072 7682 131076
rect 7698 131132 7762 131136
rect 7698 131076 7702 131132
rect 7702 131076 7758 131132
rect 7758 131076 7762 131132
rect 7698 131072 7762 131076
rect 7778 131132 7842 131136
rect 7778 131076 7782 131132
rect 7782 131076 7838 131132
rect 7838 131076 7842 131132
rect 7778 131072 7842 131076
rect 7858 131132 7922 131136
rect 7858 131076 7862 131132
rect 7862 131076 7918 131132
rect 7918 131076 7922 131132
rect 7858 131072 7922 131076
rect 2618 130588 2682 130592
rect 2618 130532 2622 130588
rect 2622 130532 2678 130588
rect 2678 130532 2682 130588
rect 2618 130528 2682 130532
rect 2698 130588 2762 130592
rect 2698 130532 2702 130588
rect 2702 130532 2758 130588
rect 2758 130532 2762 130588
rect 2698 130528 2762 130532
rect 2778 130588 2842 130592
rect 2778 130532 2782 130588
rect 2782 130532 2838 130588
rect 2838 130532 2842 130588
rect 2778 130528 2842 130532
rect 2858 130588 2922 130592
rect 2858 130532 2862 130588
rect 2862 130532 2918 130588
rect 2918 130532 2922 130588
rect 2858 130528 2922 130532
rect 5952 130588 6016 130592
rect 5952 130532 5956 130588
rect 5956 130532 6012 130588
rect 6012 130532 6016 130588
rect 5952 130528 6016 130532
rect 6032 130588 6096 130592
rect 6032 130532 6036 130588
rect 6036 130532 6092 130588
rect 6092 130532 6096 130588
rect 6032 130528 6096 130532
rect 6112 130588 6176 130592
rect 6112 130532 6116 130588
rect 6116 130532 6172 130588
rect 6172 130532 6176 130588
rect 6112 130528 6176 130532
rect 6192 130588 6256 130592
rect 6192 130532 6196 130588
rect 6196 130532 6252 130588
rect 6252 130532 6256 130588
rect 6192 130528 6256 130532
rect 4285 130044 4349 130048
rect 4285 129988 4289 130044
rect 4289 129988 4345 130044
rect 4345 129988 4349 130044
rect 4285 129984 4349 129988
rect 4365 130044 4429 130048
rect 4365 129988 4369 130044
rect 4369 129988 4425 130044
rect 4425 129988 4429 130044
rect 4365 129984 4429 129988
rect 4445 130044 4509 130048
rect 4445 129988 4449 130044
rect 4449 129988 4505 130044
rect 4505 129988 4509 130044
rect 4445 129984 4509 129988
rect 4525 130044 4589 130048
rect 4525 129988 4529 130044
rect 4529 129988 4585 130044
rect 4585 129988 4589 130044
rect 4525 129984 4589 129988
rect 7618 130044 7682 130048
rect 7618 129988 7622 130044
rect 7622 129988 7678 130044
rect 7678 129988 7682 130044
rect 7618 129984 7682 129988
rect 7698 130044 7762 130048
rect 7698 129988 7702 130044
rect 7702 129988 7758 130044
rect 7758 129988 7762 130044
rect 7698 129984 7762 129988
rect 7778 130044 7842 130048
rect 7778 129988 7782 130044
rect 7782 129988 7838 130044
rect 7838 129988 7842 130044
rect 7778 129984 7842 129988
rect 7858 130044 7922 130048
rect 7858 129988 7862 130044
rect 7862 129988 7918 130044
rect 7918 129988 7922 130044
rect 7858 129984 7922 129988
rect 2618 129500 2682 129504
rect 2618 129444 2622 129500
rect 2622 129444 2678 129500
rect 2678 129444 2682 129500
rect 2618 129440 2682 129444
rect 2698 129500 2762 129504
rect 2698 129444 2702 129500
rect 2702 129444 2758 129500
rect 2758 129444 2762 129500
rect 2698 129440 2762 129444
rect 2778 129500 2842 129504
rect 2778 129444 2782 129500
rect 2782 129444 2838 129500
rect 2838 129444 2842 129500
rect 2778 129440 2842 129444
rect 2858 129500 2922 129504
rect 2858 129444 2862 129500
rect 2862 129444 2918 129500
rect 2918 129444 2922 129500
rect 2858 129440 2922 129444
rect 5952 129500 6016 129504
rect 5952 129444 5956 129500
rect 5956 129444 6012 129500
rect 6012 129444 6016 129500
rect 5952 129440 6016 129444
rect 6032 129500 6096 129504
rect 6032 129444 6036 129500
rect 6036 129444 6092 129500
rect 6092 129444 6096 129500
rect 6032 129440 6096 129444
rect 6112 129500 6176 129504
rect 6112 129444 6116 129500
rect 6116 129444 6172 129500
rect 6172 129444 6176 129500
rect 6112 129440 6176 129444
rect 6192 129500 6256 129504
rect 6192 129444 6196 129500
rect 6196 129444 6252 129500
rect 6252 129444 6256 129500
rect 6192 129440 6256 129444
rect 4285 128956 4349 128960
rect 4285 128900 4289 128956
rect 4289 128900 4345 128956
rect 4345 128900 4349 128956
rect 4285 128896 4349 128900
rect 4365 128956 4429 128960
rect 4365 128900 4369 128956
rect 4369 128900 4425 128956
rect 4425 128900 4429 128956
rect 4365 128896 4429 128900
rect 4445 128956 4509 128960
rect 4445 128900 4449 128956
rect 4449 128900 4505 128956
rect 4505 128900 4509 128956
rect 4445 128896 4509 128900
rect 4525 128956 4589 128960
rect 4525 128900 4529 128956
rect 4529 128900 4585 128956
rect 4585 128900 4589 128956
rect 4525 128896 4589 128900
rect 7618 128956 7682 128960
rect 7618 128900 7622 128956
rect 7622 128900 7678 128956
rect 7678 128900 7682 128956
rect 7618 128896 7682 128900
rect 7698 128956 7762 128960
rect 7698 128900 7702 128956
rect 7702 128900 7758 128956
rect 7758 128900 7762 128956
rect 7698 128896 7762 128900
rect 7778 128956 7842 128960
rect 7778 128900 7782 128956
rect 7782 128900 7838 128956
rect 7838 128900 7842 128956
rect 7778 128896 7842 128900
rect 7858 128956 7922 128960
rect 7858 128900 7862 128956
rect 7862 128900 7918 128956
rect 7918 128900 7922 128956
rect 7858 128896 7922 128900
rect 2618 128412 2682 128416
rect 2618 128356 2622 128412
rect 2622 128356 2678 128412
rect 2678 128356 2682 128412
rect 2618 128352 2682 128356
rect 2698 128412 2762 128416
rect 2698 128356 2702 128412
rect 2702 128356 2758 128412
rect 2758 128356 2762 128412
rect 2698 128352 2762 128356
rect 2778 128412 2842 128416
rect 2778 128356 2782 128412
rect 2782 128356 2838 128412
rect 2838 128356 2842 128412
rect 2778 128352 2842 128356
rect 2858 128412 2922 128416
rect 2858 128356 2862 128412
rect 2862 128356 2918 128412
rect 2918 128356 2922 128412
rect 2858 128352 2922 128356
rect 5952 128412 6016 128416
rect 5952 128356 5956 128412
rect 5956 128356 6012 128412
rect 6012 128356 6016 128412
rect 5952 128352 6016 128356
rect 6032 128412 6096 128416
rect 6032 128356 6036 128412
rect 6036 128356 6092 128412
rect 6092 128356 6096 128412
rect 6032 128352 6096 128356
rect 6112 128412 6176 128416
rect 6112 128356 6116 128412
rect 6116 128356 6172 128412
rect 6172 128356 6176 128412
rect 6112 128352 6176 128356
rect 6192 128412 6256 128416
rect 6192 128356 6196 128412
rect 6196 128356 6252 128412
rect 6252 128356 6256 128412
rect 6192 128352 6256 128356
rect 4285 127868 4349 127872
rect 4285 127812 4289 127868
rect 4289 127812 4345 127868
rect 4345 127812 4349 127868
rect 4285 127808 4349 127812
rect 4365 127868 4429 127872
rect 4365 127812 4369 127868
rect 4369 127812 4425 127868
rect 4425 127812 4429 127868
rect 4365 127808 4429 127812
rect 4445 127868 4509 127872
rect 4445 127812 4449 127868
rect 4449 127812 4505 127868
rect 4505 127812 4509 127868
rect 4445 127808 4509 127812
rect 4525 127868 4589 127872
rect 4525 127812 4529 127868
rect 4529 127812 4585 127868
rect 4585 127812 4589 127868
rect 4525 127808 4589 127812
rect 7618 127868 7682 127872
rect 7618 127812 7622 127868
rect 7622 127812 7678 127868
rect 7678 127812 7682 127868
rect 7618 127808 7682 127812
rect 7698 127868 7762 127872
rect 7698 127812 7702 127868
rect 7702 127812 7758 127868
rect 7758 127812 7762 127868
rect 7698 127808 7762 127812
rect 7778 127868 7842 127872
rect 7778 127812 7782 127868
rect 7782 127812 7838 127868
rect 7838 127812 7842 127868
rect 7778 127808 7842 127812
rect 7858 127868 7922 127872
rect 7858 127812 7862 127868
rect 7862 127812 7918 127868
rect 7918 127812 7922 127868
rect 7858 127808 7922 127812
rect 2618 127324 2682 127328
rect 2618 127268 2622 127324
rect 2622 127268 2678 127324
rect 2678 127268 2682 127324
rect 2618 127264 2682 127268
rect 2698 127324 2762 127328
rect 2698 127268 2702 127324
rect 2702 127268 2758 127324
rect 2758 127268 2762 127324
rect 2698 127264 2762 127268
rect 2778 127324 2842 127328
rect 2778 127268 2782 127324
rect 2782 127268 2838 127324
rect 2838 127268 2842 127324
rect 2778 127264 2842 127268
rect 2858 127324 2922 127328
rect 2858 127268 2862 127324
rect 2862 127268 2918 127324
rect 2918 127268 2922 127324
rect 2858 127264 2922 127268
rect 5952 127324 6016 127328
rect 5952 127268 5956 127324
rect 5956 127268 6012 127324
rect 6012 127268 6016 127324
rect 5952 127264 6016 127268
rect 6032 127324 6096 127328
rect 6032 127268 6036 127324
rect 6036 127268 6092 127324
rect 6092 127268 6096 127324
rect 6032 127264 6096 127268
rect 6112 127324 6176 127328
rect 6112 127268 6116 127324
rect 6116 127268 6172 127324
rect 6172 127268 6176 127324
rect 6112 127264 6176 127268
rect 6192 127324 6256 127328
rect 6192 127268 6196 127324
rect 6196 127268 6252 127324
rect 6252 127268 6256 127324
rect 6192 127264 6256 127268
rect 4285 126780 4349 126784
rect 4285 126724 4289 126780
rect 4289 126724 4345 126780
rect 4345 126724 4349 126780
rect 4285 126720 4349 126724
rect 4365 126780 4429 126784
rect 4365 126724 4369 126780
rect 4369 126724 4425 126780
rect 4425 126724 4429 126780
rect 4365 126720 4429 126724
rect 4445 126780 4509 126784
rect 4445 126724 4449 126780
rect 4449 126724 4505 126780
rect 4505 126724 4509 126780
rect 4445 126720 4509 126724
rect 4525 126780 4589 126784
rect 4525 126724 4529 126780
rect 4529 126724 4585 126780
rect 4585 126724 4589 126780
rect 4525 126720 4589 126724
rect 7618 126780 7682 126784
rect 7618 126724 7622 126780
rect 7622 126724 7678 126780
rect 7678 126724 7682 126780
rect 7618 126720 7682 126724
rect 7698 126780 7762 126784
rect 7698 126724 7702 126780
rect 7702 126724 7758 126780
rect 7758 126724 7762 126780
rect 7698 126720 7762 126724
rect 7778 126780 7842 126784
rect 7778 126724 7782 126780
rect 7782 126724 7838 126780
rect 7838 126724 7842 126780
rect 7778 126720 7842 126724
rect 7858 126780 7922 126784
rect 7858 126724 7862 126780
rect 7862 126724 7918 126780
rect 7918 126724 7922 126780
rect 7858 126720 7922 126724
rect 2618 126236 2682 126240
rect 2618 126180 2622 126236
rect 2622 126180 2678 126236
rect 2678 126180 2682 126236
rect 2618 126176 2682 126180
rect 2698 126236 2762 126240
rect 2698 126180 2702 126236
rect 2702 126180 2758 126236
rect 2758 126180 2762 126236
rect 2698 126176 2762 126180
rect 2778 126236 2842 126240
rect 2778 126180 2782 126236
rect 2782 126180 2838 126236
rect 2838 126180 2842 126236
rect 2778 126176 2842 126180
rect 2858 126236 2922 126240
rect 2858 126180 2862 126236
rect 2862 126180 2918 126236
rect 2918 126180 2922 126236
rect 2858 126176 2922 126180
rect 5952 126236 6016 126240
rect 5952 126180 5956 126236
rect 5956 126180 6012 126236
rect 6012 126180 6016 126236
rect 5952 126176 6016 126180
rect 6032 126236 6096 126240
rect 6032 126180 6036 126236
rect 6036 126180 6092 126236
rect 6092 126180 6096 126236
rect 6032 126176 6096 126180
rect 6112 126236 6176 126240
rect 6112 126180 6116 126236
rect 6116 126180 6172 126236
rect 6172 126180 6176 126236
rect 6112 126176 6176 126180
rect 6192 126236 6256 126240
rect 6192 126180 6196 126236
rect 6196 126180 6252 126236
rect 6252 126180 6256 126236
rect 6192 126176 6256 126180
rect 4285 125692 4349 125696
rect 4285 125636 4289 125692
rect 4289 125636 4345 125692
rect 4345 125636 4349 125692
rect 4285 125632 4349 125636
rect 4365 125692 4429 125696
rect 4365 125636 4369 125692
rect 4369 125636 4425 125692
rect 4425 125636 4429 125692
rect 4365 125632 4429 125636
rect 4445 125692 4509 125696
rect 4445 125636 4449 125692
rect 4449 125636 4505 125692
rect 4505 125636 4509 125692
rect 4445 125632 4509 125636
rect 4525 125692 4589 125696
rect 4525 125636 4529 125692
rect 4529 125636 4585 125692
rect 4585 125636 4589 125692
rect 4525 125632 4589 125636
rect 7618 125692 7682 125696
rect 7618 125636 7622 125692
rect 7622 125636 7678 125692
rect 7678 125636 7682 125692
rect 7618 125632 7682 125636
rect 7698 125692 7762 125696
rect 7698 125636 7702 125692
rect 7702 125636 7758 125692
rect 7758 125636 7762 125692
rect 7698 125632 7762 125636
rect 7778 125692 7842 125696
rect 7778 125636 7782 125692
rect 7782 125636 7838 125692
rect 7838 125636 7842 125692
rect 7778 125632 7842 125636
rect 7858 125692 7922 125696
rect 7858 125636 7862 125692
rect 7862 125636 7918 125692
rect 7918 125636 7922 125692
rect 7858 125632 7922 125636
rect 2618 125148 2682 125152
rect 2618 125092 2622 125148
rect 2622 125092 2678 125148
rect 2678 125092 2682 125148
rect 2618 125088 2682 125092
rect 2698 125148 2762 125152
rect 2698 125092 2702 125148
rect 2702 125092 2758 125148
rect 2758 125092 2762 125148
rect 2698 125088 2762 125092
rect 2778 125148 2842 125152
rect 2778 125092 2782 125148
rect 2782 125092 2838 125148
rect 2838 125092 2842 125148
rect 2778 125088 2842 125092
rect 2858 125148 2922 125152
rect 2858 125092 2862 125148
rect 2862 125092 2918 125148
rect 2918 125092 2922 125148
rect 2858 125088 2922 125092
rect 5952 125148 6016 125152
rect 5952 125092 5956 125148
rect 5956 125092 6012 125148
rect 6012 125092 6016 125148
rect 5952 125088 6016 125092
rect 6032 125148 6096 125152
rect 6032 125092 6036 125148
rect 6036 125092 6092 125148
rect 6092 125092 6096 125148
rect 6032 125088 6096 125092
rect 6112 125148 6176 125152
rect 6112 125092 6116 125148
rect 6116 125092 6172 125148
rect 6172 125092 6176 125148
rect 6112 125088 6176 125092
rect 6192 125148 6256 125152
rect 6192 125092 6196 125148
rect 6196 125092 6252 125148
rect 6252 125092 6256 125148
rect 6192 125088 6256 125092
rect 4285 124604 4349 124608
rect 4285 124548 4289 124604
rect 4289 124548 4345 124604
rect 4345 124548 4349 124604
rect 4285 124544 4349 124548
rect 4365 124604 4429 124608
rect 4365 124548 4369 124604
rect 4369 124548 4425 124604
rect 4425 124548 4429 124604
rect 4365 124544 4429 124548
rect 4445 124604 4509 124608
rect 4445 124548 4449 124604
rect 4449 124548 4505 124604
rect 4505 124548 4509 124604
rect 4445 124544 4509 124548
rect 4525 124604 4589 124608
rect 4525 124548 4529 124604
rect 4529 124548 4585 124604
rect 4585 124548 4589 124604
rect 4525 124544 4589 124548
rect 7618 124604 7682 124608
rect 7618 124548 7622 124604
rect 7622 124548 7678 124604
rect 7678 124548 7682 124604
rect 7618 124544 7682 124548
rect 7698 124604 7762 124608
rect 7698 124548 7702 124604
rect 7702 124548 7758 124604
rect 7758 124548 7762 124604
rect 7698 124544 7762 124548
rect 7778 124604 7842 124608
rect 7778 124548 7782 124604
rect 7782 124548 7838 124604
rect 7838 124548 7842 124604
rect 7778 124544 7842 124548
rect 7858 124604 7922 124608
rect 7858 124548 7862 124604
rect 7862 124548 7918 124604
rect 7918 124548 7922 124604
rect 7858 124544 7922 124548
rect 2618 124060 2682 124064
rect 2618 124004 2622 124060
rect 2622 124004 2678 124060
rect 2678 124004 2682 124060
rect 2618 124000 2682 124004
rect 2698 124060 2762 124064
rect 2698 124004 2702 124060
rect 2702 124004 2758 124060
rect 2758 124004 2762 124060
rect 2698 124000 2762 124004
rect 2778 124060 2842 124064
rect 2778 124004 2782 124060
rect 2782 124004 2838 124060
rect 2838 124004 2842 124060
rect 2778 124000 2842 124004
rect 2858 124060 2922 124064
rect 2858 124004 2862 124060
rect 2862 124004 2918 124060
rect 2918 124004 2922 124060
rect 2858 124000 2922 124004
rect 5952 124060 6016 124064
rect 5952 124004 5956 124060
rect 5956 124004 6012 124060
rect 6012 124004 6016 124060
rect 5952 124000 6016 124004
rect 6032 124060 6096 124064
rect 6032 124004 6036 124060
rect 6036 124004 6092 124060
rect 6092 124004 6096 124060
rect 6032 124000 6096 124004
rect 6112 124060 6176 124064
rect 6112 124004 6116 124060
rect 6116 124004 6172 124060
rect 6172 124004 6176 124060
rect 6112 124000 6176 124004
rect 6192 124060 6256 124064
rect 6192 124004 6196 124060
rect 6196 124004 6252 124060
rect 6252 124004 6256 124060
rect 6192 124000 6256 124004
rect 4285 123516 4349 123520
rect 4285 123460 4289 123516
rect 4289 123460 4345 123516
rect 4345 123460 4349 123516
rect 4285 123456 4349 123460
rect 4365 123516 4429 123520
rect 4365 123460 4369 123516
rect 4369 123460 4425 123516
rect 4425 123460 4429 123516
rect 4365 123456 4429 123460
rect 4445 123516 4509 123520
rect 4445 123460 4449 123516
rect 4449 123460 4505 123516
rect 4505 123460 4509 123516
rect 4445 123456 4509 123460
rect 4525 123516 4589 123520
rect 4525 123460 4529 123516
rect 4529 123460 4585 123516
rect 4585 123460 4589 123516
rect 4525 123456 4589 123460
rect 7618 123516 7682 123520
rect 7618 123460 7622 123516
rect 7622 123460 7678 123516
rect 7678 123460 7682 123516
rect 7618 123456 7682 123460
rect 7698 123516 7762 123520
rect 7698 123460 7702 123516
rect 7702 123460 7758 123516
rect 7758 123460 7762 123516
rect 7698 123456 7762 123460
rect 7778 123516 7842 123520
rect 7778 123460 7782 123516
rect 7782 123460 7838 123516
rect 7838 123460 7842 123516
rect 7778 123456 7842 123460
rect 7858 123516 7922 123520
rect 7858 123460 7862 123516
rect 7862 123460 7918 123516
rect 7918 123460 7922 123516
rect 7858 123456 7922 123460
rect 2618 122972 2682 122976
rect 2618 122916 2622 122972
rect 2622 122916 2678 122972
rect 2678 122916 2682 122972
rect 2618 122912 2682 122916
rect 2698 122972 2762 122976
rect 2698 122916 2702 122972
rect 2702 122916 2758 122972
rect 2758 122916 2762 122972
rect 2698 122912 2762 122916
rect 2778 122972 2842 122976
rect 2778 122916 2782 122972
rect 2782 122916 2838 122972
rect 2838 122916 2842 122972
rect 2778 122912 2842 122916
rect 2858 122972 2922 122976
rect 2858 122916 2862 122972
rect 2862 122916 2918 122972
rect 2918 122916 2922 122972
rect 2858 122912 2922 122916
rect 5952 122972 6016 122976
rect 5952 122916 5956 122972
rect 5956 122916 6012 122972
rect 6012 122916 6016 122972
rect 5952 122912 6016 122916
rect 6032 122972 6096 122976
rect 6032 122916 6036 122972
rect 6036 122916 6092 122972
rect 6092 122916 6096 122972
rect 6032 122912 6096 122916
rect 6112 122972 6176 122976
rect 6112 122916 6116 122972
rect 6116 122916 6172 122972
rect 6172 122916 6176 122972
rect 6112 122912 6176 122916
rect 6192 122972 6256 122976
rect 6192 122916 6196 122972
rect 6196 122916 6252 122972
rect 6252 122916 6256 122972
rect 6192 122912 6256 122916
rect 4285 122428 4349 122432
rect 4285 122372 4289 122428
rect 4289 122372 4345 122428
rect 4345 122372 4349 122428
rect 4285 122368 4349 122372
rect 4365 122428 4429 122432
rect 4365 122372 4369 122428
rect 4369 122372 4425 122428
rect 4425 122372 4429 122428
rect 4365 122368 4429 122372
rect 4445 122428 4509 122432
rect 4445 122372 4449 122428
rect 4449 122372 4505 122428
rect 4505 122372 4509 122428
rect 4445 122368 4509 122372
rect 4525 122428 4589 122432
rect 4525 122372 4529 122428
rect 4529 122372 4585 122428
rect 4585 122372 4589 122428
rect 4525 122368 4589 122372
rect 7618 122428 7682 122432
rect 7618 122372 7622 122428
rect 7622 122372 7678 122428
rect 7678 122372 7682 122428
rect 7618 122368 7682 122372
rect 7698 122428 7762 122432
rect 7698 122372 7702 122428
rect 7702 122372 7758 122428
rect 7758 122372 7762 122428
rect 7698 122368 7762 122372
rect 7778 122428 7842 122432
rect 7778 122372 7782 122428
rect 7782 122372 7838 122428
rect 7838 122372 7842 122428
rect 7778 122368 7842 122372
rect 7858 122428 7922 122432
rect 7858 122372 7862 122428
rect 7862 122372 7918 122428
rect 7918 122372 7922 122428
rect 7858 122368 7922 122372
rect 2618 121884 2682 121888
rect 2618 121828 2622 121884
rect 2622 121828 2678 121884
rect 2678 121828 2682 121884
rect 2618 121824 2682 121828
rect 2698 121884 2762 121888
rect 2698 121828 2702 121884
rect 2702 121828 2758 121884
rect 2758 121828 2762 121884
rect 2698 121824 2762 121828
rect 2778 121884 2842 121888
rect 2778 121828 2782 121884
rect 2782 121828 2838 121884
rect 2838 121828 2842 121884
rect 2778 121824 2842 121828
rect 2858 121884 2922 121888
rect 2858 121828 2862 121884
rect 2862 121828 2918 121884
rect 2918 121828 2922 121884
rect 2858 121824 2922 121828
rect 5952 121884 6016 121888
rect 5952 121828 5956 121884
rect 5956 121828 6012 121884
rect 6012 121828 6016 121884
rect 5952 121824 6016 121828
rect 6032 121884 6096 121888
rect 6032 121828 6036 121884
rect 6036 121828 6092 121884
rect 6092 121828 6096 121884
rect 6032 121824 6096 121828
rect 6112 121884 6176 121888
rect 6112 121828 6116 121884
rect 6116 121828 6172 121884
rect 6172 121828 6176 121884
rect 6112 121824 6176 121828
rect 6192 121884 6256 121888
rect 6192 121828 6196 121884
rect 6196 121828 6252 121884
rect 6252 121828 6256 121884
rect 6192 121824 6256 121828
rect 4285 121340 4349 121344
rect 4285 121284 4289 121340
rect 4289 121284 4345 121340
rect 4345 121284 4349 121340
rect 4285 121280 4349 121284
rect 4365 121340 4429 121344
rect 4365 121284 4369 121340
rect 4369 121284 4425 121340
rect 4425 121284 4429 121340
rect 4365 121280 4429 121284
rect 4445 121340 4509 121344
rect 4445 121284 4449 121340
rect 4449 121284 4505 121340
rect 4505 121284 4509 121340
rect 4445 121280 4509 121284
rect 4525 121340 4589 121344
rect 4525 121284 4529 121340
rect 4529 121284 4585 121340
rect 4585 121284 4589 121340
rect 4525 121280 4589 121284
rect 7618 121340 7682 121344
rect 7618 121284 7622 121340
rect 7622 121284 7678 121340
rect 7678 121284 7682 121340
rect 7618 121280 7682 121284
rect 7698 121340 7762 121344
rect 7698 121284 7702 121340
rect 7702 121284 7758 121340
rect 7758 121284 7762 121340
rect 7698 121280 7762 121284
rect 7778 121340 7842 121344
rect 7778 121284 7782 121340
rect 7782 121284 7838 121340
rect 7838 121284 7842 121340
rect 7778 121280 7842 121284
rect 7858 121340 7922 121344
rect 7858 121284 7862 121340
rect 7862 121284 7918 121340
rect 7918 121284 7922 121340
rect 7858 121280 7922 121284
rect 2618 120796 2682 120800
rect 2618 120740 2622 120796
rect 2622 120740 2678 120796
rect 2678 120740 2682 120796
rect 2618 120736 2682 120740
rect 2698 120796 2762 120800
rect 2698 120740 2702 120796
rect 2702 120740 2758 120796
rect 2758 120740 2762 120796
rect 2698 120736 2762 120740
rect 2778 120796 2842 120800
rect 2778 120740 2782 120796
rect 2782 120740 2838 120796
rect 2838 120740 2842 120796
rect 2778 120736 2842 120740
rect 2858 120796 2922 120800
rect 2858 120740 2862 120796
rect 2862 120740 2918 120796
rect 2918 120740 2922 120796
rect 2858 120736 2922 120740
rect 5952 120796 6016 120800
rect 5952 120740 5956 120796
rect 5956 120740 6012 120796
rect 6012 120740 6016 120796
rect 5952 120736 6016 120740
rect 6032 120796 6096 120800
rect 6032 120740 6036 120796
rect 6036 120740 6092 120796
rect 6092 120740 6096 120796
rect 6032 120736 6096 120740
rect 6112 120796 6176 120800
rect 6112 120740 6116 120796
rect 6116 120740 6172 120796
rect 6172 120740 6176 120796
rect 6112 120736 6176 120740
rect 6192 120796 6256 120800
rect 6192 120740 6196 120796
rect 6196 120740 6252 120796
rect 6252 120740 6256 120796
rect 6192 120736 6256 120740
rect 4285 120252 4349 120256
rect 4285 120196 4289 120252
rect 4289 120196 4345 120252
rect 4345 120196 4349 120252
rect 4285 120192 4349 120196
rect 4365 120252 4429 120256
rect 4365 120196 4369 120252
rect 4369 120196 4425 120252
rect 4425 120196 4429 120252
rect 4365 120192 4429 120196
rect 4445 120252 4509 120256
rect 4445 120196 4449 120252
rect 4449 120196 4505 120252
rect 4505 120196 4509 120252
rect 4445 120192 4509 120196
rect 4525 120252 4589 120256
rect 4525 120196 4529 120252
rect 4529 120196 4585 120252
rect 4585 120196 4589 120252
rect 4525 120192 4589 120196
rect 7618 120252 7682 120256
rect 7618 120196 7622 120252
rect 7622 120196 7678 120252
rect 7678 120196 7682 120252
rect 7618 120192 7682 120196
rect 7698 120252 7762 120256
rect 7698 120196 7702 120252
rect 7702 120196 7758 120252
rect 7758 120196 7762 120252
rect 7698 120192 7762 120196
rect 7778 120252 7842 120256
rect 7778 120196 7782 120252
rect 7782 120196 7838 120252
rect 7838 120196 7842 120252
rect 7778 120192 7842 120196
rect 7858 120252 7922 120256
rect 7858 120196 7862 120252
rect 7862 120196 7918 120252
rect 7918 120196 7922 120252
rect 7858 120192 7922 120196
rect 2618 119708 2682 119712
rect 2618 119652 2622 119708
rect 2622 119652 2678 119708
rect 2678 119652 2682 119708
rect 2618 119648 2682 119652
rect 2698 119708 2762 119712
rect 2698 119652 2702 119708
rect 2702 119652 2758 119708
rect 2758 119652 2762 119708
rect 2698 119648 2762 119652
rect 2778 119708 2842 119712
rect 2778 119652 2782 119708
rect 2782 119652 2838 119708
rect 2838 119652 2842 119708
rect 2778 119648 2842 119652
rect 2858 119708 2922 119712
rect 2858 119652 2862 119708
rect 2862 119652 2918 119708
rect 2918 119652 2922 119708
rect 2858 119648 2922 119652
rect 5952 119708 6016 119712
rect 5952 119652 5956 119708
rect 5956 119652 6012 119708
rect 6012 119652 6016 119708
rect 5952 119648 6016 119652
rect 6032 119708 6096 119712
rect 6032 119652 6036 119708
rect 6036 119652 6092 119708
rect 6092 119652 6096 119708
rect 6032 119648 6096 119652
rect 6112 119708 6176 119712
rect 6112 119652 6116 119708
rect 6116 119652 6172 119708
rect 6172 119652 6176 119708
rect 6112 119648 6176 119652
rect 6192 119708 6256 119712
rect 6192 119652 6196 119708
rect 6196 119652 6252 119708
rect 6252 119652 6256 119708
rect 6192 119648 6256 119652
rect 4285 119164 4349 119168
rect 4285 119108 4289 119164
rect 4289 119108 4345 119164
rect 4345 119108 4349 119164
rect 4285 119104 4349 119108
rect 4365 119164 4429 119168
rect 4365 119108 4369 119164
rect 4369 119108 4425 119164
rect 4425 119108 4429 119164
rect 4365 119104 4429 119108
rect 4445 119164 4509 119168
rect 4445 119108 4449 119164
rect 4449 119108 4505 119164
rect 4505 119108 4509 119164
rect 4445 119104 4509 119108
rect 4525 119164 4589 119168
rect 4525 119108 4529 119164
rect 4529 119108 4585 119164
rect 4585 119108 4589 119164
rect 4525 119104 4589 119108
rect 7618 119164 7682 119168
rect 7618 119108 7622 119164
rect 7622 119108 7678 119164
rect 7678 119108 7682 119164
rect 7618 119104 7682 119108
rect 7698 119164 7762 119168
rect 7698 119108 7702 119164
rect 7702 119108 7758 119164
rect 7758 119108 7762 119164
rect 7698 119104 7762 119108
rect 7778 119164 7842 119168
rect 7778 119108 7782 119164
rect 7782 119108 7838 119164
rect 7838 119108 7842 119164
rect 7778 119104 7842 119108
rect 7858 119164 7922 119168
rect 7858 119108 7862 119164
rect 7862 119108 7918 119164
rect 7918 119108 7922 119164
rect 7858 119104 7922 119108
rect 2618 118620 2682 118624
rect 2618 118564 2622 118620
rect 2622 118564 2678 118620
rect 2678 118564 2682 118620
rect 2618 118560 2682 118564
rect 2698 118620 2762 118624
rect 2698 118564 2702 118620
rect 2702 118564 2758 118620
rect 2758 118564 2762 118620
rect 2698 118560 2762 118564
rect 2778 118620 2842 118624
rect 2778 118564 2782 118620
rect 2782 118564 2838 118620
rect 2838 118564 2842 118620
rect 2778 118560 2842 118564
rect 2858 118620 2922 118624
rect 2858 118564 2862 118620
rect 2862 118564 2918 118620
rect 2918 118564 2922 118620
rect 2858 118560 2922 118564
rect 5952 118620 6016 118624
rect 5952 118564 5956 118620
rect 5956 118564 6012 118620
rect 6012 118564 6016 118620
rect 5952 118560 6016 118564
rect 6032 118620 6096 118624
rect 6032 118564 6036 118620
rect 6036 118564 6092 118620
rect 6092 118564 6096 118620
rect 6032 118560 6096 118564
rect 6112 118620 6176 118624
rect 6112 118564 6116 118620
rect 6116 118564 6172 118620
rect 6172 118564 6176 118620
rect 6112 118560 6176 118564
rect 6192 118620 6256 118624
rect 6192 118564 6196 118620
rect 6196 118564 6252 118620
rect 6252 118564 6256 118620
rect 6192 118560 6256 118564
rect 4285 118076 4349 118080
rect 4285 118020 4289 118076
rect 4289 118020 4345 118076
rect 4345 118020 4349 118076
rect 4285 118016 4349 118020
rect 4365 118076 4429 118080
rect 4365 118020 4369 118076
rect 4369 118020 4425 118076
rect 4425 118020 4429 118076
rect 4365 118016 4429 118020
rect 4445 118076 4509 118080
rect 4445 118020 4449 118076
rect 4449 118020 4505 118076
rect 4505 118020 4509 118076
rect 4445 118016 4509 118020
rect 4525 118076 4589 118080
rect 4525 118020 4529 118076
rect 4529 118020 4585 118076
rect 4585 118020 4589 118076
rect 4525 118016 4589 118020
rect 7618 118076 7682 118080
rect 7618 118020 7622 118076
rect 7622 118020 7678 118076
rect 7678 118020 7682 118076
rect 7618 118016 7682 118020
rect 7698 118076 7762 118080
rect 7698 118020 7702 118076
rect 7702 118020 7758 118076
rect 7758 118020 7762 118076
rect 7698 118016 7762 118020
rect 7778 118076 7842 118080
rect 7778 118020 7782 118076
rect 7782 118020 7838 118076
rect 7838 118020 7842 118076
rect 7778 118016 7842 118020
rect 7858 118076 7922 118080
rect 7858 118020 7862 118076
rect 7862 118020 7918 118076
rect 7918 118020 7922 118076
rect 7858 118016 7922 118020
rect 2618 117532 2682 117536
rect 2618 117476 2622 117532
rect 2622 117476 2678 117532
rect 2678 117476 2682 117532
rect 2618 117472 2682 117476
rect 2698 117532 2762 117536
rect 2698 117476 2702 117532
rect 2702 117476 2758 117532
rect 2758 117476 2762 117532
rect 2698 117472 2762 117476
rect 2778 117532 2842 117536
rect 2778 117476 2782 117532
rect 2782 117476 2838 117532
rect 2838 117476 2842 117532
rect 2778 117472 2842 117476
rect 2858 117532 2922 117536
rect 2858 117476 2862 117532
rect 2862 117476 2918 117532
rect 2918 117476 2922 117532
rect 2858 117472 2922 117476
rect 5952 117532 6016 117536
rect 5952 117476 5956 117532
rect 5956 117476 6012 117532
rect 6012 117476 6016 117532
rect 5952 117472 6016 117476
rect 6032 117532 6096 117536
rect 6032 117476 6036 117532
rect 6036 117476 6092 117532
rect 6092 117476 6096 117532
rect 6032 117472 6096 117476
rect 6112 117532 6176 117536
rect 6112 117476 6116 117532
rect 6116 117476 6172 117532
rect 6172 117476 6176 117532
rect 6112 117472 6176 117476
rect 6192 117532 6256 117536
rect 6192 117476 6196 117532
rect 6196 117476 6252 117532
rect 6252 117476 6256 117532
rect 6192 117472 6256 117476
rect 4285 116988 4349 116992
rect 4285 116932 4289 116988
rect 4289 116932 4345 116988
rect 4345 116932 4349 116988
rect 4285 116928 4349 116932
rect 4365 116988 4429 116992
rect 4365 116932 4369 116988
rect 4369 116932 4425 116988
rect 4425 116932 4429 116988
rect 4365 116928 4429 116932
rect 4445 116988 4509 116992
rect 4445 116932 4449 116988
rect 4449 116932 4505 116988
rect 4505 116932 4509 116988
rect 4445 116928 4509 116932
rect 4525 116988 4589 116992
rect 4525 116932 4529 116988
rect 4529 116932 4585 116988
rect 4585 116932 4589 116988
rect 4525 116928 4589 116932
rect 7618 116988 7682 116992
rect 7618 116932 7622 116988
rect 7622 116932 7678 116988
rect 7678 116932 7682 116988
rect 7618 116928 7682 116932
rect 7698 116988 7762 116992
rect 7698 116932 7702 116988
rect 7702 116932 7758 116988
rect 7758 116932 7762 116988
rect 7698 116928 7762 116932
rect 7778 116988 7842 116992
rect 7778 116932 7782 116988
rect 7782 116932 7838 116988
rect 7838 116932 7842 116988
rect 7778 116928 7842 116932
rect 7858 116988 7922 116992
rect 7858 116932 7862 116988
rect 7862 116932 7918 116988
rect 7918 116932 7922 116988
rect 7858 116928 7922 116932
rect 2618 116444 2682 116448
rect 2618 116388 2622 116444
rect 2622 116388 2678 116444
rect 2678 116388 2682 116444
rect 2618 116384 2682 116388
rect 2698 116444 2762 116448
rect 2698 116388 2702 116444
rect 2702 116388 2758 116444
rect 2758 116388 2762 116444
rect 2698 116384 2762 116388
rect 2778 116444 2842 116448
rect 2778 116388 2782 116444
rect 2782 116388 2838 116444
rect 2838 116388 2842 116444
rect 2778 116384 2842 116388
rect 2858 116444 2922 116448
rect 2858 116388 2862 116444
rect 2862 116388 2918 116444
rect 2918 116388 2922 116444
rect 2858 116384 2922 116388
rect 5952 116444 6016 116448
rect 5952 116388 5956 116444
rect 5956 116388 6012 116444
rect 6012 116388 6016 116444
rect 5952 116384 6016 116388
rect 6032 116444 6096 116448
rect 6032 116388 6036 116444
rect 6036 116388 6092 116444
rect 6092 116388 6096 116444
rect 6032 116384 6096 116388
rect 6112 116444 6176 116448
rect 6112 116388 6116 116444
rect 6116 116388 6172 116444
rect 6172 116388 6176 116444
rect 6112 116384 6176 116388
rect 6192 116444 6256 116448
rect 6192 116388 6196 116444
rect 6196 116388 6252 116444
rect 6252 116388 6256 116444
rect 6192 116384 6256 116388
rect 4285 115900 4349 115904
rect 4285 115844 4289 115900
rect 4289 115844 4345 115900
rect 4345 115844 4349 115900
rect 4285 115840 4349 115844
rect 4365 115900 4429 115904
rect 4365 115844 4369 115900
rect 4369 115844 4425 115900
rect 4425 115844 4429 115900
rect 4365 115840 4429 115844
rect 4445 115900 4509 115904
rect 4445 115844 4449 115900
rect 4449 115844 4505 115900
rect 4505 115844 4509 115900
rect 4445 115840 4509 115844
rect 4525 115900 4589 115904
rect 4525 115844 4529 115900
rect 4529 115844 4585 115900
rect 4585 115844 4589 115900
rect 4525 115840 4589 115844
rect 7618 115900 7682 115904
rect 7618 115844 7622 115900
rect 7622 115844 7678 115900
rect 7678 115844 7682 115900
rect 7618 115840 7682 115844
rect 7698 115900 7762 115904
rect 7698 115844 7702 115900
rect 7702 115844 7758 115900
rect 7758 115844 7762 115900
rect 7698 115840 7762 115844
rect 7778 115900 7842 115904
rect 7778 115844 7782 115900
rect 7782 115844 7838 115900
rect 7838 115844 7842 115900
rect 7778 115840 7842 115844
rect 7858 115900 7922 115904
rect 7858 115844 7862 115900
rect 7862 115844 7918 115900
rect 7918 115844 7922 115900
rect 7858 115840 7922 115844
rect 2618 115356 2682 115360
rect 2618 115300 2622 115356
rect 2622 115300 2678 115356
rect 2678 115300 2682 115356
rect 2618 115296 2682 115300
rect 2698 115356 2762 115360
rect 2698 115300 2702 115356
rect 2702 115300 2758 115356
rect 2758 115300 2762 115356
rect 2698 115296 2762 115300
rect 2778 115356 2842 115360
rect 2778 115300 2782 115356
rect 2782 115300 2838 115356
rect 2838 115300 2842 115356
rect 2778 115296 2842 115300
rect 2858 115356 2922 115360
rect 2858 115300 2862 115356
rect 2862 115300 2918 115356
rect 2918 115300 2922 115356
rect 2858 115296 2922 115300
rect 5952 115356 6016 115360
rect 5952 115300 5956 115356
rect 5956 115300 6012 115356
rect 6012 115300 6016 115356
rect 5952 115296 6016 115300
rect 6032 115356 6096 115360
rect 6032 115300 6036 115356
rect 6036 115300 6092 115356
rect 6092 115300 6096 115356
rect 6032 115296 6096 115300
rect 6112 115356 6176 115360
rect 6112 115300 6116 115356
rect 6116 115300 6172 115356
rect 6172 115300 6176 115356
rect 6112 115296 6176 115300
rect 6192 115356 6256 115360
rect 6192 115300 6196 115356
rect 6196 115300 6252 115356
rect 6252 115300 6256 115356
rect 6192 115296 6256 115300
rect 4285 114812 4349 114816
rect 4285 114756 4289 114812
rect 4289 114756 4345 114812
rect 4345 114756 4349 114812
rect 4285 114752 4349 114756
rect 4365 114812 4429 114816
rect 4365 114756 4369 114812
rect 4369 114756 4425 114812
rect 4425 114756 4429 114812
rect 4365 114752 4429 114756
rect 4445 114812 4509 114816
rect 4445 114756 4449 114812
rect 4449 114756 4505 114812
rect 4505 114756 4509 114812
rect 4445 114752 4509 114756
rect 4525 114812 4589 114816
rect 4525 114756 4529 114812
rect 4529 114756 4585 114812
rect 4585 114756 4589 114812
rect 4525 114752 4589 114756
rect 7618 114812 7682 114816
rect 7618 114756 7622 114812
rect 7622 114756 7678 114812
rect 7678 114756 7682 114812
rect 7618 114752 7682 114756
rect 7698 114812 7762 114816
rect 7698 114756 7702 114812
rect 7702 114756 7758 114812
rect 7758 114756 7762 114812
rect 7698 114752 7762 114756
rect 7778 114812 7842 114816
rect 7778 114756 7782 114812
rect 7782 114756 7838 114812
rect 7838 114756 7842 114812
rect 7778 114752 7842 114756
rect 7858 114812 7922 114816
rect 7858 114756 7862 114812
rect 7862 114756 7918 114812
rect 7918 114756 7922 114812
rect 7858 114752 7922 114756
rect 2618 114268 2682 114272
rect 2618 114212 2622 114268
rect 2622 114212 2678 114268
rect 2678 114212 2682 114268
rect 2618 114208 2682 114212
rect 2698 114268 2762 114272
rect 2698 114212 2702 114268
rect 2702 114212 2758 114268
rect 2758 114212 2762 114268
rect 2698 114208 2762 114212
rect 2778 114268 2842 114272
rect 2778 114212 2782 114268
rect 2782 114212 2838 114268
rect 2838 114212 2842 114268
rect 2778 114208 2842 114212
rect 2858 114268 2922 114272
rect 2858 114212 2862 114268
rect 2862 114212 2918 114268
rect 2918 114212 2922 114268
rect 2858 114208 2922 114212
rect 5952 114268 6016 114272
rect 5952 114212 5956 114268
rect 5956 114212 6012 114268
rect 6012 114212 6016 114268
rect 5952 114208 6016 114212
rect 6032 114268 6096 114272
rect 6032 114212 6036 114268
rect 6036 114212 6092 114268
rect 6092 114212 6096 114268
rect 6032 114208 6096 114212
rect 6112 114268 6176 114272
rect 6112 114212 6116 114268
rect 6116 114212 6172 114268
rect 6172 114212 6176 114268
rect 6112 114208 6176 114212
rect 6192 114268 6256 114272
rect 6192 114212 6196 114268
rect 6196 114212 6252 114268
rect 6252 114212 6256 114268
rect 6192 114208 6256 114212
rect 4285 113724 4349 113728
rect 4285 113668 4289 113724
rect 4289 113668 4345 113724
rect 4345 113668 4349 113724
rect 4285 113664 4349 113668
rect 4365 113724 4429 113728
rect 4365 113668 4369 113724
rect 4369 113668 4425 113724
rect 4425 113668 4429 113724
rect 4365 113664 4429 113668
rect 4445 113724 4509 113728
rect 4445 113668 4449 113724
rect 4449 113668 4505 113724
rect 4505 113668 4509 113724
rect 4445 113664 4509 113668
rect 4525 113724 4589 113728
rect 4525 113668 4529 113724
rect 4529 113668 4585 113724
rect 4585 113668 4589 113724
rect 4525 113664 4589 113668
rect 7618 113724 7682 113728
rect 7618 113668 7622 113724
rect 7622 113668 7678 113724
rect 7678 113668 7682 113724
rect 7618 113664 7682 113668
rect 7698 113724 7762 113728
rect 7698 113668 7702 113724
rect 7702 113668 7758 113724
rect 7758 113668 7762 113724
rect 7698 113664 7762 113668
rect 7778 113724 7842 113728
rect 7778 113668 7782 113724
rect 7782 113668 7838 113724
rect 7838 113668 7842 113724
rect 7778 113664 7842 113668
rect 7858 113724 7922 113728
rect 7858 113668 7862 113724
rect 7862 113668 7918 113724
rect 7918 113668 7922 113724
rect 7858 113664 7922 113668
rect 2618 113180 2682 113184
rect 2618 113124 2622 113180
rect 2622 113124 2678 113180
rect 2678 113124 2682 113180
rect 2618 113120 2682 113124
rect 2698 113180 2762 113184
rect 2698 113124 2702 113180
rect 2702 113124 2758 113180
rect 2758 113124 2762 113180
rect 2698 113120 2762 113124
rect 2778 113180 2842 113184
rect 2778 113124 2782 113180
rect 2782 113124 2838 113180
rect 2838 113124 2842 113180
rect 2778 113120 2842 113124
rect 2858 113180 2922 113184
rect 2858 113124 2862 113180
rect 2862 113124 2918 113180
rect 2918 113124 2922 113180
rect 2858 113120 2922 113124
rect 5952 113180 6016 113184
rect 5952 113124 5956 113180
rect 5956 113124 6012 113180
rect 6012 113124 6016 113180
rect 5952 113120 6016 113124
rect 6032 113180 6096 113184
rect 6032 113124 6036 113180
rect 6036 113124 6092 113180
rect 6092 113124 6096 113180
rect 6032 113120 6096 113124
rect 6112 113180 6176 113184
rect 6112 113124 6116 113180
rect 6116 113124 6172 113180
rect 6172 113124 6176 113180
rect 6112 113120 6176 113124
rect 6192 113180 6256 113184
rect 6192 113124 6196 113180
rect 6196 113124 6252 113180
rect 6252 113124 6256 113180
rect 6192 113120 6256 113124
rect 4285 112636 4349 112640
rect 4285 112580 4289 112636
rect 4289 112580 4345 112636
rect 4345 112580 4349 112636
rect 4285 112576 4349 112580
rect 4365 112636 4429 112640
rect 4365 112580 4369 112636
rect 4369 112580 4425 112636
rect 4425 112580 4429 112636
rect 4365 112576 4429 112580
rect 4445 112636 4509 112640
rect 4445 112580 4449 112636
rect 4449 112580 4505 112636
rect 4505 112580 4509 112636
rect 4445 112576 4509 112580
rect 4525 112636 4589 112640
rect 4525 112580 4529 112636
rect 4529 112580 4585 112636
rect 4585 112580 4589 112636
rect 4525 112576 4589 112580
rect 7618 112636 7682 112640
rect 7618 112580 7622 112636
rect 7622 112580 7678 112636
rect 7678 112580 7682 112636
rect 7618 112576 7682 112580
rect 7698 112636 7762 112640
rect 7698 112580 7702 112636
rect 7702 112580 7758 112636
rect 7758 112580 7762 112636
rect 7698 112576 7762 112580
rect 7778 112636 7842 112640
rect 7778 112580 7782 112636
rect 7782 112580 7838 112636
rect 7838 112580 7842 112636
rect 7778 112576 7842 112580
rect 7858 112636 7922 112640
rect 7858 112580 7862 112636
rect 7862 112580 7918 112636
rect 7918 112580 7922 112636
rect 7858 112576 7922 112580
rect 2618 112092 2682 112096
rect 2618 112036 2622 112092
rect 2622 112036 2678 112092
rect 2678 112036 2682 112092
rect 2618 112032 2682 112036
rect 2698 112092 2762 112096
rect 2698 112036 2702 112092
rect 2702 112036 2758 112092
rect 2758 112036 2762 112092
rect 2698 112032 2762 112036
rect 2778 112092 2842 112096
rect 2778 112036 2782 112092
rect 2782 112036 2838 112092
rect 2838 112036 2842 112092
rect 2778 112032 2842 112036
rect 2858 112092 2922 112096
rect 2858 112036 2862 112092
rect 2862 112036 2918 112092
rect 2918 112036 2922 112092
rect 2858 112032 2922 112036
rect 5952 112092 6016 112096
rect 5952 112036 5956 112092
rect 5956 112036 6012 112092
rect 6012 112036 6016 112092
rect 5952 112032 6016 112036
rect 6032 112092 6096 112096
rect 6032 112036 6036 112092
rect 6036 112036 6092 112092
rect 6092 112036 6096 112092
rect 6032 112032 6096 112036
rect 6112 112092 6176 112096
rect 6112 112036 6116 112092
rect 6116 112036 6172 112092
rect 6172 112036 6176 112092
rect 6112 112032 6176 112036
rect 6192 112092 6256 112096
rect 6192 112036 6196 112092
rect 6196 112036 6252 112092
rect 6252 112036 6256 112092
rect 6192 112032 6256 112036
rect 4285 111548 4349 111552
rect 4285 111492 4289 111548
rect 4289 111492 4345 111548
rect 4345 111492 4349 111548
rect 4285 111488 4349 111492
rect 4365 111548 4429 111552
rect 4365 111492 4369 111548
rect 4369 111492 4425 111548
rect 4425 111492 4429 111548
rect 4365 111488 4429 111492
rect 4445 111548 4509 111552
rect 4445 111492 4449 111548
rect 4449 111492 4505 111548
rect 4505 111492 4509 111548
rect 4445 111488 4509 111492
rect 4525 111548 4589 111552
rect 4525 111492 4529 111548
rect 4529 111492 4585 111548
rect 4585 111492 4589 111548
rect 4525 111488 4589 111492
rect 7618 111548 7682 111552
rect 7618 111492 7622 111548
rect 7622 111492 7678 111548
rect 7678 111492 7682 111548
rect 7618 111488 7682 111492
rect 7698 111548 7762 111552
rect 7698 111492 7702 111548
rect 7702 111492 7758 111548
rect 7758 111492 7762 111548
rect 7698 111488 7762 111492
rect 7778 111548 7842 111552
rect 7778 111492 7782 111548
rect 7782 111492 7838 111548
rect 7838 111492 7842 111548
rect 7778 111488 7842 111492
rect 7858 111548 7922 111552
rect 7858 111492 7862 111548
rect 7862 111492 7918 111548
rect 7918 111492 7922 111548
rect 7858 111488 7922 111492
rect 2618 111004 2682 111008
rect 2618 110948 2622 111004
rect 2622 110948 2678 111004
rect 2678 110948 2682 111004
rect 2618 110944 2682 110948
rect 2698 111004 2762 111008
rect 2698 110948 2702 111004
rect 2702 110948 2758 111004
rect 2758 110948 2762 111004
rect 2698 110944 2762 110948
rect 2778 111004 2842 111008
rect 2778 110948 2782 111004
rect 2782 110948 2838 111004
rect 2838 110948 2842 111004
rect 2778 110944 2842 110948
rect 2858 111004 2922 111008
rect 2858 110948 2862 111004
rect 2862 110948 2918 111004
rect 2918 110948 2922 111004
rect 2858 110944 2922 110948
rect 5952 111004 6016 111008
rect 5952 110948 5956 111004
rect 5956 110948 6012 111004
rect 6012 110948 6016 111004
rect 5952 110944 6016 110948
rect 6032 111004 6096 111008
rect 6032 110948 6036 111004
rect 6036 110948 6092 111004
rect 6092 110948 6096 111004
rect 6032 110944 6096 110948
rect 6112 111004 6176 111008
rect 6112 110948 6116 111004
rect 6116 110948 6172 111004
rect 6172 110948 6176 111004
rect 6112 110944 6176 110948
rect 6192 111004 6256 111008
rect 6192 110948 6196 111004
rect 6196 110948 6252 111004
rect 6252 110948 6256 111004
rect 6192 110944 6256 110948
rect 4285 110460 4349 110464
rect 4285 110404 4289 110460
rect 4289 110404 4345 110460
rect 4345 110404 4349 110460
rect 4285 110400 4349 110404
rect 4365 110460 4429 110464
rect 4365 110404 4369 110460
rect 4369 110404 4425 110460
rect 4425 110404 4429 110460
rect 4365 110400 4429 110404
rect 4445 110460 4509 110464
rect 4445 110404 4449 110460
rect 4449 110404 4505 110460
rect 4505 110404 4509 110460
rect 4445 110400 4509 110404
rect 4525 110460 4589 110464
rect 4525 110404 4529 110460
rect 4529 110404 4585 110460
rect 4585 110404 4589 110460
rect 4525 110400 4589 110404
rect 7618 110460 7682 110464
rect 7618 110404 7622 110460
rect 7622 110404 7678 110460
rect 7678 110404 7682 110460
rect 7618 110400 7682 110404
rect 7698 110460 7762 110464
rect 7698 110404 7702 110460
rect 7702 110404 7758 110460
rect 7758 110404 7762 110460
rect 7698 110400 7762 110404
rect 7778 110460 7842 110464
rect 7778 110404 7782 110460
rect 7782 110404 7838 110460
rect 7838 110404 7842 110460
rect 7778 110400 7842 110404
rect 7858 110460 7922 110464
rect 7858 110404 7862 110460
rect 7862 110404 7918 110460
rect 7918 110404 7922 110460
rect 7858 110400 7922 110404
rect 2618 109916 2682 109920
rect 2618 109860 2622 109916
rect 2622 109860 2678 109916
rect 2678 109860 2682 109916
rect 2618 109856 2682 109860
rect 2698 109916 2762 109920
rect 2698 109860 2702 109916
rect 2702 109860 2758 109916
rect 2758 109860 2762 109916
rect 2698 109856 2762 109860
rect 2778 109916 2842 109920
rect 2778 109860 2782 109916
rect 2782 109860 2838 109916
rect 2838 109860 2842 109916
rect 2778 109856 2842 109860
rect 2858 109916 2922 109920
rect 2858 109860 2862 109916
rect 2862 109860 2918 109916
rect 2918 109860 2922 109916
rect 2858 109856 2922 109860
rect 5952 109916 6016 109920
rect 5952 109860 5956 109916
rect 5956 109860 6012 109916
rect 6012 109860 6016 109916
rect 5952 109856 6016 109860
rect 6032 109916 6096 109920
rect 6032 109860 6036 109916
rect 6036 109860 6092 109916
rect 6092 109860 6096 109916
rect 6032 109856 6096 109860
rect 6112 109916 6176 109920
rect 6112 109860 6116 109916
rect 6116 109860 6172 109916
rect 6172 109860 6176 109916
rect 6112 109856 6176 109860
rect 6192 109916 6256 109920
rect 6192 109860 6196 109916
rect 6196 109860 6252 109916
rect 6252 109860 6256 109916
rect 6192 109856 6256 109860
rect 4285 109372 4349 109376
rect 4285 109316 4289 109372
rect 4289 109316 4345 109372
rect 4345 109316 4349 109372
rect 4285 109312 4349 109316
rect 4365 109372 4429 109376
rect 4365 109316 4369 109372
rect 4369 109316 4425 109372
rect 4425 109316 4429 109372
rect 4365 109312 4429 109316
rect 4445 109372 4509 109376
rect 4445 109316 4449 109372
rect 4449 109316 4505 109372
rect 4505 109316 4509 109372
rect 4445 109312 4509 109316
rect 4525 109372 4589 109376
rect 4525 109316 4529 109372
rect 4529 109316 4585 109372
rect 4585 109316 4589 109372
rect 4525 109312 4589 109316
rect 7618 109372 7682 109376
rect 7618 109316 7622 109372
rect 7622 109316 7678 109372
rect 7678 109316 7682 109372
rect 7618 109312 7682 109316
rect 7698 109372 7762 109376
rect 7698 109316 7702 109372
rect 7702 109316 7758 109372
rect 7758 109316 7762 109372
rect 7698 109312 7762 109316
rect 7778 109372 7842 109376
rect 7778 109316 7782 109372
rect 7782 109316 7838 109372
rect 7838 109316 7842 109372
rect 7778 109312 7842 109316
rect 7858 109372 7922 109376
rect 7858 109316 7862 109372
rect 7862 109316 7918 109372
rect 7918 109316 7922 109372
rect 7858 109312 7922 109316
rect 2618 108828 2682 108832
rect 2618 108772 2622 108828
rect 2622 108772 2678 108828
rect 2678 108772 2682 108828
rect 2618 108768 2682 108772
rect 2698 108828 2762 108832
rect 2698 108772 2702 108828
rect 2702 108772 2758 108828
rect 2758 108772 2762 108828
rect 2698 108768 2762 108772
rect 2778 108828 2842 108832
rect 2778 108772 2782 108828
rect 2782 108772 2838 108828
rect 2838 108772 2842 108828
rect 2778 108768 2842 108772
rect 2858 108828 2922 108832
rect 2858 108772 2862 108828
rect 2862 108772 2918 108828
rect 2918 108772 2922 108828
rect 2858 108768 2922 108772
rect 5952 108828 6016 108832
rect 5952 108772 5956 108828
rect 5956 108772 6012 108828
rect 6012 108772 6016 108828
rect 5952 108768 6016 108772
rect 6032 108828 6096 108832
rect 6032 108772 6036 108828
rect 6036 108772 6092 108828
rect 6092 108772 6096 108828
rect 6032 108768 6096 108772
rect 6112 108828 6176 108832
rect 6112 108772 6116 108828
rect 6116 108772 6172 108828
rect 6172 108772 6176 108828
rect 6112 108768 6176 108772
rect 6192 108828 6256 108832
rect 6192 108772 6196 108828
rect 6196 108772 6252 108828
rect 6252 108772 6256 108828
rect 6192 108768 6256 108772
rect 4285 108284 4349 108288
rect 4285 108228 4289 108284
rect 4289 108228 4345 108284
rect 4345 108228 4349 108284
rect 4285 108224 4349 108228
rect 4365 108284 4429 108288
rect 4365 108228 4369 108284
rect 4369 108228 4425 108284
rect 4425 108228 4429 108284
rect 4365 108224 4429 108228
rect 4445 108284 4509 108288
rect 4445 108228 4449 108284
rect 4449 108228 4505 108284
rect 4505 108228 4509 108284
rect 4445 108224 4509 108228
rect 4525 108284 4589 108288
rect 4525 108228 4529 108284
rect 4529 108228 4585 108284
rect 4585 108228 4589 108284
rect 4525 108224 4589 108228
rect 7618 108284 7682 108288
rect 7618 108228 7622 108284
rect 7622 108228 7678 108284
rect 7678 108228 7682 108284
rect 7618 108224 7682 108228
rect 7698 108284 7762 108288
rect 7698 108228 7702 108284
rect 7702 108228 7758 108284
rect 7758 108228 7762 108284
rect 7698 108224 7762 108228
rect 7778 108284 7842 108288
rect 7778 108228 7782 108284
rect 7782 108228 7838 108284
rect 7838 108228 7842 108284
rect 7778 108224 7842 108228
rect 7858 108284 7922 108288
rect 7858 108228 7862 108284
rect 7862 108228 7918 108284
rect 7918 108228 7922 108284
rect 7858 108224 7922 108228
rect 2618 107740 2682 107744
rect 2618 107684 2622 107740
rect 2622 107684 2678 107740
rect 2678 107684 2682 107740
rect 2618 107680 2682 107684
rect 2698 107740 2762 107744
rect 2698 107684 2702 107740
rect 2702 107684 2758 107740
rect 2758 107684 2762 107740
rect 2698 107680 2762 107684
rect 2778 107740 2842 107744
rect 2778 107684 2782 107740
rect 2782 107684 2838 107740
rect 2838 107684 2842 107740
rect 2778 107680 2842 107684
rect 2858 107740 2922 107744
rect 2858 107684 2862 107740
rect 2862 107684 2918 107740
rect 2918 107684 2922 107740
rect 2858 107680 2922 107684
rect 5952 107740 6016 107744
rect 5952 107684 5956 107740
rect 5956 107684 6012 107740
rect 6012 107684 6016 107740
rect 5952 107680 6016 107684
rect 6032 107740 6096 107744
rect 6032 107684 6036 107740
rect 6036 107684 6092 107740
rect 6092 107684 6096 107740
rect 6032 107680 6096 107684
rect 6112 107740 6176 107744
rect 6112 107684 6116 107740
rect 6116 107684 6172 107740
rect 6172 107684 6176 107740
rect 6112 107680 6176 107684
rect 6192 107740 6256 107744
rect 6192 107684 6196 107740
rect 6196 107684 6252 107740
rect 6252 107684 6256 107740
rect 6192 107680 6256 107684
rect 4285 107196 4349 107200
rect 4285 107140 4289 107196
rect 4289 107140 4345 107196
rect 4345 107140 4349 107196
rect 4285 107136 4349 107140
rect 4365 107196 4429 107200
rect 4365 107140 4369 107196
rect 4369 107140 4425 107196
rect 4425 107140 4429 107196
rect 4365 107136 4429 107140
rect 4445 107196 4509 107200
rect 4445 107140 4449 107196
rect 4449 107140 4505 107196
rect 4505 107140 4509 107196
rect 4445 107136 4509 107140
rect 4525 107196 4589 107200
rect 4525 107140 4529 107196
rect 4529 107140 4585 107196
rect 4585 107140 4589 107196
rect 4525 107136 4589 107140
rect 7618 107196 7682 107200
rect 7618 107140 7622 107196
rect 7622 107140 7678 107196
rect 7678 107140 7682 107196
rect 7618 107136 7682 107140
rect 7698 107196 7762 107200
rect 7698 107140 7702 107196
rect 7702 107140 7758 107196
rect 7758 107140 7762 107196
rect 7698 107136 7762 107140
rect 7778 107196 7842 107200
rect 7778 107140 7782 107196
rect 7782 107140 7838 107196
rect 7838 107140 7842 107196
rect 7778 107136 7842 107140
rect 7858 107196 7922 107200
rect 7858 107140 7862 107196
rect 7862 107140 7918 107196
rect 7918 107140 7922 107196
rect 7858 107136 7922 107140
rect 2618 106652 2682 106656
rect 2618 106596 2622 106652
rect 2622 106596 2678 106652
rect 2678 106596 2682 106652
rect 2618 106592 2682 106596
rect 2698 106652 2762 106656
rect 2698 106596 2702 106652
rect 2702 106596 2758 106652
rect 2758 106596 2762 106652
rect 2698 106592 2762 106596
rect 2778 106652 2842 106656
rect 2778 106596 2782 106652
rect 2782 106596 2838 106652
rect 2838 106596 2842 106652
rect 2778 106592 2842 106596
rect 2858 106652 2922 106656
rect 2858 106596 2862 106652
rect 2862 106596 2918 106652
rect 2918 106596 2922 106652
rect 2858 106592 2922 106596
rect 5952 106652 6016 106656
rect 5952 106596 5956 106652
rect 5956 106596 6012 106652
rect 6012 106596 6016 106652
rect 5952 106592 6016 106596
rect 6032 106652 6096 106656
rect 6032 106596 6036 106652
rect 6036 106596 6092 106652
rect 6092 106596 6096 106652
rect 6032 106592 6096 106596
rect 6112 106652 6176 106656
rect 6112 106596 6116 106652
rect 6116 106596 6172 106652
rect 6172 106596 6176 106652
rect 6112 106592 6176 106596
rect 6192 106652 6256 106656
rect 6192 106596 6196 106652
rect 6196 106596 6252 106652
rect 6252 106596 6256 106652
rect 6192 106592 6256 106596
rect 4285 106108 4349 106112
rect 4285 106052 4289 106108
rect 4289 106052 4345 106108
rect 4345 106052 4349 106108
rect 4285 106048 4349 106052
rect 4365 106108 4429 106112
rect 4365 106052 4369 106108
rect 4369 106052 4425 106108
rect 4425 106052 4429 106108
rect 4365 106048 4429 106052
rect 4445 106108 4509 106112
rect 4445 106052 4449 106108
rect 4449 106052 4505 106108
rect 4505 106052 4509 106108
rect 4445 106048 4509 106052
rect 4525 106108 4589 106112
rect 4525 106052 4529 106108
rect 4529 106052 4585 106108
rect 4585 106052 4589 106108
rect 4525 106048 4589 106052
rect 7618 106108 7682 106112
rect 7618 106052 7622 106108
rect 7622 106052 7678 106108
rect 7678 106052 7682 106108
rect 7618 106048 7682 106052
rect 7698 106108 7762 106112
rect 7698 106052 7702 106108
rect 7702 106052 7758 106108
rect 7758 106052 7762 106108
rect 7698 106048 7762 106052
rect 7778 106108 7842 106112
rect 7778 106052 7782 106108
rect 7782 106052 7838 106108
rect 7838 106052 7842 106108
rect 7778 106048 7842 106052
rect 7858 106108 7922 106112
rect 7858 106052 7862 106108
rect 7862 106052 7918 106108
rect 7918 106052 7922 106108
rect 7858 106048 7922 106052
rect 2618 105564 2682 105568
rect 2618 105508 2622 105564
rect 2622 105508 2678 105564
rect 2678 105508 2682 105564
rect 2618 105504 2682 105508
rect 2698 105564 2762 105568
rect 2698 105508 2702 105564
rect 2702 105508 2758 105564
rect 2758 105508 2762 105564
rect 2698 105504 2762 105508
rect 2778 105564 2842 105568
rect 2778 105508 2782 105564
rect 2782 105508 2838 105564
rect 2838 105508 2842 105564
rect 2778 105504 2842 105508
rect 2858 105564 2922 105568
rect 2858 105508 2862 105564
rect 2862 105508 2918 105564
rect 2918 105508 2922 105564
rect 2858 105504 2922 105508
rect 5952 105564 6016 105568
rect 5952 105508 5956 105564
rect 5956 105508 6012 105564
rect 6012 105508 6016 105564
rect 5952 105504 6016 105508
rect 6032 105564 6096 105568
rect 6032 105508 6036 105564
rect 6036 105508 6092 105564
rect 6092 105508 6096 105564
rect 6032 105504 6096 105508
rect 6112 105564 6176 105568
rect 6112 105508 6116 105564
rect 6116 105508 6172 105564
rect 6172 105508 6176 105564
rect 6112 105504 6176 105508
rect 6192 105564 6256 105568
rect 6192 105508 6196 105564
rect 6196 105508 6252 105564
rect 6252 105508 6256 105564
rect 6192 105504 6256 105508
rect 4285 105020 4349 105024
rect 4285 104964 4289 105020
rect 4289 104964 4345 105020
rect 4345 104964 4349 105020
rect 4285 104960 4349 104964
rect 4365 105020 4429 105024
rect 4365 104964 4369 105020
rect 4369 104964 4425 105020
rect 4425 104964 4429 105020
rect 4365 104960 4429 104964
rect 4445 105020 4509 105024
rect 4445 104964 4449 105020
rect 4449 104964 4505 105020
rect 4505 104964 4509 105020
rect 4445 104960 4509 104964
rect 4525 105020 4589 105024
rect 4525 104964 4529 105020
rect 4529 104964 4585 105020
rect 4585 104964 4589 105020
rect 4525 104960 4589 104964
rect 7618 105020 7682 105024
rect 7618 104964 7622 105020
rect 7622 104964 7678 105020
rect 7678 104964 7682 105020
rect 7618 104960 7682 104964
rect 7698 105020 7762 105024
rect 7698 104964 7702 105020
rect 7702 104964 7758 105020
rect 7758 104964 7762 105020
rect 7698 104960 7762 104964
rect 7778 105020 7842 105024
rect 7778 104964 7782 105020
rect 7782 104964 7838 105020
rect 7838 104964 7842 105020
rect 7778 104960 7842 104964
rect 7858 105020 7922 105024
rect 7858 104964 7862 105020
rect 7862 104964 7918 105020
rect 7918 104964 7922 105020
rect 7858 104960 7922 104964
rect 2618 104476 2682 104480
rect 2618 104420 2622 104476
rect 2622 104420 2678 104476
rect 2678 104420 2682 104476
rect 2618 104416 2682 104420
rect 2698 104476 2762 104480
rect 2698 104420 2702 104476
rect 2702 104420 2758 104476
rect 2758 104420 2762 104476
rect 2698 104416 2762 104420
rect 2778 104476 2842 104480
rect 2778 104420 2782 104476
rect 2782 104420 2838 104476
rect 2838 104420 2842 104476
rect 2778 104416 2842 104420
rect 2858 104476 2922 104480
rect 2858 104420 2862 104476
rect 2862 104420 2918 104476
rect 2918 104420 2922 104476
rect 2858 104416 2922 104420
rect 5952 104476 6016 104480
rect 5952 104420 5956 104476
rect 5956 104420 6012 104476
rect 6012 104420 6016 104476
rect 5952 104416 6016 104420
rect 6032 104476 6096 104480
rect 6032 104420 6036 104476
rect 6036 104420 6092 104476
rect 6092 104420 6096 104476
rect 6032 104416 6096 104420
rect 6112 104476 6176 104480
rect 6112 104420 6116 104476
rect 6116 104420 6172 104476
rect 6172 104420 6176 104476
rect 6112 104416 6176 104420
rect 6192 104476 6256 104480
rect 6192 104420 6196 104476
rect 6196 104420 6252 104476
rect 6252 104420 6256 104476
rect 6192 104416 6256 104420
rect 4285 103932 4349 103936
rect 4285 103876 4289 103932
rect 4289 103876 4345 103932
rect 4345 103876 4349 103932
rect 4285 103872 4349 103876
rect 4365 103932 4429 103936
rect 4365 103876 4369 103932
rect 4369 103876 4425 103932
rect 4425 103876 4429 103932
rect 4365 103872 4429 103876
rect 4445 103932 4509 103936
rect 4445 103876 4449 103932
rect 4449 103876 4505 103932
rect 4505 103876 4509 103932
rect 4445 103872 4509 103876
rect 4525 103932 4589 103936
rect 4525 103876 4529 103932
rect 4529 103876 4585 103932
rect 4585 103876 4589 103932
rect 4525 103872 4589 103876
rect 7618 103932 7682 103936
rect 7618 103876 7622 103932
rect 7622 103876 7678 103932
rect 7678 103876 7682 103932
rect 7618 103872 7682 103876
rect 7698 103932 7762 103936
rect 7698 103876 7702 103932
rect 7702 103876 7758 103932
rect 7758 103876 7762 103932
rect 7698 103872 7762 103876
rect 7778 103932 7842 103936
rect 7778 103876 7782 103932
rect 7782 103876 7838 103932
rect 7838 103876 7842 103932
rect 7778 103872 7842 103876
rect 7858 103932 7922 103936
rect 7858 103876 7862 103932
rect 7862 103876 7918 103932
rect 7918 103876 7922 103932
rect 7858 103872 7922 103876
rect 2618 103388 2682 103392
rect 2618 103332 2622 103388
rect 2622 103332 2678 103388
rect 2678 103332 2682 103388
rect 2618 103328 2682 103332
rect 2698 103388 2762 103392
rect 2698 103332 2702 103388
rect 2702 103332 2758 103388
rect 2758 103332 2762 103388
rect 2698 103328 2762 103332
rect 2778 103388 2842 103392
rect 2778 103332 2782 103388
rect 2782 103332 2838 103388
rect 2838 103332 2842 103388
rect 2778 103328 2842 103332
rect 2858 103388 2922 103392
rect 2858 103332 2862 103388
rect 2862 103332 2918 103388
rect 2918 103332 2922 103388
rect 2858 103328 2922 103332
rect 5952 103388 6016 103392
rect 5952 103332 5956 103388
rect 5956 103332 6012 103388
rect 6012 103332 6016 103388
rect 5952 103328 6016 103332
rect 6032 103388 6096 103392
rect 6032 103332 6036 103388
rect 6036 103332 6092 103388
rect 6092 103332 6096 103388
rect 6032 103328 6096 103332
rect 6112 103388 6176 103392
rect 6112 103332 6116 103388
rect 6116 103332 6172 103388
rect 6172 103332 6176 103388
rect 6112 103328 6176 103332
rect 6192 103388 6256 103392
rect 6192 103332 6196 103388
rect 6196 103332 6252 103388
rect 6252 103332 6256 103388
rect 6192 103328 6256 103332
rect 4285 102844 4349 102848
rect 4285 102788 4289 102844
rect 4289 102788 4345 102844
rect 4345 102788 4349 102844
rect 4285 102784 4349 102788
rect 4365 102844 4429 102848
rect 4365 102788 4369 102844
rect 4369 102788 4425 102844
rect 4425 102788 4429 102844
rect 4365 102784 4429 102788
rect 4445 102844 4509 102848
rect 4445 102788 4449 102844
rect 4449 102788 4505 102844
rect 4505 102788 4509 102844
rect 4445 102784 4509 102788
rect 4525 102844 4589 102848
rect 4525 102788 4529 102844
rect 4529 102788 4585 102844
rect 4585 102788 4589 102844
rect 4525 102784 4589 102788
rect 7618 102844 7682 102848
rect 7618 102788 7622 102844
rect 7622 102788 7678 102844
rect 7678 102788 7682 102844
rect 7618 102784 7682 102788
rect 7698 102844 7762 102848
rect 7698 102788 7702 102844
rect 7702 102788 7758 102844
rect 7758 102788 7762 102844
rect 7698 102784 7762 102788
rect 7778 102844 7842 102848
rect 7778 102788 7782 102844
rect 7782 102788 7838 102844
rect 7838 102788 7842 102844
rect 7778 102784 7842 102788
rect 7858 102844 7922 102848
rect 7858 102788 7862 102844
rect 7862 102788 7918 102844
rect 7918 102788 7922 102844
rect 7858 102784 7922 102788
rect 2618 102300 2682 102304
rect 2618 102244 2622 102300
rect 2622 102244 2678 102300
rect 2678 102244 2682 102300
rect 2618 102240 2682 102244
rect 2698 102300 2762 102304
rect 2698 102244 2702 102300
rect 2702 102244 2758 102300
rect 2758 102244 2762 102300
rect 2698 102240 2762 102244
rect 2778 102300 2842 102304
rect 2778 102244 2782 102300
rect 2782 102244 2838 102300
rect 2838 102244 2842 102300
rect 2778 102240 2842 102244
rect 2858 102300 2922 102304
rect 2858 102244 2862 102300
rect 2862 102244 2918 102300
rect 2918 102244 2922 102300
rect 2858 102240 2922 102244
rect 5952 102300 6016 102304
rect 5952 102244 5956 102300
rect 5956 102244 6012 102300
rect 6012 102244 6016 102300
rect 5952 102240 6016 102244
rect 6032 102300 6096 102304
rect 6032 102244 6036 102300
rect 6036 102244 6092 102300
rect 6092 102244 6096 102300
rect 6032 102240 6096 102244
rect 6112 102300 6176 102304
rect 6112 102244 6116 102300
rect 6116 102244 6172 102300
rect 6172 102244 6176 102300
rect 6112 102240 6176 102244
rect 6192 102300 6256 102304
rect 6192 102244 6196 102300
rect 6196 102244 6252 102300
rect 6252 102244 6256 102300
rect 6192 102240 6256 102244
rect 4285 101756 4349 101760
rect 4285 101700 4289 101756
rect 4289 101700 4345 101756
rect 4345 101700 4349 101756
rect 4285 101696 4349 101700
rect 4365 101756 4429 101760
rect 4365 101700 4369 101756
rect 4369 101700 4425 101756
rect 4425 101700 4429 101756
rect 4365 101696 4429 101700
rect 4445 101756 4509 101760
rect 4445 101700 4449 101756
rect 4449 101700 4505 101756
rect 4505 101700 4509 101756
rect 4445 101696 4509 101700
rect 4525 101756 4589 101760
rect 4525 101700 4529 101756
rect 4529 101700 4585 101756
rect 4585 101700 4589 101756
rect 4525 101696 4589 101700
rect 7618 101756 7682 101760
rect 7618 101700 7622 101756
rect 7622 101700 7678 101756
rect 7678 101700 7682 101756
rect 7618 101696 7682 101700
rect 7698 101756 7762 101760
rect 7698 101700 7702 101756
rect 7702 101700 7758 101756
rect 7758 101700 7762 101756
rect 7698 101696 7762 101700
rect 7778 101756 7842 101760
rect 7778 101700 7782 101756
rect 7782 101700 7838 101756
rect 7838 101700 7842 101756
rect 7778 101696 7842 101700
rect 7858 101756 7922 101760
rect 7858 101700 7862 101756
rect 7862 101700 7918 101756
rect 7918 101700 7922 101756
rect 7858 101696 7922 101700
rect 2618 101212 2682 101216
rect 2618 101156 2622 101212
rect 2622 101156 2678 101212
rect 2678 101156 2682 101212
rect 2618 101152 2682 101156
rect 2698 101212 2762 101216
rect 2698 101156 2702 101212
rect 2702 101156 2758 101212
rect 2758 101156 2762 101212
rect 2698 101152 2762 101156
rect 2778 101212 2842 101216
rect 2778 101156 2782 101212
rect 2782 101156 2838 101212
rect 2838 101156 2842 101212
rect 2778 101152 2842 101156
rect 2858 101212 2922 101216
rect 2858 101156 2862 101212
rect 2862 101156 2918 101212
rect 2918 101156 2922 101212
rect 2858 101152 2922 101156
rect 5952 101212 6016 101216
rect 5952 101156 5956 101212
rect 5956 101156 6012 101212
rect 6012 101156 6016 101212
rect 5952 101152 6016 101156
rect 6032 101212 6096 101216
rect 6032 101156 6036 101212
rect 6036 101156 6092 101212
rect 6092 101156 6096 101212
rect 6032 101152 6096 101156
rect 6112 101212 6176 101216
rect 6112 101156 6116 101212
rect 6116 101156 6172 101212
rect 6172 101156 6176 101212
rect 6112 101152 6176 101156
rect 6192 101212 6256 101216
rect 6192 101156 6196 101212
rect 6196 101156 6252 101212
rect 6252 101156 6256 101212
rect 6192 101152 6256 101156
rect 4285 100668 4349 100672
rect 4285 100612 4289 100668
rect 4289 100612 4345 100668
rect 4345 100612 4349 100668
rect 4285 100608 4349 100612
rect 4365 100668 4429 100672
rect 4365 100612 4369 100668
rect 4369 100612 4425 100668
rect 4425 100612 4429 100668
rect 4365 100608 4429 100612
rect 4445 100668 4509 100672
rect 4445 100612 4449 100668
rect 4449 100612 4505 100668
rect 4505 100612 4509 100668
rect 4445 100608 4509 100612
rect 4525 100668 4589 100672
rect 4525 100612 4529 100668
rect 4529 100612 4585 100668
rect 4585 100612 4589 100668
rect 4525 100608 4589 100612
rect 7618 100668 7682 100672
rect 7618 100612 7622 100668
rect 7622 100612 7678 100668
rect 7678 100612 7682 100668
rect 7618 100608 7682 100612
rect 7698 100668 7762 100672
rect 7698 100612 7702 100668
rect 7702 100612 7758 100668
rect 7758 100612 7762 100668
rect 7698 100608 7762 100612
rect 7778 100668 7842 100672
rect 7778 100612 7782 100668
rect 7782 100612 7838 100668
rect 7838 100612 7842 100668
rect 7778 100608 7842 100612
rect 7858 100668 7922 100672
rect 7858 100612 7862 100668
rect 7862 100612 7918 100668
rect 7918 100612 7922 100668
rect 7858 100608 7922 100612
rect 2618 100124 2682 100128
rect 2618 100068 2622 100124
rect 2622 100068 2678 100124
rect 2678 100068 2682 100124
rect 2618 100064 2682 100068
rect 2698 100124 2762 100128
rect 2698 100068 2702 100124
rect 2702 100068 2758 100124
rect 2758 100068 2762 100124
rect 2698 100064 2762 100068
rect 2778 100124 2842 100128
rect 2778 100068 2782 100124
rect 2782 100068 2838 100124
rect 2838 100068 2842 100124
rect 2778 100064 2842 100068
rect 2858 100124 2922 100128
rect 2858 100068 2862 100124
rect 2862 100068 2918 100124
rect 2918 100068 2922 100124
rect 2858 100064 2922 100068
rect 5952 100124 6016 100128
rect 5952 100068 5956 100124
rect 5956 100068 6012 100124
rect 6012 100068 6016 100124
rect 5952 100064 6016 100068
rect 6032 100124 6096 100128
rect 6032 100068 6036 100124
rect 6036 100068 6092 100124
rect 6092 100068 6096 100124
rect 6032 100064 6096 100068
rect 6112 100124 6176 100128
rect 6112 100068 6116 100124
rect 6116 100068 6172 100124
rect 6172 100068 6176 100124
rect 6112 100064 6176 100068
rect 6192 100124 6256 100128
rect 6192 100068 6196 100124
rect 6196 100068 6252 100124
rect 6252 100068 6256 100124
rect 6192 100064 6256 100068
rect 4285 99580 4349 99584
rect 4285 99524 4289 99580
rect 4289 99524 4345 99580
rect 4345 99524 4349 99580
rect 4285 99520 4349 99524
rect 4365 99580 4429 99584
rect 4365 99524 4369 99580
rect 4369 99524 4425 99580
rect 4425 99524 4429 99580
rect 4365 99520 4429 99524
rect 4445 99580 4509 99584
rect 4445 99524 4449 99580
rect 4449 99524 4505 99580
rect 4505 99524 4509 99580
rect 4445 99520 4509 99524
rect 4525 99580 4589 99584
rect 4525 99524 4529 99580
rect 4529 99524 4585 99580
rect 4585 99524 4589 99580
rect 4525 99520 4589 99524
rect 7618 99580 7682 99584
rect 7618 99524 7622 99580
rect 7622 99524 7678 99580
rect 7678 99524 7682 99580
rect 7618 99520 7682 99524
rect 7698 99580 7762 99584
rect 7698 99524 7702 99580
rect 7702 99524 7758 99580
rect 7758 99524 7762 99580
rect 7698 99520 7762 99524
rect 7778 99580 7842 99584
rect 7778 99524 7782 99580
rect 7782 99524 7838 99580
rect 7838 99524 7842 99580
rect 7778 99520 7842 99524
rect 7858 99580 7922 99584
rect 7858 99524 7862 99580
rect 7862 99524 7918 99580
rect 7918 99524 7922 99580
rect 7858 99520 7922 99524
rect 2618 99036 2682 99040
rect 2618 98980 2622 99036
rect 2622 98980 2678 99036
rect 2678 98980 2682 99036
rect 2618 98976 2682 98980
rect 2698 99036 2762 99040
rect 2698 98980 2702 99036
rect 2702 98980 2758 99036
rect 2758 98980 2762 99036
rect 2698 98976 2762 98980
rect 2778 99036 2842 99040
rect 2778 98980 2782 99036
rect 2782 98980 2838 99036
rect 2838 98980 2842 99036
rect 2778 98976 2842 98980
rect 2858 99036 2922 99040
rect 2858 98980 2862 99036
rect 2862 98980 2918 99036
rect 2918 98980 2922 99036
rect 2858 98976 2922 98980
rect 5952 99036 6016 99040
rect 5952 98980 5956 99036
rect 5956 98980 6012 99036
rect 6012 98980 6016 99036
rect 5952 98976 6016 98980
rect 6032 99036 6096 99040
rect 6032 98980 6036 99036
rect 6036 98980 6092 99036
rect 6092 98980 6096 99036
rect 6032 98976 6096 98980
rect 6112 99036 6176 99040
rect 6112 98980 6116 99036
rect 6116 98980 6172 99036
rect 6172 98980 6176 99036
rect 6112 98976 6176 98980
rect 6192 99036 6256 99040
rect 6192 98980 6196 99036
rect 6196 98980 6252 99036
rect 6252 98980 6256 99036
rect 6192 98976 6256 98980
rect 4285 98492 4349 98496
rect 4285 98436 4289 98492
rect 4289 98436 4345 98492
rect 4345 98436 4349 98492
rect 4285 98432 4349 98436
rect 4365 98492 4429 98496
rect 4365 98436 4369 98492
rect 4369 98436 4425 98492
rect 4425 98436 4429 98492
rect 4365 98432 4429 98436
rect 4445 98492 4509 98496
rect 4445 98436 4449 98492
rect 4449 98436 4505 98492
rect 4505 98436 4509 98492
rect 4445 98432 4509 98436
rect 4525 98492 4589 98496
rect 4525 98436 4529 98492
rect 4529 98436 4585 98492
rect 4585 98436 4589 98492
rect 4525 98432 4589 98436
rect 7618 98492 7682 98496
rect 7618 98436 7622 98492
rect 7622 98436 7678 98492
rect 7678 98436 7682 98492
rect 7618 98432 7682 98436
rect 7698 98492 7762 98496
rect 7698 98436 7702 98492
rect 7702 98436 7758 98492
rect 7758 98436 7762 98492
rect 7698 98432 7762 98436
rect 7778 98492 7842 98496
rect 7778 98436 7782 98492
rect 7782 98436 7838 98492
rect 7838 98436 7842 98492
rect 7778 98432 7842 98436
rect 7858 98492 7922 98496
rect 7858 98436 7862 98492
rect 7862 98436 7918 98492
rect 7918 98436 7922 98492
rect 7858 98432 7922 98436
rect 2618 97948 2682 97952
rect 2618 97892 2622 97948
rect 2622 97892 2678 97948
rect 2678 97892 2682 97948
rect 2618 97888 2682 97892
rect 2698 97948 2762 97952
rect 2698 97892 2702 97948
rect 2702 97892 2758 97948
rect 2758 97892 2762 97948
rect 2698 97888 2762 97892
rect 2778 97948 2842 97952
rect 2778 97892 2782 97948
rect 2782 97892 2838 97948
rect 2838 97892 2842 97948
rect 2778 97888 2842 97892
rect 2858 97948 2922 97952
rect 2858 97892 2862 97948
rect 2862 97892 2918 97948
rect 2918 97892 2922 97948
rect 2858 97888 2922 97892
rect 5952 97948 6016 97952
rect 5952 97892 5956 97948
rect 5956 97892 6012 97948
rect 6012 97892 6016 97948
rect 5952 97888 6016 97892
rect 6032 97948 6096 97952
rect 6032 97892 6036 97948
rect 6036 97892 6092 97948
rect 6092 97892 6096 97948
rect 6032 97888 6096 97892
rect 6112 97948 6176 97952
rect 6112 97892 6116 97948
rect 6116 97892 6172 97948
rect 6172 97892 6176 97948
rect 6112 97888 6176 97892
rect 6192 97948 6256 97952
rect 6192 97892 6196 97948
rect 6196 97892 6252 97948
rect 6252 97892 6256 97948
rect 6192 97888 6256 97892
rect 4285 97404 4349 97408
rect 4285 97348 4289 97404
rect 4289 97348 4345 97404
rect 4345 97348 4349 97404
rect 4285 97344 4349 97348
rect 4365 97404 4429 97408
rect 4365 97348 4369 97404
rect 4369 97348 4425 97404
rect 4425 97348 4429 97404
rect 4365 97344 4429 97348
rect 4445 97404 4509 97408
rect 4445 97348 4449 97404
rect 4449 97348 4505 97404
rect 4505 97348 4509 97404
rect 4445 97344 4509 97348
rect 4525 97404 4589 97408
rect 4525 97348 4529 97404
rect 4529 97348 4585 97404
rect 4585 97348 4589 97404
rect 4525 97344 4589 97348
rect 7618 97404 7682 97408
rect 7618 97348 7622 97404
rect 7622 97348 7678 97404
rect 7678 97348 7682 97404
rect 7618 97344 7682 97348
rect 7698 97404 7762 97408
rect 7698 97348 7702 97404
rect 7702 97348 7758 97404
rect 7758 97348 7762 97404
rect 7698 97344 7762 97348
rect 7778 97404 7842 97408
rect 7778 97348 7782 97404
rect 7782 97348 7838 97404
rect 7838 97348 7842 97404
rect 7778 97344 7842 97348
rect 7858 97404 7922 97408
rect 7858 97348 7862 97404
rect 7862 97348 7918 97404
rect 7918 97348 7922 97404
rect 7858 97344 7922 97348
rect 2618 96860 2682 96864
rect 2618 96804 2622 96860
rect 2622 96804 2678 96860
rect 2678 96804 2682 96860
rect 2618 96800 2682 96804
rect 2698 96860 2762 96864
rect 2698 96804 2702 96860
rect 2702 96804 2758 96860
rect 2758 96804 2762 96860
rect 2698 96800 2762 96804
rect 2778 96860 2842 96864
rect 2778 96804 2782 96860
rect 2782 96804 2838 96860
rect 2838 96804 2842 96860
rect 2778 96800 2842 96804
rect 2858 96860 2922 96864
rect 2858 96804 2862 96860
rect 2862 96804 2918 96860
rect 2918 96804 2922 96860
rect 2858 96800 2922 96804
rect 5952 96860 6016 96864
rect 5952 96804 5956 96860
rect 5956 96804 6012 96860
rect 6012 96804 6016 96860
rect 5952 96800 6016 96804
rect 6032 96860 6096 96864
rect 6032 96804 6036 96860
rect 6036 96804 6092 96860
rect 6092 96804 6096 96860
rect 6032 96800 6096 96804
rect 6112 96860 6176 96864
rect 6112 96804 6116 96860
rect 6116 96804 6172 96860
rect 6172 96804 6176 96860
rect 6112 96800 6176 96804
rect 6192 96860 6256 96864
rect 6192 96804 6196 96860
rect 6196 96804 6252 96860
rect 6252 96804 6256 96860
rect 6192 96800 6256 96804
rect 4285 96316 4349 96320
rect 4285 96260 4289 96316
rect 4289 96260 4345 96316
rect 4345 96260 4349 96316
rect 4285 96256 4349 96260
rect 4365 96316 4429 96320
rect 4365 96260 4369 96316
rect 4369 96260 4425 96316
rect 4425 96260 4429 96316
rect 4365 96256 4429 96260
rect 4445 96316 4509 96320
rect 4445 96260 4449 96316
rect 4449 96260 4505 96316
rect 4505 96260 4509 96316
rect 4445 96256 4509 96260
rect 4525 96316 4589 96320
rect 4525 96260 4529 96316
rect 4529 96260 4585 96316
rect 4585 96260 4589 96316
rect 4525 96256 4589 96260
rect 7618 96316 7682 96320
rect 7618 96260 7622 96316
rect 7622 96260 7678 96316
rect 7678 96260 7682 96316
rect 7618 96256 7682 96260
rect 7698 96316 7762 96320
rect 7698 96260 7702 96316
rect 7702 96260 7758 96316
rect 7758 96260 7762 96316
rect 7698 96256 7762 96260
rect 7778 96316 7842 96320
rect 7778 96260 7782 96316
rect 7782 96260 7838 96316
rect 7838 96260 7842 96316
rect 7778 96256 7842 96260
rect 7858 96316 7922 96320
rect 7858 96260 7862 96316
rect 7862 96260 7918 96316
rect 7918 96260 7922 96316
rect 7858 96256 7922 96260
rect 2618 95772 2682 95776
rect 2618 95716 2622 95772
rect 2622 95716 2678 95772
rect 2678 95716 2682 95772
rect 2618 95712 2682 95716
rect 2698 95772 2762 95776
rect 2698 95716 2702 95772
rect 2702 95716 2758 95772
rect 2758 95716 2762 95772
rect 2698 95712 2762 95716
rect 2778 95772 2842 95776
rect 2778 95716 2782 95772
rect 2782 95716 2838 95772
rect 2838 95716 2842 95772
rect 2778 95712 2842 95716
rect 2858 95772 2922 95776
rect 2858 95716 2862 95772
rect 2862 95716 2918 95772
rect 2918 95716 2922 95772
rect 2858 95712 2922 95716
rect 5952 95772 6016 95776
rect 5952 95716 5956 95772
rect 5956 95716 6012 95772
rect 6012 95716 6016 95772
rect 5952 95712 6016 95716
rect 6032 95772 6096 95776
rect 6032 95716 6036 95772
rect 6036 95716 6092 95772
rect 6092 95716 6096 95772
rect 6032 95712 6096 95716
rect 6112 95772 6176 95776
rect 6112 95716 6116 95772
rect 6116 95716 6172 95772
rect 6172 95716 6176 95772
rect 6112 95712 6176 95716
rect 6192 95772 6256 95776
rect 6192 95716 6196 95772
rect 6196 95716 6252 95772
rect 6252 95716 6256 95772
rect 6192 95712 6256 95716
rect 4285 95228 4349 95232
rect 4285 95172 4289 95228
rect 4289 95172 4345 95228
rect 4345 95172 4349 95228
rect 4285 95168 4349 95172
rect 4365 95228 4429 95232
rect 4365 95172 4369 95228
rect 4369 95172 4425 95228
rect 4425 95172 4429 95228
rect 4365 95168 4429 95172
rect 4445 95228 4509 95232
rect 4445 95172 4449 95228
rect 4449 95172 4505 95228
rect 4505 95172 4509 95228
rect 4445 95168 4509 95172
rect 4525 95228 4589 95232
rect 4525 95172 4529 95228
rect 4529 95172 4585 95228
rect 4585 95172 4589 95228
rect 4525 95168 4589 95172
rect 7618 95228 7682 95232
rect 7618 95172 7622 95228
rect 7622 95172 7678 95228
rect 7678 95172 7682 95228
rect 7618 95168 7682 95172
rect 7698 95228 7762 95232
rect 7698 95172 7702 95228
rect 7702 95172 7758 95228
rect 7758 95172 7762 95228
rect 7698 95168 7762 95172
rect 7778 95228 7842 95232
rect 7778 95172 7782 95228
rect 7782 95172 7838 95228
rect 7838 95172 7842 95228
rect 7778 95168 7842 95172
rect 7858 95228 7922 95232
rect 7858 95172 7862 95228
rect 7862 95172 7918 95228
rect 7918 95172 7922 95228
rect 7858 95168 7922 95172
rect 2618 94684 2682 94688
rect 2618 94628 2622 94684
rect 2622 94628 2678 94684
rect 2678 94628 2682 94684
rect 2618 94624 2682 94628
rect 2698 94684 2762 94688
rect 2698 94628 2702 94684
rect 2702 94628 2758 94684
rect 2758 94628 2762 94684
rect 2698 94624 2762 94628
rect 2778 94684 2842 94688
rect 2778 94628 2782 94684
rect 2782 94628 2838 94684
rect 2838 94628 2842 94684
rect 2778 94624 2842 94628
rect 2858 94684 2922 94688
rect 2858 94628 2862 94684
rect 2862 94628 2918 94684
rect 2918 94628 2922 94684
rect 2858 94624 2922 94628
rect 5952 94684 6016 94688
rect 5952 94628 5956 94684
rect 5956 94628 6012 94684
rect 6012 94628 6016 94684
rect 5952 94624 6016 94628
rect 6032 94684 6096 94688
rect 6032 94628 6036 94684
rect 6036 94628 6092 94684
rect 6092 94628 6096 94684
rect 6032 94624 6096 94628
rect 6112 94684 6176 94688
rect 6112 94628 6116 94684
rect 6116 94628 6172 94684
rect 6172 94628 6176 94684
rect 6112 94624 6176 94628
rect 6192 94684 6256 94688
rect 6192 94628 6196 94684
rect 6196 94628 6252 94684
rect 6252 94628 6256 94684
rect 6192 94624 6256 94628
rect 4285 94140 4349 94144
rect 4285 94084 4289 94140
rect 4289 94084 4345 94140
rect 4345 94084 4349 94140
rect 4285 94080 4349 94084
rect 4365 94140 4429 94144
rect 4365 94084 4369 94140
rect 4369 94084 4425 94140
rect 4425 94084 4429 94140
rect 4365 94080 4429 94084
rect 4445 94140 4509 94144
rect 4445 94084 4449 94140
rect 4449 94084 4505 94140
rect 4505 94084 4509 94140
rect 4445 94080 4509 94084
rect 4525 94140 4589 94144
rect 4525 94084 4529 94140
rect 4529 94084 4585 94140
rect 4585 94084 4589 94140
rect 4525 94080 4589 94084
rect 7618 94140 7682 94144
rect 7618 94084 7622 94140
rect 7622 94084 7678 94140
rect 7678 94084 7682 94140
rect 7618 94080 7682 94084
rect 7698 94140 7762 94144
rect 7698 94084 7702 94140
rect 7702 94084 7758 94140
rect 7758 94084 7762 94140
rect 7698 94080 7762 94084
rect 7778 94140 7842 94144
rect 7778 94084 7782 94140
rect 7782 94084 7838 94140
rect 7838 94084 7842 94140
rect 7778 94080 7842 94084
rect 7858 94140 7922 94144
rect 7858 94084 7862 94140
rect 7862 94084 7918 94140
rect 7918 94084 7922 94140
rect 7858 94080 7922 94084
rect 2618 93596 2682 93600
rect 2618 93540 2622 93596
rect 2622 93540 2678 93596
rect 2678 93540 2682 93596
rect 2618 93536 2682 93540
rect 2698 93596 2762 93600
rect 2698 93540 2702 93596
rect 2702 93540 2758 93596
rect 2758 93540 2762 93596
rect 2698 93536 2762 93540
rect 2778 93596 2842 93600
rect 2778 93540 2782 93596
rect 2782 93540 2838 93596
rect 2838 93540 2842 93596
rect 2778 93536 2842 93540
rect 2858 93596 2922 93600
rect 2858 93540 2862 93596
rect 2862 93540 2918 93596
rect 2918 93540 2922 93596
rect 2858 93536 2922 93540
rect 5952 93596 6016 93600
rect 5952 93540 5956 93596
rect 5956 93540 6012 93596
rect 6012 93540 6016 93596
rect 5952 93536 6016 93540
rect 6032 93596 6096 93600
rect 6032 93540 6036 93596
rect 6036 93540 6092 93596
rect 6092 93540 6096 93596
rect 6032 93536 6096 93540
rect 6112 93596 6176 93600
rect 6112 93540 6116 93596
rect 6116 93540 6172 93596
rect 6172 93540 6176 93596
rect 6112 93536 6176 93540
rect 6192 93596 6256 93600
rect 6192 93540 6196 93596
rect 6196 93540 6252 93596
rect 6252 93540 6256 93596
rect 6192 93536 6256 93540
rect 4285 93052 4349 93056
rect 4285 92996 4289 93052
rect 4289 92996 4345 93052
rect 4345 92996 4349 93052
rect 4285 92992 4349 92996
rect 4365 93052 4429 93056
rect 4365 92996 4369 93052
rect 4369 92996 4425 93052
rect 4425 92996 4429 93052
rect 4365 92992 4429 92996
rect 4445 93052 4509 93056
rect 4445 92996 4449 93052
rect 4449 92996 4505 93052
rect 4505 92996 4509 93052
rect 4445 92992 4509 92996
rect 4525 93052 4589 93056
rect 4525 92996 4529 93052
rect 4529 92996 4585 93052
rect 4585 92996 4589 93052
rect 4525 92992 4589 92996
rect 7618 93052 7682 93056
rect 7618 92996 7622 93052
rect 7622 92996 7678 93052
rect 7678 92996 7682 93052
rect 7618 92992 7682 92996
rect 7698 93052 7762 93056
rect 7698 92996 7702 93052
rect 7702 92996 7758 93052
rect 7758 92996 7762 93052
rect 7698 92992 7762 92996
rect 7778 93052 7842 93056
rect 7778 92996 7782 93052
rect 7782 92996 7838 93052
rect 7838 92996 7842 93052
rect 7778 92992 7842 92996
rect 7858 93052 7922 93056
rect 7858 92996 7862 93052
rect 7862 92996 7918 93052
rect 7918 92996 7922 93052
rect 7858 92992 7922 92996
rect 2618 92508 2682 92512
rect 2618 92452 2622 92508
rect 2622 92452 2678 92508
rect 2678 92452 2682 92508
rect 2618 92448 2682 92452
rect 2698 92508 2762 92512
rect 2698 92452 2702 92508
rect 2702 92452 2758 92508
rect 2758 92452 2762 92508
rect 2698 92448 2762 92452
rect 2778 92508 2842 92512
rect 2778 92452 2782 92508
rect 2782 92452 2838 92508
rect 2838 92452 2842 92508
rect 2778 92448 2842 92452
rect 2858 92508 2922 92512
rect 2858 92452 2862 92508
rect 2862 92452 2918 92508
rect 2918 92452 2922 92508
rect 2858 92448 2922 92452
rect 5952 92508 6016 92512
rect 5952 92452 5956 92508
rect 5956 92452 6012 92508
rect 6012 92452 6016 92508
rect 5952 92448 6016 92452
rect 6032 92508 6096 92512
rect 6032 92452 6036 92508
rect 6036 92452 6092 92508
rect 6092 92452 6096 92508
rect 6032 92448 6096 92452
rect 6112 92508 6176 92512
rect 6112 92452 6116 92508
rect 6116 92452 6172 92508
rect 6172 92452 6176 92508
rect 6112 92448 6176 92452
rect 6192 92508 6256 92512
rect 6192 92452 6196 92508
rect 6196 92452 6252 92508
rect 6252 92452 6256 92508
rect 6192 92448 6256 92452
rect 4285 91964 4349 91968
rect 4285 91908 4289 91964
rect 4289 91908 4345 91964
rect 4345 91908 4349 91964
rect 4285 91904 4349 91908
rect 4365 91964 4429 91968
rect 4365 91908 4369 91964
rect 4369 91908 4425 91964
rect 4425 91908 4429 91964
rect 4365 91904 4429 91908
rect 4445 91964 4509 91968
rect 4445 91908 4449 91964
rect 4449 91908 4505 91964
rect 4505 91908 4509 91964
rect 4445 91904 4509 91908
rect 4525 91964 4589 91968
rect 4525 91908 4529 91964
rect 4529 91908 4585 91964
rect 4585 91908 4589 91964
rect 4525 91904 4589 91908
rect 7618 91964 7682 91968
rect 7618 91908 7622 91964
rect 7622 91908 7678 91964
rect 7678 91908 7682 91964
rect 7618 91904 7682 91908
rect 7698 91964 7762 91968
rect 7698 91908 7702 91964
rect 7702 91908 7758 91964
rect 7758 91908 7762 91964
rect 7698 91904 7762 91908
rect 7778 91964 7842 91968
rect 7778 91908 7782 91964
rect 7782 91908 7838 91964
rect 7838 91908 7842 91964
rect 7778 91904 7842 91908
rect 7858 91964 7922 91968
rect 7858 91908 7862 91964
rect 7862 91908 7918 91964
rect 7918 91908 7922 91964
rect 7858 91904 7922 91908
rect 2618 91420 2682 91424
rect 2618 91364 2622 91420
rect 2622 91364 2678 91420
rect 2678 91364 2682 91420
rect 2618 91360 2682 91364
rect 2698 91420 2762 91424
rect 2698 91364 2702 91420
rect 2702 91364 2758 91420
rect 2758 91364 2762 91420
rect 2698 91360 2762 91364
rect 2778 91420 2842 91424
rect 2778 91364 2782 91420
rect 2782 91364 2838 91420
rect 2838 91364 2842 91420
rect 2778 91360 2842 91364
rect 2858 91420 2922 91424
rect 2858 91364 2862 91420
rect 2862 91364 2918 91420
rect 2918 91364 2922 91420
rect 2858 91360 2922 91364
rect 5952 91420 6016 91424
rect 5952 91364 5956 91420
rect 5956 91364 6012 91420
rect 6012 91364 6016 91420
rect 5952 91360 6016 91364
rect 6032 91420 6096 91424
rect 6032 91364 6036 91420
rect 6036 91364 6092 91420
rect 6092 91364 6096 91420
rect 6032 91360 6096 91364
rect 6112 91420 6176 91424
rect 6112 91364 6116 91420
rect 6116 91364 6172 91420
rect 6172 91364 6176 91420
rect 6112 91360 6176 91364
rect 6192 91420 6256 91424
rect 6192 91364 6196 91420
rect 6196 91364 6252 91420
rect 6252 91364 6256 91420
rect 6192 91360 6256 91364
rect 4285 90876 4349 90880
rect 4285 90820 4289 90876
rect 4289 90820 4345 90876
rect 4345 90820 4349 90876
rect 4285 90816 4349 90820
rect 4365 90876 4429 90880
rect 4365 90820 4369 90876
rect 4369 90820 4425 90876
rect 4425 90820 4429 90876
rect 4365 90816 4429 90820
rect 4445 90876 4509 90880
rect 4445 90820 4449 90876
rect 4449 90820 4505 90876
rect 4505 90820 4509 90876
rect 4445 90816 4509 90820
rect 4525 90876 4589 90880
rect 4525 90820 4529 90876
rect 4529 90820 4585 90876
rect 4585 90820 4589 90876
rect 4525 90816 4589 90820
rect 7618 90876 7682 90880
rect 7618 90820 7622 90876
rect 7622 90820 7678 90876
rect 7678 90820 7682 90876
rect 7618 90816 7682 90820
rect 7698 90876 7762 90880
rect 7698 90820 7702 90876
rect 7702 90820 7758 90876
rect 7758 90820 7762 90876
rect 7698 90816 7762 90820
rect 7778 90876 7842 90880
rect 7778 90820 7782 90876
rect 7782 90820 7838 90876
rect 7838 90820 7842 90876
rect 7778 90816 7842 90820
rect 7858 90876 7922 90880
rect 7858 90820 7862 90876
rect 7862 90820 7918 90876
rect 7918 90820 7922 90876
rect 7858 90816 7922 90820
rect 2618 90332 2682 90336
rect 2618 90276 2622 90332
rect 2622 90276 2678 90332
rect 2678 90276 2682 90332
rect 2618 90272 2682 90276
rect 2698 90332 2762 90336
rect 2698 90276 2702 90332
rect 2702 90276 2758 90332
rect 2758 90276 2762 90332
rect 2698 90272 2762 90276
rect 2778 90332 2842 90336
rect 2778 90276 2782 90332
rect 2782 90276 2838 90332
rect 2838 90276 2842 90332
rect 2778 90272 2842 90276
rect 2858 90332 2922 90336
rect 2858 90276 2862 90332
rect 2862 90276 2918 90332
rect 2918 90276 2922 90332
rect 2858 90272 2922 90276
rect 5952 90332 6016 90336
rect 5952 90276 5956 90332
rect 5956 90276 6012 90332
rect 6012 90276 6016 90332
rect 5952 90272 6016 90276
rect 6032 90332 6096 90336
rect 6032 90276 6036 90332
rect 6036 90276 6092 90332
rect 6092 90276 6096 90332
rect 6032 90272 6096 90276
rect 6112 90332 6176 90336
rect 6112 90276 6116 90332
rect 6116 90276 6172 90332
rect 6172 90276 6176 90332
rect 6112 90272 6176 90276
rect 6192 90332 6256 90336
rect 6192 90276 6196 90332
rect 6196 90276 6252 90332
rect 6252 90276 6256 90332
rect 6192 90272 6256 90276
rect 4285 89788 4349 89792
rect 4285 89732 4289 89788
rect 4289 89732 4345 89788
rect 4345 89732 4349 89788
rect 4285 89728 4349 89732
rect 4365 89788 4429 89792
rect 4365 89732 4369 89788
rect 4369 89732 4425 89788
rect 4425 89732 4429 89788
rect 4365 89728 4429 89732
rect 4445 89788 4509 89792
rect 4445 89732 4449 89788
rect 4449 89732 4505 89788
rect 4505 89732 4509 89788
rect 4445 89728 4509 89732
rect 4525 89788 4589 89792
rect 4525 89732 4529 89788
rect 4529 89732 4585 89788
rect 4585 89732 4589 89788
rect 4525 89728 4589 89732
rect 7618 89788 7682 89792
rect 7618 89732 7622 89788
rect 7622 89732 7678 89788
rect 7678 89732 7682 89788
rect 7618 89728 7682 89732
rect 7698 89788 7762 89792
rect 7698 89732 7702 89788
rect 7702 89732 7758 89788
rect 7758 89732 7762 89788
rect 7698 89728 7762 89732
rect 7778 89788 7842 89792
rect 7778 89732 7782 89788
rect 7782 89732 7838 89788
rect 7838 89732 7842 89788
rect 7778 89728 7842 89732
rect 7858 89788 7922 89792
rect 7858 89732 7862 89788
rect 7862 89732 7918 89788
rect 7918 89732 7922 89788
rect 7858 89728 7922 89732
rect 2618 89244 2682 89248
rect 2618 89188 2622 89244
rect 2622 89188 2678 89244
rect 2678 89188 2682 89244
rect 2618 89184 2682 89188
rect 2698 89244 2762 89248
rect 2698 89188 2702 89244
rect 2702 89188 2758 89244
rect 2758 89188 2762 89244
rect 2698 89184 2762 89188
rect 2778 89244 2842 89248
rect 2778 89188 2782 89244
rect 2782 89188 2838 89244
rect 2838 89188 2842 89244
rect 2778 89184 2842 89188
rect 2858 89244 2922 89248
rect 2858 89188 2862 89244
rect 2862 89188 2918 89244
rect 2918 89188 2922 89244
rect 2858 89184 2922 89188
rect 5952 89244 6016 89248
rect 5952 89188 5956 89244
rect 5956 89188 6012 89244
rect 6012 89188 6016 89244
rect 5952 89184 6016 89188
rect 6032 89244 6096 89248
rect 6032 89188 6036 89244
rect 6036 89188 6092 89244
rect 6092 89188 6096 89244
rect 6032 89184 6096 89188
rect 6112 89244 6176 89248
rect 6112 89188 6116 89244
rect 6116 89188 6172 89244
rect 6172 89188 6176 89244
rect 6112 89184 6176 89188
rect 6192 89244 6256 89248
rect 6192 89188 6196 89244
rect 6196 89188 6252 89244
rect 6252 89188 6256 89244
rect 6192 89184 6256 89188
rect 4285 88700 4349 88704
rect 4285 88644 4289 88700
rect 4289 88644 4345 88700
rect 4345 88644 4349 88700
rect 4285 88640 4349 88644
rect 4365 88700 4429 88704
rect 4365 88644 4369 88700
rect 4369 88644 4425 88700
rect 4425 88644 4429 88700
rect 4365 88640 4429 88644
rect 4445 88700 4509 88704
rect 4445 88644 4449 88700
rect 4449 88644 4505 88700
rect 4505 88644 4509 88700
rect 4445 88640 4509 88644
rect 4525 88700 4589 88704
rect 4525 88644 4529 88700
rect 4529 88644 4585 88700
rect 4585 88644 4589 88700
rect 4525 88640 4589 88644
rect 7618 88700 7682 88704
rect 7618 88644 7622 88700
rect 7622 88644 7678 88700
rect 7678 88644 7682 88700
rect 7618 88640 7682 88644
rect 7698 88700 7762 88704
rect 7698 88644 7702 88700
rect 7702 88644 7758 88700
rect 7758 88644 7762 88700
rect 7698 88640 7762 88644
rect 7778 88700 7842 88704
rect 7778 88644 7782 88700
rect 7782 88644 7838 88700
rect 7838 88644 7842 88700
rect 7778 88640 7842 88644
rect 7858 88700 7922 88704
rect 7858 88644 7862 88700
rect 7862 88644 7918 88700
rect 7918 88644 7922 88700
rect 7858 88640 7922 88644
rect 2618 88156 2682 88160
rect 2618 88100 2622 88156
rect 2622 88100 2678 88156
rect 2678 88100 2682 88156
rect 2618 88096 2682 88100
rect 2698 88156 2762 88160
rect 2698 88100 2702 88156
rect 2702 88100 2758 88156
rect 2758 88100 2762 88156
rect 2698 88096 2762 88100
rect 2778 88156 2842 88160
rect 2778 88100 2782 88156
rect 2782 88100 2838 88156
rect 2838 88100 2842 88156
rect 2778 88096 2842 88100
rect 2858 88156 2922 88160
rect 2858 88100 2862 88156
rect 2862 88100 2918 88156
rect 2918 88100 2922 88156
rect 2858 88096 2922 88100
rect 5952 88156 6016 88160
rect 5952 88100 5956 88156
rect 5956 88100 6012 88156
rect 6012 88100 6016 88156
rect 5952 88096 6016 88100
rect 6032 88156 6096 88160
rect 6032 88100 6036 88156
rect 6036 88100 6092 88156
rect 6092 88100 6096 88156
rect 6032 88096 6096 88100
rect 6112 88156 6176 88160
rect 6112 88100 6116 88156
rect 6116 88100 6172 88156
rect 6172 88100 6176 88156
rect 6112 88096 6176 88100
rect 6192 88156 6256 88160
rect 6192 88100 6196 88156
rect 6196 88100 6252 88156
rect 6252 88100 6256 88156
rect 6192 88096 6256 88100
rect 4285 87612 4349 87616
rect 4285 87556 4289 87612
rect 4289 87556 4345 87612
rect 4345 87556 4349 87612
rect 4285 87552 4349 87556
rect 4365 87612 4429 87616
rect 4365 87556 4369 87612
rect 4369 87556 4425 87612
rect 4425 87556 4429 87612
rect 4365 87552 4429 87556
rect 4445 87612 4509 87616
rect 4445 87556 4449 87612
rect 4449 87556 4505 87612
rect 4505 87556 4509 87612
rect 4445 87552 4509 87556
rect 4525 87612 4589 87616
rect 4525 87556 4529 87612
rect 4529 87556 4585 87612
rect 4585 87556 4589 87612
rect 4525 87552 4589 87556
rect 7618 87612 7682 87616
rect 7618 87556 7622 87612
rect 7622 87556 7678 87612
rect 7678 87556 7682 87612
rect 7618 87552 7682 87556
rect 7698 87612 7762 87616
rect 7698 87556 7702 87612
rect 7702 87556 7758 87612
rect 7758 87556 7762 87612
rect 7698 87552 7762 87556
rect 7778 87612 7842 87616
rect 7778 87556 7782 87612
rect 7782 87556 7838 87612
rect 7838 87556 7842 87612
rect 7778 87552 7842 87556
rect 7858 87612 7922 87616
rect 7858 87556 7862 87612
rect 7862 87556 7918 87612
rect 7918 87556 7922 87612
rect 7858 87552 7922 87556
rect 2618 87068 2682 87072
rect 2618 87012 2622 87068
rect 2622 87012 2678 87068
rect 2678 87012 2682 87068
rect 2618 87008 2682 87012
rect 2698 87068 2762 87072
rect 2698 87012 2702 87068
rect 2702 87012 2758 87068
rect 2758 87012 2762 87068
rect 2698 87008 2762 87012
rect 2778 87068 2842 87072
rect 2778 87012 2782 87068
rect 2782 87012 2838 87068
rect 2838 87012 2842 87068
rect 2778 87008 2842 87012
rect 2858 87068 2922 87072
rect 2858 87012 2862 87068
rect 2862 87012 2918 87068
rect 2918 87012 2922 87068
rect 2858 87008 2922 87012
rect 5952 87068 6016 87072
rect 5952 87012 5956 87068
rect 5956 87012 6012 87068
rect 6012 87012 6016 87068
rect 5952 87008 6016 87012
rect 6032 87068 6096 87072
rect 6032 87012 6036 87068
rect 6036 87012 6092 87068
rect 6092 87012 6096 87068
rect 6032 87008 6096 87012
rect 6112 87068 6176 87072
rect 6112 87012 6116 87068
rect 6116 87012 6172 87068
rect 6172 87012 6176 87068
rect 6112 87008 6176 87012
rect 6192 87068 6256 87072
rect 6192 87012 6196 87068
rect 6196 87012 6252 87068
rect 6252 87012 6256 87068
rect 6192 87008 6256 87012
rect 4285 86524 4349 86528
rect 4285 86468 4289 86524
rect 4289 86468 4345 86524
rect 4345 86468 4349 86524
rect 4285 86464 4349 86468
rect 4365 86524 4429 86528
rect 4365 86468 4369 86524
rect 4369 86468 4425 86524
rect 4425 86468 4429 86524
rect 4365 86464 4429 86468
rect 4445 86524 4509 86528
rect 4445 86468 4449 86524
rect 4449 86468 4505 86524
rect 4505 86468 4509 86524
rect 4445 86464 4509 86468
rect 4525 86524 4589 86528
rect 4525 86468 4529 86524
rect 4529 86468 4585 86524
rect 4585 86468 4589 86524
rect 4525 86464 4589 86468
rect 7618 86524 7682 86528
rect 7618 86468 7622 86524
rect 7622 86468 7678 86524
rect 7678 86468 7682 86524
rect 7618 86464 7682 86468
rect 7698 86524 7762 86528
rect 7698 86468 7702 86524
rect 7702 86468 7758 86524
rect 7758 86468 7762 86524
rect 7698 86464 7762 86468
rect 7778 86524 7842 86528
rect 7778 86468 7782 86524
rect 7782 86468 7838 86524
rect 7838 86468 7842 86524
rect 7778 86464 7842 86468
rect 7858 86524 7922 86528
rect 7858 86468 7862 86524
rect 7862 86468 7918 86524
rect 7918 86468 7922 86524
rect 7858 86464 7922 86468
rect 2618 85980 2682 85984
rect 2618 85924 2622 85980
rect 2622 85924 2678 85980
rect 2678 85924 2682 85980
rect 2618 85920 2682 85924
rect 2698 85980 2762 85984
rect 2698 85924 2702 85980
rect 2702 85924 2758 85980
rect 2758 85924 2762 85980
rect 2698 85920 2762 85924
rect 2778 85980 2842 85984
rect 2778 85924 2782 85980
rect 2782 85924 2838 85980
rect 2838 85924 2842 85980
rect 2778 85920 2842 85924
rect 2858 85980 2922 85984
rect 2858 85924 2862 85980
rect 2862 85924 2918 85980
rect 2918 85924 2922 85980
rect 2858 85920 2922 85924
rect 5952 85980 6016 85984
rect 5952 85924 5956 85980
rect 5956 85924 6012 85980
rect 6012 85924 6016 85980
rect 5952 85920 6016 85924
rect 6032 85980 6096 85984
rect 6032 85924 6036 85980
rect 6036 85924 6092 85980
rect 6092 85924 6096 85980
rect 6032 85920 6096 85924
rect 6112 85980 6176 85984
rect 6112 85924 6116 85980
rect 6116 85924 6172 85980
rect 6172 85924 6176 85980
rect 6112 85920 6176 85924
rect 6192 85980 6256 85984
rect 6192 85924 6196 85980
rect 6196 85924 6252 85980
rect 6252 85924 6256 85980
rect 6192 85920 6256 85924
rect 4285 85436 4349 85440
rect 4285 85380 4289 85436
rect 4289 85380 4345 85436
rect 4345 85380 4349 85436
rect 4285 85376 4349 85380
rect 4365 85436 4429 85440
rect 4365 85380 4369 85436
rect 4369 85380 4425 85436
rect 4425 85380 4429 85436
rect 4365 85376 4429 85380
rect 4445 85436 4509 85440
rect 4445 85380 4449 85436
rect 4449 85380 4505 85436
rect 4505 85380 4509 85436
rect 4445 85376 4509 85380
rect 4525 85436 4589 85440
rect 4525 85380 4529 85436
rect 4529 85380 4585 85436
rect 4585 85380 4589 85436
rect 4525 85376 4589 85380
rect 7618 85436 7682 85440
rect 7618 85380 7622 85436
rect 7622 85380 7678 85436
rect 7678 85380 7682 85436
rect 7618 85376 7682 85380
rect 7698 85436 7762 85440
rect 7698 85380 7702 85436
rect 7702 85380 7758 85436
rect 7758 85380 7762 85436
rect 7698 85376 7762 85380
rect 7778 85436 7842 85440
rect 7778 85380 7782 85436
rect 7782 85380 7838 85436
rect 7838 85380 7842 85436
rect 7778 85376 7842 85380
rect 7858 85436 7922 85440
rect 7858 85380 7862 85436
rect 7862 85380 7918 85436
rect 7918 85380 7922 85436
rect 7858 85376 7922 85380
rect 2618 84892 2682 84896
rect 2618 84836 2622 84892
rect 2622 84836 2678 84892
rect 2678 84836 2682 84892
rect 2618 84832 2682 84836
rect 2698 84892 2762 84896
rect 2698 84836 2702 84892
rect 2702 84836 2758 84892
rect 2758 84836 2762 84892
rect 2698 84832 2762 84836
rect 2778 84892 2842 84896
rect 2778 84836 2782 84892
rect 2782 84836 2838 84892
rect 2838 84836 2842 84892
rect 2778 84832 2842 84836
rect 2858 84892 2922 84896
rect 2858 84836 2862 84892
rect 2862 84836 2918 84892
rect 2918 84836 2922 84892
rect 2858 84832 2922 84836
rect 5952 84892 6016 84896
rect 5952 84836 5956 84892
rect 5956 84836 6012 84892
rect 6012 84836 6016 84892
rect 5952 84832 6016 84836
rect 6032 84892 6096 84896
rect 6032 84836 6036 84892
rect 6036 84836 6092 84892
rect 6092 84836 6096 84892
rect 6032 84832 6096 84836
rect 6112 84892 6176 84896
rect 6112 84836 6116 84892
rect 6116 84836 6172 84892
rect 6172 84836 6176 84892
rect 6112 84832 6176 84836
rect 6192 84892 6256 84896
rect 6192 84836 6196 84892
rect 6196 84836 6252 84892
rect 6252 84836 6256 84892
rect 6192 84832 6256 84836
rect 4285 84348 4349 84352
rect 4285 84292 4289 84348
rect 4289 84292 4345 84348
rect 4345 84292 4349 84348
rect 4285 84288 4349 84292
rect 4365 84348 4429 84352
rect 4365 84292 4369 84348
rect 4369 84292 4425 84348
rect 4425 84292 4429 84348
rect 4365 84288 4429 84292
rect 4445 84348 4509 84352
rect 4445 84292 4449 84348
rect 4449 84292 4505 84348
rect 4505 84292 4509 84348
rect 4445 84288 4509 84292
rect 4525 84348 4589 84352
rect 4525 84292 4529 84348
rect 4529 84292 4585 84348
rect 4585 84292 4589 84348
rect 4525 84288 4589 84292
rect 7618 84348 7682 84352
rect 7618 84292 7622 84348
rect 7622 84292 7678 84348
rect 7678 84292 7682 84348
rect 7618 84288 7682 84292
rect 7698 84348 7762 84352
rect 7698 84292 7702 84348
rect 7702 84292 7758 84348
rect 7758 84292 7762 84348
rect 7698 84288 7762 84292
rect 7778 84348 7842 84352
rect 7778 84292 7782 84348
rect 7782 84292 7838 84348
rect 7838 84292 7842 84348
rect 7778 84288 7842 84292
rect 7858 84348 7922 84352
rect 7858 84292 7862 84348
rect 7862 84292 7918 84348
rect 7918 84292 7922 84348
rect 7858 84288 7922 84292
rect 2618 83804 2682 83808
rect 2618 83748 2622 83804
rect 2622 83748 2678 83804
rect 2678 83748 2682 83804
rect 2618 83744 2682 83748
rect 2698 83804 2762 83808
rect 2698 83748 2702 83804
rect 2702 83748 2758 83804
rect 2758 83748 2762 83804
rect 2698 83744 2762 83748
rect 2778 83804 2842 83808
rect 2778 83748 2782 83804
rect 2782 83748 2838 83804
rect 2838 83748 2842 83804
rect 2778 83744 2842 83748
rect 2858 83804 2922 83808
rect 2858 83748 2862 83804
rect 2862 83748 2918 83804
rect 2918 83748 2922 83804
rect 2858 83744 2922 83748
rect 5952 83804 6016 83808
rect 5952 83748 5956 83804
rect 5956 83748 6012 83804
rect 6012 83748 6016 83804
rect 5952 83744 6016 83748
rect 6032 83804 6096 83808
rect 6032 83748 6036 83804
rect 6036 83748 6092 83804
rect 6092 83748 6096 83804
rect 6032 83744 6096 83748
rect 6112 83804 6176 83808
rect 6112 83748 6116 83804
rect 6116 83748 6172 83804
rect 6172 83748 6176 83804
rect 6112 83744 6176 83748
rect 6192 83804 6256 83808
rect 6192 83748 6196 83804
rect 6196 83748 6252 83804
rect 6252 83748 6256 83804
rect 6192 83744 6256 83748
rect 4285 83260 4349 83264
rect 4285 83204 4289 83260
rect 4289 83204 4345 83260
rect 4345 83204 4349 83260
rect 4285 83200 4349 83204
rect 4365 83260 4429 83264
rect 4365 83204 4369 83260
rect 4369 83204 4425 83260
rect 4425 83204 4429 83260
rect 4365 83200 4429 83204
rect 4445 83260 4509 83264
rect 4445 83204 4449 83260
rect 4449 83204 4505 83260
rect 4505 83204 4509 83260
rect 4445 83200 4509 83204
rect 4525 83260 4589 83264
rect 4525 83204 4529 83260
rect 4529 83204 4585 83260
rect 4585 83204 4589 83260
rect 4525 83200 4589 83204
rect 7618 83260 7682 83264
rect 7618 83204 7622 83260
rect 7622 83204 7678 83260
rect 7678 83204 7682 83260
rect 7618 83200 7682 83204
rect 7698 83260 7762 83264
rect 7698 83204 7702 83260
rect 7702 83204 7758 83260
rect 7758 83204 7762 83260
rect 7698 83200 7762 83204
rect 7778 83260 7842 83264
rect 7778 83204 7782 83260
rect 7782 83204 7838 83260
rect 7838 83204 7842 83260
rect 7778 83200 7842 83204
rect 7858 83260 7922 83264
rect 7858 83204 7862 83260
rect 7862 83204 7918 83260
rect 7918 83204 7922 83260
rect 7858 83200 7922 83204
rect 2618 82716 2682 82720
rect 2618 82660 2622 82716
rect 2622 82660 2678 82716
rect 2678 82660 2682 82716
rect 2618 82656 2682 82660
rect 2698 82716 2762 82720
rect 2698 82660 2702 82716
rect 2702 82660 2758 82716
rect 2758 82660 2762 82716
rect 2698 82656 2762 82660
rect 2778 82716 2842 82720
rect 2778 82660 2782 82716
rect 2782 82660 2838 82716
rect 2838 82660 2842 82716
rect 2778 82656 2842 82660
rect 2858 82716 2922 82720
rect 2858 82660 2862 82716
rect 2862 82660 2918 82716
rect 2918 82660 2922 82716
rect 2858 82656 2922 82660
rect 5952 82716 6016 82720
rect 5952 82660 5956 82716
rect 5956 82660 6012 82716
rect 6012 82660 6016 82716
rect 5952 82656 6016 82660
rect 6032 82716 6096 82720
rect 6032 82660 6036 82716
rect 6036 82660 6092 82716
rect 6092 82660 6096 82716
rect 6032 82656 6096 82660
rect 6112 82716 6176 82720
rect 6112 82660 6116 82716
rect 6116 82660 6172 82716
rect 6172 82660 6176 82716
rect 6112 82656 6176 82660
rect 6192 82716 6256 82720
rect 6192 82660 6196 82716
rect 6196 82660 6252 82716
rect 6252 82660 6256 82716
rect 6192 82656 6256 82660
rect 4285 82172 4349 82176
rect 4285 82116 4289 82172
rect 4289 82116 4345 82172
rect 4345 82116 4349 82172
rect 4285 82112 4349 82116
rect 4365 82172 4429 82176
rect 4365 82116 4369 82172
rect 4369 82116 4425 82172
rect 4425 82116 4429 82172
rect 4365 82112 4429 82116
rect 4445 82172 4509 82176
rect 4445 82116 4449 82172
rect 4449 82116 4505 82172
rect 4505 82116 4509 82172
rect 4445 82112 4509 82116
rect 4525 82172 4589 82176
rect 4525 82116 4529 82172
rect 4529 82116 4585 82172
rect 4585 82116 4589 82172
rect 4525 82112 4589 82116
rect 7618 82172 7682 82176
rect 7618 82116 7622 82172
rect 7622 82116 7678 82172
rect 7678 82116 7682 82172
rect 7618 82112 7682 82116
rect 7698 82172 7762 82176
rect 7698 82116 7702 82172
rect 7702 82116 7758 82172
rect 7758 82116 7762 82172
rect 7698 82112 7762 82116
rect 7778 82172 7842 82176
rect 7778 82116 7782 82172
rect 7782 82116 7838 82172
rect 7838 82116 7842 82172
rect 7778 82112 7842 82116
rect 7858 82172 7922 82176
rect 7858 82116 7862 82172
rect 7862 82116 7918 82172
rect 7918 82116 7922 82172
rect 7858 82112 7922 82116
rect 2618 81628 2682 81632
rect 2618 81572 2622 81628
rect 2622 81572 2678 81628
rect 2678 81572 2682 81628
rect 2618 81568 2682 81572
rect 2698 81628 2762 81632
rect 2698 81572 2702 81628
rect 2702 81572 2758 81628
rect 2758 81572 2762 81628
rect 2698 81568 2762 81572
rect 2778 81628 2842 81632
rect 2778 81572 2782 81628
rect 2782 81572 2838 81628
rect 2838 81572 2842 81628
rect 2778 81568 2842 81572
rect 2858 81628 2922 81632
rect 2858 81572 2862 81628
rect 2862 81572 2918 81628
rect 2918 81572 2922 81628
rect 2858 81568 2922 81572
rect 5952 81628 6016 81632
rect 5952 81572 5956 81628
rect 5956 81572 6012 81628
rect 6012 81572 6016 81628
rect 5952 81568 6016 81572
rect 6032 81628 6096 81632
rect 6032 81572 6036 81628
rect 6036 81572 6092 81628
rect 6092 81572 6096 81628
rect 6032 81568 6096 81572
rect 6112 81628 6176 81632
rect 6112 81572 6116 81628
rect 6116 81572 6172 81628
rect 6172 81572 6176 81628
rect 6112 81568 6176 81572
rect 6192 81628 6256 81632
rect 6192 81572 6196 81628
rect 6196 81572 6252 81628
rect 6252 81572 6256 81628
rect 6192 81568 6256 81572
rect 4285 81084 4349 81088
rect 4285 81028 4289 81084
rect 4289 81028 4345 81084
rect 4345 81028 4349 81084
rect 4285 81024 4349 81028
rect 4365 81084 4429 81088
rect 4365 81028 4369 81084
rect 4369 81028 4425 81084
rect 4425 81028 4429 81084
rect 4365 81024 4429 81028
rect 4445 81084 4509 81088
rect 4445 81028 4449 81084
rect 4449 81028 4505 81084
rect 4505 81028 4509 81084
rect 4445 81024 4509 81028
rect 4525 81084 4589 81088
rect 4525 81028 4529 81084
rect 4529 81028 4585 81084
rect 4585 81028 4589 81084
rect 4525 81024 4589 81028
rect 7618 81084 7682 81088
rect 7618 81028 7622 81084
rect 7622 81028 7678 81084
rect 7678 81028 7682 81084
rect 7618 81024 7682 81028
rect 7698 81084 7762 81088
rect 7698 81028 7702 81084
rect 7702 81028 7758 81084
rect 7758 81028 7762 81084
rect 7698 81024 7762 81028
rect 7778 81084 7842 81088
rect 7778 81028 7782 81084
rect 7782 81028 7838 81084
rect 7838 81028 7842 81084
rect 7778 81024 7842 81028
rect 7858 81084 7922 81088
rect 7858 81028 7862 81084
rect 7862 81028 7918 81084
rect 7918 81028 7922 81084
rect 7858 81024 7922 81028
rect 2618 80540 2682 80544
rect 2618 80484 2622 80540
rect 2622 80484 2678 80540
rect 2678 80484 2682 80540
rect 2618 80480 2682 80484
rect 2698 80540 2762 80544
rect 2698 80484 2702 80540
rect 2702 80484 2758 80540
rect 2758 80484 2762 80540
rect 2698 80480 2762 80484
rect 2778 80540 2842 80544
rect 2778 80484 2782 80540
rect 2782 80484 2838 80540
rect 2838 80484 2842 80540
rect 2778 80480 2842 80484
rect 2858 80540 2922 80544
rect 2858 80484 2862 80540
rect 2862 80484 2918 80540
rect 2918 80484 2922 80540
rect 2858 80480 2922 80484
rect 5952 80540 6016 80544
rect 5952 80484 5956 80540
rect 5956 80484 6012 80540
rect 6012 80484 6016 80540
rect 5952 80480 6016 80484
rect 6032 80540 6096 80544
rect 6032 80484 6036 80540
rect 6036 80484 6092 80540
rect 6092 80484 6096 80540
rect 6032 80480 6096 80484
rect 6112 80540 6176 80544
rect 6112 80484 6116 80540
rect 6116 80484 6172 80540
rect 6172 80484 6176 80540
rect 6112 80480 6176 80484
rect 6192 80540 6256 80544
rect 6192 80484 6196 80540
rect 6196 80484 6252 80540
rect 6252 80484 6256 80540
rect 6192 80480 6256 80484
rect 4285 79996 4349 80000
rect 4285 79940 4289 79996
rect 4289 79940 4345 79996
rect 4345 79940 4349 79996
rect 4285 79936 4349 79940
rect 4365 79996 4429 80000
rect 4365 79940 4369 79996
rect 4369 79940 4425 79996
rect 4425 79940 4429 79996
rect 4365 79936 4429 79940
rect 4445 79996 4509 80000
rect 4445 79940 4449 79996
rect 4449 79940 4505 79996
rect 4505 79940 4509 79996
rect 4445 79936 4509 79940
rect 4525 79996 4589 80000
rect 4525 79940 4529 79996
rect 4529 79940 4585 79996
rect 4585 79940 4589 79996
rect 4525 79936 4589 79940
rect 7618 79996 7682 80000
rect 7618 79940 7622 79996
rect 7622 79940 7678 79996
rect 7678 79940 7682 79996
rect 7618 79936 7682 79940
rect 7698 79996 7762 80000
rect 7698 79940 7702 79996
rect 7702 79940 7758 79996
rect 7758 79940 7762 79996
rect 7698 79936 7762 79940
rect 7778 79996 7842 80000
rect 7778 79940 7782 79996
rect 7782 79940 7838 79996
rect 7838 79940 7842 79996
rect 7778 79936 7842 79940
rect 7858 79996 7922 80000
rect 7858 79940 7862 79996
rect 7862 79940 7918 79996
rect 7918 79940 7922 79996
rect 7858 79936 7922 79940
rect 2618 79452 2682 79456
rect 2618 79396 2622 79452
rect 2622 79396 2678 79452
rect 2678 79396 2682 79452
rect 2618 79392 2682 79396
rect 2698 79452 2762 79456
rect 2698 79396 2702 79452
rect 2702 79396 2758 79452
rect 2758 79396 2762 79452
rect 2698 79392 2762 79396
rect 2778 79452 2842 79456
rect 2778 79396 2782 79452
rect 2782 79396 2838 79452
rect 2838 79396 2842 79452
rect 2778 79392 2842 79396
rect 2858 79452 2922 79456
rect 2858 79396 2862 79452
rect 2862 79396 2918 79452
rect 2918 79396 2922 79452
rect 2858 79392 2922 79396
rect 5952 79452 6016 79456
rect 5952 79396 5956 79452
rect 5956 79396 6012 79452
rect 6012 79396 6016 79452
rect 5952 79392 6016 79396
rect 6032 79452 6096 79456
rect 6032 79396 6036 79452
rect 6036 79396 6092 79452
rect 6092 79396 6096 79452
rect 6032 79392 6096 79396
rect 6112 79452 6176 79456
rect 6112 79396 6116 79452
rect 6116 79396 6172 79452
rect 6172 79396 6176 79452
rect 6112 79392 6176 79396
rect 6192 79452 6256 79456
rect 6192 79396 6196 79452
rect 6196 79396 6252 79452
rect 6252 79396 6256 79452
rect 6192 79392 6256 79396
rect 4285 78908 4349 78912
rect 4285 78852 4289 78908
rect 4289 78852 4345 78908
rect 4345 78852 4349 78908
rect 4285 78848 4349 78852
rect 4365 78908 4429 78912
rect 4365 78852 4369 78908
rect 4369 78852 4425 78908
rect 4425 78852 4429 78908
rect 4365 78848 4429 78852
rect 4445 78908 4509 78912
rect 4445 78852 4449 78908
rect 4449 78852 4505 78908
rect 4505 78852 4509 78908
rect 4445 78848 4509 78852
rect 4525 78908 4589 78912
rect 4525 78852 4529 78908
rect 4529 78852 4585 78908
rect 4585 78852 4589 78908
rect 4525 78848 4589 78852
rect 7618 78908 7682 78912
rect 7618 78852 7622 78908
rect 7622 78852 7678 78908
rect 7678 78852 7682 78908
rect 7618 78848 7682 78852
rect 7698 78908 7762 78912
rect 7698 78852 7702 78908
rect 7702 78852 7758 78908
rect 7758 78852 7762 78908
rect 7698 78848 7762 78852
rect 7778 78908 7842 78912
rect 7778 78852 7782 78908
rect 7782 78852 7838 78908
rect 7838 78852 7842 78908
rect 7778 78848 7842 78852
rect 7858 78908 7922 78912
rect 7858 78852 7862 78908
rect 7862 78852 7918 78908
rect 7918 78852 7922 78908
rect 7858 78848 7922 78852
rect 2618 78364 2682 78368
rect 2618 78308 2622 78364
rect 2622 78308 2678 78364
rect 2678 78308 2682 78364
rect 2618 78304 2682 78308
rect 2698 78364 2762 78368
rect 2698 78308 2702 78364
rect 2702 78308 2758 78364
rect 2758 78308 2762 78364
rect 2698 78304 2762 78308
rect 2778 78364 2842 78368
rect 2778 78308 2782 78364
rect 2782 78308 2838 78364
rect 2838 78308 2842 78364
rect 2778 78304 2842 78308
rect 2858 78364 2922 78368
rect 2858 78308 2862 78364
rect 2862 78308 2918 78364
rect 2918 78308 2922 78364
rect 2858 78304 2922 78308
rect 5952 78364 6016 78368
rect 5952 78308 5956 78364
rect 5956 78308 6012 78364
rect 6012 78308 6016 78364
rect 5952 78304 6016 78308
rect 6032 78364 6096 78368
rect 6032 78308 6036 78364
rect 6036 78308 6092 78364
rect 6092 78308 6096 78364
rect 6032 78304 6096 78308
rect 6112 78364 6176 78368
rect 6112 78308 6116 78364
rect 6116 78308 6172 78364
rect 6172 78308 6176 78364
rect 6112 78304 6176 78308
rect 6192 78364 6256 78368
rect 6192 78308 6196 78364
rect 6196 78308 6252 78364
rect 6252 78308 6256 78364
rect 6192 78304 6256 78308
rect 4285 77820 4349 77824
rect 4285 77764 4289 77820
rect 4289 77764 4345 77820
rect 4345 77764 4349 77820
rect 4285 77760 4349 77764
rect 4365 77820 4429 77824
rect 4365 77764 4369 77820
rect 4369 77764 4425 77820
rect 4425 77764 4429 77820
rect 4365 77760 4429 77764
rect 4445 77820 4509 77824
rect 4445 77764 4449 77820
rect 4449 77764 4505 77820
rect 4505 77764 4509 77820
rect 4445 77760 4509 77764
rect 4525 77820 4589 77824
rect 4525 77764 4529 77820
rect 4529 77764 4585 77820
rect 4585 77764 4589 77820
rect 4525 77760 4589 77764
rect 7618 77820 7682 77824
rect 7618 77764 7622 77820
rect 7622 77764 7678 77820
rect 7678 77764 7682 77820
rect 7618 77760 7682 77764
rect 7698 77820 7762 77824
rect 7698 77764 7702 77820
rect 7702 77764 7758 77820
rect 7758 77764 7762 77820
rect 7698 77760 7762 77764
rect 7778 77820 7842 77824
rect 7778 77764 7782 77820
rect 7782 77764 7838 77820
rect 7838 77764 7842 77820
rect 7778 77760 7842 77764
rect 7858 77820 7922 77824
rect 7858 77764 7862 77820
rect 7862 77764 7918 77820
rect 7918 77764 7922 77820
rect 7858 77760 7922 77764
rect 2618 77276 2682 77280
rect 2618 77220 2622 77276
rect 2622 77220 2678 77276
rect 2678 77220 2682 77276
rect 2618 77216 2682 77220
rect 2698 77276 2762 77280
rect 2698 77220 2702 77276
rect 2702 77220 2758 77276
rect 2758 77220 2762 77276
rect 2698 77216 2762 77220
rect 2778 77276 2842 77280
rect 2778 77220 2782 77276
rect 2782 77220 2838 77276
rect 2838 77220 2842 77276
rect 2778 77216 2842 77220
rect 2858 77276 2922 77280
rect 2858 77220 2862 77276
rect 2862 77220 2918 77276
rect 2918 77220 2922 77276
rect 2858 77216 2922 77220
rect 5952 77276 6016 77280
rect 5952 77220 5956 77276
rect 5956 77220 6012 77276
rect 6012 77220 6016 77276
rect 5952 77216 6016 77220
rect 6032 77276 6096 77280
rect 6032 77220 6036 77276
rect 6036 77220 6092 77276
rect 6092 77220 6096 77276
rect 6032 77216 6096 77220
rect 6112 77276 6176 77280
rect 6112 77220 6116 77276
rect 6116 77220 6172 77276
rect 6172 77220 6176 77276
rect 6112 77216 6176 77220
rect 6192 77276 6256 77280
rect 6192 77220 6196 77276
rect 6196 77220 6252 77276
rect 6252 77220 6256 77276
rect 6192 77216 6256 77220
rect 4285 76732 4349 76736
rect 4285 76676 4289 76732
rect 4289 76676 4345 76732
rect 4345 76676 4349 76732
rect 4285 76672 4349 76676
rect 4365 76732 4429 76736
rect 4365 76676 4369 76732
rect 4369 76676 4425 76732
rect 4425 76676 4429 76732
rect 4365 76672 4429 76676
rect 4445 76732 4509 76736
rect 4445 76676 4449 76732
rect 4449 76676 4505 76732
rect 4505 76676 4509 76732
rect 4445 76672 4509 76676
rect 4525 76732 4589 76736
rect 4525 76676 4529 76732
rect 4529 76676 4585 76732
rect 4585 76676 4589 76732
rect 4525 76672 4589 76676
rect 7618 76732 7682 76736
rect 7618 76676 7622 76732
rect 7622 76676 7678 76732
rect 7678 76676 7682 76732
rect 7618 76672 7682 76676
rect 7698 76732 7762 76736
rect 7698 76676 7702 76732
rect 7702 76676 7758 76732
rect 7758 76676 7762 76732
rect 7698 76672 7762 76676
rect 7778 76732 7842 76736
rect 7778 76676 7782 76732
rect 7782 76676 7838 76732
rect 7838 76676 7842 76732
rect 7778 76672 7842 76676
rect 7858 76732 7922 76736
rect 7858 76676 7862 76732
rect 7862 76676 7918 76732
rect 7918 76676 7922 76732
rect 7858 76672 7922 76676
rect 2618 76188 2682 76192
rect 2618 76132 2622 76188
rect 2622 76132 2678 76188
rect 2678 76132 2682 76188
rect 2618 76128 2682 76132
rect 2698 76188 2762 76192
rect 2698 76132 2702 76188
rect 2702 76132 2758 76188
rect 2758 76132 2762 76188
rect 2698 76128 2762 76132
rect 2778 76188 2842 76192
rect 2778 76132 2782 76188
rect 2782 76132 2838 76188
rect 2838 76132 2842 76188
rect 2778 76128 2842 76132
rect 2858 76188 2922 76192
rect 2858 76132 2862 76188
rect 2862 76132 2918 76188
rect 2918 76132 2922 76188
rect 2858 76128 2922 76132
rect 5952 76188 6016 76192
rect 5952 76132 5956 76188
rect 5956 76132 6012 76188
rect 6012 76132 6016 76188
rect 5952 76128 6016 76132
rect 6032 76188 6096 76192
rect 6032 76132 6036 76188
rect 6036 76132 6092 76188
rect 6092 76132 6096 76188
rect 6032 76128 6096 76132
rect 6112 76188 6176 76192
rect 6112 76132 6116 76188
rect 6116 76132 6172 76188
rect 6172 76132 6176 76188
rect 6112 76128 6176 76132
rect 6192 76188 6256 76192
rect 6192 76132 6196 76188
rect 6196 76132 6252 76188
rect 6252 76132 6256 76188
rect 6192 76128 6256 76132
rect 4285 75644 4349 75648
rect 4285 75588 4289 75644
rect 4289 75588 4345 75644
rect 4345 75588 4349 75644
rect 4285 75584 4349 75588
rect 4365 75644 4429 75648
rect 4365 75588 4369 75644
rect 4369 75588 4425 75644
rect 4425 75588 4429 75644
rect 4365 75584 4429 75588
rect 4445 75644 4509 75648
rect 4445 75588 4449 75644
rect 4449 75588 4505 75644
rect 4505 75588 4509 75644
rect 4445 75584 4509 75588
rect 4525 75644 4589 75648
rect 4525 75588 4529 75644
rect 4529 75588 4585 75644
rect 4585 75588 4589 75644
rect 4525 75584 4589 75588
rect 7618 75644 7682 75648
rect 7618 75588 7622 75644
rect 7622 75588 7678 75644
rect 7678 75588 7682 75644
rect 7618 75584 7682 75588
rect 7698 75644 7762 75648
rect 7698 75588 7702 75644
rect 7702 75588 7758 75644
rect 7758 75588 7762 75644
rect 7698 75584 7762 75588
rect 7778 75644 7842 75648
rect 7778 75588 7782 75644
rect 7782 75588 7838 75644
rect 7838 75588 7842 75644
rect 7778 75584 7842 75588
rect 7858 75644 7922 75648
rect 7858 75588 7862 75644
rect 7862 75588 7918 75644
rect 7918 75588 7922 75644
rect 7858 75584 7922 75588
rect 2618 75100 2682 75104
rect 2618 75044 2622 75100
rect 2622 75044 2678 75100
rect 2678 75044 2682 75100
rect 2618 75040 2682 75044
rect 2698 75100 2762 75104
rect 2698 75044 2702 75100
rect 2702 75044 2758 75100
rect 2758 75044 2762 75100
rect 2698 75040 2762 75044
rect 2778 75100 2842 75104
rect 2778 75044 2782 75100
rect 2782 75044 2838 75100
rect 2838 75044 2842 75100
rect 2778 75040 2842 75044
rect 2858 75100 2922 75104
rect 2858 75044 2862 75100
rect 2862 75044 2918 75100
rect 2918 75044 2922 75100
rect 2858 75040 2922 75044
rect 5952 75100 6016 75104
rect 5952 75044 5956 75100
rect 5956 75044 6012 75100
rect 6012 75044 6016 75100
rect 5952 75040 6016 75044
rect 6032 75100 6096 75104
rect 6032 75044 6036 75100
rect 6036 75044 6092 75100
rect 6092 75044 6096 75100
rect 6032 75040 6096 75044
rect 6112 75100 6176 75104
rect 6112 75044 6116 75100
rect 6116 75044 6172 75100
rect 6172 75044 6176 75100
rect 6112 75040 6176 75044
rect 6192 75100 6256 75104
rect 6192 75044 6196 75100
rect 6196 75044 6252 75100
rect 6252 75044 6256 75100
rect 6192 75040 6256 75044
rect 4285 74556 4349 74560
rect 4285 74500 4289 74556
rect 4289 74500 4345 74556
rect 4345 74500 4349 74556
rect 4285 74496 4349 74500
rect 4365 74556 4429 74560
rect 4365 74500 4369 74556
rect 4369 74500 4425 74556
rect 4425 74500 4429 74556
rect 4365 74496 4429 74500
rect 4445 74556 4509 74560
rect 4445 74500 4449 74556
rect 4449 74500 4505 74556
rect 4505 74500 4509 74556
rect 4445 74496 4509 74500
rect 4525 74556 4589 74560
rect 4525 74500 4529 74556
rect 4529 74500 4585 74556
rect 4585 74500 4589 74556
rect 4525 74496 4589 74500
rect 7618 74556 7682 74560
rect 7618 74500 7622 74556
rect 7622 74500 7678 74556
rect 7678 74500 7682 74556
rect 7618 74496 7682 74500
rect 7698 74556 7762 74560
rect 7698 74500 7702 74556
rect 7702 74500 7758 74556
rect 7758 74500 7762 74556
rect 7698 74496 7762 74500
rect 7778 74556 7842 74560
rect 7778 74500 7782 74556
rect 7782 74500 7838 74556
rect 7838 74500 7842 74556
rect 7778 74496 7842 74500
rect 7858 74556 7922 74560
rect 7858 74500 7862 74556
rect 7862 74500 7918 74556
rect 7918 74500 7922 74556
rect 7858 74496 7922 74500
rect 2618 74012 2682 74016
rect 2618 73956 2622 74012
rect 2622 73956 2678 74012
rect 2678 73956 2682 74012
rect 2618 73952 2682 73956
rect 2698 74012 2762 74016
rect 2698 73956 2702 74012
rect 2702 73956 2758 74012
rect 2758 73956 2762 74012
rect 2698 73952 2762 73956
rect 2778 74012 2842 74016
rect 2778 73956 2782 74012
rect 2782 73956 2838 74012
rect 2838 73956 2842 74012
rect 2778 73952 2842 73956
rect 2858 74012 2922 74016
rect 2858 73956 2862 74012
rect 2862 73956 2918 74012
rect 2918 73956 2922 74012
rect 2858 73952 2922 73956
rect 5952 74012 6016 74016
rect 5952 73956 5956 74012
rect 5956 73956 6012 74012
rect 6012 73956 6016 74012
rect 5952 73952 6016 73956
rect 6032 74012 6096 74016
rect 6032 73956 6036 74012
rect 6036 73956 6092 74012
rect 6092 73956 6096 74012
rect 6032 73952 6096 73956
rect 6112 74012 6176 74016
rect 6112 73956 6116 74012
rect 6116 73956 6172 74012
rect 6172 73956 6176 74012
rect 6112 73952 6176 73956
rect 6192 74012 6256 74016
rect 6192 73956 6196 74012
rect 6196 73956 6252 74012
rect 6252 73956 6256 74012
rect 6192 73952 6256 73956
rect 4285 73468 4349 73472
rect 4285 73412 4289 73468
rect 4289 73412 4345 73468
rect 4345 73412 4349 73468
rect 4285 73408 4349 73412
rect 4365 73468 4429 73472
rect 4365 73412 4369 73468
rect 4369 73412 4425 73468
rect 4425 73412 4429 73468
rect 4365 73408 4429 73412
rect 4445 73468 4509 73472
rect 4445 73412 4449 73468
rect 4449 73412 4505 73468
rect 4505 73412 4509 73468
rect 4445 73408 4509 73412
rect 4525 73468 4589 73472
rect 4525 73412 4529 73468
rect 4529 73412 4585 73468
rect 4585 73412 4589 73468
rect 4525 73408 4589 73412
rect 7618 73468 7682 73472
rect 7618 73412 7622 73468
rect 7622 73412 7678 73468
rect 7678 73412 7682 73468
rect 7618 73408 7682 73412
rect 7698 73468 7762 73472
rect 7698 73412 7702 73468
rect 7702 73412 7758 73468
rect 7758 73412 7762 73468
rect 7698 73408 7762 73412
rect 7778 73468 7842 73472
rect 7778 73412 7782 73468
rect 7782 73412 7838 73468
rect 7838 73412 7842 73468
rect 7778 73408 7842 73412
rect 7858 73468 7922 73472
rect 7858 73412 7862 73468
rect 7862 73412 7918 73468
rect 7918 73412 7922 73468
rect 7858 73408 7922 73412
rect 2618 72924 2682 72928
rect 2618 72868 2622 72924
rect 2622 72868 2678 72924
rect 2678 72868 2682 72924
rect 2618 72864 2682 72868
rect 2698 72924 2762 72928
rect 2698 72868 2702 72924
rect 2702 72868 2758 72924
rect 2758 72868 2762 72924
rect 2698 72864 2762 72868
rect 2778 72924 2842 72928
rect 2778 72868 2782 72924
rect 2782 72868 2838 72924
rect 2838 72868 2842 72924
rect 2778 72864 2842 72868
rect 2858 72924 2922 72928
rect 2858 72868 2862 72924
rect 2862 72868 2918 72924
rect 2918 72868 2922 72924
rect 2858 72864 2922 72868
rect 5952 72924 6016 72928
rect 5952 72868 5956 72924
rect 5956 72868 6012 72924
rect 6012 72868 6016 72924
rect 5952 72864 6016 72868
rect 6032 72924 6096 72928
rect 6032 72868 6036 72924
rect 6036 72868 6092 72924
rect 6092 72868 6096 72924
rect 6032 72864 6096 72868
rect 6112 72924 6176 72928
rect 6112 72868 6116 72924
rect 6116 72868 6172 72924
rect 6172 72868 6176 72924
rect 6112 72864 6176 72868
rect 6192 72924 6256 72928
rect 6192 72868 6196 72924
rect 6196 72868 6252 72924
rect 6252 72868 6256 72924
rect 6192 72864 6256 72868
rect 4285 72380 4349 72384
rect 4285 72324 4289 72380
rect 4289 72324 4345 72380
rect 4345 72324 4349 72380
rect 4285 72320 4349 72324
rect 4365 72380 4429 72384
rect 4365 72324 4369 72380
rect 4369 72324 4425 72380
rect 4425 72324 4429 72380
rect 4365 72320 4429 72324
rect 4445 72380 4509 72384
rect 4445 72324 4449 72380
rect 4449 72324 4505 72380
rect 4505 72324 4509 72380
rect 4445 72320 4509 72324
rect 4525 72380 4589 72384
rect 4525 72324 4529 72380
rect 4529 72324 4585 72380
rect 4585 72324 4589 72380
rect 4525 72320 4589 72324
rect 7618 72380 7682 72384
rect 7618 72324 7622 72380
rect 7622 72324 7678 72380
rect 7678 72324 7682 72380
rect 7618 72320 7682 72324
rect 7698 72380 7762 72384
rect 7698 72324 7702 72380
rect 7702 72324 7758 72380
rect 7758 72324 7762 72380
rect 7698 72320 7762 72324
rect 7778 72380 7842 72384
rect 7778 72324 7782 72380
rect 7782 72324 7838 72380
rect 7838 72324 7842 72380
rect 7778 72320 7842 72324
rect 7858 72380 7922 72384
rect 7858 72324 7862 72380
rect 7862 72324 7918 72380
rect 7918 72324 7922 72380
rect 7858 72320 7922 72324
rect 2618 71836 2682 71840
rect 2618 71780 2622 71836
rect 2622 71780 2678 71836
rect 2678 71780 2682 71836
rect 2618 71776 2682 71780
rect 2698 71836 2762 71840
rect 2698 71780 2702 71836
rect 2702 71780 2758 71836
rect 2758 71780 2762 71836
rect 2698 71776 2762 71780
rect 2778 71836 2842 71840
rect 2778 71780 2782 71836
rect 2782 71780 2838 71836
rect 2838 71780 2842 71836
rect 2778 71776 2842 71780
rect 2858 71836 2922 71840
rect 2858 71780 2862 71836
rect 2862 71780 2918 71836
rect 2918 71780 2922 71836
rect 2858 71776 2922 71780
rect 5952 71836 6016 71840
rect 5952 71780 5956 71836
rect 5956 71780 6012 71836
rect 6012 71780 6016 71836
rect 5952 71776 6016 71780
rect 6032 71836 6096 71840
rect 6032 71780 6036 71836
rect 6036 71780 6092 71836
rect 6092 71780 6096 71836
rect 6032 71776 6096 71780
rect 6112 71836 6176 71840
rect 6112 71780 6116 71836
rect 6116 71780 6172 71836
rect 6172 71780 6176 71836
rect 6112 71776 6176 71780
rect 6192 71836 6256 71840
rect 6192 71780 6196 71836
rect 6196 71780 6252 71836
rect 6252 71780 6256 71836
rect 6192 71776 6256 71780
rect 4285 71292 4349 71296
rect 4285 71236 4289 71292
rect 4289 71236 4345 71292
rect 4345 71236 4349 71292
rect 4285 71232 4349 71236
rect 4365 71292 4429 71296
rect 4365 71236 4369 71292
rect 4369 71236 4425 71292
rect 4425 71236 4429 71292
rect 4365 71232 4429 71236
rect 4445 71292 4509 71296
rect 4445 71236 4449 71292
rect 4449 71236 4505 71292
rect 4505 71236 4509 71292
rect 4445 71232 4509 71236
rect 4525 71292 4589 71296
rect 4525 71236 4529 71292
rect 4529 71236 4585 71292
rect 4585 71236 4589 71292
rect 4525 71232 4589 71236
rect 7618 71292 7682 71296
rect 7618 71236 7622 71292
rect 7622 71236 7678 71292
rect 7678 71236 7682 71292
rect 7618 71232 7682 71236
rect 7698 71292 7762 71296
rect 7698 71236 7702 71292
rect 7702 71236 7758 71292
rect 7758 71236 7762 71292
rect 7698 71232 7762 71236
rect 7778 71292 7842 71296
rect 7778 71236 7782 71292
rect 7782 71236 7838 71292
rect 7838 71236 7842 71292
rect 7778 71232 7842 71236
rect 7858 71292 7922 71296
rect 7858 71236 7862 71292
rect 7862 71236 7918 71292
rect 7918 71236 7922 71292
rect 7858 71232 7922 71236
rect 2618 70748 2682 70752
rect 2618 70692 2622 70748
rect 2622 70692 2678 70748
rect 2678 70692 2682 70748
rect 2618 70688 2682 70692
rect 2698 70748 2762 70752
rect 2698 70692 2702 70748
rect 2702 70692 2758 70748
rect 2758 70692 2762 70748
rect 2698 70688 2762 70692
rect 2778 70748 2842 70752
rect 2778 70692 2782 70748
rect 2782 70692 2838 70748
rect 2838 70692 2842 70748
rect 2778 70688 2842 70692
rect 2858 70748 2922 70752
rect 2858 70692 2862 70748
rect 2862 70692 2918 70748
rect 2918 70692 2922 70748
rect 2858 70688 2922 70692
rect 5952 70748 6016 70752
rect 5952 70692 5956 70748
rect 5956 70692 6012 70748
rect 6012 70692 6016 70748
rect 5952 70688 6016 70692
rect 6032 70748 6096 70752
rect 6032 70692 6036 70748
rect 6036 70692 6092 70748
rect 6092 70692 6096 70748
rect 6032 70688 6096 70692
rect 6112 70748 6176 70752
rect 6112 70692 6116 70748
rect 6116 70692 6172 70748
rect 6172 70692 6176 70748
rect 6112 70688 6176 70692
rect 6192 70748 6256 70752
rect 6192 70692 6196 70748
rect 6196 70692 6252 70748
rect 6252 70692 6256 70748
rect 6192 70688 6256 70692
rect 4285 70204 4349 70208
rect 4285 70148 4289 70204
rect 4289 70148 4345 70204
rect 4345 70148 4349 70204
rect 4285 70144 4349 70148
rect 4365 70204 4429 70208
rect 4365 70148 4369 70204
rect 4369 70148 4425 70204
rect 4425 70148 4429 70204
rect 4365 70144 4429 70148
rect 4445 70204 4509 70208
rect 4445 70148 4449 70204
rect 4449 70148 4505 70204
rect 4505 70148 4509 70204
rect 4445 70144 4509 70148
rect 4525 70204 4589 70208
rect 4525 70148 4529 70204
rect 4529 70148 4585 70204
rect 4585 70148 4589 70204
rect 4525 70144 4589 70148
rect 7618 70204 7682 70208
rect 7618 70148 7622 70204
rect 7622 70148 7678 70204
rect 7678 70148 7682 70204
rect 7618 70144 7682 70148
rect 7698 70204 7762 70208
rect 7698 70148 7702 70204
rect 7702 70148 7758 70204
rect 7758 70148 7762 70204
rect 7698 70144 7762 70148
rect 7778 70204 7842 70208
rect 7778 70148 7782 70204
rect 7782 70148 7838 70204
rect 7838 70148 7842 70204
rect 7778 70144 7842 70148
rect 7858 70204 7922 70208
rect 7858 70148 7862 70204
rect 7862 70148 7918 70204
rect 7918 70148 7922 70204
rect 7858 70144 7922 70148
rect 2618 69660 2682 69664
rect 2618 69604 2622 69660
rect 2622 69604 2678 69660
rect 2678 69604 2682 69660
rect 2618 69600 2682 69604
rect 2698 69660 2762 69664
rect 2698 69604 2702 69660
rect 2702 69604 2758 69660
rect 2758 69604 2762 69660
rect 2698 69600 2762 69604
rect 2778 69660 2842 69664
rect 2778 69604 2782 69660
rect 2782 69604 2838 69660
rect 2838 69604 2842 69660
rect 2778 69600 2842 69604
rect 2858 69660 2922 69664
rect 2858 69604 2862 69660
rect 2862 69604 2918 69660
rect 2918 69604 2922 69660
rect 2858 69600 2922 69604
rect 5952 69660 6016 69664
rect 5952 69604 5956 69660
rect 5956 69604 6012 69660
rect 6012 69604 6016 69660
rect 5952 69600 6016 69604
rect 6032 69660 6096 69664
rect 6032 69604 6036 69660
rect 6036 69604 6092 69660
rect 6092 69604 6096 69660
rect 6032 69600 6096 69604
rect 6112 69660 6176 69664
rect 6112 69604 6116 69660
rect 6116 69604 6172 69660
rect 6172 69604 6176 69660
rect 6112 69600 6176 69604
rect 6192 69660 6256 69664
rect 6192 69604 6196 69660
rect 6196 69604 6252 69660
rect 6252 69604 6256 69660
rect 6192 69600 6256 69604
rect 4285 69116 4349 69120
rect 4285 69060 4289 69116
rect 4289 69060 4345 69116
rect 4345 69060 4349 69116
rect 4285 69056 4349 69060
rect 4365 69116 4429 69120
rect 4365 69060 4369 69116
rect 4369 69060 4425 69116
rect 4425 69060 4429 69116
rect 4365 69056 4429 69060
rect 4445 69116 4509 69120
rect 4445 69060 4449 69116
rect 4449 69060 4505 69116
rect 4505 69060 4509 69116
rect 4445 69056 4509 69060
rect 4525 69116 4589 69120
rect 4525 69060 4529 69116
rect 4529 69060 4585 69116
rect 4585 69060 4589 69116
rect 4525 69056 4589 69060
rect 7618 69116 7682 69120
rect 7618 69060 7622 69116
rect 7622 69060 7678 69116
rect 7678 69060 7682 69116
rect 7618 69056 7682 69060
rect 7698 69116 7762 69120
rect 7698 69060 7702 69116
rect 7702 69060 7758 69116
rect 7758 69060 7762 69116
rect 7698 69056 7762 69060
rect 7778 69116 7842 69120
rect 7778 69060 7782 69116
rect 7782 69060 7838 69116
rect 7838 69060 7842 69116
rect 7778 69056 7842 69060
rect 7858 69116 7922 69120
rect 7858 69060 7862 69116
rect 7862 69060 7918 69116
rect 7918 69060 7922 69116
rect 7858 69056 7922 69060
rect 2618 68572 2682 68576
rect 2618 68516 2622 68572
rect 2622 68516 2678 68572
rect 2678 68516 2682 68572
rect 2618 68512 2682 68516
rect 2698 68572 2762 68576
rect 2698 68516 2702 68572
rect 2702 68516 2758 68572
rect 2758 68516 2762 68572
rect 2698 68512 2762 68516
rect 2778 68572 2842 68576
rect 2778 68516 2782 68572
rect 2782 68516 2838 68572
rect 2838 68516 2842 68572
rect 2778 68512 2842 68516
rect 2858 68572 2922 68576
rect 2858 68516 2862 68572
rect 2862 68516 2918 68572
rect 2918 68516 2922 68572
rect 2858 68512 2922 68516
rect 5952 68572 6016 68576
rect 5952 68516 5956 68572
rect 5956 68516 6012 68572
rect 6012 68516 6016 68572
rect 5952 68512 6016 68516
rect 6032 68572 6096 68576
rect 6032 68516 6036 68572
rect 6036 68516 6092 68572
rect 6092 68516 6096 68572
rect 6032 68512 6096 68516
rect 6112 68572 6176 68576
rect 6112 68516 6116 68572
rect 6116 68516 6172 68572
rect 6172 68516 6176 68572
rect 6112 68512 6176 68516
rect 6192 68572 6256 68576
rect 6192 68516 6196 68572
rect 6196 68516 6252 68572
rect 6252 68516 6256 68572
rect 6192 68512 6256 68516
rect 4285 68028 4349 68032
rect 4285 67972 4289 68028
rect 4289 67972 4345 68028
rect 4345 67972 4349 68028
rect 4285 67968 4349 67972
rect 4365 68028 4429 68032
rect 4365 67972 4369 68028
rect 4369 67972 4425 68028
rect 4425 67972 4429 68028
rect 4365 67968 4429 67972
rect 4445 68028 4509 68032
rect 4445 67972 4449 68028
rect 4449 67972 4505 68028
rect 4505 67972 4509 68028
rect 4445 67968 4509 67972
rect 4525 68028 4589 68032
rect 4525 67972 4529 68028
rect 4529 67972 4585 68028
rect 4585 67972 4589 68028
rect 4525 67968 4589 67972
rect 7618 68028 7682 68032
rect 7618 67972 7622 68028
rect 7622 67972 7678 68028
rect 7678 67972 7682 68028
rect 7618 67968 7682 67972
rect 7698 68028 7762 68032
rect 7698 67972 7702 68028
rect 7702 67972 7758 68028
rect 7758 67972 7762 68028
rect 7698 67968 7762 67972
rect 7778 68028 7842 68032
rect 7778 67972 7782 68028
rect 7782 67972 7838 68028
rect 7838 67972 7842 68028
rect 7778 67968 7842 67972
rect 7858 68028 7922 68032
rect 7858 67972 7862 68028
rect 7862 67972 7918 68028
rect 7918 67972 7922 68028
rect 7858 67968 7922 67972
rect 2618 67484 2682 67488
rect 2618 67428 2622 67484
rect 2622 67428 2678 67484
rect 2678 67428 2682 67484
rect 2618 67424 2682 67428
rect 2698 67484 2762 67488
rect 2698 67428 2702 67484
rect 2702 67428 2758 67484
rect 2758 67428 2762 67484
rect 2698 67424 2762 67428
rect 2778 67484 2842 67488
rect 2778 67428 2782 67484
rect 2782 67428 2838 67484
rect 2838 67428 2842 67484
rect 2778 67424 2842 67428
rect 2858 67484 2922 67488
rect 2858 67428 2862 67484
rect 2862 67428 2918 67484
rect 2918 67428 2922 67484
rect 2858 67424 2922 67428
rect 5952 67484 6016 67488
rect 5952 67428 5956 67484
rect 5956 67428 6012 67484
rect 6012 67428 6016 67484
rect 5952 67424 6016 67428
rect 6032 67484 6096 67488
rect 6032 67428 6036 67484
rect 6036 67428 6092 67484
rect 6092 67428 6096 67484
rect 6032 67424 6096 67428
rect 6112 67484 6176 67488
rect 6112 67428 6116 67484
rect 6116 67428 6172 67484
rect 6172 67428 6176 67484
rect 6112 67424 6176 67428
rect 6192 67484 6256 67488
rect 6192 67428 6196 67484
rect 6196 67428 6252 67484
rect 6252 67428 6256 67484
rect 6192 67424 6256 67428
rect 4285 66940 4349 66944
rect 4285 66884 4289 66940
rect 4289 66884 4345 66940
rect 4345 66884 4349 66940
rect 4285 66880 4349 66884
rect 4365 66940 4429 66944
rect 4365 66884 4369 66940
rect 4369 66884 4425 66940
rect 4425 66884 4429 66940
rect 4365 66880 4429 66884
rect 4445 66940 4509 66944
rect 4445 66884 4449 66940
rect 4449 66884 4505 66940
rect 4505 66884 4509 66940
rect 4445 66880 4509 66884
rect 4525 66940 4589 66944
rect 4525 66884 4529 66940
rect 4529 66884 4585 66940
rect 4585 66884 4589 66940
rect 4525 66880 4589 66884
rect 7618 66940 7682 66944
rect 7618 66884 7622 66940
rect 7622 66884 7678 66940
rect 7678 66884 7682 66940
rect 7618 66880 7682 66884
rect 7698 66940 7762 66944
rect 7698 66884 7702 66940
rect 7702 66884 7758 66940
rect 7758 66884 7762 66940
rect 7698 66880 7762 66884
rect 7778 66940 7842 66944
rect 7778 66884 7782 66940
rect 7782 66884 7838 66940
rect 7838 66884 7842 66940
rect 7778 66880 7842 66884
rect 7858 66940 7922 66944
rect 7858 66884 7862 66940
rect 7862 66884 7918 66940
rect 7918 66884 7922 66940
rect 7858 66880 7922 66884
rect 2618 66396 2682 66400
rect 2618 66340 2622 66396
rect 2622 66340 2678 66396
rect 2678 66340 2682 66396
rect 2618 66336 2682 66340
rect 2698 66396 2762 66400
rect 2698 66340 2702 66396
rect 2702 66340 2758 66396
rect 2758 66340 2762 66396
rect 2698 66336 2762 66340
rect 2778 66396 2842 66400
rect 2778 66340 2782 66396
rect 2782 66340 2838 66396
rect 2838 66340 2842 66396
rect 2778 66336 2842 66340
rect 2858 66396 2922 66400
rect 2858 66340 2862 66396
rect 2862 66340 2918 66396
rect 2918 66340 2922 66396
rect 2858 66336 2922 66340
rect 5952 66396 6016 66400
rect 5952 66340 5956 66396
rect 5956 66340 6012 66396
rect 6012 66340 6016 66396
rect 5952 66336 6016 66340
rect 6032 66396 6096 66400
rect 6032 66340 6036 66396
rect 6036 66340 6092 66396
rect 6092 66340 6096 66396
rect 6032 66336 6096 66340
rect 6112 66396 6176 66400
rect 6112 66340 6116 66396
rect 6116 66340 6172 66396
rect 6172 66340 6176 66396
rect 6112 66336 6176 66340
rect 6192 66396 6256 66400
rect 6192 66340 6196 66396
rect 6196 66340 6252 66396
rect 6252 66340 6256 66396
rect 6192 66336 6256 66340
rect 4285 65852 4349 65856
rect 4285 65796 4289 65852
rect 4289 65796 4345 65852
rect 4345 65796 4349 65852
rect 4285 65792 4349 65796
rect 4365 65852 4429 65856
rect 4365 65796 4369 65852
rect 4369 65796 4425 65852
rect 4425 65796 4429 65852
rect 4365 65792 4429 65796
rect 4445 65852 4509 65856
rect 4445 65796 4449 65852
rect 4449 65796 4505 65852
rect 4505 65796 4509 65852
rect 4445 65792 4509 65796
rect 4525 65852 4589 65856
rect 4525 65796 4529 65852
rect 4529 65796 4585 65852
rect 4585 65796 4589 65852
rect 4525 65792 4589 65796
rect 7618 65852 7682 65856
rect 7618 65796 7622 65852
rect 7622 65796 7678 65852
rect 7678 65796 7682 65852
rect 7618 65792 7682 65796
rect 7698 65852 7762 65856
rect 7698 65796 7702 65852
rect 7702 65796 7758 65852
rect 7758 65796 7762 65852
rect 7698 65792 7762 65796
rect 7778 65852 7842 65856
rect 7778 65796 7782 65852
rect 7782 65796 7838 65852
rect 7838 65796 7842 65852
rect 7778 65792 7842 65796
rect 7858 65852 7922 65856
rect 7858 65796 7862 65852
rect 7862 65796 7918 65852
rect 7918 65796 7922 65852
rect 7858 65792 7922 65796
rect 2618 65308 2682 65312
rect 2618 65252 2622 65308
rect 2622 65252 2678 65308
rect 2678 65252 2682 65308
rect 2618 65248 2682 65252
rect 2698 65308 2762 65312
rect 2698 65252 2702 65308
rect 2702 65252 2758 65308
rect 2758 65252 2762 65308
rect 2698 65248 2762 65252
rect 2778 65308 2842 65312
rect 2778 65252 2782 65308
rect 2782 65252 2838 65308
rect 2838 65252 2842 65308
rect 2778 65248 2842 65252
rect 2858 65308 2922 65312
rect 2858 65252 2862 65308
rect 2862 65252 2918 65308
rect 2918 65252 2922 65308
rect 2858 65248 2922 65252
rect 5952 65308 6016 65312
rect 5952 65252 5956 65308
rect 5956 65252 6012 65308
rect 6012 65252 6016 65308
rect 5952 65248 6016 65252
rect 6032 65308 6096 65312
rect 6032 65252 6036 65308
rect 6036 65252 6092 65308
rect 6092 65252 6096 65308
rect 6032 65248 6096 65252
rect 6112 65308 6176 65312
rect 6112 65252 6116 65308
rect 6116 65252 6172 65308
rect 6172 65252 6176 65308
rect 6112 65248 6176 65252
rect 6192 65308 6256 65312
rect 6192 65252 6196 65308
rect 6196 65252 6252 65308
rect 6252 65252 6256 65308
rect 6192 65248 6256 65252
rect 4285 64764 4349 64768
rect 4285 64708 4289 64764
rect 4289 64708 4345 64764
rect 4345 64708 4349 64764
rect 4285 64704 4349 64708
rect 4365 64764 4429 64768
rect 4365 64708 4369 64764
rect 4369 64708 4425 64764
rect 4425 64708 4429 64764
rect 4365 64704 4429 64708
rect 4445 64764 4509 64768
rect 4445 64708 4449 64764
rect 4449 64708 4505 64764
rect 4505 64708 4509 64764
rect 4445 64704 4509 64708
rect 4525 64764 4589 64768
rect 4525 64708 4529 64764
rect 4529 64708 4585 64764
rect 4585 64708 4589 64764
rect 4525 64704 4589 64708
rect 7618 64764 7682 64768
rect 7618 64708 7622 64764
rect 7622 64708 7678 64764
rect 7678 64708 7682 64764
rect 7618 64704 7682 64708
rect 7698 64764 7762 64768
rect 7698 64708 7702 64764
rect 7702 64708 7758 64764
rect 7758 64708 7762 64764
rect 7698 64704 7762 64708
rect 7778 64764 7842 64768
rect 7778 64708 7782 64764
rect 7782 64708 7838 64764
rect 7838 64708 7842 64764
rect 7778 64704 7842 64708
rect 7858 64764 7922 64768
rect 7858 64708 7862 64764
rect 7862 64708 7918 64764
rect 7918 64708 7922 64764
rect 7858 64704 7922 64708
rect 2618 64220 2682 64224
rect 2618 64164 2622 64220
rect 2622 64164 2678 64220
rect 2678 64164 2682 64220
rect 2618 64160 2682 64164
rect 2698 64220 2762 64224
rect 2698 64164 2702 64220
rect 2702 64164 2758 64220
rect 2758 64164 2762 64220
rect 2698 64160 2762 64164
rect 2778 64220 2842 64224
rect 2778 64164 2782 64220
rect 2782 64164 2838 64220
rect 2838 64164 2842 64220
rect 2778 64160 2842 64164
rect 2858 64220 2922 64224
rect 2858 64164 2862 64220
rect 2862 64164 2918 64220
rect 2918 64164 2922 64220
rect 2858 64160 2922 64164
rect 5952 64220 6016 64224
rect 5952 64164 5956 64220
rect 5956 64164 6012 64220
rect 6012 64164 6016 64220
rect 5952 64160 6016 64164
rect 6032 64220 6096 64224
rect 6032 64164 6036 64220
rect 6036 64164 6092 64220
rect 6092 64164 6096 64220
rect 6032 64160 6096 64164
rect 6112 64220 6176 64224
rect 6112 64164 6116 64220
rect 6116 64164 6172 64220
rect 6172 64164 6176 64220
rect 6112 64160 6176 64164
rect 6192 64220 6256 64224
rect 6192 64164 6196 64220
rect 6196 64164 6252 64220
rect 6252 64164 6256 64220
rect 6192 64160 6256 64164
rect 4285 63676 4349 63680
rect 4285 63620 4289 63676
rect 4289 63620 4345 63676
rect 4345 63620 4349 63676
rect 4285 63616 4349 63620
rect 4365 63676 4429 63680
rect 4365 63620 4369 63676
rect 4369 63620 4425 63676
rect 4425 63620 4429 63676
rect 4365 63616 4429 63620
rect 4445 63676 4509 63680
rect 4445 63620 4449 63676
rect 4449 63620 4505 63676
rect 4505 63620 4509 63676
rect 4445 63616 4509 63620
rect 4525 63676 4589 63680
rect 4525 63620 4529 63676
rect 4529 63620 4585 63676
rect 4585 63620 4589 63676
rect 4525 63616 4589 63620
rect 7618 63676 7682 63680
rect 7618 63620 7622 63676
rect 7622 63620 7678 63676
rect 7678 63620 7682 63676
rect 7618 63616 7682 63620
rect 7698 63676 7762 63680
rect 7698 63620 7702 63676
rect 7702 63620 7758 63676
rect 7758 63620 7762 63676
rect 7698 63616 7762 63620
rect 7778 63676 7842 63680
rect 7778 63620 7782 63676
rect 7782 63620 7838 63676
rect 7838 63620 7842 63676
rect 7778 63616 7842 63620
rect 7858 63676 7922 63680
rect 7858 63620 7862 63676
rect 7862 63620 7918 63676
rect 7918 63620 7922 63676
rect 7858 63616 7922 63620
rect 2618 63132 2682 63136
rect 2618 63076 2622 63132
rect 2622 63076 2678 63132
rect 2678 63076 2682 63132
rect 2618 63072 2682 63076
rect 2698 63132 2762 63136
rect 2698 63076 2702 63132
rect 2702 63076 2758 63132
rect 2758 63076 2762 63132
rect 2698 63072 2762 63076
rect 2778 63132 2842 63136
rect 2778 63076 2782 63132
rect 2782 63076 2838 63132
rect 2838 63076 2842 63132
rect 2778 63072 2842 63076
rect 2858 63132 2922 63136
rect 2858 63076 2862 63132
rect 2862 63076 2918 63132
rect 2918 63076 2922 63132
rect 2858 63072 2922 63076
rect 5952 63132 6016 63136
rect 5952 63076 5956 63132
rect 5956 63076 6012 63132
rect 6012 63076 6016 63132
rect 5952 63072 6016 63076
rect 6032 63132 6096 63136
rect 6032 63076 6036 63132
rect 6036 63076 6092 63132
rect 6092 63076 6096 63132
rect 6032 63072 6096 63076
rect 6112 63132 6176 63136
rect 6112 63076 6116 63132
rect 6116 63076 6172 63132
rect 6172 63076 6176 63132
rect 6112 63072 6176 63076
rect 6192 63132 6256 63136
rect 6192 63076 6196 63132
rect 6196 63076 6252 63132
rect 6252 63076 6256 63132
rect 6192 63072 6256 63076
rect 4285 62588 4349 62592
rect 4285 62532 4289 62588
rect 4289 62532 4345 62588
rect 4345 62532 4349 62588
rect 4285 62528 4349 62532
rect 4365 62588 4429 62592
rect 4365 62532 4369 62588
rect 4369 62532 4425 62588
rect 4425 62532 4429 62588
rect 4365 62528 4429 62532
rect 4445 62588 4509 62592
rect 4445 62532 4449 62588
rect 4449 62532 4505 62588
rect 4505 62532 4509 62588
rect 4445 62528 4509 62532
rect 4525 62588 4589 62592
rect 4525 62532 4529 62588
rect 4529 62532 4585 62588
rect 4585 62532 4589 62588
rect 4525 62528 4589 62532
rect 7618 62588 7682 62592
rect 7618 62532 7622 62588
rect 7622 62532 7678 62588
rect 7678 62532 7682 62588
rect 7618 62528 7682 62532
rect 7698 62588 7762 62592
rect 7698 62532 7702 62588
rect 7702 62532 7758 62588
rect 7758 62532 7762 62588
rect 7698 62528 7762 62532
rect 7778 62588 7842 62592
rect 7778 62532 7782 62588
rect 7782 62532 7838 62588
rect 7838 62532 7842 62588
rect 7778 62528 7842 62532
rect 7858 62588 7922 62592
rect 7858 62532 7862 62588
rect 7862 62532 7918 62588
rect 7918 62532 7922 62588
rect 7858 62528 7922 62532
rect 2618 62044 2682 62048
rect 2618 61988 2622 62044
rect 2622 61988 2678 62044
rect 2678 61988 2682 62044
rect 2618 61984 2682 61988
rect 2698 62044 2762 62048
rect 2698 61988 2702 62044
rect 2702 61988 2758 62044
rect 2758 61988 2762 62044
rect 2698 61984 2762 61988
rect 2778 62044 2842 62048
rect 2778 61988 2782 62044
rect 2782 61988 2838 62044
rect 2838 61988 2842 62044
rect 2778 61984 2842 61988
rect 2858 62044 2922 62048
rect 2858 61988 2862 62044
rect 2862 61988 2918 62044
rect 2918 61988 2922 62044
rect 2858 61984 2922 61988
rect 5952 62044 6016 62048
rect 5952 61988 5956 62044
rect 5956 61988 6012 62044
rect 6012 61988 6016 62044
rect 5952 61984 6016 61988
rect 6032 62044 6096 62048
rect 6032 61988 6036 62044
rect 6036 61988 6092 62044
rect 6092 61988 6096 62044
rect 6032 61984 6096 61988
rect 6112 62044 6176 62048
rect 6112 61988 6116 62044
rect 6116 61988 6172 62044
rect 6172 61988 6176 62044
rect 6112 61984 6176 61988
rect 6192 62044 6256 62048
rect 6192 61988 6196 62044
rect 6196 61988 6252 62044
rect 6252 61988 6256 62044
rect 6192 61984 6256 61988
rect 4285 61500 4349 61504
rect 4285 61444 4289 61500
rect 4289 61444 4345 61500
rect 4345 61444 4349 61500
rect 4285 61440 4349 61444
rect 4365 61500 4429 61504
rect 4365 61444 4369 61500
rect 4369 61444 4425 61500
rect 4425 61444 4429 61500
rect 4365 61440 4429 61444
rect 4445 61500 4509 61504
rect 4445 61444 4449 61500
rect 4449 61444 4505 61500
rect 4505 61444 4509 61500
rect 4445 61440 4509 61444
rect 4525 61500 4589 61504
rect 4525 61444 4529 61500
rect 4529 61444 4585 61500
rect 4585 61444 4589 61500
rect 4525 61440 4589 61444
rect 7618 61500 7682 61504
rect 7618 61444 7622 61500
rect 7622 61444 7678 61500
rect 7678 61444 7682 61500
rect 7618 61440 7682 61444
rect 7698 61500 7762 61504
rect 7698 61444 7702 61500
rect 7702 61444 7758 61500
rect 7758 61444 7762 61500
rect 7698 61440 7762 61444
rect 7778 61500 7842 61504
rect 7778 61444 7782 61500
rect 7782 61444 7838 61500
rect 7838 61444 7842 61500
rect 7778 61440 7842 61444
rect 7858 61500 7922 61504
rect 7858 61444 7862 61500
rect 7862 61444 7918 61500
rect 7918 61444 7922 61500
rect 7858 61440 7922 61444
rect 2618 60956 2682 60960
rect 2618 60900 2622 60956
rect 2622 60900 2678 60956
rect 2678 60900 2682 60956
rect 2618 60896 2682 60900
rect 2698 60956 2762 60960
rect 2698 60900 2702 60956
rect 2702 60900 2758 60956
rect 2758 60900 2762 60956
rect 2698 60896 2762 60900
rect 2778 60956 2842 60960
rect 2778 60900 2782 60956
rect 2782 60900 2838 60956
rect 2838 60900 2842 60956
rect 2778 60896 2842 60900
rect 2858 60956 2922 60960
rect 2858 60900 2862 60956
rect 2862 60900 2918 60956
rect 2918 60900 2922 60956
rect 2858 60896 2922 60900
rect 5952 60956 6016 60960
rect 5952 60900 5956 60956
rect 5956 60900 6012 60956
rect 6012 60900 6016 60956
rect 5952 60896 6016 60900
rect 6032 60956 6096 60960
rect 6032 60900 6036 60956
rect 6036 60900 6092 60956
rect 6092 60900 6096 60956
rect 6032 60896 6096 60900
rect 6112 60956 6176 60960
rect 6112 60900 6116 60956
rect 6116 60900 6172 60956
rect 6172 60900 6176 60956
rect 6112 60896 6176 60900
rect 6192 60956 6256 60960
rect 6192 60900 6196 60956
rect 6196 60900 6252 60956
rect 6252 60900 6256 60956
rect 6192 60896 6256 60900
rect 4285 60412 4349 60416
rect 4285 60356 4289 60412
rect 4289 60356 4345 60412
rect 4345 60356 4349 60412
rect 4285 60352 4349 60356
rect 4365 60412 4429 60416
rect 4365 60356 4369 60412
rect 4369 60356 4425 60412
rect 4425 60356 4429 60412
rect 4365 60352 4429 60356
rect 4445 60412 4509 60416
rect 4445 60356 4449 60412
rect 4449 60356 4505 60412
rect 4505 60356 4509 60412
rect 4445 60352 4509 60356
rect 4525 60412 4589 60416
rect 4525 60356 4529 60412
rect 4529 60356 4585 60412
rect 4585 60356 4589 60412
rect 4525 60352 4589 60356
rect 7618 60412 7682 60416
rect 7618 60356 7622 60412
rect 7622 60356 7678 60412
rect 7678 60356 7682 60412
rect 7618 60352 7682 60356
rect 7698 60412 7762 60416
rect 7698 60356 7702 60412
rect 7702 60356 7758 60412
rect 7758 60356 7762 60412
rect 7698 60352 7762 60356
rect 7778 60412 7842 60416
rect 7778 60356 7782 60412
rect 7782 60356 7838 60412
rect 7838 60356 7842 60412
rect 7778 60352 7842 60356
rect 7858 60412 7922 60416
rect 7858 60356 7862 60412
rect 7862 60356 7918 60412
rect 7918 60356 7922 60412
rect 7858 60352 7922 60356
rect 2618 59868 2682 59872
rect 2618 59812 2622 59868
rect 2622 59812 2678 59868
rect 2678 59812 2682 59868
rect 2618 59808 2682 59812
rect 2698 59868 2762 59872
rect 2698 59812 2702 59868
rect 2702 59812 2758 59868
rect 2758 59812 2762 59868
rect 2698 59808 2762 59812
rect 2778 59868 2842 59872
rect 2778 59812 2782 59868
rect 2782 59812 2838 59868
rect 2838 59812 2842 59868
rect 2778 59808 2842 59812
rect 2858 59868 2922 59872
rect 2858 59812 2862 59868
rect 2862 59812 2918 59868
rect 2918 59812 2922 59868
rect 2858 59808 2922 59812
rect 5952 59868 6016 59872
rect 5952 59812 5956 59868
rect 5956 59812 6012 59868
rect 6012 59812 6016 59868
rect 5952 59808 6016 59812
rect 6032 59868 6096 59872
rect 6032 59812 6036 59868
rect 6036 59812 6092 59868
rect 6092 59812 6096 59868
rect 6032 59808 6096 59812
rect 6112 59868 6176 59872
rect 6112 59812 6116 59868
rect 6116 59812 6172 59868
rect 6172 59812 6176 59868
rect 6112 59808 6176 59812
rect 6192 59868 6256 59872
rect 6192 59812 6196 59868
rect 6196 59812 6252 59868
rect 6252 59812 6256 59868
rect 6192 59808 6256 59812
rect 4285 59324 4349 59328
rect 4285 59268 4289 59324
rect 4289 59268 4345 59324
rect 4345 59268 4349 59324
rect 4285 59264 4349 59268
rect 4365 59324 4429 59328
rect 4365 59268 4369 59324
rect 4369 59268 4425 59324
rect 4425 59268 4429 59324
rect 4365 59264 4429 59268
rect 4445 59324 4509 59328
rect 4445 59268 4449 59324
rect 4449 59268 4505 59324
rect 4505 59268 4509 59324
rect 4445 59264 4509 59268
rect 4525 59324 4589 59328
rect 4525 59268 4529 59324
rect 4529 59268 4585 59324
rect 4585 59268 4589 59324
rect 4525 59264 4589 59268
rect 7618 59324 7682 59328
rect 7618 59268 7622 59324
rect 7622 59268 7678 59324
rect 7678 59268 7682 59324
rect 7618 59264 7682 59268
rect 7698 59324 7762 59328
rect 7698 59268 7702 59324
rect 7702 59268 7758 59324
rect 7758 59268 7762 59324
rect 7698 59264 7762 59268
rect 7778 59324 7842 59328
rect 7778 59268 7782 59324
rect 7782 59268 7838 59324
rect 7838 59268 7842 59324
rect 7778 59264 7842 59268
rect 7858 59324 7922 59328
rect 7858 59268 7862 59324
rect 7862 59268 7918 59324
rect 7918 59268 7922 59324
rect 7858 59264 7922 59268
rect 2618 58780 2682 58784
rect 2618 58724 2622 58780
rect 2622 58724 2678 58780
rect 2678 58724 2682 58780
rect 2618 58720 2682 58724
rect 2698 58780 2762 58784
rect 2698 58724 2702 58780
rect 2702 58724 2758 58780
rect 2758 58724 2762 58780
rect 2698 58720 2762 58724
rect 2778 58780 2842 58784
rect 2778 58724 2782 58780
rect 2782 58724 2838 58780
rect 2838 58724 2842 58780
rect 2778 58720 2842 58724
rect 2858 58780 2922 58784
rect 2858 58724 2862 58780
rect 2862 58724 2918 58780
rect 2918 58724 2922 58780
rect 2858 58720 2922 58724
rect 5952 58780 6016 58784
rect 5952 58724 5956 58780
rect 5956 58724 6012 58780
rect 6012 58724 6016 58780
rect 5952 58720 6016 58724
rect 6032 58780 6096 58784
rect 6032 58724 6036 58780
rect 6036 58724 6092 58780
rect 6092 58724 6096 58780
rect 6032 58720 6096 58724
rect 6112 58780 6176 58784
rect 6112 58724 6116 58780
rect 6116 58724 6172 58780
rect 6172 58724 6176 58780
rect 6112 58720 6176 58724
rect 6192 58780 6256 58784
rect 6192 58724 6196 58780
rect 6196 58724 6252 58780
rect 6252 58724 6256 58780
rect 6192 58720 6256 58724
rect 4285 58236 4349 58240
rect 4285 58180 4289 58236
rect 4289 58180 4345 58236
rect 4345 58180 4349 58236
rect 4285 58176 4349 58180
rect 4365 58236 4429 58240
rect 4365 58180 4369 58236
rect 4369 58180 4425 58236
rect 4425 58180 4429 58236
rect 4365 58176 4429 58180
rect 4445 58236 4509 58240
rect 4445 58180 4449 58236
rect 4449 58180 4505 58236
rect 4505 58180 4509 58236
rect 4445 58176 4509 58180
rect 4525 58236 4589 58240
rect 4525 58180 4529 58236
rect 4529 58180 4585 58236
rect 4585 58180 4589 58236
rect 4525 58176 4589 58180
rect 7618 58236 7682 58240
rect 7618 58180 7622 58236
rect 7622 58180 7678 58236
rect 7678 58180 7682 58236
rect 7618 58176 7682 58180
rect 7698 58236 7762 58240
rect 7698 58180 7702 58236
rect 7702 58180 7758 58236
rect 7758 58180 7762 58236
rect 7698 58176 7762 58180
rect 7778 58236 7842 58240
rect 7778 58180 7782 58236
rect 7782 58180 7838 58236
rect 7838 58180 7842 58236
rect 7778 58176 7842 58180
rect 7858 58236 7922 58240
rect 7858 58180 7862 58236
rect 7862 58180 7918 58236
rect 7918 58180 7922 58236
rect 7858 58176 7922 58180
rect 2618 57692 2682 57696
rect 2618 57636 2622 57692
rect 2622 57636 2678 57692
rect 2678 57636 2682 57692
rect 2618 57632 2682 57636
rect 2698 57692 2762 57696
rect 2698 57636 2702 57692
rect 2702 57636 2758 57692
rect 2758 57636 2762 57692
rect 2698 57632 2762 57636
rect 2778 57692 2842 57696
rect 2778 57636 2782 57692
rect 2782 57636 2838 57692
rect 2838 57636 2842 57692
rect 2778 57632 2842 57636
rect 2858 57692 2922 57696
rect 2858 57636 2862 57692
rect 2862 57636 2918 57692
rect 2918 57636 2922 57692
rect 2858 57632 2922 57636
rect 5952 57692 6016 57696
rect 5952 57636 5956 57692
rect 5956 57636 6012 57692
rect 6012 57636 6016 57692
rect 5952 57632 6016 57636
rect 6032 57692 6096 57696
rect 6032 57636 6036 57692
rect 6036 57636 6092 57692
rect 6092 57636 6096 57692
rect 6032 57632 6096 57636
rect 6112 57692 6176 57696
rect 6112 57636 6116 57692
rect 6116 57636 6172 57692
rect 6172 57636 6176 57692
rect 6112 57632 6176 57636
rect 6192 57692 6256 57696
rect 6192 57636 6196 57692
rect 6196 57636 6252 57692
rect 6252 57636 6256 57692
rect 6192 57632 6256 57636
rect 4285 57148 4349 57152
rect 4285 57092 4289 57148
rect 4289 57092 4345 57148
rect 4345 57092 4349 57148
rect 4285 57088 4349 57092
rect 4365 57148 4429 57152
rect 4365 57092 4369 57148
rect 4369 57092 4425 57148
rect 4425 57092 4429 57148
rect 4365 57088 4429 57092
rect 4445 57148 4509 57152
rect 4445 57092 4449 57148
rect 4449 57092 4505 57148
rect 4505 57092 4509 57148
rect 4445 57088 4509 57092
rect 4525 57148 4589 57152
rect 4525 57092 4529 57148
rect 4529 57092 4585 57148
rect 4585 57092 4589 57148
rect 4525 57088 4589 57092
rect 7618 57148 7682 57152
rect 7618 57092 7622 57148
rect 7622 57092 7678 57148
rect 7678 57092 7682 57148
rect 7618 57088 7682 57092
rect 7698 57148 7762 57152
rect 7698 57092 7702 57148
rect 7702 57092 7758 57148
rect 7758 57092 7762 57148
rect 7698 57088 7762 57092
rect 7778 57148 7842 57152
rect 7778 57092 7782 57148
rect 7782 57092 7838 57148
rect 7838 57092 7842 57148
rect 7778 57088 7842 57092
rect 7858 57148 7922 57152
rect 7858 57092 7862 57148
rect 7862 57092 7918 57148
rect 7918 57092 7922 57148
rect 7858 57088 7922 57092
rect 2618 56604 2682 56608
rect 2618 56548 2622 56604
rect 2622 56548 2678 56604
rect 2678 56548 2682 56604
rect 2618 56544 2682 56548
rect 2698 56604 2762 56608
rect 2698 56548 2702 56604
rect 2702 56548 2758 56604
rect 2758 56548 2762 56604
rect 2698 56544 2762 56548
rect 2778 56604 2842 56608
rect 2778 56548 2782 56604
rect 2782 56548 2838 56604
rect 2838 56548 2842 56604
rect 2778 56544 2842 56548
rect 2858 56604 2922 56608
rect 2858 56548 2862 56604
rect 2862 56548 2918 56604
rect 2918 56548 2922 56604
rect 2858 56544 2922 56548
rect 5952 56604 6016 56608
rect 5952 56548 5956 56604
rect 5956 56548 6012 56604
rect 6012 56548 6016 56604
rect 5952 56544 6016 56548
rect 6032 56604 6096 56608
rect 6032 56548 6036 56604
rect 6036 56548 6092 56604
rect 6092 56548 6096 56604
rect 6032 56544 6096 56548
rect 6112 56604 6176 56608
rect 6112 56548 6116 56604
rect 6116 56548 6172 56604
rect 6172 56548 6176 56604
rect 6112 56544 6176 56548
rect 6192 56604 6256 56608
rect 6192 56548 6196 56604
rect 6196 56548 6252 56604
rect 6252 56548 6256 56604
rect 6192 56544 6256 56548
rect 4285 56060 4349 56064
rect 4285 56004 4289 56060
rect 4289 56004 4345 56060
rect 4345 56004 4349 56060
rect 4285 56000 4349 56004
rect 4365 56060 4429 56064
rect 4365 56004 4369 56060
rect 4369 56004 4425 56060
rect 4425 56004 4429 56060
rect 4365 56000 4429 56004
rect 4445 56060 4509 56064
rect 4445 56004 4449 56060
rect 4449 56004 4505 56060
rect 4505 56004 4509 56060
rect 4445 56000 4509 56004
rect 4525 56060 4589 56064
rect 4525 56004 4529 56060
rect 4529 56004 4585 56060
rect 4585 56004 4589 56060
rect 4525 56000 4589 56004
rect 7618 56060 7682 56064
rect 7618 56004 7622 56060
rect 7622 56004 7678 56060
rect 7678 56004 7682 56060
rect 7618 56000 7682 56004
rect 7698 56060 7762 56064
rect 7698 56004 7702 56060
rect 7702 56004 7758 56060
rect 7758 56004 7762 56060
rect 7698 56000 7762 56004
rect 7778 56060 7842 56064
rect 7778 56004 7782 56060
rect 7782 56004 7838 56060
rect 7838 56004 7842 56060
rect 7778 56000 7842 56004
rect 7858 56060 7922 56064
rect 7858 56004 7862 56060
rect 7862 56004 7918 56060
rect 7918 56004 7922 56060
rect 7858 56000 7922 56004
rect 2618 55516 2682 55520
rect 2618 55460 2622 55516
rect 2622 55460 2678 55516
rect 2678 55460 2682 55516
rect 2618 55456 2682 55460
rect 2698 55516 2762 55520
rect 2698 55460 2702 55516
rect 2702 55460 2758 55516
rect 2758 55460 2762 55516
rect 2698 55456 2762 55460
rect 2778 55516 2842 55520
rect 2778 55460 2782 55516
rect 2782 55460 2838 55516
rect 2838 55460 2842 55516
rect 2778 55456 2842 55460
rect 2858 55516 2922 55520
rect 2858 55460 2862 55516
rect 2862 55460 2918 55516
rect 2918 55460 2922 55516
rect 2858 55456 2922 55460
rect 5952 55516 6016 55520
rect 5952 55460 5956 55516
rect 5956 55460 6012 55516
rect 6012 55460 6016 55516
rect 5952 55456 6016 55460
rect 6032 55516 6096 55520
rect 6032 55460 6036 55516
rect 6036 55460 6092 55516
rect 6092 55460 6096 55516
rect 6032 55456 6096 55460
rect 6112 55516 6176 55520
rect 6112 55460 6116 55516
rect 6116 55460 6172 55516
rect 6172 55460 6176 55516
rect 6112 55456 6176 55460
rect 6192 55516 6256 55520
rect 6192 55460 6196 55516
rect 6196 55460 6252 55516
rect 6252 55460 6256 55516
rect 6192 55456 6256 55460
rect 4285 54972 4349 54976
rect 4285 54916 4289 54972
rect 4289 54916 4345 54972
rect 4345 54916 4349 54972
rect 4285 54912 4349 54916
rect 4365 54972 4429 54976
rect 4365 54916 4369 54972
rect 4369 54916 4425 54972
rect 4425 54916 4429 54972
rect 4365 54912 4429 54916
rect 4445 54972 4509 54976
rect 4445 54916 4449 54972
rect 4449 54916 4505 54972
rect 4505 54916 4509 54972
rect 4445 54912 4509 54916
rect 4525 54972 4589 54976
rect 4525 54916 4529 54972
rect 4529 54916 4585 54972
rect 4585 54916 4589 54972
rect 4525 54912 4589 54916
rect 7618 54972 7682 54976
rect 7618 54916 7622 54972
rect 7622 54916 7678 54972
rect 7678 54916 7682 54972
rect 7618 54912 7682 54916
rect 7698 54972 7762 54976
rect 7698 54916 7702 54972
rect 7702 54916 7758 54972
rect 7758 54916 7762 54972
rect 7698 54912 7762 54916
rect 7778 54972 7842 54976
rect 7778 54916 7782 54972
rect 7782 54916 7838 54972
rect 7838 54916 7842 54972
rect 7778 54912 7842 54916
rect 7858 54972 7922 54976
rect 7858 54916 7862 54972
rect 7862 54916 7918 54972
rect 7918 54916 7922 54972
rect 7858 54912 7922 54916
rect 2618 54428 2682 54432
rect 2618 54372 2622 54428
rect 2622 54372 2678 54428
rect 2678 54372 2682 54428
rect 2618 54368 2682 54372
rect 2698 54428 2762 54432
rect 2698 54372 2702 54428
rect 2702 54372 2758 54428
rect 2758 54372 2762 54428
rect 2698 54368 2762 54372
rect 2778 54428 2842 54432
rect 2778 54372 2782 54428
rect 2782 54372 2838 54428
rect 2838 54372 2842 54428
rect 2778 54368 2842 54372
rect 2858 54428 2922 54432
rect 2858 54372 2862 54428
rect 2862 54372 2918 54428
rect 2918 54372 2922 54428
rect 2858 54368 2922 54372
rect 5952 54428 6016 54432
rect 5952 54372 5956 54428
rect 5956 54372 6012 54428
rect 6012 54372 6016 54428
rect 5952 54368 6016 54372
rect 6032 54428 6096 54432
rect 6032 54372 6036 54428
rect 6036 54372 6092 54428
rect 6092 54372 6096 54428
rect 6032 54368 6096 54372
rect 6112 54428 6176 54432
rect 6112 54372 6116 54428
rect 6116 54372 6172 54428
rect 6172 54372 6176 54428
rect 6112 54368 6176 54372
rect 6192 54428 6256 54432
rect 6192 54372 6196 54428
rect 6196 54372 6252 54428
rect 6252 54372 6256 54428
rect 6192 54368 6256 54372
rect 4285 53884 4349 53888
rect 4285 53828 4289 53884
rect 4289 53828 4345 53884
rect 4345 53828 4349 53884
rect 4285 53824 4349 53828
rect 4365 53884 4429 53888
rect 4365 53828 4369 53884
rect 4369 53828 4425 53884
rect 4425 53828 4429 53884
rect 4365 53824 4429 53828
rect 4445 53884 4509 53888
rect 4445 53828 4449 53884
rect 4449 53828 4505 53884
rect 4505 53828 4509 53884
rect 4445 53824 4509 53828
rect 4525 53884 4589 53888
rect 4525 53828 4529 53884
rect 4529 53828 4585 53884
rect 4585 53828 4589 53884
rect 4525 53824 4589 53828
rect 7618 53884 7682 53888
rect 7618 53828 7622 53884
rect 7622 53828 7678 53884
rect 7678 53828 7682 53884
rect 7618 53824 7682 53828
rect 7698 53884 7762 53888
rect 7698 53828 7702 53884
rect 7702 53828 7758 53884
rect 7758 53828 7762 53884
rect 7698 53824 7762 53828
rect 7778 53884 7842 53888
rect 7778 53828 7782 53884
rect 7782 53828 7838 53884
rect 7838 53828 7842 53884
rect 7778 53824 7842 53828
rect 7858 53884 7922 53888
rect 7858 53828 7862 53884
rect 7862 53828 7918 53884
rect 7918 53828 7922 53884
rect 7858 53824 7922 53828
rect 2618 53340 2682 53344
rect 2618 53284 2622 53340
rect 2622 53284 2678 53340
rect 2678 53284 2682 53340
rect 2618 53280 2682 53284
rect 2698 53340 2762 53344
rect 2698 53284 2702 53340
rect 2702 53284 2758 53340
rect 2758 53284 2762 53340
rect 2698 53280 2762 53284
rect 2778 53340 2842 53344
rect 2778 53284 2782 53340
rect 2782 53284 2838 53340
rect 2838 53284 2842 53340
rect 2778 53280 2842 53284
rect 2858 53340 2922 53344
rect 2858 53284 2862 53340
rect 2862 53284 2918 53340
rect 2918 53284 2922 53340
rect 2858 53280 2922 53284
rect 5952 53340 6016 53344
rect 5952 53284 5956 53340
rect 5956 53284 6012 53340
rect 6012 53284 6016 53340
rect 5952 53280 6016 53284
rect 6032 53340 6096 53344
rect 6032 53284 6036 53340
rect 6036 53284 6092 53340
rect 6092 53284 6096 53340
rect 6032 53280 6096 53284
rect 6112 53340 6176 53344
rect 6112 53284 6116 53340
rect 6116 53284 6172 53340
rect 6172 53284 6176 53340
rect 6112 53280 6176 53284
rect 6192 53340 6256 53344
rect 6192 53284 6196 53340
rect 6196 53284 6252 53340
rect 6252 53284 6256 53340
rect 6192 53280 6256 53284
rect 4285 52796 4349 52800
rect 4285 52740 4289 52796
rect 4289 52740 4345 52796
rect 4345 52740 4349 52796
rect 4285 52736 4349 52740
rect 4365 52796 4429 52800
rect 4365 52740 4369 52796
rect 4369 52740 4425 52796
rect 4425 52740 4429 52796
rect 4365 52736 4429 52740
rect 4445 52796 4509 52800
rect 4445 52740 4449 52796
rect 4449 52740 4505 52796
rect 4505 52740 4509 52796
rect 4445 52736 4509 52740
rect 4525 52796 4589 52800
rect 4525 52740 4529 52796
rect 4529 52740 4585 52796
rect 4585 52740 4589 52796
rect 4525 52736 4589 52740
rect 7618 52796 7682 52800
rect 7618 52740 7622 52796
rect 7622 52740 7678 52796
rect 7678 52740 7682 52796
rect 7618 52736 7682 52740
rect 7698 52796 7762 52800
rect 7698 52740 7702 52796
rect 7702 52740 7758 52796
rect 7758 52740 7762 52796
rect 7698 52736 7762 52740
rect 7778 52796 7842 52800
rect 7778 52740 7782 52796
rect 7782 52740 7838 52796
rect 7838 52740 7842 52796
rect 7778 52736 7842 52740
rect 7858 52796 7922 52800
rect 7858 52740 7862 52796
rect 7862 52740 7918 52796
rect 7918 52740 7922 52796
rect 7858 52736 7922 52740
rect 2618 52252 2682 52256
rect 2618 52196 2622 52252
rect 2622 52196 2678 52252
rect 2678 52196 2682 52252
rect 2618 52192 2682 52196
rect 2698 52252 2762 52256
rect 2698 52196 2702 52252
rect 2702 52196 2758 52252
rect 2758 52196 2762 52252
rect 2698 52192 2762 52196
rect 2778 52252 2842 52256
rect 2778 52196 2782 52252
rect 2782 52196 2838 52252
rect 2838 52196 2842 52252
rect 2778 52192 2842 52196
rect 2858 52252 2922 52256
rect 2858 52196 2862 52252
rect 2862 52196 2918 52252
rect 2918 52196 2922 52252
rect 2858 52192 2922 52196
rect 5952 52252 6016 52256
rect 5952 52196 5956 52252
rect 5956 52196 6012 52252
rect 6012 52196 6016 52252
rect 5952 52192 6016 52196
rect 6032 52252 6096 52256
rect 6032 52196 6036 52252
rect 6036 52196 6092 52252
rect 6092 52196 6096 52252
rect 6032 52192 6096 52196
rect 6112 52252 6176 52256
rect 6112 52196 6116 52252
rect 6116 52196 6172 52252
rect 6172 52196 6176 52252
rect 6112 52192 6176 52196
rect 6192 52252 6256 52256
rect 6192 52196 6196 52252
rect 6196 52196 6252 52252
rect 6252 52196 6256 52252
rect 6192 52192 6256 52196
rect 4285 51708 4349 51712
rect 4285 51652 4289 51708
rect 4289 51652 4345 51708
rect 4345 51652 4349 51708
rect 4285 51648 4349 51652
rect 4365 51708 4429 51712
rect 4365 51652 4369 51708
rect 4369 51652 4425 51708
rect 4425 51652 4429 51708
rect 4365 51648 4429 51652
rect 4445 51708 4509 51712
rect 4445 51652 4449 51708
rect 4449 51652 4505 51708
rect 4505 51652 4509 51708
rect 4445 51648 4509 51652
rect 4525 51708 4589 51712
rect 4525 51652 4529 51708
rect 4529 51652 4585 51708
rect 4585 51652 4589 51708
rect 4525 51648 4589 51652
rect 7618 51708 7682 51712
rect 7618 51652 7622 51708
rect 7622 51652 7678 51708
rect 7678 51652 7682 51708
rect 7618 51648 7682 51652
rect 7698 51708 7762 51712
rect 7698 51652 7702 51708
rect 7702 51652 7758 51708
rect 7758 51652 7762 51708
rect 7698 51648 7762 51652
rect 7778 51708 7842 51712
rect 7778 51652 7782 51708
rect 7782 51652 7838 51708
rect 7838 51652 7842 51708
rect 7778 51648 7842 51652
rect 7858 51708 7922 51712
rect 7858 51652 7862 51708
rect 7862 51652 7918 51708
rect 7918 51652 7922 51708
rect 7858 51648 7922 51652
rect 2618 51164 2682 51168
rect 2618 51108 2622 51164
rect 2622 51108 2678 51164
rect 2678 51108 2682 51164
rect 2618 51104 2682 51108
rect 2698 51164 2762 51168
rect 2698 51108 2702 51164
rect 2702 51108 2758 51164
rect 2758 51108 2762 51164
rect 2698 51104 2762 51108
rect 2778 51164 2842 51168
rect 2778 51108 2782 51164
rect 2782 51108 2838 51164
rect 2838 51108 2842 51164
rect 2778 51104 2842 51108
rect 2858 51164 2922 51168
rect 2858 51108 2862 51164
rect 2862 51108 2918 51164
rect 2918 51108 2922 51164
rect 2858 51104 2922 51108
rect 5952 51164 6016 51168
rect 5952 51108 5956 51164
rect 5956 51108 6012 51164
rect 6012 51108 6016 51164
rect 5952 51104 6016 51108
rect 6032 51164 6096 51168
rect 6032 51108 6036 51164
rect 6036 51108 6092 51164
rect 6092 51108 6096 51164
rect 6032 51104 6096 51108
rect 6112 51164 6176 51168
rect 6112 51108 6116 51164
rect 6116 51108 6172 51164
rect 6172 51108 6176 51164
rect 6112 51104 6176 51108
rect 6192 51164 6256 51168
rect 6192 51108 6196 51164
rect 6196 51108 6252 51164
rect 6252 51108 6256 51164
rect 6192 51104 6256 51108
rect 4285 50620 4349 50624
rect 4285 50564 4289 50620
rect 4289 50564 4345 50620
rect 4345 50564 4349 50620
rect 4285 50560 4349 50564
rect 4365 50620 4429 50624
rect 4365 50564 4369 50620
rect 4369 50564 4425 50620
rect 4425 50564 4429 50620
rect 4365 50560 4429 50564
rect 4445 50620 4509 50624
rect 4445 50564 4449 50620
rect 4449 50564 4505 50620
rect 4505 50564 4509 50620
rect 4445 50560 4509 50564
rect 4525 50620 4589 50624
rect 4525 50564 4529 50620
rect 4529 50564 4585 50620
rect 4585 50564 4589 50620
rect 4525 50560 4589 50564
rect 7618 50620 7682 50624
rect 7618 50564 7622 50620
rect 7622 50564 7678 50620
rect 7678 50564 7682 50620
rect 7618 50560 7682 50564
rect 7698 50620 7762 50624
rect 7698 50564 7702 50620
rect 7702 50564 7758 50620
rect 7758 50564 7762 50620
rect 7698 50560 7762 50564
rect 7778 50620 7842 50624
rect 7778 50564 7782 50620
rect 7782 50564 7838 50620
rect 7838 50564 7842 50620
rect 7778 50560 7842 50564
rect 7858 50620 7922 50624
rect 7858 50564 7862 50620
rect 7862 50564 7918 50620
rect 7918 50564 7922 50620
rect 7858 50560 7922 50564
rect 2618 50076 2682 50080
rect 2618 50020 2622 50076
rect 2622 50020 2678 50076
rect 2678 50020 2682 50076
rect 2618 50016 2682 50020
rect 2698 50076 2762 50080
rect 2698 50020 2702 50076
rect 2702 50020 2758 50076
rect 2758 50020 2762 50076
rect 2698 50016 2762 50020
rect 2778 50076 2842 50080
rect 2778 50020 2782 50076
rect 2782 50020 2838 50076
rect 2838 50020 2842 50076
rect 2778 50016 2842 50020
rect 2858 50076 2922 50080
rect 2858 50020 2862 50076
rect 2862 50020 2918 50076
rect 2918 50020 2922 50076
rect 2858 50016 2922 50020
rect 5952 50076 6016 50080
rect 5952 50020 5956 50076
rect 5956 50020 6012 50076
rect 6012 50020 6016 50076
rect 5952 50016 6016 50020
rect 6032 50076 6096 50080
rect 6032 50020 6036 50076
rect 6036 50020 6092 50076
rect 6092 50020 6096 50076
rect 6032 50016 6096 50020
rect 6112 50076 6176 50080
rect 6112 50020 6116 50076
rect 6116 50020 6172 50076
rect 6172 50020 6176 50076
rect 6112 50016 6176 50020
rect 6192 50076 6256 50080
rect 6192 50020 6196 50076
rect 6196 50020 6252 50076
rect 6252 50020 6256 50076
rect 6192 50016 6256 50020
rect 4285 49532 4349 49536
rect 4285 49476 4289 49532
rect 4289 49476 4345 49532
rect 4345 49476 4349 49532
rect 4285 49472 4349 49476
rect 4365 49532 4429 49536
rect 4365 49476 4369 49532
rect 4369 49476 4425 49532
rect 4425 49476 4429 49532
rect 4365 49472 4429 49476
rect 4445 49532 4509 49536
rect 4445 49476 4449 49532
rect 4449 49476 4505 49532
rect 4505 49476 4509 49532
rect 4445 49472 4509 49476
rect 4525 49532 4589 49536
rect 4525 49476 4529 49532
rect 4529 49476 4585 49532
rect 4585 49476 4589 49532
rect 4525 49472 4589 49476
rect 7618 49532 7682 49536
rect 7618 49476 7622 49532
rect 7622 49476 7678 49532
rect 7678 49476 7682 49532
rect 7618 49472 7682 49476
rect 7698 49532 7762 49536
rect 7698 49476 7702 49532
rect 7702 49476 7758 49532
rect 7758 49476 7762 49532
rect 7698 49472 7762 49476
rect 7778 49532 7842 49536
rect 7778 49476 7782 49532
rect 7782 49476 7838 49532
rect 7838 49476 7842 49532
rect 7778 49472 7842 49476
rect 7858 49532 7922 49536
rect 7858 49476 7862 49532
rect 7862 49476 7918 49532
rect 7918 49476 7922 49532
rect 7858 49472 7922 49476
rect 2618 48988 2682 48992
rect 2618 48932 2622 48988
rect 2622 48932 2678 48988
rect 2678 48932 2682 48988
rect 2618 48928 2682 48932
rect 2698 48988 2762 48992
rect 2698 48932 2702 48988
rect 2702 48932 2758 48988
rect 2758 48932 2762 48988
rect 2698 48928 2762 48932
rect 2778 48988 2842 48992
rect 2778 48932 2782 48988
rect 2782 48932 2838 48988
rect 2838 48932 2842 48988
rect 2778 48928 2842 48932
rect 2858 48988 2922 48992
rect 2858 48932 2862 48988
rect 2862 48932 2918 48988
rect 2918 48932 2922 48988
rect 2858 48928 2922 48932
rect 5952 48988 6016 48992
rect 5952 48932 5956 48988
rect 5956 48932 6012 48988
rect 6012 48932 6016 48988
rect 5952 48928 6016 48932
rect 6032 48988 6096 48992
rect 6032 48932 6036 48988
rect 6036 48932 6092 48988
rect 6092 48932 6096 48988
rect 6032 48928 6096 48932
rect 6112 48988 6176 48992
rect 6112 48932 6116 48988
rect 6116 48932 6172 48988
rect 6172 48932 6176 48988
rect 6112 48928 6176 48932
rect 6192 48988 6256 48992
rect 6192 48932 6196 48988
rect 6196 48932 6252 48988
rect 6252 48932 6256 48988
rect 6192 48928 6256 48932
rect 4285 48444 4349 48448
rect 4285 48388 4289 48444
rect 4289 48388 4345 48444
rect 4345 48388 4349 48444
rect 4285 48384 4349 48388
rect 4365 48444 4429 48448
rect 4365 48388 4369 48444
rect 4369 48388 4425 48444
rect 4425 48388 4429 48444
rect 4365 48384 4429 48388
rect 4445 48444 4509 48448
rect 4445 48388 4449 48444
rect 4449 48388 4505 48444
rect 4505 48388 4509 48444
rect 4445 48384 4509 48388
rect 4525 48444 4589 48448
rect 4525 48388 4529 48444
rect 4529 48388 4585 48444
rect 4585 48388 4589 48444
rect 4525 48384 4589 48388
rect 7618 48444 7682 48448
rect 7618 48388 7622 48444
rect 7622 48388 7678 48444
rect 7678 48388 7682 48444
rect 7618 48384 7682 48388
rect 7698 48444 7762 48448
rect 7698 48388 7702 48444
rect 7702 48388 7758 48444
rect 7758 48388 7762 48444
rect 7698 48384 7762 48388
rect 7778 48444 7842 48448
rect 7778 48388 7782 48444
rect 7782 48388 7838 48444
rect 7838 48388 7842 48444
rect 7778 48384 7842 48388
rect 7858 48444 7922 48448
rect 7858 48388 7862 48444
rect 7862 48388 7918 48444
rect 7918 48388 7922 48444
rect 7858 48384 7922 48388
rect 2618 47900 2682 47904
rect 2618 47844 2622 47900
rect 2622 47844 2678 47900
rect 2678 47844 2682 47900
rect 2618 47840 2682 47844
rect 2698 47900 2762 47904
rect 2698 47844 2702 47900
rect 2702 47844 2758 47900
rect 2758 47844 2762 47900
rect 2698 47840 2762 47844
rect 2778 47900 2842 47904
rect 2778 47844 2782 47900
rect 2782 47844 2838 47900
rect 2838 47844 2842 47900
rect 2778 47840 2842 47844
rect 2858 47900 2922 47904
rect 2858 47844 2862 47900
rect 2862 47844 2918 47900
rect 2918 47844 2922 47900
rect 2858 47840 2922 47844
rect 5952 47900 6016 47904
rect 5952 47844 5956 47900
rect 5956 47844 6012 47900
rect 6012 47844 6016 47900
rect 5952 47840 6016 47844
rect 6032 47900 6096 47904
rect 6032 47844 6036 47900
rect 6036 47844 6092 47900
rect 6092 47844 6096 47900
rect 6032 47840 6096 47844
rect 6112 47900 6176 47904
rect 6112 47844 6116 47900
rect 6116 47844 6172 47900
rect 6172 47844 6176 47900
rect 6112 47840 6176 47844
rect 6192 47900 6256 47904
rect 6192 47844 6196 47900
rect 6196 47844 6252 47900
rect 6252 47844 6256 47900
rect 6192 47840 6256 47844
rect 4285 47356 4349 47360
rect 4285 47300 4289 47356
rect 4289 47300 4345 47356
rect 4345 47300 4349 47356
rect 4285 47296 4349 47300
rect 4365 47356 4429 47360
rect 4365 47300 4369 47356
rect 4369 47300 4425 47356
rect 4425 47300 4429 47356
rect 4365 47296 4429 47300
rect 4445 47356 4509 47360
rect 4445 47300 4449 47356
rect 4449 47300 4505 47356
rect 4505 47300 4509 47356
rect 4445 47296 4509 47300
rect 4525 47356 4589 47360
rect 4525 47300 4529 47356
rect 4529 47300 4585 47356
rect 4585 47300 4589 47356
rect 4525 47296 4589 47300
rect 7618 47356 7682 47360
rect 7618 47300 7622 47356
rect 7622 47300 7678 47356
rect 7678 47300 7682 47356
rect 7618 47296 7682 47300
rect 7698 47356 7762 47360
rect 7698 47300 7702 47356
rect 7702 47300 7758 47356
rect 7758 47300 7762 47356
rect 7698 47296 7762 47300
rect 7778 47356 7842 47360
rect 7778 47300 7782 47356
rect 7782 47300 7838 47356
rect 7838 47300 7842 47356
rect 7778 47296 7842 47300
rect 7858 47356 7922 47360
rect 7858 47300 7862 47356
rect 7862 47300 7918 47356
rect 7918 47300 7922 47356
rect 7858 47296 7922 47300
rect 2618 46812 2682 46816
rect 2618 46756 2622 46812
rect 2622 46756 2678 46812
rect 2678 46756 2682 46812
rect 2618 46752 2682 46756
rect 2698 46812 2762 46816
rect 2698 46756 2702 46812
rect 2702 46756 2758 46812
rect 2758 46756 2762 46812
rect 2698 46752 2762 46756
rect 2778 46812 2842 46816
rect 2778 46756 2782 46812
rect 2782 46756 2838 46812
rect 2838 46756 2842 46812
rect 2778 46752 2842 46756
rect 2858 46812 2922 46816
rect 2858 46756 2862 46812
rect 2862 46756 2918 46812
rect 2918 46756 2922 46812
rect 2858 46752 2922 46756
rect 5952 46812 6016 46816
rect 5952 46756 5956 46812
rect 5956 46756 6012 46812
rect 6012 46756 6016 46812
rect 5952 46752 6016 46756
rect 6032 46812 6096 46816
rect 6032 46756 6036 46812
rect 6036 46756 6092 46812
rect 6092 46756 6096 46812
rect 6032 46752 6096 46756
rect 6112 46812 6176 46816
rect 6112 46756 6116 46812
rect 6116 46756 6172 46812
rect 6172 46756 6176 46812
rect 6112 46752 6176 46756
rect 6192 46812 6256 46816
rect 6192 46756 6196 46812
rect 6196 46756 6252 46812
rect 6252 46756 6256 46812
rect 6192 46752 6256 46756
rect 4285 46268 4349 46272
rect 4285 46212 4289 46268
rect 4289 46212 4345 46268
rect 4345 46212 4349 46268
rect 4285 46208 4349 46212
rect 4365 46268 4429 46272
rect 4365 46212 4369 46268
rect 4369 46212 4425 46268
rect 4425 46212 4429 46268
rect 4365 46208 4429 46212
rect 4445 46268 4509 46272
rect 4445 46212 4449 46268
rect 4449 46212 4505 46268
rect 4505 46212 4509 46268
rect 4445 46208 4509 46212
rect 4525 46268 4589 46272
rect 4525 46212 4529 46268
rect 4529 46212 4585 46268
rect 4585 46212 4589 46268
rect 4525 46208 4589 46212
rect 7618 46268 7682 46272
rect 7618 46212 7622 46268
rect 7622 46212 7678 46268
rect 7678 46212 7682 46268
rect 7618 46208 7682 46212
rect 7698 46268 7762 46272
rect 7698 46212 7702 46268
rect 7702 46212 7758 46268
rect 7758 46212 7762 46268
rect 7698 46208 7762 46212
rect 7778 46268 7842 46272
rect 7778 46212 7782 46268
rect 7782 46212 7838 46268
rect 7838 46212 7842 46268
rect 7778 46208 7842 46212
rect 7858 46268 7922 46272
rect 7858 46212 7862 46268
rect 7862 46212 7918 46268
rect 7918 46212 7922 46268
rect 7858 46208 7922 46212
rect 2618 45724 2682 45728
rect 2618 45668 2622 45724
rect 2622 45668 2678 45724
rect 2678 45668 2682 45724
rect 2618 45664 2682 45668
rect 2698 45724 2762 45728
rect 2698 45668 2702 45724
rect 2702 45668 2758 45724
rect 2758 45668 2762 45724
rect 2698 45664 2762 45668
rect 2778 45724 2842 45728
rect 2778 45668 2782 45724
rect 2782 45668 2838 45724
rect 2838 45668 2842 45724
rect 2778 45664 2842 45668
rect 2858 45724 2922 45728
rect 2858 45668 2862 45724
rect 2862 45668 2918 45724
rect 2918 45668 2922 45724
rect 2858 45664 2922 45668
rect 5952 45724 6016 45728
rect 5952 45668 5956 45724
rect 5956 45668 6012 45724
rect 6012 45668 6016 45724
rect 5952 45664 6016 45668
rect 6032 45724 6096 45728
rect 6032 45668 6036 45724
rect 6036 45668 6092 45724
rect 6092 45668 6096 45724
rect 6032 45664 6096 45668
rect 6112 45724 6176 45728
rect 6112 45668 6116 45724
rect 6116 45668 6172 45724
rect 6172 45668 6176 45724
rect 6112 45664 6176 45668
rect 6192 45724 6256 45728
rect 6192 45668 6196 45724
rect 6196 45668 6252 45724
rect 6252 45668 6256 45724
rect 6192 45664 6256 45668
rect 4285 45180 4349 45184
rect 4285 45124 4289 45180
rect 4289 45124 4345 45180
rect 4345 45124 4349 45180
rect 4285 45120 4349 45124
rect 4365 45180 4429 45184
rect 4365 45124 4369 45180
rect 4369 45124 4425 45180
rect 4425 45124 4429 45180
rect 4365 45120 4429 45124
rect 4445 45180 4509 45184
rect 4445 45124 4449 45180
rect 4449 45124 4505 45180
rect 4505 45124 4509 45180
rect 4445 45120 4509 45124
rect 4525 45180 4589 45184
rect 4525 45124 4529 45180
rect 4529 45124 4585 45180
rect 4585 45124 4589 45180
rect 4525 45120 4589 45124
rect 7618 45180 7682 45184
rect 7618 45124 7622 45180
rect 7622 45124 7678 45180
rect 7678 45124 7682 45180
rect 7618 45120 7682 45124
rect 7698 45180 7762 45184
rect 7698 45124 7702 45180
rect 7702 45124 7758 45180
rect 7758 45124 7762 45180
rect 7698 45120 7762 45124
rect 7778 45180 7842 45184
rect 7778 45124 7782 45180
rect 7782 45124 7838 45180
rect 7838 45124 7842 45180
rect 7778 45120 7842 45124
rect 7858 45180 7922 45184
rect 7858 45124 7862 45180
rect 7862 45124 7918 45180
rect 7918 45124 7922 45180
rect 7858 45120 7922 45124
rect 2618 44636 2682 44640
rect 2618 44580 2622 44636
rect 2622 44580 2678 44636
rect 2678 44580 2682 44636
rect 2618 44576 2682 44580
rect 2698 44636 2762 44640
rect 2698 44580 2702 44636
rect 2702 44580 2758 44636
rect 2758 44580 2762 44636
rect 2698 44576 2762 44580
rect 2778 44636 2842 44640
rect 2778 44580 2782 44636
rect 2782 44580 2838 44636
rect 2838 44580 2842 44636
rect 2778 44576 2842 44580
rect 2858 44636 2922 44640
rect 2858 44580 2862 44636
rect 2862 44580 2918 44636
rect 2918 44580 2922 44636
rect 2858 44576 2922 44580
rect 5952 44636 6016 44640
rect 5952 44580 5956 44636
rect 5956 44580 6012 44636
rect 6012 44580 6016 44636
rect 5952 44576 6016 44580
rect 6032 44636 6096 44640
rect 6032 44580 6036 44636
rect 6036 44580 6092 44636
rect 6092 44580 6096 44636
rect 6032 44576 6096 44580
rect 6112 44636 6176 44640
rect 6112 44580 6116 44636
rect 6116 44580 6172 44636
rect 6172 44580 6176 44636
rect 6112 44576 6176 44580
rect 6192 44636 6256 44640
rect 6192 44580 6196 44636
rect 6196 44580 6252 44636
rect 6252 44580 6256 44636
rect 6192 44576 6256 44580
rect 4285 44092 4349 44096
rect 4285 44036 4289 44092
rect 4289 44036 4345 44092
rect 4345 44036 4349 44092
rect 4285 44032 4349 44036
rect 4365 44092 4429 44096
rect 4365 44036 4369 44092
rect 4369 44036 4425 44092
rect 4425 44036 4429 44092
rect 4365 44032 4429 44036
rect 4445 44092 4509 44096
rect 4445 44036 4449 44092
rect 4449 44036 4505 44092
rect 4505 44036 4509 44092
rect 4445 44032 4509 44036
rect 4525 44092 4589 44096
rect 4525 44036 4529 44092
rect 4529 44036 4585 44092
rect 4585 44036 4589 44092
rect 4525 44032 4589 44036
rect 7618 44092 7682 44096
rect 7618 44036 7622 44092
rect 7622 44036 7678 44092
rect 7678 44036 7682 44092
rect 7618 44032 7682 44036
rect 7698 44092 7762 44096
rect 7698 44036 7702 44092
rect 7702 44036 7758 44092
rect 7758 44036 7762 44092
rect 7698 44032 7762 44036
rect 7778 44092 7842 44096
rect 7778 44036 7782 44092
rect 7782 44036 7838 44092
rect 7838 44036 7842 44092
rect 7778 44032 7842 44036
rect 7858 44092 7922 44096
rect 7858 44036 7862 44092
rect 7862 44036 7918 44092
rect 7918 44036 7922 44092
rect 7858 44032 7922 44036
rect 2618 43548 2682 43552
rect 2618 43492 2622 43548
rect 2622 43492 2678 43548
rect 2678 43492 2682 43548
rect 2618 43488 2682 43492
rect 2698 43548 2762 43552
rect 2698 43492 2702 43548
rect 2702 43492 2758 43548
rect 2758 43492 2762 43548
rect 2698 43488 2762 43492
rect 2778 43548 2842 43552
rect 2778 43492 2782 43548
rect 2782 43492 2838 43548
rect 2838 43492 2842 43548
rect 2778 43488 2842 43492
rect 2858 43548 2922 43552
rect 2858 43492 2862 43548
rect 2862 43492 2918 43548
rect 2918 43492 2922 43548
rect 2858 43488 2922 43492
rect 5952 43548 6016 43552
rect 5952 43492 5956 43548
rect 5956 43492 6012 43548
rect 6012 43492 6016 43548
rect 5952 43488 6016 43492
rect 6032 43548 6096 43552
rect 6032 43492 6036 43548
rect 6036 43492 6092 43548
rect 6092 43492 6096 43548
rect 6032 43488 6096 43492
rect 6112 43548 6176 43552
rect 6112 43492 6116 43548
rect 6116 43492 6172 43548
rect 6172 43492 6176 43548
rect 6112 43488 6176 43492
rect 6192 43548 6256 43552
rect 6192 43492 6196 43548
rect 6196 43492 6252 43548
rect 6252 43492 6256 43548
rect 6192 43488 6256 43492
rect 4285 43004 4349 43008
rect 4285 42948 4289 43004
rect 4289 42948 4345 43004
rect 4345 42948 4349 43004
rect 4285 42944 4349 42948
rect 4365 43004 4429 43008
rect 4365 42948 4369 43004
rect 4369 42948 4425 43004
rect 4425 42948 4429 43004
rect 4365 42944 4429 42948
rect 4445 43004 4509 43008
rect 4445 42948 4449 43004
rect 4449 42948 4505 43004
rect 4505 42948 4509 43004
rect 4445 42944 4509 42948
rect 4525 43004 4589 43008
rect 4525 42948 4529 43004
rect 4529 42948 4585 43004
rect 4585 42948 4589 43004
rect 4525 42944 4589 42948
rect 7618 43004 7682 43008
rect 7618 42948 7622 43004
rect 7622 42948 7678 43004
rect 7678 42948 7682 43004
rect 7618 42944 7682 42948
rect 7698 43004 7762 43008
rect 7698 42948 7702 43004
rect 7702 42948 7758 43004
rect 7758 42948 7762 43004
rect 7698 42944 7762 42948
rect 7778 43004 7842 43008
rect 7778 42948 7782 43004
rect 7782 42948 7838 43004
rect 7838 42948 7842 43004
rect 7778 42944 7842 42948
rect 7858 43004 7922 43008
rect 7858 42948 7862 43004
rect 7862 42948 7918 43004
rect 7918 42948 7922 43004
rect 7858 42944 7922 42948
rect 2618 42460 2682 42464
rect 2618 42404 2622 42460
rect 2622 42404 2678 42460
rect 2678 42404 2682 42460
rect 2618 42400 2682 42404
rect 2698 42460 2762 42464
rect 2698 42404 2702 42460
rect 2702 42404 2758 42460
rect 2758 42404 2762 42460
rect 2698 42400 2762 42404
rect 2778 42460 2842 42464
rect 2778 42404 2782 42460
rect 2782 42404 2838 42460
rect 2838 42404 2842 42460
rect 2778 42400 2842 42404
rect 2858 42460 2922 42464
rect 2858 42404 2862 42460
rect 2862 42404 2918 42460
rect 2918 42404 2922 42460
rect 2858 42400 2922 42404
rect 5952 42460 6016 42464
rect 5952 42404 5956 42460
rect 5956 42404 6012 42460
rect 6012 42404 6016 42460
rect 5952 42400 6016 42404
rect 6032 42460 6096 42464
rect 6032 42404 6036 42460
rect 6036 42404 6092 42460
rect 6092 42404 6096 42460
rect 6032 42400 6096 42404
rect 6112 42460 6176 42464
rect 6112 42404 6116 42460
rect 6116 42404 6172 42460
rect 6172 42404 6176 42460
rect 6112 42400 6176 42404
rect 6192 42460 6256 42464
rect 6192 42404 6196 42460
rect 6196 42404 6252 42460
rect 6252 42404 6256 42460
rect 6192 42400 6256 42404
rect 4285 41916 4349 41920
rect 4285 41860 4289 41916
rect 4289 41860 4345 41916
rect 4345 41860 4349 41916
rect 4285 41856 4349 41860
rect 4365 41916 4429 41920
rect 4365 41860 4369 41916
rect 4369 41860 4425 41916
rect 4425 41860 4429 41916
rect 4365 41856 4429 41860
rect 4445 41916 4509 41920
rect 4445 41860 4449 41916
rect 4449 41860 4505 41916
rect 4505 41860 4509 41916
rect 4445 41856 4509 41860
rect 4525 41916 4589 41920
rect 4525 41860 4529 41916
rect 4529 41860 4585 41916
rect 4585 41860 4589 41916
rect 4525 41856 4589 41860
rect 7618 41916 7682 41920
rect 7618 41860 7622 41916
rect 7622 41860 7678 41916
rect 7678 41860 7682 41916
rect 7618 41856 7682 41860
rect 7698 41916 7762 41920
rect 7698 41860 7702 41916
rect 7702 41860 7758 41916
rect 7758 41860 7762 41916
rect 7698 41856 7762 41860
rect 7778 41916 7842 41920
rect 7778 41860 7782 41916
rect 7782 41860 7838 41916
rect 7838 41860 7842 41916
rect 7778 41856 7842 41860
rect 7858 41916 7922 41920
rect 7858 41860 7862 41916
rect 7862 41860 7918 41916
rect 7918 41860 7922 41916
rect 7858 41856 7922 41860
rect 2618 41372 2682 41376
rect 2618 41316 2622 41372
rect 2622 41316 2678 41372
rect 2678 41316 2682 41372
rect 2618 41312 2682 41316
rect 2698 41372 2762 41376
rect 2698 41316 2702 41372
rect 2702 41316 2758 41372
rect 2758 41316 2762 41372
rect 2698 41312 2762 41316
rect 2778 41372 2842 41376
rect 2778 41316 2782 41372
rect 2782 41316 2838 41372
rect 2838 41316 2842 41372
rect 2778 41312 2842 41316
rect 2858 41372 2922 41376
rect 2858 41316 2862 41372
rect 2862 41316 2918 41372
rect 2918 41316 2922 41372
rect 2858 41312 2922 41316
rect 5952 41372 6016 41376
rect 5952 41316 5956 41372
rect 5956 41316 6012 41372
rect 6012 41316 6016 41372
rect 5952 41312 6016 41316
rect 6032 41372 6096 41376
rect 6032 41316 6036 41372
rect 6036 41316 6092 41372
rect 6092 41316 6096 41372
rect 6032 41312 6096 41316
rect 6112 41372 6176 41376
rect 6112 41316 6116 41372
rect 6116 41316 6172 41372
rect 6172 41316 6176 41372
rect 6112 41312 6176 41316
rect 6192 41372 6256 41376
rect 6192 41316 6196 41372
rect 6196 41316 6252 41372
rect 6252 41316 6256 41372
rect 6192 41312 6256 41316
rect 4285 40828 4349 40832
rect 4285 40772 4289 40828
rect 4289 40772 4345 40828
rect 4345 40772 4349 40828
rect 4285 40768 4349 40772
rect 4365 40828 4429 40832
rect 4365 40772 4369 40828
rect 4369 40772 4425 40828
rect 4425 40772 4429 40828
rect 4365 40768 4429 40772
rect 4445 40828 4509 40832
rect 4445 40772 4449 40828
rect 4449 40772 4505 40828
rect 4505 40772 4509 40828
rect 4445 40768 4509 40772
rect 4525 40828 4589 40832
rect 4525 40772 4529 40828
rect 4529 40772 4585 40828
rect 4585 40772 4589 40828
rect 4525 40768 4589 40772
rect 7618 40828 7682 40832
rect 7618 40772 7622 40828
rect 7622 40772 7678 40828
rect 7678 40772 7682 40828
rect 7618 40768 7682 40772
rect 7698 40828 7762 40832
rect 7698 40772 7702 40828
rect 7702 40772 7758 40828
rect 7758 40772 7762 40828
rect 7698 40768 7762 40772
rect 7778 40828 7842 40832
rect 7778 40772 7782 40828
rect 7782 40772 7838 40828
rect 7838 40772 7842 40828
rect 7778 40768 7842 40772
rect 7858 40828 7922 40832
rect 7858 40772 7862 40828
rect 7862 40772 7918 40828
rect 7918 40772 7922 40828
rect 7858 40768 7922 40772
rect 2618 40284 2682 40288
rect 2618 40228 2622 40284
rect 2622 40228 2678 40284
rect 2678 40228 2682 40284
rect 2618 40224 2682 40228
rect 2698 40284 2762 40288
rect 2698 40228 2702 40284
rect 2702 40228 2758 40284
rect 2758 40228 2762 40284
rect 2698 40224 2762 40228
rect 2778 40284 2842 40288
rect 2778 40228 2782 40284
rect 2782 40228 2838 40284
rect 2838 40228 2842 40284
rect 2778 40224 2842 40228
rect 2858 40284 2922 40288
rect 2858 40228 2862 40284
rect 2862 40228 2918 40284
rect 2918 40228 2922 40284
rect 2858 40224 2922 40228
rect 5952 40284 6016 40288
rect 5952 40228 5956 40284
rect 5956 40228 6012 40284
rect 6012 40228 6016 40284
rect 5952 40224 6016 40228
rect 6032 40284 6096 40288
rect 6032 40228 6036 40284
rect 6036 40228 6092 40284
rect 6092 40228 6096 40284
rect 6032 40224 6096 40228
rect 6112 40284 6176 40288
rect 6112 40228 6116 40284
rect 6116 40228 6172 40284
rect 6172 40228 6176 40284
rect 6112 40224 6176 40228
rect 6192 40284 6256 40288
rect 6192 40228 6196 40284
rect 6196 40228 6252 40284
rect 6252 40228 6256 40284
rect 6192 40224 6256 40228
rect 4285 39740 4349 39744
rect 4285 39684 4289 39740
rect 4289 39684 4345 39740
rect 4345 39684 4349 39740
rect 4285 39680 4349 39684
rect 4365 39740 4429 39744
rect 4365 39684 4369 39740
rect 4369 39684 4425 39740
rect 4425 39684 4429 39740
rect 4365 39680 4429 39684
rect 4445 39740 4509 39744
rect 4445 39684 4449 39740
rect 4449 39684 4505 39740
rect 4505 39684 4509 39740
rect 4445 39680 4509 39684
rect 4525 39740 4589 39744
rect 4525 39684 4529 39740
rect 4529 39684 4585 39740
rect 4585 39684 4589 39740
rect 4525 39680 4589 39684
rect 7618 39740 7682 39744
rect 7618 39684 7622 39740
rect 7622 39684 7678 39740
rect 7678 39684 7682 39740
rect 7618 39680 7682 39684
rect 7698 39740 7762 39744
rect 7698 39684 7702 39740
rect 7702 39684 7758 39740
rect 7758 39684 7762 39740
rect 7698 39680 7762 39684
rect 7778 39740 7842 39744
rect 7778 39684 7782 39740
rect 7782 39684 7838 39740
rect 7838 39684 7842 39740
rect 7778 39680 7842 39684
rect 7858 39740 7922 39744
rect 7858 39684 7862 39740
rect 7862 39684 7918 39740
rect 7918 39684 7922 39740
rect 7858 39680 7922 39684
rect 2618 39196 2682 39200
rect 2618 39140 2622 39196
rect 2622 39140 2678 39196
rect 2678 39140 2682 39196
rect 2618 39136 2682 39140
rect 2698 39196 2762 39200
rect 2698 39140 2702 39196
rect 2702 39140 2758 39196
rect 2758 39140 2762 39196
rect 2698 39136 2762 39140
rect 2778 39196 2842 39200
rect 2778 39140 2782 39196
rect 2782 39140 2838 39196
rect 2838 39140 2842 39196
rect 2778 39136 2842 39140
rect 2858 39196 2922 39200
rect 2858 39140 2862 39196
rect 2862 39140 2918 39196
rect 2918 39140 2922 39196
rect 2858 39136 2922 39140
rect 5952 39196 6016 39200
rect 5952 39140 5956 39196
rect 5956 39140 6012 39196
rect 6012 39140 6016 39196
rect 5952 39136 6016 39140
rect 6032 39196 6096 39200
rect 6032 39140 6036 39196
rect 6036 39140 6092 39196
rect 6092 39140 6096 39196
rect 6032 39136 6096 39140
rect 6112 39196 6176 39200
rect 6112 39140 6116 39196
rect 6116 39140 6172 39196
rect 6172 39140 6176 39196
rect 6112 39136 6176 39140
rect 6192 39196 6256 39200
rect 6192 39140 6196 39196
rect 6196 39140 6252 39196
rect 6252 39140 6256 39196
rect 6192 39136 6256 39140
rect 4285 38652 4349 38656
rect 4285 38596 4289 38652
rect 4289 38596 4345 38652
rect 4345 38596 4349 38652
rect 4285 38592 4349 38596
rect 4365 38652 4429 38656
rect 4365 38596 4369 38652
rect 4369 38596 4425 38652
rect 4425 38596 4429 38652
rect 4365 38592 4429 38596
rect 4445 38652 4509 38656
rect 4445 38596 4449 38652
rect 4449 38596 4505 38652
rect 4505 38596 4509 38652
rect 4445 38592 4509 38596
rect 4525 38652 4589 38656
rect 4525 38596 4529 38652
rect 4529 38596 4585 38652
rect 4585 38596 4589 38652
rect 4525 38592 4589 38596
rect 7618 38652 7682 38656
rect 7618 38596 7622 38652
rect 7622 38596 7678 38652
rect 7678 38596 7682 38652
rect 7618 38592 7682 38596
rect 7698 38652 7762 38656
rect 7698 38596 7702 38652
rect 7702 38596 7758 38652
rect 7758 38596 7762 38652
rect 7698 38592 7762 38596
rect 7778 38652 7842 38656
rect 7778 38596 7782 38652
rect 7782 38596 7838 38652
rect 7838 38596 7842 38652
rect 7778 38592 7842 38596
rect 7858 38652 7922 38656
rect 7858 38596 7862 38652
rect 7862 38596 7918 38652
rect 7918 38596 7922 38652
rect 7858 38592 7922 38596
rect 2618 38108 2682 38112
rect 2618 38052 2622 38108
rect 2622 38052 2678 38108
rect 2678 38052 2682 38108
rect 2618 38048 2682 38052
rect 2698 38108 2762 38112
rect 2698 38052 2702 38108
rect 2702 38052 2758 38108
rect 2758 38052 2762 38108
rect 2698 38048 2762 38052
rect 2778 38108 2842 38112
rect 2778 38052 2782 38108
rect 2782 38052 2838 38108
rect 2838 38052 2842 38108
rect 2778 38048 2842 38052
rect 2858 38108 2922 38112
rect 2858 38052 2862 38108
rect 2862 38052 2918 38108
rect 2918 38052 2922 38108
rect 2858 38048 2922 38052
rect 5952 38108 6016 38112
rect 5952 38052 5956 38108
rect 5956 38052 6012 38108
rect 6012 38052 6016 38108
rect 5952 38048 6016 38052
rect 6032 38108 6096 38112
rect 6032 38052 6036 38108
rect 6036 38052 6092 38108
rect 6092 38052 6096 38108
rect 6032 38048 6096 38052
rect 6112 38108 6176 38112
rect 6112 38052 6116 38108
rect 6116 38052 6172 38108
rect 6172 38052 6176 38108
rect 6112 38048 6176 38052
rect 6192 38108 6256 38112
rect 6192 38052 6196 38108
rect 6196 38052 6252 38108
rect 6252 38052 6256 38108
rect 6192 38048 6256 38052
rect 4285 37564 4349 37568
rect 4285 37508 4289 37564
rect 4289 37508 4345 37564
rect 4345 37508 4349 37564
rect 4285 37504 4349 37508
rect 4365 37564 4429 37568
rect 4365 37508 4369 37564
rect 4369 37508 4425 37564
rect 4425 37508 4429 37564
rect 4365 37504 4429 37508
rect 4445 37564 4509 37568
rect 4445 37508 4449 37564
rect 4449 37508 4505 37564
rect 4505 37508 4509 37564
rect 4445 37504 4509 37508
rect 4525 37564 4589 37568
rect 4525 37508 4529 37564
rect 4529 37508 4585 37564
rect 4585 37508 4589 37564
rect 4525 37504 4589 37508
rect 7618 37564 7682 37568
rect 7618 37508 7622 37564
rect 7622 37508 7678 37564
rect 7678 37508 7682 37564
rect 7618 37504 7682 37508
rect 7698 37564 7762 37568
rect 7698 37508 7702 37564
rect 7702 37508 7758 37564
rect 7758 37508 7762 37564
rect 7698 37504 7762 37508
rect 7778 37564 7842 37568
rect 7778 37508 7782 37564
rect 7782 37508 7838 37564
rect 7838 37508 7842 37564
rect 7778 37504 7842 37508
rect 7858 37564 7922 37568
rect 7858 37508 7862 37564
rect 7862 37508 7918 37564
rect 7918 37508 7922 37564
rect 7858 37504 7922 37508
rect 2618 37020 2682 37024
rect 2618 36964 2622 37020
rect 2622 36964 2678 37020
rect 2678 36964 2682 37020
rect 2618 36960 2682 36964
rect 2698 37020 2762 37024
rect 2698 36964 2702 37020
rect 2702 36964 2758 37020
rect 2758 36964 2762 37020
rect 2698 36960 2762 36964
rect 2778 37020 2842 37024
rect 2778 36964 2782 37020
rect 2782 36964 2838 37020
rect 2838 36964 2842 37020
rect 2778 36960 2842 36964
rect 2858 37020 2922 37024
rect 2858 36964 2862 37020
rect 2862 36964 2918 37020
rect 2918 36964 2922 37020
rect 2858 36960 2922 36964
rect 5952 37020 6016 37024
rect 5952 36964 5956 37020
rect 5956 36964 6012 37020
rect 6012 36964 6016 37020
rect 5952 36960 6016 36964
rect 6032 37020 6096 37024
rect 6032 36964 6036 37020
rect 6036 36964 6092 37020
rect 6092 36964 6096 37020
rect 6032 36960 6096 36964
rect 6112 37020 6176 37024
rect 6112 36964 6116 37020
rect 6116 36964 6172 37020
rect 6172 36964 6176 37020
rect 6112 36960 6176 36964
rect 6192 37020 6256 37024
rect 6192 36964 6196 37020
rect 6196 36964 6252 37020
rect 6252 36964 6256 37020
rect 6192 36960 6256 36964
rect 4285 36476 4349 36480
rect 4285 36420 4289 36476
rect 4289 36420 4345 36476
rect 4345 36420 4349 36476
rect 4285 36416 4349 36420
rect 4365 36476 4429 36480
rect 4365 36420 4369 36476
rect 4369 36420 4425 36476
rect 4425 36420 4429 36476
rect 4365 36416 4429 36420
rect 4445 36476 4509 36480
rect 4445 36420 4449 36476
rect 4449 36420 4505 36476
rect 4505 36420 4509 36476
rect 4445 36416 4509 36420
rect 4525 36476 4589 36480
rect 4525 36420 4529 36476
rect 4529 36420 4585 36476
rect 4585 36420 4589 36476
rect 4525 36416 4589 36420
rect 7618 36476 7682 36480
rect 7618 36420 7622 36476
rect 7622 36420 7678 36476
rect 7678 36420 7682 36476
rect 7618 36416 7682 36420
rect 7698 36476 7762 36480
rect 7698 36420 7702 36476
rect 7702 36420 7758 36476
rect 7758 36420 7762 36476
rect 7698 36416 7762 36420
rect 7778 36476 7842 36480
rect 7778 36420 7782 36476
rect 7782 36420 7838 36476
rect 7838 36420 7842 36476
rect 7778 36416 7842 36420
rect 7858 36476 7922 36480
rect 7858 36420 7862 36476
rect 7862 36420 7918 36476
rect 7918 36420 7922 36476
rect 7858 36416 7922 36420
rect 2618 35932 2682 35936
rect 2618 35876 2622 35932
rect 2622 35876 2678 35932
rect 2678 35876 2682 35932
rect 2618 35872 2682 35876
rect 2698 35932 2762 35936
rect 2698 35876 2702 35932
rect 2702 35876 2758 35932
rect 2758 35876 2762 35932
rect 2698 35872 2762 35876
rect 2778 35932 2842 35936
rect 2778 35876 2782 35932
rect 2782 35876 2838 35932
rect 2838 35876 2842 35932
rect 2778 35872 2842 35876
rect 2858 35932 2922 35936
rect 2858 35876 2862 35932
rect 2862 35876 2918 35932
rect 2918 35876 2922 35932
rect 2858 35872 2922 35876
rect 5952 35932 6016 35936
rect 5952 35876 5956 35932
rect 5956 35876 6012 35932
rect 6012 35876 6016 35932
rect 5952 35872 6016 35876
rect 6032 35932 6096 35936
rect 6032 35876 6036 35932
rect 6036 35876 6092 35932
rect 6092 35876 6096 35932
rect 6032 35872 6096 35876
rect 6112 35932 6176 35936
rect 6112 35876 6116 35932
rect 6116 35876 6172 35932
rect 6172 35876 6176 35932
rect 6112 35872 6176 35876
rect 6192 35932 6256 35936
rect 6192 35876 6196 35932
rect 6196 35876 6252 35932
rect 6252 35876 6256 35932
rect 6192 35872 6256 35876
rect 4285 35388 4349 35392
rect 4285 35332 4289 35388
rect 4289 35332 4345 35388
rect 4345 35332 4349 35388
rect 4285 35328 4349 35332
rect 4365 35388 4429 35392
rect 4365 35332 4369 35388
rect 4369 35332 4425 35388
rect 4425 35332 4429 35388
rect 4365 35328 4429 35332
rect 4445 35388 4509 35392
rect 4445 35332 4449 35388
rect 4449 35332 4505 35388
rect 4505 35332 4509 35388
rect 4445 35328 4509 35332
rect 4525 35388 4589 35392
rect 4525 35332 4529 35388
rect 4529 35332 4585 35388
rect 4585 35332 4589 35388
rect 4525 35328 4589 35332
rect 7618 35388 7682 35392
rect 7618 35332 7622 35388
rect 7622 35332 7678 35388
rect 7678 35332 7682 35388
rect 7618 35328 7682 35332
rect 7698 35388 7762 35392
rect 7698 35332 7702 35388
rect 7702 35332 7758 35388
rect 7758 35332 7762 35388
rect 7698 35328 7762 35332
rect 7778 35388 7842 35392
rect 7778 35332 7782 35388
rect 7782 35332 7838 35388
rect 7838 35332 7842 35388
rect 7778 35328 7842 35332
rect 7858 35388 7922 35392
rect 7858 35332 7862 35388
rect 7862 35332 7918 35388
rect 7918 35332 7922 35388
rect 7858 35328 7922 35332
rect 2618 34844 2682 34848
rect 2618 34788 2622 34844
rect 2622 34788 2678 34844
rect 2678 34788 2682 34844
rect 2618 34784 2682 34788
rect 2698 34844 2762 34848
rect 2698 34788 2702 34844
rect 2702 34788 2758 34844
rect 2758 34788 2762 34844
rect 2698 34784 2762 34788
rect 2778 34844 2842 34848
rect 2778 34788 2782 34844
rect 2782 34788 2838 34844
rect 2838 34788 2842 34844
rect 2778 34784 2842 34788
rect 2858 34844 2922 34848
rect 2858 34788 2862 34844
rect 2862 34788 2918 34844
rect 2918 34788 2922 34844
rect 2858 34784 2922 34788
rect 5952 34844 6016 34848
rect 5952 34788 5956 34844
rect 5956 34788 6012 34844
rect 6012 34788 6016 34844
rect 5952 34784 6016 34788
rect 6032 34844 6096 34848
rect 6032 34788 6036 34844
rect 6036 34788 6092 34844
rect 6092 34788 6096 34844
rect 6032 34784 6096 34788
rect 6112 34844 6176 34848
rect 6112 34788 6116 34844
rect 6116 34788 6172 34844
rect 6172 34788 6176 34844
rect 6112 34784 6176 34788
rect 6192 34844 6256 34848
rect 6192 34788 6196 34844
rect 6196 34788 6252 34844
rect 6252 34788 6256 34844
rect 6192 34784 6256 34788
rect 4285 34300 4349 34304
rect 4285 34244 4289 34300
rect 4289 34244 4345 34300
rect 4345 34244 4349 34300
rect 4285 34240 4349 34244
rect 4365 34300 4429 34304
rect 4365 34244 4369 34300
rect 4369 34244 4425 34300
rect 4425 34244 4429 34300
rect 4365 34240 4429 34244
rect 4445 34300 4509 34304
rect 4445 34244 4449 34300
rect 4449 34244 4505 34300
rect 4505 34244 4509 34300
rect 4445 34240 4509 34244
rect 4525 34300 4589 34304
rect 4525 34244 4529 34300
rect 4529 34244 4585 34300
rect 4585 34244 4589 34300
rect 4525 34240 4589 34244
rect 7618 34300 7682 34304
rect 7618 34244 7622 34300
rect 7622 34244 7678 34300
rect 7678 34244 7682 34300
rect 7618 34240 7682 34244
rect 7698 34300 7762 34304
rect 7698 34244 7702 34300
rect 7702 34244 7758 34300
rect 7758 34244 7762 34300
rect 7698 34240 7762 34244
rect 7778 34300 7842 34304
rect 7778 34244 7782 34300
rect 7782 34244 7838 34300
rect 7838 34244 7842 34300
rect 7778 34240 7842 34244
rect 7858 34300 7922 34304
rect 7858 34244 7862 34300
rect 7862 34244 7918 34300
rect 7918 34244 7922 34300
rect 7858 34240 7922 34244
rect 2618 33756 2682 33760
rect 2618 33700 2622 33756
rect 2622 33700 2678 33756
rect 2678 33700 2682 33756
rect 2618 33696 2682 33700
rect 2698 33756 2762 33760
rect 2698 33700 2702 33756
rect 2702 33700 2758 33756
rect 2758 33700 2762 33756
rect 2698 33696 2762 33700
rect 2778 33756 2842 33760
rect 2778 33700 2782 33756
rect 2782 33700 2838 33756
rect 2838 33700 2842 33756
rect 2778 33696 2842 33700
rect 2858 33756 2922 33760
rect 2858 33700 2862 33756
rect 2862 33700 2918 33756
rect 2918 33700 2922 33756
rect 2858 33696 2922 33700
rect 5952 33756 6016 33760
rect 5952 33700 5956 33756
rect 5956 33700 6012 33756
rect 6012 33700 6016 33756
rect 5952 33696 6016 33700
rect 6032 33756 6096 33760
rect 6032 33700 6036 33756
rect 6036 33700 6092 33756
rect 6092 33700 6096 33756
rect 6032 33696 6096 33700
rect 6112 33756 6176 33760
rect 6112 33700 6116 33756
rect 6116 33700 6172 33756
rect 6172 33700 6176 33756
rect 6112 33696 6176 33700
rect 6192 33756 6256 33760
rect 6192 33700 6196 33756
rect 6196 33700 6252 33756
rect 6252 33700 6256 33756
rect 6192 33696 6256 33700
rect 4285 33212 4349 33216
rect 4285 33156 4289 33212
rect 4289 33156 4345 33212
rect 4345 33156 4349 33212
rect 4285 33152 4349 33156
rect 4365 33212 4429 33216
rect 4365 33156 4369 33212
rect 4369 33156 4425 33212
rect 4425 33156 4429 33212
rect 4365 33152 4429 33156
rect 4445 33212 4509 33216
rect 4445 33156 4449 33212
rect 4449 33156 4505 33212
rect 4505 33156 4509 33212
rect 4445 33152 4509 33156
rect 4525 33212 4589 33216
rect 4525 33156 4529 33212
rect 4529 33156 4585 33212
rect 4585 33156 4589 33212
rect 4525 33152 4589 33156
rect 7618 33212 7682 33216
rect 7618 33156 7622 33212
rect 7622 33156 7678 33212
rect 7678 33156 7682 33212
rect 7618 33152 7682 33156
rect 7698 33212 7762 33216
rect 7698 33156 7702 33212
rect 7702 33156 7758 33212
rect 7758 33156 7762 33212
rect 7698 33152 7762 33156
rect 7778 33212 7842 33216
rect 7778 33156 7782 33212
rect 7782 33156 7838 33212
rect 7838 33156 7842 33212
rect 7778 33152 7842 33156
rect 7858 33212 7922 33216
rect 7858 33156 7862 33212
rect 7862 33156 7918 33212
rect 7918 33156 7922 33212
rect 7858 33152 7922 33156
rect 2618 32668 2682 32672
rect 2618 32612 2622 32668
rect 2622 32612 2678 32668
rect 2678 32612 2682 32668
rect 2618 32608 2682 32612
rect 2698 32668 2762 32672
rect 2698 32612 2702 32668
rect 2702 32612 2758 32668
rect 2758 32612 2762 32668
rect 2698 32608 2762 32612
rect 2778 32668 2842 32672
rect 2778 32612 2782 32668
rect 2782 32612 2838 32668
rect 2838 32612 2842 32668
rect 2778 32608 2842 32612
rect 2858 32668 2922 32672
rect 2858 32612 2862 32668
rect 2862 32612 2918 32668
rect 2918 32612 2922 32668
rect 2858 32608 2922 32612
rect 5952 32668 6016 32672
rect 5952 32612 5956 32668
rect 5956 32612 6012 32668
rect 6012 32612 6016 32668
rect 5952 32608 6016 32612
rect 6032 32668 6096 32672
rect 6032 32612 6036 32668
rect 6036 32612 6092 32668
rect 6092 32612 6096 32668
rect 6032 32608 6096 32612
rect 6112 32668 6176 32672
rect 6112 32612 6116 32668
rect 6116 32612 6172 32668
rect 6172 32612 6176 32668
rect 6112 32608 6176 32612
rect 6192 32668 6256 32672
rect 6192 32612 6196 32668
rect 6196 32612 6252 32668
rect 6252 32612 6256 32668
rect 6192 32608 6256 32612
rect 4285 32124 4349 32128
rect 4285 32068 4289 32124
rect 4289 32068 4345 32124
rect 4345 32068 4349 32124
rect 4285 32064 4349 32068
rect 4365 32124 4429 32128
rect 4365 32068 4369 32124
rect 4369 32068 4425 32124
rect 4425 32068 4429 32124
rect 4365 32064 4429 32068
rect 4445 32124 4509 32128
rect 4445 32068 4449 32124
rect 4449 32068 4505 32124
rect 4505 32068 4509 32124
rect 4445 32064 4509 32068
rect 4525 32124 4589 32128
rect 4525 32068 4529 32124
rect 4529 32068 4585 32124
rect 4585 32068 4589 32124
rect 4525 32064 4589 32068
rect 7618 32124 7682 32128
rect 7618 32068 7622 32124
rect 7622 32068 7678 32124
rect 7678 32068 7682 32124
rect 7618 32064 7682 32068
rect 7698 32124 7762 32128
rect 7698 32068 7702 32124
rect 7702 32068 7758 32124
rect 7758 32068 7762 32124
rect 7698 32064 7762 32068
rect 7778 32124 7842 32128
rect 7778 32068 7782 32124
rect 7782 32068 7838 32124
rect 7838 32068 7842 32124
rect 7778 32064 7842 32068
rect 7858 32124 7922 32128
rect 7858 32068 7862 32124
rect 7862 32068 7918 32124
rect 7918 32068 7922 32124
rect 7858 32064 7922 32068
rect 2618 31580 2682 31584
rect 2618 31524 2622 31580
rect 2622 31524 2678 31580
rect 2678 31524 2682 31580
rect 2618 31520 2682 31524
rect 2698 31580 2762 31584
rect 2698 31524 2702 31580
rect 2702 31524 2758 31580
rect 2758 31524 2762 31580
rect 2698 31520 2762 31524
rect 2778 31580 2842 31584
rect 2778 31524 2782 31580
rect 2782 31524 2838 31580
rect 2838 31524 2842 31580
rect 2778 31520 2842 31524
rect 2858 31580 2922 31584
rect 2858 31524 2862 31580
rect 2862 31524 2918 31580
rect 2918 31524 2922 31580
rect 2858 31520 2922 31524
rect 5952 31580 6016 31584
rect 5952 31524 5956 31580
rect 5956 31524 6012 31580
rect 6012 31524 6016 31580
rect 5952 31520 6016 31524
rect 6032 31580 6096 31584
rect 6032 31524 6036 31580
rect 6036 31524 6092 31580
rect 6092 31524 6096 31580
rect 6032 31520 6096 31524
rect 6112 31580 6176 31584
rect 6112 31524 6116 31580
rect 6116 31524 6172 31580
rect 6172 31524 6176 31580
rect 6112 31520 6176 31524
rect 6192 31580 6256 31584
rect 6192 31524 6196 31580
rect 6196 31524 6252 31580
rect 6252 31524 6256 31580
rect 6192 31520 6256 31524
rect 4285 31036 4349 31040
rect 4285 30980 4289 31036
rect 4289 30980 4345 31036
rect 4345 30980 4349 31036
rect 4285 30976 4349 30980
rect 4365 31036 4429 31040
rect 4365 30980 4369 31036
rect 4369 30980 4425 31036
rect 4425 30980 4429 31036
rect 4365 30976 4429 30980
rect 4445 31036 4509 31040
rect 4445 30980 4449 31036
rect 4449 30980 4505 31036
rect 4505 30980 4509 31036
rect 4445 30976 4509 30980
rect 4525 31036 4589 31040
rect 4525 30980 4529 31036
rect 4529 30980 4585 31036
rect 4585 30980 4589 31036
rect 4525 30976 4589 30980
rect 7618 31036 7682 31040
rect 7618 30980 7622 31036
rect 7622 30980 7678 31036
rect 7678 30980 7682 31036
rect 7618 30976 7682 30980
rect 7698 31036 7762 31040
rect 7698 30980 7702 31036
rect 7702 30980 7758 31036
rect 7758 30980 7762 31036
rect 7698 30976 7762 30980
rect 7778 31036 7842 31040
rect 7778 30980 7782 31036
rect 7782 30980 7838 31036
rect 7838 30980 7842 31036
rect 7778 30976 7842 30980
rect 7858 31036 7922 31040
rect 7858 30980 7862 31036
rect 7862 30980 7918 31036
rect 7918 30980 7922 31036
rect 7858 30976 7922 30980
rect 2618 30492 2682 30496
rect 2618 30436 2622 30492
rect 2622 30436 2678 30492
rect 2678 30436 2682 30492
rect 2618 30432 2682 30436
rect 2698 30492 2762 30496
rect 2698 30436 2702 30492
rect 2702 30436 2758 30492
rect 2758 30436 2762 30492
rect 2698 30432 2762 30436
rect 2778 30492 2842 30496
rect 2778 30436 2782 30492
rect 2782 30436 2838 30492
rect 2838 30436 2842 30492
rect 2778 30432 2842 30436
rect 2858 30492 2922 30496
rect 2858 30436 2862 30492
rect 2862 30436 2918 30492
rect 2918 30436 2922 30492
rect 2858 30432 2922 30436
rect 5952 30492 6016 30496
rect 5952 30436 5956 30492
rect 5956 30436 6012 30492
rect 6012 30436 6016 30492
rect 5952 30432 6016 30436
rect 6032 30492 6096 30496
rect 6032 30436 6036 30492
rect 6036 30436 6092 30492
rect 6092 30436 6096 30492
rect 6032 30432 6096 30436
rect 6112 30492 6176 30496
rect 6112 30436 6116 30492
rect 6116 30436 6172 30492
rect 6172 30436 6176 30492
rect 6112 30432 6176 30436
rect 6192 30492 6256 30496
rect 6192 30436 6196 30492
rect 6196 30436 6252 30492
rect 6252 30436 6256 30492
rect 6192 30432 6256 30436
rect 4285 29948 4349 29952
rect 4285 29892 4289 29948
rect 4289 29892 4345 29948
rect 4345 29892 4349 29948
rect 4285 29888 4349 29892
rect 4365 29948 4429 29952
rect 4365 29892 4369 29948
rect 4369 29892 4425 29948
rect 4425 29892 4429 29948
rect 4365 29888 4429 29892
rect 4445 29948 4509 29952
rect 4445 29892 4449 29948
rect 4449 29892 4505 29948
rect 4505 29892 4509 29948
rect 4445 29888 4509 29892
rect 4525 29948 4589 29952
rect 4525 29892 4529 29948
rect 4529 29892 4585 29948
rect 4585 29892 4589 29948
rect 4525 29888 4589 29892
rect 7618 29948 7682 29952
rect 7618 29892 7622 29948
rect 7622 29892 7678 29948
rect 7678 29892 7682 29948
rect 7618 29888 7682 29892
rect 7698 29948 7762 29952
rect 7698 29892 7702 29948
rect 7702 29892 7758 29948
rect 7758 29892 7762 29948
rect 7698 29888 7762 29892
rect 7778 29948 7842 29952
rect 7778 29892 7782 29948
rect 7782 29892 7838 29948
rect 7838 29892 7842 29948
rect 7778 29888 7842 29892
rect 7858 29948 7922 29952
rect 7858 29892 7862 29948
rect 7862 29892 7918 29948
rect 7918 29892 7922 29948
rect 7858 29888 7922 29892
rect 2618 29404 2682 29408
rect 2618 29348 2622 29404
rect 2622 29348 2678 29404
rect 2678 29348 2682 29404
rect 2618 29344 2682 29348
rect 2698 29404 2762 29408
rect 2698 29348 2702 29404
rect 2702 29348 2758 29404
rect 2758 29348 2762 29404
rect 2698 29344 2762 29348
rect 2778 29404 2842 29408
rect 2778 29348 2782 29404
rect 2782 29348 2838 29404
rect 2838 29348 2842 29404
rect 2778 29344 2842 29348
rect 2858 29404 2922 29408
rect 2858 29348 2862 29404
rect 2862 29348 2918 29404
rect 2918 29348 2922 29404
rect 2858 29344 2922 29348
rect 5952 29404 6016 29408
rect 5952 29348 5956 29404
rect 5956 29348 6012 29404
rect 6012 29348 6016 29404
rect 5952 29344 6016 29348
rect 6032 29404 6096 29408
rect 6032 29348 6036 29404
rect 6036 29348 6092 29404
rect 6092 29348 6096 29404
rect 6032 29344 6096 29348
rect 6112 29404 6176 29408
rect 6112 29348 6116 29404
rect 6116 29348 6172 29404
rect 6172 29348 6176 29404
rect 6112 29344 6176 29348
rect 6192 29404 6256 29408
rect 6192 29348 6196 29404
rect 6196 29348 6252 29404
rect 6252 29348 6256 29404
rect 6192 29344 6256 29348
rect 4285 28860 4349 28864
rect 4285 28804 4289 28860
rect 4289 28804 4345 28860
rect 4345 28804 4349 28860
rect 4285 28800 4349 28804
rect 4365 28860 4429 28864
rect 4365 28804 4369 28860
rect 4369 28804 4425 28860
rect 4425 28804 4429 28860
rect 4365 28800 4429 28804
rect 4445 28860 4509 28864
rect 4445 28804 4449 28860
rect 4449 28804 4505 28860
rect 4505 28804 4509 28860
rect 4445 28800 4509 28804
rect 4525 28860 4589 28864
rect 4525 28804 4529 28860
rect 4529 28804 4585 28860
rect 4585 28804 4589 28860
rect 4525 28800 4589 28804
rect 7618 28860 7682 28864
rect 7618 28804 7622 28860
rect 7622 28804 7678 28860
rect 7678 28804 7682 28860
rect 7618 28800 7682 28804
rect 7698 28860 7762 28864
rect 7698 28804 7702 28860
rect 7702 28804 7758 28860
rect 7758 28804 7762 28860
rect 7698 28800 7762 28804
rect 7778 28860 7842 28864
rect 7778 28804 7782 28860
rect 7782 28804 7838 28860
rect 7838 28804 7842 28860
rect 7778 28800 7842 28804
rect 7858 28860 7922 28864
rect 7858 28804 7862 28860
rect 7862 28804 7918 28860
rect 7918 28804 7922 28860
rect 7858 28800 7922 28804
rect 2618 28316 2682 28320
rect 2618 28260 2622 28316
rect 2622 28260 2678 28316
rect 2678 28260 2682 28316
rect 2618 28256 2682 28260
rect 2698 28316 2762 28320
rect 2698 28260 2702 28316
rect 2702 28260 2758 28316
rect 2758 28260 2762 28316
rect 2698 28256 2762 28260
rect 2778 28316 2842 28320
rect 2778 28260 2782 28316
rect 2782 28260 2838 28316
rect 2838 28260 2842 28316
rect 2778 28256 2842 28260
rect 2858 28316 2922 28320
rect 2858 28260 2862 28316
rect 2862 28260 2918 28316
rect 2918 28260 2922 28316
rect 2858 28256 2922 28260
rect 5952 28316 6016 28320
rect 5952 28260 5956 28316
rect 5956 28260 6012 28316
rect 6012 28260 6016 28316
rect 5952 28256 6016 28260
rect 6032 28316 6096 28320
rect 6032 28260 6036 28316
rect 6036 28260 6092 28316
rect 6092 28260 6096 28316
rect 6032 28256 6096 28260
rect 6112 28316 6176 28320
rect 6112 28260 6116 28316
rect 6116 28260 6172 28316
rect 6172 28260 6176 28316
rect 6112 28256 6176 28260
rect 6192 28316 6256 28320
rect 6192 28260 6196 28316
rect 6196 28260 6252 28316
rect 6252 28260 6256 28316
rect 6192 28256 6256 28260
rect 4285 27772 4349 27776
rect 4285 27716 4289 27772
rect 4289 27716 4345 27772
rect 4345 27716 4349 27772
rect 4285 27712 4349 27716
rect 4365 27772 4429 27776
rect 4365 27716 4369 27772
rect 4369 27716 4425 27772
rect 4425 27716 4429 27772
rect 4365 27712 4429 27716
rect 4445 27772 4509 27776
rect 4445 27716 4449 27772
rect 4449 27716 4505 27772
rect 4505 27716 4509 27772
rect 4445 27712 4509 27716
rect 4525 27772 4589 27776
rect 4525 27716 4529 27772
rect 4529 27716 4585 27772
rect 4585 27716 4589 27772
rect 4525 27712 4589 27716
rect 7618 27772 7682 27776
rect 7618 27716 7622 27772
rect 7622 27716 7678 27772
rect 7678 27716 7682 27772
rect 7618 27712 7682 27716
rect 7698 27772 7762 27776
rect 7698 27716 7702 27772
rect 7702 27716 7758 27772
rect 7758 27716 7762 27772
rect 7698 27712 7762 27716
rect 7778 27772 7842 27776
rect 7778 27716 7782 27772
rect 7782 27716 7838 27772
rect 7838 27716 7842 27772
rect 7778 27712 7842 27716
rect 7858 27772 7922 27776
rect 7858 27716 7862 27772
rect 7862 27716 7918 27772
rect 7918 27716 7922 27772
rect 7858 27712 7922 27716
rect 2618 27228 2682 27232
rect 2618 27172 2622 27228
rect 2622 27172 2678 27228
rect 2678 27172 2682 27228
rect 2618 27168 2682 27172
rect 2698 27228 2762 27232
rect 2698 27172 2702 27228
rect 2702 27172 2758 27228
rect 2758 27172 2762 27228
rect 2698 27168 2762 27172
rect 2778 27228 2842 27232
rect 2778 27172 2782 27228
rect 2782 27172 2838 27228
rect 2838 27172 2842 27228
rect 2778 27168 2842 27172
rect 2858 27228 2922 27232
rect 2858 27172 2862 27228
rect 2862 27172 2918 27228
rect 2918 27172 2922 27228
rect 2858 27168 2922 27172
rect 5952 27228 6016 27232
rect 5952 27172 5956 27228
rect 5956 27172 6012 27228
rect 6012 27172 6016 27228
rect 5952 27168 6016 27172
rect 6032 27228 6096 27232
rect 6032 27172 6036 27228
rect 6036 27172 6092 27228
rect 6092 27172 6096 27228
rect 6032 27168 6096 27172
rect 6112 27228 6176 27232
rect 6112 27172 6116 27228
rect 6116 27172 6172 27228
rect 6172 27172 6176 27228
rect 6112 27168 6176 27172
rect 6192 27228 6256 27232
rect 6192 27172 6196 27228
rect 6196 27172 6252 27228
rect 6252 27172 6256 27228
rect 6192 27168 6256 27172
rect 4285 26684 4349 26688
rect 4285 26628 4289 26684
rect 4289 26628 4345 26684
rect 4345 26628 4349 26684
rect 4285 26624 4349 26628
rect 4365 26684 4429 26688
rect 4365 26628 4369 26684
rect 4369 26628 4425 26684
rect 4425 26628 4429 26684
rect 4365 26624 4429 26628
rect 4445 26684 4509 26688
rect 4445 26628 4449 26684
rect 4449 26628 4505 26684
rect 4505 26628 4509 26684
rect 4445 26624 4509 26628
rect 4525 26684 4589 26688
rect 4525 26628 4529 26684
rect 4529 26628 4585 26684
rect 4585 26628 4589 26684
rect 4525 26624 4589 26628
rect 7618 26684 7682 26688
rect 7618 26628 7622 26684
rect 7622 26628 7678 26684
rect 7678 26628 7682 26684
rect 7618 26624 7682 26628
rect 7698 26684 7762 26688
rect 7698 26628 7702 26684
rect 7702 26628 7758 26684
rect 7758 26628 7762 26684
rect 7698 26624 7762 26628
rect 7778 26684 7842 26688
rect 7778 26628 7782 26684
rect 7782 26628 7838 26684
rect 7838 26628 7842 26684
rect 7778 26624 7842 26628
rect 7858 26684 7922 26688
rect 7858 26628 7862 26684
rect 7862 26628 7918 26684
rect 7918 26628 7922 26684
rect 7858 26624 7922 26628
rect 2618 26140 2682 26144
rect 2618 26084 2622 26140
rect 2622 26084 2678 26140
rect 2678 26084 2682 26140
rect 2618 26080 2682 26084
rect 2698 26140 2762 26144
rect 2698 26084 2702 26140
rect 2702 26084 2758 26140
rect 2758 26084 2762 26140
rect 2698 26080 2762 26084
rect 2778 26140 2842 26144
rect 2778 26084 2782 26140
rect 2782 26084 2838 26140
rect 2838 26084 2842 26140
rect 2778 26080 2842 26084
rect 2858 26140 2922 26144
rect 2858 26084 2862 26140
rect 2862 26084 2918 26140
rect 2918 26084 2922 26140
rect 2858 26080 2922 26084
rect 5952 26140 6016 26144
rect 5952 26084 5956 26140
rect 5956 26084 6012 26140
rect 6012 26084 6016 26140
rect 5952 26080 6016 26084
rect 6032 26140 6096 26144
rect 6032 26084 6036 26140
rect 6036 26084 6092 26140
rect 6092 26084 6096 26140
rect 6032 26080 6096 26084
rect 6112 26140 6176 26144
rect 6112 26084 6116 26140
rect 6116 26084 6172 26140
rect 6172 26084 6176 26140
rect 6112 26080 6176 26084
rect 6192 26140 6256 26144
rect 6192 26084 6196 26140
rect 6196 26084 6252 26140
rect 6252 26084 6256 26140
rect 6192 26080 6256 26084
rect 4285 25596 4349 25600
rect 4285 25540 4289 25596
rect 4289 25540 4345 25596
rect 4345 25540 4349 25596
rect 4285 25536 4349 25540
rect 4365 25596 4429 25600
rect 4365 25540 4369 25596
rect 4369 25540 4425 25596
rect 4425 25540 4429 25596
rect 4365 25536 4429 25540
rect 4445 25596 4509 25600
rect 4445 25540 4449 25596
rect 4449 25540 4505 25596
rect 4505 25540 4509 25596
rect 4445 25536 4509 25540
rect 4525 25596 4589 25600
rect 4525 25540 4529 25596
rect 4529 25540 4585 25596
rect 4585 25540 4589 25596
rect 4525 25536 4589 25540
rect 7618 25596 7682 25600
rect 7618 25540 7622 25596
rect 7622 25540 7678 25596
rect 7678 25540 7682 25596
rect 7618 25536 7682 25540
rect 7698 25596 7762 25600
rect 7698 25540 7702 25596
rect 7702 25540 7758 25596
rect 7758 25540 7762 25596
rect 7698 25536 7762 25540
rect 7778 25596 7842 25600
rect 7778 25540 7782 25596
rect 7782 25540 7838 25596
rect 7838 25540 7842 25596
rect 7778 25536 7842 25540
rect 7858 25596 7922 25600
rect 7858 25540 7862 25596
rect 7862 25540 7918 25596
rect 7918 25540 7922 25596
rect 7858 25536 7922 25540
rect 2618 25052 2682 25056
rect 2618 24996 2622 25052
rect 2622 24996 2678 25052
rect 2678 24996 2682 25052
rect 2618 24992 2682 24996
rect 2698 25052 2762 25056
rect 2698 24996 2702 25052
rect 2702 24996 2758 25052
rect 2758 24996 2762 25052
rect 2698 24992 2762 24996
rect 2778 25052 2842 25056
rect 2778 24996 2782 25052
rect 2782 24996 2838 25052
rect 2838 24996 2842 25052
rect 2778 24992 2842 24996
rect 2858 25052 2922 25056
rect 2858 24996 2862 25052
rect 2862 24996 2918 25052
rect 2918 24996 2922 25052
rect 2858 24992 2922 24996
rect 5952 25052 6016 25056
rect 5952 24996 5956 25052
rect 5956 24996 6012 25052
rect 6012 24996 6016 25052
rect 5952 24992 6016 24996
rect 6032 25052 6096 25056
rect 6032 24996 6036 25052
rect 6036 24996 6092 25052
rect 6092 24996 6096 25052
rect 6032 24992 6096 24996
rect 6112 25052 6176 25056
rect 6112 24996 6116 25052
rect 6116 24996 6172 25052
rect 6172 24996 6176 25052
rect 6112 24992 6176 24996
rect 6192 25052 6256 25056
rect 6192 24996 6196 25052
rect 6196 24996 6252 25052
rect 6252 24996 6256 25052
rect 6192 24992 6256 24996
rect 4285 24508 4349 24512
rect 4285 24452 4289 24508
rect 4289 24452 4345 24508
rect 4345 24452 4349 24508
rect 4285 24448 4349 24452
rect 4365 24508 4429 24512
rect 4365 24452 4369 24508
rect 4369 24452 4425 24508
rect 4425 24452 4429 24508
rect 4365 24448 4429 24452
rect 4445 24508 4509 24512
rect 4445 24452 4449 24508
rect 4449 24452 4505 24508
rect 4505 24452 4509 24508
rect 4445 24448 4509 24452
rect 4525 24508 4589 24512
rect 4525 24452 4529 24508
rect 4529 24452 4585 24508
rect 4585 24452 4589 24508
rect 4525 24448 4589 24452
rect 7618 24508 7682 24512
rect 7618 24452 7622 24508
rect 7622 24452 7678 24508
rect 7678 24452 7682 24508
rect 7618 24448 7682 24452
rect 7698 24508 7762 24512
rect 7698 24452 7702 24508
rect 7702 24452 7758 24508
rect 7758 24452 7762 24508
rect 7698 24448 7762 24452
rect 7778 24508 7842 24512
rect 7778 24452 7782 24508
rect 7782 24452 7838 24508
rect 7838 24452 7842 24508
rect 7778 24448 7842 24452
rect 7858 24508 7922 24512
rect 7858 24452 7862 24508
rect 7862 24452 7918 24508
rect 7918 24452 7922 24508
rect 7858 24448 7922 24452
rect 2618 23964 2682 23968
rect 2618 23908 2622 23964
rect 2622 23908 2678 23964
rect 2678 23908 2682 23964
rect 2618 23904 2682 23908
rect 2698 23964 2762 23968
rect 2698 23908 2702 23964
rect 2702 23908 2758 23964
rect 2758 23908 2762 23964
rect 2698 23904 2762 23908
rect 2778 23964 2842 23968
rect 2778 23908 2782 23964
rect 2782 23908 2838 23964
rect 2838 23908 2842 23964
rect 2778 23904 2842 23908
rect 2858 23964 2922 23968
rect 2858 23908 2862 23964
rect 2862 23908 2918 23964
rect 2918 23908 2922 23964
rect 2858 23904 2922 23908
rect 5952 23964 6016 23968
rect 5952 23908 5956 23964
rect 5956 23908 6012 23964
rect 6012 23908 6016 23964
rect 5952 23904 6016 23908
rect 6032 23964 6096 23968
rect 6032 23908 6036 23964
rect 6036 23908 6092 23964
rect 6092 23908 6096 23964
rect 6032 23904 6096 23908
rect 6112 23964 6176 23968
rect 6112 23908 6116 23964
rect 6116 23908 6172 23964
rect 6172 23908 6176 23964
rect 6112 23904 6176 23908
rect 6192 23964 6256 23968
rect 6192 23908 6196 23964
rect 6196 23908 6252 23964
rect 6252 23908 6256 23964
rect 6192 23904 6256 23908
rect 4285 23420 4349 23424
rect 4285 23364 4289 23420
rect 4289 23364 4345 23420
rect 4345 23364 4349 23420
rect 4285 23360 4349 23364
rect 4365 23420 4429 23424
rect 4365 23364 4369 23420
rect 4369 23364 4425 23420
rect 4425 23364 4429 23420
rect 4365 23360 4429 23364
rect 4445 23420 4509 23424
rect 4445 23364 4449 23420
rect 4449 23364 4505 23420
rect 4505 23364 4509 23420
rect 4445 23360 4509 23364
rect 4525 23420 4589 23424
rect 4525 23364 4529 23420
rect 4529 23364 4585 23420
rect 4585 23364 4589 23420
rect 4525 23360 4589 23364
rect 7618 23420 7682 23424
rect 7618 23364 7622 23420
rect 7622 23364 7678 23420
rect 7678 23364 7682 23420
rect 7618 23360 7682 23364
rect 7698 23420 7762 23424
rect 7698 23364 7702 23420
rect 7702 23364 7758 23420
rect 7758 23364 7762 23420
rect 7698 23360 7762 23364
rect 7778 23420 7842 23424
rect 7778 23364 7782 23420
rect 7782 23364 7838 23420
rect 7838 23364 7842 23420
rect 7778 23360 7842 23364
rect 7858 23420 7922 23424
rect 7858 23364 7862 23420
rect 7862 23364 7918 23420
rect 7918 23364 7922 23420
rect 7858 23360 7922 23364
rect 2618 22876 2682 22880
rect 2618 22820 2622 22876
rect 2622 22820 2678 22876
rect 2678 22820 2682 22876
rect 2618 22816 2682 22820
rect 2698 22876 2762 22880
rect 2698 22820 2702 22876
rect 2702 22820 2758 22876
rect 2758 22820 2762 22876
rect 2698 22816 2762 22820
rect 2778 22876 2842 22880
rect 2778 22820 2782 22876
rect 2782 22820 2838 22876
rect 2838 22820 2842 22876
rect 2778 22816 2842 22820
rect 2858 22876 2922 22880
rect 2858 22820 2862 22876
rect 2862 22820 2918 22876
rect 2918 22820 2922 22876
rect 2858 22816 2922 22820
rect 5952 22876 6016 22880
rect 5952 22820 5956 22876
rect 5956 22820 6012 22876
rect 6012 22820 6016 22876
rect 5952 22816 6016 22820
rect 6032 22876 6096 22880
rect 6032 22820 6036 22876
rect 6036 22820 6092 22876
rect 6092 22820 6096 22876
rect 6032 22816 6096 22820
rect 6112 22876 6176 22880
rect 6112 22820 6116 22876
rect 6116 22820 6172 22876
rect 6172 22820 6176 22876
rect 6112 22816 6176 22820
rect 6192 22876 6256 22880
rect 6192 22820 6196 22876
rect 6196 22820 6252 22876
rect 6252 22820 6256 22876
rect 6192 22816 6256 22820
rect 4285 22332 4349 22336
rect 4285 22276 4289 22332
rect 4289 22276 4345 22332
rect 4345 22276 4349 22332
rect 4285 22272 4349 22276
rect 4365 22332 4429 22336
rect 4365 22276 4369 22332
rect 4369 22276 4425 22332
rect 4425 22276 4429 22332
rect 4365 22272 4429 22276
rect 4445 22332 4509 22336
rect 4445 22276 4449 22332
rect 4449 22276 4505 22332
rect 4505 22276 4509 22332
rect 4445 22272 4509 22276
rect 4525 22332 4589 22336
rect 4525 22276 4529 22332
rect 4529 22276 4585 22332
rect 4585 22276 4589 22332
rect 4525 22272 4589 22276
rect 7618 22332 7682 22336
rect 7618 22276 7622 22332
rect 7622 22276 7678 22332
rect 7678 22276 7682 22332
rect 7618 22272 7682 22276
rect 7698 22332 7762 22336
rect 7698 22276 7702 22332
rect 7702 22276 7758 22332
rect 7758 22276 7762 22332
rect 7698 22272 7762 22276
rect 7778 22332 7842 22336
rect 7778 22276 7782 22332
rect 7782 22276 7838 22332
rect 7838 22276 7842 22332
rect 7778 22272 7842 22276
rect 7858 22332 7922 22336
rect 7858 22276 7862 22332
rect 7862 22276 7918 22332
rect 7918 22276 7922 22332
rect 7858 22272 7922 22276
rect 2618 21788 2682 21792
rect 2618 21732 2622 21788
rect 2622 21732 2678 21788
rect 2678 21732 2682 21788
rect 2618 21728 2682 21732
rect 2698 21788 2762 21792
rect 2698 21732 2702 21788
rect 2702 21732 2758 21788
rect 2758 21732 2762 21788
rect 2698 21728 2762 21732
rect 2778 21788 2842 21792
rect 2778 21732 2782 21788
rect 2782 21732 2838 21788
rect 2838 21732 2842 21788
rect 2778 21728 2842 21732
rect 2858 21788 2922 21792
rect 2858 21732 2862 21788
rect 2862 21732 2918 21788
rect 2918 21732 2922 21788
rect 2858 21728 2922 21732
rect 5952 21788 6016 21792
rect 5952 21732 5956 21788
rect 5956 21732 6012 21788
rect 6012 21732 6016 21788
rect 5952 21728 6016 21732
rect 6032 21788 6096 21792
rect 6032 21732 6036 21788
rect 6036 21732 6092 21788
rect 6092 21732 6096 21788
rect 6032 21728 6096 21732
rect 6112 21788 6176 21792
rect 6112 21732 6116 21788
rect 6116 21732 6172 21788
rect 6172 21732 6176 21788
rect 6112 21728 6176 21732
rect 6192 21788 6256 21792
rect 6192 21732 6196 21788
rect 6196 21732 6252 21788
rect 6252 21732 6256 21788
rect 6192 21728 6256 21732
rect 4285 21244 4349 21248
rect 4285 21188 4289 21244
rect 4289 21188 4345 21244
rect 4345 21188 4349 21244
rect 4285 21184 4349 21188
rect 4365 21244 4429 21248
rect 4365 21188 4369 21244
rect 4369 21188 4425 21244
rect 4425 21188 4429 21244
rect 4365 21184 4429 21188
rect 4445 21244 4509 21248
rect 4445 21188 4449 21244
rect 4449 21188 4505 21244
rect 4505 21188 4509 21244
rect 4445 21184 4509 21188
rect 4525 21244 4589 21248
rect 4525 21188 4529 21244
rect 4529 21188 4585 21244
rect 4585 21188 4589 21244
rect 4525 21184 4589 21188
rect 7618 21244 7682 21248
rect 7618 21188 7622 21244
rect 7622 21188 7678 21244
rect 7678 21188 7682 21244
rect 7618 21184 7682 21188
rect 7698 21244 7762 21248
rect 7698 21188 7702 21244
rect 7702 21188 7758 21244
rect 7758 21188 7762 21244
rect 7698 21184 7762 21188
rect 7778 21244 7842 21248
rect 7778 21188 7782 21244
rect 7782 21188 7838 21244
rect 7838 21188 7842 21244
rect 7778 21184 7842 21188
rect 7858 21244 7922 21248
rect 7858 21188 7862 21244
rect 7862 21188 7918 21244
rect 7918 21188 7922 21244
rect 7858 21184 7922 21188
rect 2618 20700 2682 20704
rect 2618 20644 2622 20700
rect 2622 20644 2678 20700
rect 2678 20644 2682 20700
rect 2618 20640 2682 20644
rect 2698 20700 2762 20704
rect 2698 20644 2702 20700
rect 2702 20644 2758 20700
rect 2758 20644 2762 20700
rect 2698 20640 2762 20644
rect 2778 20700 2842 20704
rect 2778 20644 2782 20700
rect 2782 20644 2838 20700
rect 2838 20644 2842 20700
rect 2778 20640 2842 20644
rect 2858 20700 2922 20704
rect 2858 20644 2862 20700
rect 2862 20644 2918 20700
rect 2918 20644 2922 20700
rect 2858 20640 2922 20644
rect 5952 20700 6016 20704
rect 5952 20644 5956 20700
rect 5956 20644 6012 20700
rect 6012 20644 6016 20700
rect 5952 20640 6016 20644
rect 6032 20700 6096 20704
rect 6032 20644 6036 20700
rect 6036 20644 6092 20700
rect 6092 20644 6096 20700
rect 6032 20640 6096 20644
rect 6112 20700 6176 20704
rect 6112 20644 6116 20700
rect 6116 20644 6172 20700
rect 6172 20644 6176 20700
rect 6112 20640 6176 20644
rect 6192 20700 6256 20704
rect 6192 20644 6196 20700
rect 6196 20644 6252 20700
rect 6252 20644 6256 20700
rect 6192 20640 6256 20644
rect 4285 20156 4349 20160
rect 4285 20100 4289 20156
rect 4289 20100 4345 20156
rect 4345 20100 4349 20156
rect 4285 20096 4349 20100
rect 4365 20156 4429 20160
rect 4365 20100 4369 20156
rect 4369 20100 4425 20156
rect 4425 20100 4429 20156
rect 4365 20096 4429 20100
rect 4445 20156 4509 20160
rect 4445 20100 4449 20156
rect 4449 20100 4505 20156
rect 4505 20100 4509 20156
rect 4445 20096 4509 20100
rect 4525 20156 4589 20160
rect 4525 20100 4529 20156
rect 4529 20100 4585 20156
rect 4585 20100 4589 20156
rect 4525 20096 4589 20100
rect 7618 20156 7682 20160
rect 7618 20100 7622 20156
rect 7622 20100 7678 20156
rect 7678 20100 7682 20156
rect 7618 20096 7682 20100
rect 7698 20156 7762 20160
rect 7698 20100 7702 20156
rect 7702 20100 7758 20156
rect 7758 20100 7762 20156
rect 7698 20096 7762 20100
rect 7778 20156 7842 20160
rect 7778 20100 7782 20156
rect 7782 20100 7838 20156
rect 7838 20100 7842 20156
rect 7778 20096 7842 20100
rect 7858 20156 7922 20160
rect 7858 20100 7862 20156
rect 7862 20100 7918 20156
rect 7918 20100 7922 20156
rect 7858 20096 7922 20100
rect 2618 19612 2682 19616
rect 2618 19556 2622 19612
rect 2622 19556 2678 19612
rect 2678 19556 2682 19612
rect 2618 19552 2682 19556
rect 2698 19612 2762 19616
rect 2698 19556 2702 19612
rect 2702 19556 2758 19612
rect 2758 19556 2762 19612
rect 2698 19552 2762 19556
rect 2778 19612 2842 19616
rect 2778 19556 2782 19612
rect 2782 19556 2838 19612
rect 2838 19556 2842 19612
rect 2778 19552 2842 19556
rect 2858 19612 2922 19616
rect 2858 19556 2862 19612
rect 2862 19556 2918 19612
rect 2918 19556 2922 19612
rect 2858 19552 2922 19556
rect 5952 19612 6016 19616
rect 5952 19556 5956 19612
rect 5956 19556 6012 19612
rect 6012 19556 6016 19612
rect 5952 19552 6016 19556
rect 6032 19612 6096 19616
rect 6032 19556 6036 19612
rect 6036 19556 6092 19612
rect 6092 19556 6096 19612
rect 6032 19552 6096 19556
rect 6112 19612 6176 19616
rect 6112 19556 6116 19612
rect 6116 19556 6172 19612
rect 6172 19556 6176 19612
rect 6112 19552 6176 19556
rect 6192 19612 6256 19616
rect 6192 19556 6196 19612
rect 6196 19556 6252 19612
rect 6252 19556 6256 19612
rect 6192 19552 6256 19556
rect 4285 19068 4349 19072
rect 4285 19012 4289 19068
rect 4289 19012 4345 19068
rect 4345 19012 4349 19068
rect 4285 19008 4349 19012
rect 4365 19068 4429 19072
rect 4365 19012 4369 19068
rect 4369 19012 4425 19068
rect 4425 19012 4429 19068
rect 4365 19008 4429 19012
rect 4445 19068 4509 19072
rect 4445 19012 4449 19068
rect 4449 19012 4505 19068
rect 4505 19012 4509 19068
rect 4445 19008 4509 19012
rect 4525 19068 4589 19072
rect 4525 19012 4529 19068
rect 4529 19012 4585 19068
rect 4585 19012 4589 19068
rect 4525 19008 4589 19012
rect 7618 19068 7682 19072
rect 7618 19012 7622 19068
rect 7622 19012 7678 19068
rect 7678 19012 7682 19068
rect 7618 19008 7682 19012
rect 7698 19068 7762 19072
rect 7698 19012 7702 19068
rect 7702 19012 7758 19068
rect 7758 19012 7762 19068
rect 7698 19008 7762 19012
rect 7778 19068 7842 19072
rect 7778 19012 7782 19068
rect 7782 19012 7838 19068
rect 7838 19012 7842 19068
rect 7778 19008 7842 19012
rect 7858 19068 7922 19072
rect 7858 19012 7862 19068
rect 7862 19012 7918 19068
rect 7918 19012 7922 19068
rect 7858 19008 7922 19012
rect 2618 18524 2682 18528
rect 2618 18468 2622 18524
rect 2622 18468 2678 18524
rect 2678 18468 2682 18524
rect 2618 18464 2682 18468
rect 2698 18524 2762 18528
rect 2698 18468 2702 18524
rect 2702 18468 2758 18524
rect 2758 18468 2762 18524
rect 2698 18464 2762 18468
rect 2778 18524 2842 18528
rect 2778 18468 2782 18524
rect 2782 18468 2838 18524
rect 2838 18468 2842 18524
rect 2778 18464 2842 18468
rect 2858 18524 2922 18528
rect 2858 18468 2862 18524
rect 2862 18468 2918 18524
rect 2918 18468 2922 18524
rect 2858 18464 2922 18468
rect 5952 18524 6016 18528
rect 5952 18468 5956 18524
rect 5956 18468 6012 18524
rect 6012 18468 6016 18524
rect 5952 18464 6016 18468
rect 6032 18524 6096 18528
rect 6032 18468 6036 18524
rect 6036 18468 6092 18524
rect 6092 18468 6096 18524
rect 6032 18464 6096 18468
rect 6112 18524 6176 18528
rect 6112 18468 6116 18524
rect 6116 18468 6172 18524
rect 6172 18468 6176 18524
rect 6112 18464 6176 18468
rect 6192 18524 6256 18528
rect 6192 18468 6196 18524
rect 6196 18468 6252 18524
rect 6252 18468 6256 18524
rect 6192 18464 6256 18468
rect 4285 17980 4349 17984
rect 4285 17924 4289 17980
rect 4289 17924 4345 17980
rect 4345 17924 4349 17980
rect 4285 17920 4349 17924
rect 4365 17980 4429 17984
rect 4365 17924 4369 17980
rect 4369 17924 4425 17980
rect 4425 17924 4429 17980
rect 4365 17920 4429 17924
rect 4445 17980 4509 17984
rect 4445 17924 4449 17980
rect 4449 17924 4505 17980
rect 4505 17924 4509 17980
rect 4445 17920 4509 17924
rect 4525 17980 4589 17984
rect 4525 17924 4529 17980
rect 4529 17924 4585 17980
rect 4585 17924 4589 17980
rect 4525 17920 4589 17924
rect 7618 17980 7682 17984
rect 7618 17924 7622 17980
rect 7622 17924 7678 17980
rect 7678 17924 7682 17980
rect 7618 17920 7682 17924
rect 7698 17980 7762 17984
rect 7698 17924 7702 17980
rect 7702 17924 7758 17980
rect 7758 17924 7762 17980
rect 7698 17920 7762 17924
rect 7778 17980 7842 17984
rect 7778 17924 7782 17980
rect 7782 17924 7838 17980
rect 7838 17924 7842 17980
rect 7778 17920 7842 17924
rect 7858 17980 7922 17984
rect 7858 17924 7862 17980
rect 7862 17924 7918 17980
rect 7918 17924 7922 17980
rect 7858 17920 7922 17924
rect 2618 17436 2682 17440
rect 2618 17380 2622 17436
rect 2622 17380 2678 17436
rect 2678 17380 2682 17436
rect 2618 17376 2682 17380
rect 2698 17436 2762 17440
rect 2698 17380 2702 17436
rect 2702 17380 2758 17436
rect 2758 17380 2762 17436
rect 2698 17376 2762 17380
rect 2778 17436 2842 17440
rect 2778 17380 2782 17436
rect 2782 17380 2838 17436
rect 2838 17380 2842 17436
rect 2778 17376 2842 17380
rect 2858 17436 2922 17440
rect 2858 17380 2862 17436
rect 2862 17380 2918 17436
rect 2918 17380 2922 17436
rect 2858 17376 2922 17380
rect 5952 17436 6016 17440
rect 5952 17380 5956 17436
rect 5956 17380 6012 17436
rect 6012 17380 6016 17436
rect 5952 17376 6016 17380
rect 6032 17436 6096 17440
rect 6032 17380 6036 17436
rect 6036 17380 6092 17436
rect 6092 17380 6096 17436
rect 6032 17376 6096 17380
rect 6112 17436 6176 17440
rect 6112 17380 6116 17436
rect 6116 17380 6172 17436
rect 6172 17380 6176 17436
rect 6112 17376 6176 17380
rect 6192 17436 6256 17440
rect 6192 17380 6196 17436
rect 6196 17380 6252 17436
rect 6252 17380 6256 17436
rect 6192 17376 6256 17380
rect 4285 16892 4349 16896
rect 4285 16836 4289 16892
rect 4289 16836 4345 16892
rect 4345 16836 4349 16892
rect 4285 16832 4349 16836
rect 4365 16892 4429 16896
rect 4365 16836 4369 16892
rect 4369 16836 4425 16892
rect 4425 16836 4429 16892
rect 4365 16832 4429 16836
rect 4445 16892 4509 16896
rect 4445 16836 4449 16892
rect 4449 16836 4505 16892
rect 4505 16836 4509 16892
rect 4445 16832 4509 16836
rect 4525 16892 4589 16896
rect 4525 16836 4529 16892
rect 4529 16836 4585 16892
rect 4585 16836 4589 16892
rect 4525 16832 4589 16836
rect 7618 16892 7682 16896
rect 7618 16836 7622 16892
rect 7622 16836 7678 16892
rect 7678 16836 7682 16892
rect 7618 16832 7682 16836
rect 7698 16892 7762 16896
rect 7698 16836 7702 16892
rect 7702 16836 7758 16892
rect 7758 16836 7762 16892
rect 7698 16832 7762 16836
rect 7778 16892 7842 16896
rect 7778 16836 7782 16892
rect 7782 16836 7838 16892
rect 7838 16836 7842 16892
rect 7778 16832 7842 16836
rect 7858 16892 7922 16896
rect 7858 16836 7862 16892
rect 7862 16836 7918 16892
rect 7918 16836 7922 16892
rect 7858 16832 7922 16836
rect 2618 16348 2682 16352
rect 2618 16292 2622 16348
rect 2622 16292 2678 16348
rect 2678 16292 2682 16348
rect 2618 16288 2682 16292
rect 2698 16348 2762 16352
rect 2698 16292 2702 16348
rect 2702 16292 2758 16348
rect 2758 16292 2762 16348
rect 2698 16288 2762 16292
rect 2778 16348 2842 16352
rect 2778 16292 2782 16348
rect 2782 16292 2838 16348
rect 2838 16292 2842 16348
rect 2778 16288 2842 16292
rect 2858 16348 2922 16352
rect 2858 16292 2862 16348
rect 2862 16292 2918 16348
rect 2918 16292 2922 16348
rect 2858 16288 2922 16292
rect 5952 16348 6016 16352
rect 5952 16292 5956 16348
rect 5956 16292 6012 16348
rect 6012 16292 6016 16348
rect 5952 16288 6016 16292
rect 6032 16348 6096 16352
rect 6032 16292 6036 16348
rect 6036 16292 6092 16348
rect 6092 16292 6096 16348
rect 6032 16288 6096 16292
rect 6112 16348 6176 16352
rect 6112 16292 6116 16348
rect 6116 16292 6172 16348
rect 6172 16292 6176 16348
rect 6112 16288 6176 16292
rect 6192 16348 6256 16352
rect 6192 16292 6196 16348
rect 6196 16292 6252 16348
rect 6252 16292 6256 16348
rect 6192 16288 6256 16292
rect 4285 15804 4349 15808
rect 4285 15748 4289 15804
rect 4289 15748 4345 15804
rect 4345 15748 4349 15804
rect 4285 15744 4349 15748
rect 4365 15804 4429 15808
rect 4365 15748 4369 15804
rect 4369 15748 4425 15804
rect 4425 15748 4429 15804
rect 4365 15744 4429 15748
rect 4445 15804 4509 15808
rect 4445 15748 4449 15804
rect 4449 15748 4505 15804
rect 4505 15748 4509 15804
rect 4445 15744 4509 15748
rect 4525 15804 4589 15808
rect 4525 15748 4529 15804
rect 4529 15748 4585 15804
rect 4585 15748 4589 15804
rect 4525 15744 4589 15748
rect 7618 15804 7682 15808
rect 7618 15748 7622 15804
rect 7622 15748 7678 15804
rect 7678 15748 7682 15804
rect 7618 15744 7682 15748
rect 7698 15804 7762 15808
rect 7698 15748 7702 15804
rect 7702 15748 7758 15804
rect 7758 15748 7762 15804
rect 7698 15744 7762 15748
rect 7778 15804 7842 15808
rect 7778 15748 7782 15804
rect 7782 15748 7838 15804
rect 7838 15748 7842 15804
rect 7778 15744 7842 15748
rect 7858 15804 7922 15808
rect 7858 15748 7862 15804
rect 7862 15748 7918 15804
rect 7918 15748 7922 15804
rect 7858 15744 7922 15748
rect 2618 15260 2682 15264
rect 2618 15204 2622 15260
rect 2622 15204 2678 15260
rect 2678 15204 2682 15260
rect 2618 15200 2682 15204
rect 2698 15260 2762 15264
rect 2698 15204 2702 15260
rect 2702 15204 2758 15260
rect 2758 15204 2762 15260
rect 2698 15200 2762 15204
rect 2778 15260 2842 15264
rect 2778 15204 2782 15260
rect 2782 15204 2838 15260
rect 2838 15204 2842 15260
rect 2778 15200 2842 15204
rect 2858 15260 2922 15264
rect 2858 15204 2862 15260
rect 2862 15204 2918 15260
rect 2918 15204 2922 15260
rect 2858 15200 2922 15204
rect 5952 15260 6016 15264
rect 5952 15204 5956 15260
rect 5956 15204 6012 15260
rect 6012 15204 6016 15260
rect 5952 15200 6016 15204
rect 6032 15260 6096 15264
rect 6032 15204 6036 15260
rect 6036 15204 6092 15260
rect 6092 15204 6096 15260
rect 6032 15200 6096 15204
rect 6112 15260 6176 15264
rect 6112 15204 6116 15260
rect 6116 15204 6172 15260
rect 6172 15204 6176 15260
rect 6112 15200 6176 15204
rect 6192 15260 6256 15264
rect 6192 15204 6196 15260
rect 6196 15204 6252 15260
rect 6252 15204 6256 15260
rect 6192 15200 6256 15204
rect 4285 14716 4349 14720
rect 4285 14660 4289 14716
rect 4289 14660 4345 14716
rect 4345 14660 4349 14716
rect 4285 14656 4349 14660
rect 4365 14716 4429 14720
rect 4365 14660 4369 14716
rect 4369 14660 4425 14716
rect 4425 14660 4429 14716
rect 4365 14656 4429 14660
rect 4445 14716 4509 14720
rect 4445 14660 4449 14716
rect 4449 14660 4505 14716
rect 4505 14660 4509 14716
rect 4445 14656 4509 14660
rect 4525 14716 4589 14720
rect 4525 14660 4529 14716
rect 4529 14660 4585 14716
rect 4585 14660 4589 14716
rect 4525 14656 4589 14660
rect 7618 14716 7682 14720
rect 7618 14660 7622 14716
rect 7622 14660 7678 14716
rect 7678 14660 7682 14716
rect 7618 14656 7682 14660
rect 7698 14716 7762 14720
rect 7698 14660 7702 14716
rect 7702 14660 7758 14716
rect 7758 14660 7762 14716
rect 7698 14656 7762 14660
rect 7778 14716 7842 14720
rect 7778 14660 7782 14716
rect 7782 14660 7838 14716
rect 7838 14660 7842 14716
rect 7778 14656 7842 14660
rect 7858 14716 7922 14720
rect 7858 14660 7862 14716
rect 7862 14660 7918 14716
rect 7918 14660 7922 14716
rect 7858 14656 7922 14660
rect 2618 14172 2682 14176
rect 2618 14116 2622 14172
rect 2622 14116 2678 14172
rect 2678 14116 2682 14172
rect 2618 14112 2682 14116
rect 2698 14172 2762 14176
rect 2698 14116 2702 14172
rect 2702 14116 2758 14172
rect 2758 14116 2762 14172
rect 2698 14112 2762 14116
rect 2778 14172 2842 14176
rect 2778 14116 2782 14172
rect 2782 14116 2838 14172
rect 2838 14116 2842 14172
rect 2778 14112 2842 14116
rect 2858 14172 2922 14176
rect 2858 14116 2862 14172
rect 2862 14116 2918 14172
rect 2918 14116 2922 14172
rect 2858 14112 2922 14116
rect 5952 14172 6016 14176
rect 5952 14116 5956 14172
rect 5956 14116 6012 14172
rect 6012 14116 6016 14172
rect 5952 14112 6016 14116
rect 6032 14172 6096 14176
rect 6032 14116 6036 14172
rect 6036 14116 6092 14172
rect 6092 14116 6096 14172
rect 6032 14112 6096 14116
rect 6112 14172 6176 14176
rect 6112 14116 6116 14172
rect 6116 14116 6172 14172
rect 6172 14116 6176 14172
rect 6112 14112 6176 14116
rect 6192 14172 6256 14176
rect 6192 14116 6196 14172
rect 6196 14116 6252 14172
rect 6252 14116 6256 14172
rect 6192 14112 6256 14116
rect 4285 13628 4349 13632
rect 4285 13572 4289 13628
rect 4289 13572 4345 13628
rect 4345 13572 4349 13628
rect 4285 13568 4349 13572
rect 4365 13628 4429 13632
rect 4365 13572 4369 13628
rect 4369 13572 4425 13628
rect 4425 13572 4429 13628
rect 4365 13568 4429 13572
rect 4445 13628 4509 13632
rect 4445 13572 4449 13628
rect 4449 13572 4505 13628
rect 4505 13572 4509 13628
rect 4445 13568 4509 13572
rect 4525 13628 4589 13632
rect 4525 13572 4529 13628
rect 4529 13572 4585 13628
rect 4585 13572 4589 13628
rect 4525 13568 4589 13572
rect 7618 13628 7682 13632
rect 7618 13572 7622 13628
rect 7622 13572 7678 13628
rect 7678 13572 7682 13628
rect 7618 13568 7682 13572
rect 7698 13628 7762 13632
rect 7698 13572 7702 13628
rect 7702 13572 7758 13628
rect 7758 13572 7762 13628
rect 7698 13568 7762 13572
rect 7778 13628 7842 13632
rect 7778 13572 7782 13628
rect 7782 13572 7838 13628
rect 7838 13572 7842 13628
rect 7778 13568 7842 13572
rect 7858 13628 7922 13632
rect 7858 13572 7862 13628
rect 7862 13572 7918 13628
rect 7918 13572 7922 13628
rect 7858 13568 7922 13572
rect 2618 13084 2682 13088
rect 2618 13028 2622 13084
rect 2622 13028 2678 13084
rect 2678 13028 2682 13084
rect 2618 13024 2682 13028
rect 2698 13084 2762 13088
rect 2698 13028 2702 13084
rect 2702 13028 2758 13084
rect 2758 13028 2762 13084
rect 2698 13024 2762 13028
rect 2778 13084 2842 13088
rect 2778 13028 2782 13084
rect 2782 13028 2838 13084
rect 2838 13028 2842 13084
rect 2778 13024 2842 13028
rect 2858 13084 2922 13088
rect 2858 13028 2862 13084
rect 2862 13028 2918 13084
rect 2918 13028 2922 13084
rect 2858 13024 2922 13028
rect 5952 13084 6016 13088
rect 5952 13028 5956 13084
rect 5956 13028 6012 13084
rect 6012 13028 6016 13084
rect 5952 13024 6016 13028
rect 6032 13084 6096 13088
rect 6032 13028 6036 13084
rect 6036 13028 6092 13084
rect 6092 13028 6096 13084
rect 6032 13024 6096 13028
rect 6112 13084 6176 13088
rect 6112 13028 6116 13084
rect 6116 13028 6172 13084
rect 6172 13028 6176 13084
rect 6112 13024 6176 13028
rect 6192 13084 6256 13088
rect 6192 13028 6196 13084
rect 6196 13028 6252 13084
rect 6252 13028 6256 13084
rect 6192 13024 6256 13028
rect 4285 12540 4349 12544
rect 4285 12484 4289 12540
rect 4289 12484 4345 12540
rect 4345 12484 4349 12540
rect 4285 12480 4349 12484
rect 4365 12540 4429 12544
rect 4365 12484 4369 12540
rect 4369 12484 4425 12540
rect 4425 12484 4429 12540
rect 4365 12480 4429 12484
rect 4445 12540 4509 12544
rect 4445 12484 4449 12540
rect 4449 12484 4505 12540
rect 4505 12484 4509 12540
rect 4445 12480 4509 12484
rect 4525 12540 4589 12544
rect 4525 12484 4529 12540
rect 4529 12484 4585 12540
rect 4585 12484 4589 12540
rect 4525 12480 4589 12484
rect 7618 12540 7682 12544
rect 7618 12484 7622 12540
rect 7622 12484 7678 12540
rect 7678 12484 7682 12540
rect 7618 12480 7682 12484
rect 7698 12540 7762 12544
rect 7698 12484 7702 12540
rect 7702 12484 7758 12540
rect 7758 12484 7762 12540
rect 7698 12480 7762 12484
rect 7778 12540 7842 12544
rect 7778 12484 7782 12540
rect 7782 12484 7838 12540
rect 7838 12484 7842 12540
rect 7778 12480 7842 12484
rect 7858 12540 7922 12544
rect 7858 12484 7862 12540
rect 7862 12484 7918 12540
rect 7918 12484 7922 12540
rect 7858 12480 7922 12484
rect 2618 11996 2682 12000
rect 2618 11940 2622 11996
rect 2622 11940 2678 11996
rect 2678 11940 2682 11996
rect 2618 11936 2682 11940
rect 2698 11996 2762 12000
rect 2698 11940 2702 11996
rect 2702 11940 2758 11996
rect 2758 11940 2762 11996
rect 2698 11936 2762 11940
rect 2778 11996 2842 12000
rect 2778 11940 2782 11996
rect 2782 11940 2838 11996
rect 2838 11940 2842 11996
rect 2778 11936 2842 11940
rect 2858 11996 2922 12000
rect 2858 11940 2862 11996
rect 2862 11940 2918 11996
rect 2918 11940 2922 11996
rect 2858 11936 2922 11940
rect 5952 11996 6016 12000
rect 5952 11940 5956 11996
rect 5956 11940 6012 11996
rect 6012 11940 6016 11996
rect 5952 11936 6016 11940
rect 6032 11996 6096 12000
rect 6032 11940 6036 11996
rect 6036 11940 6092 11996
rect 6092 11940 6096 11996
rect 6032 11936 6096 11940
rect 6112 11996 6176 12000
rect 6112 11940 6116 11996
rect 6116 11940 6172 11996
rect 6172 11940 6176 11996
rect 6112 11936 6176 11940
rect 6192 11996 6256 12000
rect 6192 11940 6196 11996
rect 6196 11940 6252 11996
rect 6252 11940 6256 11996
rect 6192 11936 6256 11940
rect 4285 11452 4349 11456
rect 4285 11396 4289 11452
rect 4289 11396 4345 11452
rect 4345 11396 4349 11452
rect 4285 11392 4349 11396
rect 4365 11452 4429 11456
rect 4365 11396 4369 11452
rect 4369 11396 4425 11452
rect 4425 11396 4429 11452
rect 4365 11392 4429 11396
rect 4445 11452 4509 11456
rect 4445 11396 4449 11452
rect 4449 11396 4505 11452
rect 4505 11396 4509 11452
rect 4445 11392 4509 11396
rect 4525 11452 4589 11456
rect 4525 11396 4529 11452
rect 4529 11396 4585 11452
rect 4585 11396 4589 11452
rect 4525 11392 4589 11396
rect 7618 11452 7682 11456
rect 7618 11396 7622 11452
rect 7622 11396 7678 11452
rect 7678 11396 7682 11452
rect 7618 11392 7682 11396
rect 7698 11452 7762 11456
rect 7698 11396 7702 11452
rect 7702 11396 7758 11452
rect 7758 11396 7762 11452
rect 7698 11392 7762 11396
rect 7778 11452 7842 11456
rect 7778 11396 7782 11452
rect 7782 11396 7838 11452
rect 7838 11396 7842 11452
rect 7778 11392 7842 11396
rect 7858 11452 7922 11456
rect 7858 11396 7862 11452
rect 7862 11396 7918 11452
rect 7918 11396 7922 11452
rect 7858 11392 7922 11396
rect 2618 10908 2682 10912
rect 2618 10852 2622 10908
rect 2622 10852 2678 10908
rect 2678 10852 2682 10908
rect 2618 10848 2682 10852
rect 2698 10908 2762 10912
rect 2698 10852 2702 10908
rect 2702 10852 2758 10908
rect 2758 10852 2762 10908
rect 2698 10848 2762 10852
rect 2778 10908 2842 10912
rect 2778 10852 2782 10908
rect 2782 10852 2838 10908
rect 2838 10852 2842 10908
rect 2778 10848 2842 10852
rect 2858 10908 2922 10912
rect 2858 10852 2862 10908
rect 2862 10852 2918 10908
rect 2918 10852 2922 10908
rect 2858 10848 2922 10852
rect 5952 10908 6016 10912
rect 5952 10852 5956 10908
rect 5956 10852 6012 10908
rect 6012 10852 6016 10908
rect 5952 10848 6016 10852
rect 6032 10908 6096 10912
rect 6032 10852 6036 10908
rect 6036 10852 6092 10908
rect 6092 10852 6096 10908
rect 6032 10848 6096 10852
rect 6112 10908 6176 10912
rect 6112 10852 6116 10908
rect 6116 10852 6172 10908
rect 6172 10852 6176 10908
rect 6112 10848 6176 10852
rect 6192 10908 6256 10912
rect 6192 10852 6196 10908
rect 6196 10852 6252 10908
rect 6252 10852 6256 10908
rect 6192 10848 6256 10852
rect 4285 10364 4349 10368
rect 4285 10308 4289 10364
rect 4289 10308 4345 10364
rect 4345 10308 4349 10364
rect 4285 10304 4349 10308
rect 4365 10364 4429 10368
rect 4365 10308 4369 10364
rect 4369 10308 4425 10364
rect 4425 10308 4429 10364
rect 4365 10304 4429 10308
rect 4445 10364 4509 10368
rect 4445 10308 4449 10364
rect 4449 10308 4505 10364
rect 4505 10308 4509 10364
rect 4445 10304 4509 10308
rect 4525 10364 4589 10368
rect 4525 10308 4529 10364
rect 4529 10308 4585 10364
rect 4585 10308 4589 10364
rect 4525 10304 4589 10308
rect 7618 10364 7682 10368
rect 7618 10308 7622 10364
rect 7622 10308 7678 10364
rect 7678 10308 7682 10364
rect 7618 10304 7682 10308
rect 7698 10364 7762 10368
rect 7698 10308 7702 10364
rect 7702 10308 7758 10364
rect 7758 10308 7762 10364
rect 7698 10304 7762 10308
rect 7778 10364 7842 10368
rect 7778 10308 7782 10364
rect 7782 10308 7838 10364
rect 7838 10308 7842 10364
rect 7778 10304 7842 10308
rect 7858 10364 7922 10368
rect 7858 10308 7862 10364
rect 7862 10308 7918 10364
rect 7918 10308 7922 10364
rect 7858 10304 7922 10308
rect 2618 9820 2682 9824
rect 2618 9764 2622 9820
rect 2622 9764 2678 9820
rect 2678 9764 2682 9820
rect 2618 9760 2682 9764
rect 2698 9820 2762 9824
rect 2698 9764 2702 9820
rect 2702 9764 2758 9820
rect 2758 9764 2762 9820
rect 2698 9760 2762 9764
rect 2778 9820 2842 9824
rect 2778 9764 2782 9820
rect 2782 9764 2838 9820
rect 2838 9764 2842 9820
rect 2778 9760 2842 9764
rect 2858 9820 2922 9824
rect 2858 9764 2862 9820
rect 2862 9764 2918 9820
rect 2918 9764 2922 9820
rect 2858 9760 2922 9764
rect 5952 9820 6016 9824
rect 5952 9764 5956 9820
rect 5956 9764 6012 9820
rect 6012 9764 6016 9820
rect 5952 9760 6016 9764
rect 6032 9820 6096 9824
rect 6032 9764 6036 9820
rect 6036 9764 6092 9820
rect 6092 9764 6096 9820
rect 6032 9760 6096 9764
rect 6112 9820 6176 9824
rect 6112 9764 6116 9820
rect 6116 9764 6172 9820
rect 6172 9764 6176 9820
rect 6112 9760 6176 9764
rect 6192 9820 6256 9824
rect 6192 9764 6196 9820
rect 6196 9764 6252 9820
rect 6252 9764 6256 9820
rect 6192 9760 6256 9764
rect 4285 9276 4349 9280
rect 4285 9220 4289 9276
rect 4289 9220 4345 9276
rect 4345 9220 4349 9276
rect 4285 9216 4349 9220
rect 4365 9276 4429 9280
rect 4365 9220 4369 9276
rect 4369 9220 4425 9276
rect 4425 9220 4429 9276
rect 4365 9216 4429 9220
rect 4445 9276 4509 9280
rect 4445 9220 4449 9276
rect 4449 9220 4505 9276
rect 4505 9220 4509 9276
rect 4445 9216 4509 9220
rect 4525 9276 4589 9280
rect 4525 9220 4529 9276
rect 4529 9220 4585 9276
rect 4585 9220 4589 9276
rect 4525 9216 4589 9220
rect 7618 9276 7682 9280
rect 7618 9220 7622 9276
rect 7622 9220 7678 9276
rect 7678 9220 7682 9276
rect 7618 9216 7682 9220
rect 7698 9276 7762 9280
rect 7698 9220 7702 9276
rect 7702 9220 7758 9276
rect 7758 9220 7762 9276
rect 7698 9216 7762 9220
rect 7778 9276 7842 9280
rect 7778 9220 7782 9276
rect 7782 9220 7838 9276
rect 7838 9220 7842 9276
rect 7778 9216 7842 9220
rect 7858 9276 7922 9280
rect 7858 9220 7862 9276
rect 7862 9220 7918 9276
rect 7918 9220 7922 9276
rect 7858 9216 7922 9220
rect 2618 8732 2682 8736
rect 2618 8676 2622 8732
rect 2622 8676 2678 8732
rect 2678 8676 2682 8732
rect 2618 8672 2682 8676
rect 2698 8732 2762 8736
rect 2698 8676 2702 8732
rect 2702 8676 2758 8732
rect 2758 8676 2762 8732
rect 2698 8672 2762 8676
rect 2778 8732 2842 8736
rect 2778 8676 2782 8732
rect 2782 8676 2838 8732
rect 2838 8676 2842 8732
rect 2778 8672 2842 8676
rect 2858 8732 2922 8736
rect 2858 8676 2862 8732
rect 2862 8676 2918 8732
rect 2918 8676 2922 8732
rect 2858 8672 2922 8676
rect 5952 8732 6016 8736
rect 5952 8676 5956 8732
rect 5956 8676 6012 8732
rect 6012 8676 6016 8732
rect 5952 8672 6016 8676
rect 6032 8732 6096 8736
rect 6032 8676 6036 8732
rect 6036 8676 6092 8732
rect 6092 8676 6096 8732
rect 6032 8672 6096 8676
rect 6112 8732 6176 8736
rect 6112 8676 6116 8732
rect 6116 8676 6172 8732
rect 6172 8676 6176 8732
rect 6112 8672 6176 8676
rect 6192 8732 6256 8736
rect 6192 8676 6196 8732
rect 6196 8676 6252 8732
rect 6252 8676 6256 8732
rect 6192 8672 6256 8676
rect 4285 8188 4349 8192
rect 4285 8132 4289 8188
rect 4289 8132 4345 8188
rect 4345 8132 4349 8188
rect 4285 8128 4349 8132
rect 4365 8188 4429 8192
rect 4365 8132 4369 8188
rect 4369 8132 4425 8188
rect 4425 8132 4429 8188
rect 4365 8128 4429 8132
rect 4445 8188 4509 8192
rect 4445 8132 4449 8188
rect 4449 8132 4505 8188
rect 4505 8132 4509 8188
rect 4445 8128 4509 8132
rect 4525 8188 4589 8192
rect 4525 8132 4529 8188
rect 4529 8132 4585 8188
rect 4585 8132 4589 8188
rect 4525 8128 4589 8132
rect 7618 8188 7682 8192
rect 7618 8132 7622 8188
rect 7622 8132 7678 8188
rect 7678 8132 7682 8188
rect 7618 8128 7682 8132
rect 7698 8188 7762 8192
rect 7698 8132 7702 8188
rect 7702 8132 7758 8188
rect 7758 8132 7762 8188
rect 7698 8128 7762 8132
rect 7778 8188 7842 8192
rect 7778 8132 7782 8188
rect 7782 8132 7838 8188
rect 7838 8132 7842 8188
rect 7778 8128 7842 8132
rect 7858 8188 7922 8192
rect 7858 8132 7862 8188
rect 7862 8132 7918 8188
rect 7918 8132 7922 8188
rect 7858 8128 7922 8132
rect 2618 7644 2682 7648
rect 2618 7588 2622 7644
rect 2622 7588 2678 7644
rect 2678 7588 2682 7644
rect 2618 7584 2682 7588
rect 2698 7644 2762 7648
rect 2698 7588 2702 7644
rect 2702 7588 2758 7644
rect 2758 7588 2762 7644
rect 2698 7584 2762 7588
rect 2778 7644 2842 7648
rect 2778 7588 2782 7644
rect 2782 7588 2838 7644
rect 2838 7588 2842 7644
rect 2778 7584 2842 7588
rect 2858 7644 2922 7648
rect 2858 7588 2862 7644
rect 2862 7588 2918 7644
rect 2918 7588 2922 7644
rect 2858 7584 2922 7588
rect 5952 7644 6016 7648
rect 5952 7588 5956 7644
rect 5956 7588 6012 7644
rect 6012 7588 6016 7644
rect 5952 7584 6016 7588
rect 6032 7644 6096 7648
rect 6032 7588 6036 7644
rect 6036 7588 6092 7644
rect 6092 7588 6096 7644
rect 6032 7584 6096 7588
rect 6112 7644 6176 7648
rect 6112 7588 6116 7644
rect 6116 7588 6172 7644
rect 6172 7588 6176 7644
rect 6112 7584 6176 7588
rect 6192 7644 6256 7648
rect 6192 7588 6196 7644
rect 6196 7588 6252 7644
rect 6252 7588 6256 7644
rect 6192 7584 6256 7588
rect 4285 7100 4349 7104
rect 4285 7044 4289 7100
rect 4289 7044 4345 7100
rect 4345 7044 4349 7100
rect 4285 7040 4349 7044
rect 4365 7100 4429 7104
rect 4365 7044 4369 7100
rect 4369 7044 4425 7100
rect 4425 7044 4429 7100
rect 4365 7040 4429 7044
rect 4445 7100 4509 7104
rect 4445 7044 4449 7100
rect 4449 7044 4505 7100
rect 4505 7044 4509 7100
rect 4445 7040 4509 7044
rect 4525 7100 4589 7104
rect 4525 7044 4529 7100
rect 4529 7044 4585 7100
rect 4585 7044 4589 7100
rect 4525 7040 4589 7044
rect 7618 7100 7682 7104
rect 7618 7044 7622 7100
rect 7622 7044 7678 7100
rect 7678 7044 7682 7100
rect 7618 7040 7682 7044
rect 7698 7100 7762 7104
rect 7698 7044 7702 7100
rect 7702 7044 7758 7100
rect 7758 7044 7762 7100
rect 7698 7040 7762 7044
rect 7778 7100 7842 7104
rect 7778 7044 7782 7100
rect 7782 7044 7838 7100
rect 7838 7044 7842 7100
rect 7778 7040 7842 7044
rect 7858 7100 7922 7104
rect 7858 7044 7862 7100
rect 7862 7044 7918 7100
rect 7918 7044 7922 7100
rect 7858 7040 7922 7044
rect 2618 6556 2682 6560
rect 2618 6500 2622 6556
rect 2622 6500 2678 6556
rect 2678 6500 2682 6556
rect 2618 6496 2682 6500
rect 2698 6556 2762 6560
rect 2698 6500 2702 6556
rect 2702 6500 2758 6556
rect 2758 6500 2762 6556
rect 2698 6496 2762 6500
rect 2778 6556 2842 6560
rect 2778 6500 2782 6556
rect 2782 6500 2838 6556
rect 2838 6500 2842 6556
rect 2778 6496 2842 6500
rect 2858 6556 2922 6560
rect 2858 6500 2862 6556
rect 2862 6500 2918 6556
rect 2918 6500 2922 6556
rect 2858 6496 2922 6500
rect 5952 6556 6016 6560
rect 5952 6500 5956 6556
rect 5956 6500 6012 6556
rect 6012 6500 6016 6556
rect 5952 6496 6016 6500
rect 6032 6556 6096 6560
rect 6032 6500 6036 6556
rect 6036 6500 6092 6556
rect 6092 6500 6096 6556
rect 6032 6496 6096 6500
rect 6112 6556 6176 6560
rect 6112 6500 6116 6556
rect 6116 6500 6172 6556
rect 6172 6500 6176 6556
rect 6112 6496 6176 6500
rect 6192 6556 6256 6560
rect 6192 6500 6196 6556
rect 6196 6500 6252 6556
rect 6252 6500 6256 6556
rect 6192 6496 6256 6500
rect 4285 6012 4349 6016
rect 4285 5956 4289 6012
rect 4289 5956 4345 6012
rect 4345 5956 4349 6012
rect 4285 5952 4349 5956
rect 4365 6012 4429 6016
rect 4365 5956 4369 6012
rect 4369 5956 4425 6012
rect 4425 5956 4429 6012
rect 4365 5952 4429 5956
rect 4445 6012 4509 6016
rect 4445 5956 4449 6012
rect 4449 5956 4505 6012
rect 4505 5956 4509 6012
rect 4445 5952 4509 5956
rect 4525 6012 4589 6016
rect 4525 5956 4529 6012
rect 4529 5956 4585 6012
rect 4585 5956 4589 6012
rect 4525 5952 4589 5956
rect 7618 6012 7682 6016
rect 7618 5956 7622 6012
rect 7622 5956 7678 6012
rect 7678 5956 7682 6012
rect 7618 5952 7682 5956
rect 7698 6012 7762 6016
rect 7698 5956 7702 6012
rect 7702 5956 7758 6012
rect 7758 5956 7762 6012
rect 7698 5952 7762 5956
rect 7778 6012 7842 6016
rect 7778 5956 7782 6012
rect 7782 5956 7838 6012
rect 7838 5956 7842 6012
rect 7778 5952 7842 5956
rect 7858 6012 7922 6016
rect 7858 5956 7862 6012
rect 7862 5956 7918 6012
rect 7918 5956 7922 6012
rect 7858 5952 7922 5956
rect 2618 5468 2682 5472
rect 2618 5412 2622 5468
rect 2622 5412 2678 5468
rect 2678 5412 2682 5468
rect 2618 5408 2682 5412
rect 2698 5468 2762 5472
rect 2698 5412 2702 5468
rect 2702 5412 2758 5468
rect 2758 5412 2762 5468
rect 2698 5408 2762 5412
rect 2778 5468 2842 5472
rect 2778 5412 2782 5468
rect 2782 5412 2838 5468
rect 2838 5412 2842 5468
rect 2778 5408 2842 5412
rect 2858 5468 2922 5472
rect 2858 5412 2862 5468
rect 2862 5412 2918 5468
rect 2918 5412 2922 5468
rect 2858 5408 2922 5412
rect 5952 5468 6016 5472
rect 5952 5412 5956 5468
rect 5956 5412 6012 5468
rect 6012 5412 6016 5468
rect 5952 5408 6016 5412
rect 6032 5468 6096 5472
rect 6032 5412 6036 5468
rect 6036 5412 6092 5468
rect 6092 5412 6096 5468
rect 6032 5408 6096 5412
rect 6112 5468 6176 5472
rect 6112 5412 6116 5468
rect 6116 5412 6172 5468
rect 6172 5412 6176 5468
rect 6112 5408 6176 5412
rect 6192 5468 6256 5472
rect 6192 5412 6196 5468
rect 6196 5412 6252 5468
rect 6252 5412 6256 5468
rect 6192 5408 6256 5412
rect 4285 4924 4349 4928
rect 4285 4868 4289 4924
rect 4289 4868 4345 4924
rect 4345 4868 4349 4924
rect 4285 4864 4349 4868
rect 4365 4924 4429 4928
rect 4365 4868 4369 4924
rect 4369 4868 4425 4924
rect 4425 4868 4429 4924
rect 4365 4864 4429 4868
rect 4445 4924 4509 4928
rect 4445 4868 4449 4924
rect 4449 4868 4505 4924
rect 4505 4868 4509 4924
rect 4445 4864 4509 4868
rect 4525 4924 4589 4928
rect 4525 4868 4529 4924
rect 4529 4868 4585 4924
rect 4585 4868 4589 4924
rect 4525 4864 4589 4868
rect 7618 4924 7682 4928
rect 7618 4868 7622 4924
rect 7622 4868 7678 4924
rect 7678 4868 7682 4924
rect 7618 4864 7682 4868
rect 7698 4924 7762 4928
rect 7698 4868 7702 4924
rect 7702 4868 7758 4924
rect 7758 4868 7762 4924
rect 7698 4864 7762 4868
rect 7778 4924 7842 4928
rect 7778 4868 7782 4924
rect 7782 4868 7838 4924
rect 7838 4868 7842 4924
rect 7778 4864 7842 4868
rect 7858 4924 7922 4928
rect 7858 4868 7862 4924
rect 7862 4868 7918 4924
rect 7918 4868 7922 4924
rect 7858 4864 7922 4868
rect 2618 4380 2682 4384
rect 2618 4324 2622 4380
rect 2622 4324 2678 4380
rect 2678 4324 2682 4380
rect 2618 4320 2682 4324
rect 2698 4380 2762 4384
rect 2698 4324 2702 4380
rect 2702 4324 2758 4380
rect 2758 4324 2762 4380
rect 2698 4320 2762 4324
rect 2778 4380 2842 4384
rect 2778 4324 2782 4380
rect 2782 4324 2838 4380
rect 2838 4324 2842 4380
rect 2778 4320 2842 4324
rect 2858 4380 2922 4384
rect 2858 4324 2862 4380
rect 2862 4324 2918 4380
rect 2918 4324 2922 4380
rect 2858 4320 2922 4324
rect 5952 4380 6016 4384
rect 5952 4324 5956 4380
rect 5956 4324 6012 4380
rect 6012 4324 6016 4380
rect 5952 4320 6016 4324
rect 6032 4380 6096 4384
rect 6032 4324 6036 4380
rect 6036 4324 6092 4380
rect 6092 4324 6096 4380
rect 6032 4320 6096 4324
rect 6112 4380 6176 4384
rect 6112 4324 6116 4380
rect 6116 4324 6172 4380
rect 6172 4324 6176 4380
rect 6112 4320 6176 4324
rect 6192 4380 6256 4384
rect 6192 4324 6196 4380
rect 6196 4324 6252 4380
rect 6252 4324 6256 4380
rect 6192 4320 6256 4324
rect 4285 3836 4349 3840
rect 4285 3780 4289 3836
rect 4289 3780 4345 3836
rect 4345 3780 4349 3836
rect 4285 3776 4349 3780
rect 4365 3836 4429 3840
rect 4365 3780 4369 3836
rect 4369 3780 4425 3836
rect 4425 3780 4429 3836
rect 4365 3776 4429 3780
rect 4445 3836 4509 3840
rect 4445 3780 4449 3836
rect 4449 3780 4505 3836
rect 4505 3780 4509 3836
rect 4445 3776 4509 3780
rect 4525 3836 4589 3840
rect 4525 3780 4529 3836
rect 4529 3780 4585 3836
rect 4585 3780 4589 3836
rect 4525 3776 4589 3780
rect 7618 3836 7682 3840
rect 7618 3780 7622 3836
rect 7622 3780 7678 3836
rect 7678 3780 7682 3836
rect 7618 3776 7682 3780
rect 7698 3836 7762 3840
rect 7698 3780 7702 3836
rect 7702 3780 7758 3836
rect 7758 3780 7762 3836
rect 7698 3776 7762 3780
rect 7778 3836 7842 3840
rect 7778 3780 7782 3836
rect 7782 3780 7838 3836
rect 7838 3780 7842 3836
rect 7778 3776 7842 3780
rect 7858 3836 7922 3840
rect 7858 3780 7862 3836
rect 7862 3780 7918 3836
rect 7918 3780 7922 3836
rect 7858 3776 7922 3780
rect 2618 3292 2682 3296
rect 2618 3236 2622 3292
rect 2622 3236 2678 3292
rect 2678 3236 2682 3292
rect 2618 3232 2682 3236
rect 2698 3292 2762 3296
rect 2698 3236 2702 3292
rect 2702 3236 2758 3292
rect 2758 3236 2762 3292
rect 2698 3232 2762 3236
rect 2778 3292 2842 3296
rect 2778 3236 2782 3292
rect 2782 3236 2838 3292
rect 2838 3236 2842 3292
rect 2778 3232 2842 3236
rect 2858 3292 2922 3296
rect 2858 3236 2862 3292
rect 2862 3236 2918 3292
rect 2918 3236 2922 3292
rect 2858 3232 2922 3236
rect 5952 3292 6016 3296
rect 5952 3236 5956 3292
rect 5956 3236 6012 3292
rect 6012 3236 6016 3292
rect 5952 3232 6016 3236
rect 6032 3292 6096 3296
rect 6032 3236 6036 3292
rect 6036 3236 6092 3292
rect 6092 3236 6096 3292
rect 6032 3232 6096 3236
rect 6112 3292 6176 3296
rect 6112 3236 6116 3292
rect 6116 3236 6172 3292
rect 6172 3236 6176 3292
rect 6112 3232 6176 3236
rect 6192 3292 6256 3296
rect 6192 3236 6196 3292
rect 6196 3236 6252 3292
rect 6252 3236 6256 3292
rect 6192 3232 6256 3236
rect 4285 2748 4349 2752
rect 4285 2692 4289 2748
rect 4289 2692 4345 2748
rect 4345 2692 4349 2748
rect 4285 2688 4349 2692
rect 4365 2748 4429 2752
rect 4365 2692 4369 2748
rect 4369 2692 4425 2748
rect 4425 2692 4429 2748
rect 4365 2688 4429 2692
rect 4445 2748 4509 2752
rect 4445 2692 4449 2748
rect 4449 2692 4505 2748
rect 4505 2692 4509 2748
rect 4445 2688 4509 2692
rect 4525 2748 4589 2752
rect 4525 2692 4529 2748
rect 4529 2692 4585 2748
rect 4585 2692 4589 2748
rect 4525 2688 4589 2692
rect 7618 2748 7682 2752
rect 7618 2692 7622 2748
rect 7622 2692 7678 2748
rect 7678 2692 7682 2748
rect 7618 2688 7682 2692
rect 7698 2748 7762 2752
rect 7698 2692 7702 2748
rect 7702 2692 7758 2748
rect 7758 2692 7762 2748
rect 7698 2688 7762 2692
rect 7778 2748 7842 2752
rect 7778 2692 7782 2748
rect 7782 2692 7838 2748
rect 7838 2692 7842 2748
rect 7778 2688 7842 2692
rect 7858 2748 7922 2752
rect 7858 2692 7862 2748
rect 7862 2692 7918 2748
rect 7918 2692 7922 2748
rect 7858 2688 7922 2692
rect 2618 2204 2682 2208
rect 2618 2148 2622 2204
rect 2622 2148 2678 2204
rect 2678 2148 2682 2204
rect 2618 2144 2682 2148
rect 2698 2204 2762 2208
rect 2698 2148 2702 2204
rect 2702 2148 2758 2204
rect 2758 2148 2762 2204
rect 2698 2144 2762 2148
rect 2778 2204 2842 2208
rect 2778 2148 2782 2204
rect 2782 2148 2838 2204
rect 2838 2148 2842 2204
rect 2778 2144 2842 2148
rect 2858 2204 2922 2208
rect 2858 2148 2862 2204
rect 2862 2148 2918 2204
rect 2918 2148 2922 2204
rect 2858 2144 2922 2148
rect 5952 2204 6016 2208
rect 5952 2148 5956 2204
rect 5956 2148 6012 2204
rect 6012 2148 6016 2204
rect 5952 2144 6016 2148
rect 6032 2204 6096 2208
rect 6032 2148 6036 2204
rect 6036 2148 6092 2204
rect 6092 2148 6096 2204
rect 6032 2144 6096 2148
rect 6112 2204 6176 2208
rect 6112 2148 6116 2204
rect 6116 2148 6172 2204
rect 6172 2148 6176 2204
rect 6112 2144 6176 2148
rect 6192 2204 6256 2208
rect 6192 2148 6196 2204
rect 6196 2148 6252 2204
rect 6252 2148 6256 2204
rect 6192 2144 6256 2148
<< metal4 >>
rect 2610 330784 2931 330800
rect 2610 330720 2618 330784
rect 2682 330720 2698 330784
rect 2762 330720 2778 330784
rect 2842 330720 2858 330784
rect 2922 330720 2931 330784
rect 2610 329696 2931 330720
rect 2610 329632 2618 329696
rect 2682 329632 2698 329696
rect 2762 329632 2778 329696
rect 2842 329632 2858 329696
rect 2922 329632 2931 329696
rect 2610 328608 2931 329632
rect 2610 328544 2618 328608
rect 2682 328544 2698 328608
rect 2762 328544 2778 328608
rect 2842 328544 2858 328608
rect 2922 328544 2931 328608
rect 2610 327520 2931 328544
rect 2610 327456 2618 327520
rect 2682 327456 2698 327520
rect 2762 327456 2778 327520
rect 2842 327456 2858 327520
rect 2922 327456 2931 327520
rect 2610 326432 2931 327456
rect 2610 326368 2618 326432
rect 2682 326368 2698 326432
rect 2762 326368 2778 326432
rect 2842 326368 2858 326432
rect 2922 326368 2931 326432
rect 2610 325344 2931 326368
rect 2610 325280 2618 325344
rect 2682 325280 2698 325344
rect 2762 325280 2778 325344
rect 2842 325280 2858 325344
rect 2922 325280 2931 325344
rect 2610 324256 2931 325280
rect 2610 324192 2618 324256
rect 2682 324192 2698 324256
rect 2762 324192 2778 324256
rect 2842 324192 2858 324256
rect 2922 324192 2931 324256
rect 2610 323168 2931 324192
rect 2610 323104 2618 323168
rect 2682 323104 2698 323168
rect 2762 323104 2778 323168
rect 2842 323104 2858 323168
rect 2922 323104 2931 323168
rect 2610 322080 2931 323104
rect 2610 322016 2618 322080
rect 2682 322016 2698 322080
rect 2762 322016 2778 322080
rect 2842 322016 2858 322080
rect 2922 322016 2931 322080
rect 2610 320992 2931 322016
rect 2610 320928 2618 320992
rect 2682 320928 2698 320992
rect 2762 320928 2778 320992
rect 2842 320928 2858 320992
rect 2922 320928 2931 320992
rect 2610 319904 2931 320928
rect 2610 319840 2618 319904
rect 2682 319840 2698 319904
rect 2762 319840 2778 319904
rect 2842 319840 2858 319904
rect 2922 319840 2931 319904
rect 2610 318816 2931 319840
rect 2610 318752 2618 318816
rect 2682 318752 2698 318816
rect 2762 318752 2778 318816
rect 2842 318752 2858 318816
rect 2922 318752 2931 318816
rect 2610 317728 2931 318752
rect 2610 317664 2618 317728
rect 2682 317664 2698 317728
rect 2762 317664 2778 317728
rect 2842 317664 2858 317728
rect 2922 317664 2931 317728
rect 2610 316640 2931 317664
rect 2610 316576 2618 316640
rect 2682 316576 2698 316640
rect 2762 316576 2778 316640
rect 2842 316576 2858 316640
rect 2922 316576 2931 316640
rect 2610 315552 2931 316576
rect 2610 315488 2618 315552
rect 2682 315488 2698 315552
rect 2762 315488 2778 315552
rect 2842 315488 2858 315552
rect 2922 315488 2931 315552
rect 2610 314464 2931 315488
rect 2610 314400 2618 314464
rect 2682 314400 2698 314464
rect 2762 314400 2778 314464
rect 2842 314400 2858 314464
rect 2922 314400 2931 314464
rect 2610 313376 2931 314400
rect 2610 313312 2618 313376
rect 2682 313312 2698 313376
rect 2762 313312 2778 313376
rect 2842 313312 2858 313376
rect 2922 313312 2931 313376
rect 2610 312288 2931 313312
rect 2610 312224 2618 312288
rect 2682 312224 2698 312288
rect 2762 312224 2778 312288
rect 2842 312224 2858 312288
rect 2922 312224 2931 312288
rect 2610 311200 2931 312224
rect 2610 311136 2618 311200
rect 2682 311136 2698 311200
rect 2762 311136 2778 311200
rect 2842 311136 2858 311200
rect 2922 311136 2931 311200
rect 2610 310112 2931 311136
rect 2610 310048 2618 310112
rect 2682 310048 2698 310112
rect 2762 310048 2778 310112
rect 2842 310048 2858 310112
rect 2922 310048 2931 310112
rect 2610 309024 2931 310048
rect 2610 308960 2618 309024
rect 2682 308960 2698 309024
rect 2762 308960 2778 309024
rect 2842 308960 2858 309024
rect 2922 308960 2931 309024
rect 2610 307936 2931 308960
rect 2610 307872 2618 307936
rect 2682 307872 2698 307936
rect 2762 307872 2778 307936
rect 2842 307872 2858 307936
rect 2922 307872 2931 307936
rect 2610 306848 2931 307872
rect 2610 306784 2618 306848
rect 2682 306784 2698 306848
rect 2762 306784 2778 306848
rect 2842 306784 2858 306848
rect 2922 306784 2931 306848
rect 2610 305760 2931 306784
rect 2610 305696 2618 305760
rect 2682 305696 2698 305760
rect 2762 305696 2778 305760
rect 2842 305696 2858 305760
rect 2922 305696 2931 305760
rect 2610 304672 2931 305696
rect 2610 304608 2618 304672
rect 2682 304608 2698 304672
rect 2762 304608 2778 304672
rect 2842 304608 2858 304672
rect 2922 304608 2931 304672
rect 2610 303584 2931 304608
rect 2610 303520 2618 303584
rect 2682 303520 2698 303584
rect 2762 303520 2778 303584
rect 2842 303520 2858 303584
rect 2922 303520 2931 303584
rect 2610 302496 2931 303520
rect 2610 302432 2618 302496
rect 2682 302432 2698 302496
rect 2762 302432 2778 302496
rect 2842 302432 2858 302496
rect 2922 302432 2931 302496
rect 2610 301408 2931 302432
rect 2610 301344 2618 301408
rect 2682 301344 2698 301408
rect 2762 301344 2778 301408
rect 2842 301344 2858 301408
rect 2922 301344 2931 301408
rect 2610 300320 2931 301344
rect 2610 300256 2618 300320
rect 2682 300256 2698 300320
rect 2762 300256 2778 300320
rect 2842 300256 2858 300320
rect 2922 300256 2931 300320
rect 2610 299232 2931 300256
rect 2610 299168 2618 299232
rect 2682 299168 2698 299232
rect 2762 299168 2778 299232
rect 2842 299168 2858 299232
rect 2922 299168 2931 299232
rect 2610 298144 2931 299168
rect 2610 298080 2618 298144
rect 2682 298080 2698 298144
rect 2762 298080 2778 298144
rect 2842 298080 2858 298144
rect 2922 298080 2931 298144
rect 2610 297056 2931 298080
rect 2610 296992 2618 297056
rect 2682 296992 2698 297056
rect 2762 296992 2778 297056
rect 2842 296992 2858 297056
rect 2922 296992 2931 297056
rect 2610 295968 2931 296992
rect 2610 295904 2618 295968
rect 2682 295904 2698 295968
rect 2762 295904 2778 295968
rect 2842 295904 2858 295968
rect 2922 295904 2931 295968
rect 2610 294880 2931 295904
rect 2610 294816 2618 294880
rect 2682 294816 2698 294880
rect 2762 294816 2778 294880
rect 2842 294816 2858 294880
rect 2922 294816 2931 294880
rect 2610 293792 2931 294816
rect 2610 293728 2618 293792
rect 2682 293728 2698 293792
rect 2762 293728 2778 293792
rect 2842 293728 2858 293792
rect 2922 293728 2931 293792
rect 2610 292704 2931 293728
rect 2610 292640 2618 292704
rect 2682 292640 2698 292704
rect 2762 292640 2778 292704
rect 2842 292640 2858 292704
rect 2922 292640 2931 292704
rect 2610 291616 2931 292640
rect 2610 291552 2618 291616
rect 2682 291552 2698 291616
rect 2762 291552 2778 291616
rect 2842 291552 2858 291616
rect 2922 291552 2931 291616
rect 2610 290528 2931 291552
rect 2610 290464 2618 290528
rect 2682 290464 2698 290528
rect 2762 290464 2778 290528
rect 2842 290464 2858 290528
rect 2922 290464 2931 290528
rect 2610 289440 2931 290464
rect 2610 289376 2618 289440
rect 2682 289376 2698 289440
rect 2762 289376 2778 289440
rect 2842 289376 2858 289440
rect 2922 289376 2931 289440
rect 2610 288352 2931 289376
rect 2610 288288 2618 288352
rect 2682 288288 2698 288352
rect 2762 288288 2778 288352
rect 2842 288288 2858 288352
rect 2922 288288 2931 288352
rect 2610 287264 2931 288288
rect 2610 287200 2618 287264
rect 2682 287200 2698 287264
rect 2762 287200 2778 287264
rect 2842 287200 2858 287264
rect 2922 287200 2931 287264
rect 2610 286176 2931 287200
rect 2610 286112 2618 286176
rect 2682 286112 2698 286176
rect 2762 286112 2778 286176
rect 2842 286112 2858 286176
rect 2922 286112 2931 286176
rect 2610 285088 2931 286112
rect 2610 285024 2618 285088
rect 2682 285024 2698 285088
rect 2762 285024 2778 285088
rect 2842 285024 2858 285088
rect 2922 285024 2931 285088
rect 2610 284000 2931 285024
rect 2610 283936 2618 284000
rect 2682 283936 2698 284000
rect 2762 283936 2778 284000
rect 2842 283936 2858 284000
rect 2922 283936 2931 284000
rect 2610 282912 2931 283936
rect 2610 282848 2618 282912
rect 2682 282848 2698 282912
rect 2762 282848 2778 282912
rect 2842 282848 2858 282912
rect 2922 282848 2931 282912
rect 2610 281824 2931 282848
rect 2610 281760 2618 281824
rect 2682 281760 2698 281824
rect 2762 281760 2778 281824
rect 2842 281760 2858 281824
rect 2922 281760 2931 281824
rect 2610 280736 2931 281760
rect 2610 280672 2618 280736
rect 2682 280672 2698 280736
rect 2762 280672 2778 280736
rect 2842 280672 2858 280736
rect 2922 280672 2931 280736
rect 2610 279648 2931 280672
rect 2610 279584 2618 279648
rect 2682 279584 2698 279648
rect 2762 279584 2778 279648
rect 2842 279584 2858 279648
rect 2922 279584 2931 279648
rect 2610 278560 2931 279584
rect 2610 278496 2618 278560
rect 2682 278496 2698 278560
rect 2762 278496 2778 278560
rect 2842 278496 2858 278560
rect 2922 278496 2931 278560
rect 2610 277472 2931 278496
rect 2610 277408 2618 277472
rect 2682 277408 2698 277472
rect 2762 277408 2778 277472
rect 2842 277408 2858 277472
rect 2922 277408 2931 277472
rect 2610 276384 2931 277408
rect 2610 276320 2618 276384
rect 2682 276320 2698 276384
rect 2762 276320 2778 276384
rect 2842 276320 2858 276384
rect 2922 276320 2931 276384
rect 2610 275296 2931 276320
rect 2610 275232 2618 275296
rect 2682 275232 2698 275296
rect 2762 275232 2778 275296
rect 2842 275232 2858 275296
rect 2922 275232 2931 275296
rect 2610 274208 2931 275232
rect 2610 274144 2618 274208
rect 2682 274144 2698 274208
rect 2762 274144 2778 274208
rect 2842 274144 2858 274208
rect 2922 274144 2931 274208
rect 2610 273120 2931 274144
rect 2610 273056 2618 273120
rect 2682 273056 2698 273120
rect 2762 273056 2778 273120
rect 2842 273056 2858 273120
rect 2922 273056 2931 273120
rect 2610 272032 2931 273056
rect 2610 271968 2618 272032
rect 2682 271968 2698 272032
rect 2762 271968 2778 272032
rect 2842 271968 2858 272032
rect 2922 271968 2931 272032
rect 2610 270944 2931 271968
rect 2610 270880 2618 270944
rect 2682 270880 2698 270944
rect 2762 270880 2778 270944
rect 2842 270880 2858 270944
rect 2922 270880 2931 270944
rect 2610 269856 2931 270880
rect 2610 269792 2618 269856
rect 2682 269792 2698 269856
rect 2762 269792 2778 269856
rect 2842 269792 2858 269856
rect 2922 269792 2931 269856
rect 2610 268768 2931 269792
rect 2610 268704 2618 268768
rect 2682 268704 2698 268768
rect 2762 268704 2778 268768
rect 2842 268704 2858 268768
rect 2922 268704 2931 268768
rect 2610 267680 2931 268704
rect 2610 267616 2618 267680
rect 2682 267616 2698 267680
rect 2762 267616 2778 267680
rect 2842 267616 2858 267680
rect 2922 267616 2931 267680
rect 2610 266592 2931 267616
rect 2610 266528 2618 266592
rect 2682 266528 2698 266592
rect 2762 266528 2778 266592
rect 2842 266528 2858 266592
rect 2922 266528 2931 266592
rect 2610 265504 2931 266528
rect 2610 265440 2618 265504
rect 2682 265440 2698 265504
rect 2762 265440 2778 265504
rect 2842 265440 2858 265504
rect 2922 265440 2931 265504
rect 2610 264416 2931 265440
rect 2610 264352 2618 264416
rect 2682 264352 2698 264416
rect 2762 264352 2778 264416
rect 2842 264352 2858 264416
rect 2922 264352 2931 264416
rect 2610 263328 2931 264352
rect 2610 263264 2618 263328
rect 2682 263264 2698 263328
rect 2762 263264 2778 263328
rect 2842 263264 2858 263328
rect 2922 263264 2931 263328
rect 2610 262240 2931 263264
rect 2610 262176 2618 262240
rect 2682 262176 2698 262240
rect 2762 262176 2778 262240
rect 2842 262176 2858 262240
rect 2922 262176 2931 262240
rect 2610 261152 2931 262176
rect 2610 261088 2618 261152
rect 2682 261088 2698 261152
rect 2762 261088 2778 261152
rect 2842 261088 2858 261152
rect 2922 261088 2931 261152
rect 2610 260064 2931 261088
rect 2610 260000 2618 260064
rect 2682 260000 2698 260064
rect 2762 260000 2778 260064
rect 2842 260000 2858 260064
rect 2922 260000 2931 260064
rect 2610 258976 2931 260000
rect 2610 258912 2618 258976
rect 2682 258912 2698 258976
rect 2762 258912 2778 258976
rect 2842 258912 2858 258976
rect 2922 258912 2931 258976
rect 2610 257888 2931 258912
rect 2610 257824 2618 257888
rect 2682 257824 2698 257888
rect 2762 257824 2778 257888
rect 2842 257824 2858 257888
rect 2922 257824 2931 257888
rect 2610 256800 2931 257824
rect 2610 256736 2618 256800
rect 2682 256736 2698 256800
rect 2762 256736 2778 256800
rect 2842 256736 2858 256800
rect 2922 256736 2931 256800
rect 2610 255712 2931 256736
rect 2610 255648 2618 255712
rect 2682 255648 2698 255712
rect 2762 255648 2778 255712
rect 2842 255648 2858 255712
rect 2922 255648 2931 255712
rect 2610 254624 2931 255648
rect 2610 254560 2618 254624
rect 2682 254560 2698 254624
rect 2762 254560 2778 254624
rect 2842 254560 2858 254624
rect 2922 254560 2931 254624
rect 2610 253536 2931 254560
rect 2610 253472 2618 253536
rect 2682 253472 2698 253536
rect 2762 253472 2778 253536
rect 2842 253472 2858 253536
rect 2922 253472 2931 253536
rect 2610 252448 2931 253472
rect 2610 252384 2618 252448
rect 2682 252384 2698 252448
rect 2762 252384 2778 252448
rect 2842 252384 2858 252448
rect 2922 252384 2931 252448
rect 2610 251360 2931 252384
rect 2610 251296 2618 251360
rect 2682 251296 2698 251360
rect 2762 251296 2778 251360
rect 2842 251296 2858 251360
rect 2922 251296 2931 251360
rect 2610 250272 2931 251296
rect 2610 250208 2618 250272
rect 2682 250208 2698 250272
rect 2762 250208 2778 250272
rect 2842 250208 2858 250272
rect 2922 250208 2931 250272
rect 2610 249184 2931 250208
rect 2610 249120 2618 249184
rect 2682 249120 2698 249184
rect 2762 249120 2778 249184
rect 2842 249120 2858 249184
rect 2922 249120 2931 249184
rect 2610 248096 2931 249120
rect 2610 248032 2618 248096
rect 2682 248032 2698 248096
rect 2762 248032 2778 248096
rect 2842 248032 2858 248096
rect 2922 248032 2931 248096
rect 2610 247008 2931 248032
rect 2610 246944 2618 247008
rect 2682 246944 2698 247008
rect 2762 246944 2778 247008
rect 2842 246944 2858 247008
rect 2922 246944 2931 247008
rect 2610 245920 2931 246944
rect 2610 245856 2618 245920
rect 2682 245856 2698 245920
rect 2762 245856 2778 245920
rect 2842 245856 2858 245920
rect 2922 245856 2931 245920
rect 2610 244832 2931 245856
rect 2610 244768 2618 244832
rect 2682 244768 2698 244832
rect 2762 244768 2778 244832
rect 2842 244768 2858 244832
rect 2922 244768 2931 244832
rect 2610 243744 2931 244768
rect 2610 243680 2618 243744
rect 2682 243680 2698 243744
rect 2762 243680 2778 243744
rect 2842 243680 2858 243744
rect 2922 243680 2931 243744
rect 2610 242656 2931 243680
rect 2610 242592 2618 242656
rect 2682 242592 2698 242656
rect 2762 242592 2778 242656
rect 2842 242592 2858 242656
rect 2922 242592 2931 242656
rect 2610 241568 2931 242592
rect 2610 241504 2618 241568
rect 2682 241504 2698 241568
rect 2762 241504 2778 241568
rect 2842 241504 2858 241568
rect 2922 241504 2931 241568
rect 2610 240480 2931 241504
rect 2610 240416 2618 240480
rect 2682 240416 2698 240480
rect 2762 240416 2778 240480
rect 2842 240416 2858 240480
rect 2922 240416 2931 240480
rect 2610 239392 2931 240416
rect 2610 239328 2618 239392
rect 2682 239328 2698 239392
rect 2762 239328 2778 239392
rect 2842 239328 2858 239392
rect 2922 239328 2931 239392
rect 2610 238304 2931 239328
rect 2610 238240 2618 238304
rect 2682 238240 2698 238304
rect 2762 238240 2778 238304
rect 2842 238240 2858 238304
rect 2922 238240 2931 238304
rect 2610 237216 2931 238240
rect 2610 237152 2618 237216
rect 2682 237152 2698 237216
rect 2762 237152 2778 237216
rect 2842 237152 2858 237216
rect 2922 237152 2931 237216
rect 2610 236128 2931 237152
rect 2610 236064 2618 236128
rect 2682 236064 2698 236128
rect 2762 236064 2778 236128
rect 2842 236064 2858 236128
rect 2922 236064 2931 236128
rect 2610 235040 2931 236064
rect 2610 234976 2618 235040
rect 2682 234976 2698 235040
rect 2762 234976 2778 235040
rect 2842 234976 2858 235040
rect 2922 234976 2931 235040
rect 2610 233952 2931 234976
rect 2610 233888 2618 233952
rect 2682 233888 2698 233952
rect 2762 233888 2778 233952
rect 2842 233888 2858 233952
rect 2922 233888 2931 233952
rect 2610 232864 2931 233888
rect 2610 232800 2618 232864
rect 2682 232800 2698 232864
rect 2762 232800 2778 232864
rect 2842 232800 2858 232864
rect 2922 232800 2931 232864
rect 2610 231776 2931 232800
rect 2610 231712 2618 231776
rect 2682 231712 2698 231776
rect 2762 231712 2778 231776
rect 2842 231712 2858 231776
rect 2922 231712 2931 231776
rect 2610 230688 2931 231712
rect 2610 230624 2618 230688
rect 2682 230624 2698 230688
rect 2762 230624 2778 230688
rect 2842 230624 2858 230688
rect 2922 230624 2931 230688
rect 2610 229600 2931 230624
rect 2610 229536 2618 229600
rect 2682 229536 2698 229600
rect 2762 229536 2778 229600
rect 2842 229536 2858 229600
rect 2922 229536 2931 229600
rect 2610 228512 2931 229536
rect 2610 228448 2618 228512
rect 2682 228448 2698 228512
rect 2762 228448 2778 228512
rect 2842 228448 2858 228512
rect 2922 228448 2931 228512
rect 2610 227424 2931 228448
rect 2610 227360 2618 227424
rect 2682 227360 2698 227424
rect 2762 227360 2778 227424
rect 2842 227360 2858 227424
rect 2922 227360 2931 227424
rect 2610 226336 2931 227360
rect 2610 226272 2618 226336
rect 2682 226272 2698 226336
rect 2762 226272 2778 226336
rect 2842 226272 2858 226336
rect 2922 226272 2931 226336
rect 2610 225248 2931 226272
rect 2610 225184 2618 225248
rect 2682 225184 2698 225248
rect 2762 225184 2778 225248
rect 2842 225184 2858 225248
rect 2922 225184 2931 225248
rect 2610 224160 2931 225184
rect 2610 224096 2618 224160
rect 2682 224096 2698 224160
rect 2762 224096 2778 224160
rect 2842 224096 2858 224160
rect 2922 224096 2931 224160
rect 2610 223072 2931 224096
rect 2610 223008 2618 223072
rect 2682 223008 2698 223072
rect 2762 223008 2778 223072
rect 2842 223008 2858 223072
rect 2922 223008 2931 223072
rect 2610 221984 2931 223008
rect 2610 221920 2618 221984
rect 2682 221920 2698 221984
rect 2762 221920 2778 221984
rect 2842 221920 2858 221984
rect 2922 221920 2931 221984
rect 2610 220896 2931 221920
rect 2610 220832 2618 220896
rect 2682 220832 2698 220896
rect 2762 220832 2778 220896
rect 2842 220832 2858 220896
rect 2922 220832 2931 220896
rect 2610 219808 2931 220832
rect 2610 219744 2618 219808
rect 2682 219744 2698 219808
rect 2762 219744 2778 219808
rect 2842 219744 2858 219808
rect 2922 219744 2931 219808
rect 2610 218720 2931 219744
rect 2610 218656 2618 218720
rect 2682 218656 2698 218720
rect 2762 218656 2778 218720
rect 2842 218656 2858 218720
rect 2922 218656 2931 218720
rect 2610 217632 2931 218656
rect 2610 217568 2618 217632
rect 2682 217568 2698 217632
rect 2762 217568 2778 217632
rect 2842 217568 2858 217632
rect 2922 217568 2931 217632
rect 2610 216544 2931 217568
rect 2610 216480 2618 216544
rect 2682 216480 2698 216544
rect 2762 216480 2778 216544
rect 2842 216480 2858 216544
rect 2922 216480 2931 216544
rect 2610 215456 2931 216480
rect 2610 215392 2618 215456
rect 2682 215392 2698 215456
rect 2762 215392 2778 215456
rect 2842 215392 2858 215456
rect 2922 215392 2931 215456
rect 2610 214368 2931 215392
rect 2610 214304 2618 214368
rect 2682 214304 2698 214368
rect 2762 214304 2778 214368
rect 2842 214304 2858 214368
rect 2922 214304 2931 214368
rect 2610 213280 2931 214304
rect 2610 213216 2618 213280
rect 2682 213216 2698 213280
rect 2762 213216 2778 213280
rect 2842 213216 2858 213280
rect 2922 213216 2931 213280
rect 2610 212192 2931 213216
rect 2610 212128 2618 212192
rect 2682 212128 2698 212192
rect 2762 212128 2778 212192
rect 2842 212128 2858 212192
rect 2922 212128 2931 212192
rect 2610 211104 2931 212128
rect 2610 211040 2618 211104
rect 2682 211040 2698 211104
rect 2762 211040 2778 211104
rect 2842 211040 2858 211104
rect 2922 211040 2931 211104
rect 2610 210016 2931 211040
rect 2610 209952 2618 210016
rect 2682 209952 2698 210016
rect 2762 209952 2778 210016
rect 2842 209952 2858 210016
rect 2922 209952 2931 210016
rect 2610 208928 2931 209952
rect 2610 208864 2618 208928
rect 2682 208864 2698 208928
rect 2762 208864 2778 208928
rect 2842 208864 2858 208928
rect 2922 208864 2931 208928
rect 2610 207840 2931 208864
rect 2610 207776 2618 207840
rect 2682 207776 2698 207840
rect 2762 207776 2778 207840
rect 2842 207776 2858 207840
rect 2922 207776 2931 207840
rect 2610 206752 2931 207776
rect 2610 206688 2618 206752
rect 2682 206688 2698 206752
rect 2762 206688 2778 206752
rect 2842 206688 2858 206752
rect 2922 206688 2931 206752
rect 2610 205664 2931 206688
rect 2610 205600 2618 205664
rect 2682 205600 2698 205664
rect 2762 205600 2778 205664
rect 2842 205600 2858 205664
rect 2922 205600 2931 205664
rect 2610 204576 2931 205600
rect 2610 204512 2618 204576
rect 2682 204512 2698 204576
rect 2762 204512 2778 204576
rect 2842 204512 2858 204576
rect 2922 204512 2931 204576
rect 2610 203488 2931 204512
rect 2610 203424 2618 203488
rect 2682 203424 2698 203488
rect 2762 203424 2778 203488
rect 2842 203424 2858 203488
rect 2922 203424 2931 203488
rect 2610 202400 2931 203424
rect 2610 202336 2618 202400
rect 2682 202336 2698 202400
rect 2762 202336 2778 202400
rect 2842 202336 2858 202400
rect 2922 202336 2931 202400
rect 2610 201312 2931 202336
rect 2610 201248 2618 201312
rect 2682 201248 2698 201312
rect 2762 201248 2778 201312
rect 2842 201248 2858 201312
rect 2922 201248 2931 201312
rect 2610 200224 2931 201248
rect 2610 200160 2618 200224
rect 2682 200160 2698 200224
rect 2762 200160 2778 200224
rect 2842 200160 2858 200224
rect 2922 200160 2931 200224
rect 2610 199136 2931 200160
rect 2610 199072 2618 199136
rect 2682 199072 2698 199136
rect 2762 199072 2778 199136
rect 2842 199072 2858 199136
rect 2922 199072 2931 199136
rect 2610 198048 2931 199072
rect 2610 197984 2618 198048
rect 2682 197984 2698 198048
rect 2762 197984 2778 198048
rect 2842 197984 2858 198048
rect 2922 197984 2931 198048
rect 2610 196960 2931 197984
rect 2610 196896 2618 196960
rect 2682 196896 2698 196960
rect 2762 196896 2778 196960
rect 2842 196896 2858 196960
rect 2922 196896 2931 196960
rect 2610 195872 2931 196896
rect 2610 195808 2618 195872
rect 2682 195808 2698 195872
rect 2762 195808 2778 195872
rect 2842 195808 2858 195872
rect 2922 195808 2931 195872
rect 2610 194784 2931 195808
rect 2610 194720 2618 194784
rect 2682 194720 2698 194784
rect 2762 194720 2778 194784
rect 2842 194720 2858 194784
rect 2922 194720 2931 194784
rect 2610 193696 2931 194720
rect 2610 193632 2618 193696
rect 2682 193632 2698 193696
rect 2762 193632 2778 193696
rect 2842 193632 2858 193696
rect 2922 193632 2931 193696
rect 2610 192608 2931 193632
rect 2610 192544 2618 192608
rect 2682 192544 2698 192608
rect 2762 192544 2778 192608
rect 2842 192544 2858 192608
rect 2922 192544 2931 192608
rect 2610 191520 2931 192544
rect 2610 191456 2618 191520
rect 2682 191456 2698 191520
rect 2762 191456 2778 191520
rect 2842 191456 2858 191520
rect 2922 191456 2931 191520
rect 2610 190432 2931 191456
rect 2610 190368 2618 190432
rect 2682 190368 2698 190432
rect 2762 190368 2778 190432
rect 2842 190368 2858 190432
rect 2922 190368 2931 190432
rect 2610 189344 2931 190368
rect 2610 189280 2618 189344
rect 2682 189280 2698 189344
rect 2762 189280 2778 189344
rect 2842 189280 2858 189344
rect 2922 189280 2931 189344
rect 2610 188256 2931 189280
rect 2610 188192 2618 188256
rect 2682 188192 2698 188256
rect 2762 188192 2778 188256
rect 2842 188192 2858 188256
rect 2922 188192 2931 188256
rect 2610 187168 2931 188192
rect 2610 187104 2618 187168
rect 2682 187104 2698 187168
rect 2762 187104 2778 187168
rect 2842 187104 2858 187168
rect 2922 187104 2931 187168
rect 2610 186080 2931 187104
rect 2610 186016 2618 186080
rect 2682 186016 2698 186080
rect 2762 186016 2778 186080
rect 2842 186016 2858 186080
rect 2922 186016 2931 186080
rect 2610 184992 2931 186016
rect 2610 184928 2618 184992
rect 2682 184928 2698 184992
rect 2762 184928 2778 184992
rect 2842 184928 2858 184992
rect 2922 184928 2931 184992
rect 2610 183904 2931 184928
rect 2610 183840 2618 183904
rect 2682 183840 2698 183904
rect 2762 183840 2778 183904
rect 2842 183840 2858 183904
rect 2922 183840 2931 183904
rect 2610 182816 2931 183840
rect 2610 182752 2618 182816
rect 2682 182752 2698 182816
rect 2762 182752 2778 182816
rect 2842 182752 2858 182816
rect 2922 182752 2931 182816
rect 2610 181728 2931 182752
rect 2610 181664 2618 181728
rect 2682 181664 2698 181728
rect 2762 181664 2778 181728
rect 2842 181664 2858 181728
rect 2922 181664 2931 181728
rect 2610 180640 2931 181664
rect 2610 180576 2618 180640
rect 2682 180576 2698 180640
rect 2762 180576 2778 180640
rect 2842 180576 2858 180640
rect 2922 180576 2931 180640
rect 2610 179552 2931 180576
rect 2610 179488 2618 179552
rect 2682 179488 2698 179552
rect 2762 179488 2778 179552
rect 2842 179488 2858 179552
rect 2922 179488 2931 179552
rect 2610 178464 2931 179488
rect 2610 178400 2618 178464
rect 2682 178400 2698 178464
rect 2762 178400 2778 178464
rect 2842 178400 2858 178464
rect 2922 178400 2931 178464
rect 2610 177376 2931 178400
rect 2610 177312 2618 177376
rect 2682 177312 2698 177376
rect 2762 177312 2778 177376
rect 2842 177312 2858 177376
rect 2922 177312 2931 177376
rect 2610 176288 2931 177312
rect 2610 176224 2618 176288
rect 2682 176224 2698 176288
rect 2762 176224 2778 176288
rect 2842 176224 2858 176288
rect 2922 176224 2931 176288
rect 2610 175200 2931 176224
rect 2610 175136 2618 175200
rect 2682 175136 2698 175200
rect 2762 175136 2778 175200
rect 2842 175136 2858 175200
rect 2922 175136 2931 175200
rect 2610 174112 2931 175136
rect 2610 174048 2618 174112
rect 2682 174048 2698 174112
rect 2762 174048 2778 174112
rect 2842 174048 2858 174112
rect 2922 174048 2931 174112
rect 2610 173024 2931 174048
rect 2610 172960 2618 173024
rect 2682 172960 2698 173024
rect 2762 172960 2778 173024
rect 2842 172960 2858 173024
rect 2922 172960 2931 173024
rect 2610 171936 2931 172960
rect 2610 171872 2618 171936
rect 2682 171872 2698 171936
rect 2762 171872 2778 171936
rect 2842 171872 2858 171936
rect 2922 171872 2931 171936
rect 2610 170848 2931 171872
rect 2610 170784 2618 170848
rect 2682 170784 2698 170848
rect 2762 170784 2778 170848
rect 2842 170784 2858 170848
rect 2922 170784 2931 170848
rect 2610 169760 2931 170784
rect 2610 169696 2618 169760
rect 2682 169696 2698 169760
rect 2762 169696 2778 169760
rect 2842 169696 2858 169760
rect 2922 169696 2931 169760
rect 2610 168672 2931 169696
rect 2610 168608 2618 168672
rect 2682 168608 2698 168672
rect 2762 168608 2778 168672
rect 2842 168608 2858 168672
rect 2922 168608 2931 168672
rect 2610 167584 2931 168608
rect 2610 167520 2618 167584
rect 2682 167520 2698 167584
rect 2762 167520 2778 167584
rect 2842 167520 2858 167584
rect 2922 167520 2931 167584
rect 2610 166496 2931 167520
rect 2610 166432 2618 166496
rect 2682 166432 2698 166496
rect 2762 166432 2778 166496
rect 2842 166432 2858 166496
rect 2922 166432 2931 166496
rect 2610 165408 2931 166432
rect 2610 165344 2618 165408
rect 2682 165344 2698 165408
rect 2762 165344 2778 165408
rect 2842 165344 2858 165408
rect 2922 165344 2931 165408
rect 2610 164320 2931 165344
rect 2610 164256 2618 164320
rect 2682 164256 2698 164320
rect 2762 164256 2778 164320
rect 2842 164256 2858 164320
rect 2922 164256 2931 164320
rect 2610 163232 2931 164256
rect 2610 163168 2618 163232
rect 2682 163168 2698 163232
rect 2762 163168 2778 163232
rect 2842 163168 2858 163232
rect 2922 163168 2931 163232
rect 2610 162144 2931 163168
rect 2610 162080 2618 162144
rect 2682 162080 2698 162144
rect 2762 162080 2778 162144
rect 2842 162080 2858 162144
rect 2922 162080 2931 162144
rect 2610 161056 2931 162080
rect 2610 160992 2618 161056
rect 2682 160992 2698 161056
rect 2762 160992 2778 161056
rect 2842 160992 2858 161056
rect 2922 160992 2931 161056
rect 2610 159968 2931 160992
rect 2610 159904 2618 159968
rect 2682 159904 2698 159968
rect 2762 159904 2778 159968
rect 2842 159904 2858 159968
rect 2922 159904 2931 159968
rect 2610 158880 2931 159904
rect 2610 158816 2618 158880
rect 2682 158816 2698 158880
rect 2762 158816 2778 158880
rect 2842 158816 2858 158880
rect 2922 158816 2931 158880
rect 2610 157792 2931 158816
rect 2610 157728 2618 157792
rect 2682 157728 2698 157792
rect 2762 157728 2778 157792
rect 2842 157728 2858 157792
rect 2922 157728 2931 157792
rect 2610 156704 2931 157728
rect 2610 156640 2618 156704
rect 2682 156640 2698 156704
rect 2762 156640 2778 156704
rect 2842 156640 2858 156704
rect 2922 156640 2931 156704
rect 2610 155616 2931 156640
rect 2610 155552 2618 155616
rect 2682 155552 2698 155616
rect 2762 155552 2778 155616
rect 2842 155552 2858 155616
rect 2922 155552 2931 155616
rect 2610 154528 2931 155552
rect 2610 154464 2618 154528
rect 2682 154464 2698 154528
rect 2762 154464 2778 154528
rect 2842 154464 2858 154528
rect 2922 154464 2931 154528
rect 2610 153440 2931 154464
rect 2610 153376 2618 153440
rect 2682 153376 2698 153440
rect 2762 153376 2778 153440
rect 2842 153376 2858 153440
rect 2922 153376 2931 153440
rect 2610 152352 2931 153376
rect 2610 152288 2618 152352
rect 2682 152288 2698 152352
rect 2762 152288 2778 152352
rect 2842 152288 2858 152352
rect 2922 152288 2931 152352
rect 2610 151264 2931 152288
rect 2610 151200 2618 151264
rect 2682 151200 2698 151264
rect 2762 151200 2778 151264
rect 2842 151200 2858 151264
rect 2922 151200 2931 151264
rect 2610 150176 2931 151200
rect 2610 150112 2618 150176
rect 2682 150112 2698 150176
rect 2762 150112 2778 150176
rect 2842 150112 2858 150176
rect 2922 150112 2931 150176
rect 2610 149088 2931 150112
rect 2610 149024 2618 149088
rect 2682 149024 2698 149088
rect 2762 149024 2778 149088
rect 2842 149024 2858 149088
rect 2922 149024 2931 149088
rect 2610 148000 2931 149024
rect 2610 147936 2618 148000
rect 2682 147936 2698 148000
rect 2762 147936 2778 148000
rect 2842 147936 2858 148000
rect 2922 147936 2931 148000
rect 2610 146912 2931 147936
rect 2610 146848 2618 146912
rect 2682 146848 2698 146912
rect 2762 146848 2778 146912
rect 2842 146848 2858 146912
rect 2922 146848 2931 146912
rect 2610 145824 2931 146848
rect 2610 145760 2618 145824
rect 2682 145760 2698 145824
rect 2762 145760 2778 145824
rect 2842 145760 2858 145824
rect 2922 145760 2931 145824
rect 2610 144736 2931 145760
rect 2610 144672 2618 144736
rect 2682 144672 2698 144736
rect 2762 144672 2778 144736
rect 2842 144672 2858 144736
rect 2922 144672 2931 144736
rect 2610 143648 2931 144672
rect 2610 143584 2618 143648
rect 2682 143584 2698 143648
rect 2762 143584 2778 143648
rect 2842 143584 2858 143648
rect 2922 143584 2931 143648
rect 2610 142560 2931 143584
rect 2610 142496 2618 142560
rect 2682 142496 2698 142560
rect 2762 142496 2778 142560
rect 2842 142496 2858 142560
rect 2922 142496 2931 142560
rect 2610 141472 2931 142496
rect 2610 141408 2618 141472
rect 2682 141408 2698 141472
rect 2762 141408 2778 141472
rect 2842 141408 2858 141472
rect 2922 141408 2931 141472
rect 2610 140384 2931 141408
rect 2610 140320 2618 140384
rect 2682 140320 2698 140384
rect 2762 140320 2778 140384
rect 2842 140320 2858 140384
rect 2922 140320 2931 140384
rect 2610 139296 2931 140320
rect 2610 139232 2618 139296
rect 2682 139232 2698 139296
rect 2762 139232 2778 139296
rect 2842 139232 2858 139296
rect 2922 139232 2931 139296
rect 2610 138208 2931 139232
rect 2610 138144 2618 138208
rect 2682 138144 2698 138208
rect 2762 138144 2778 138208
rect 2842 138144 2858 138208
rect 2922 138144 2931 138208
rect 2610 137120 2931 138144
rect 2610 137056 2618 137120
rect 2682 137056 2698 137120
rect 2762 137056 2778 137120
rect 2842 137056 2858 137120
rect 2922 137056 2931 137120
rect 2610 136032 2931 137056
rect 2610 135968 2618 136032
rect 2682 135968 2698 136032
rect 2762 135968 2778 136032
rect 2842 135968 2858 136032
rect 2922 135968 2931 136032
rect 2610 134944 2931 135968
rect 2610 134880 2618 134944
rect 2682 134880 2698 134944
rect 2762 134880 2778 134944
rect 2842 134880 2858 134944
rect 2922 134880 2931 134944
rect 2610 133856 2931 134880
rect 2610 133792 2618 133856
rect 2682 133792 2698 133856
rect 2762 133792 2778 133856
rect 2842 133792 2858 133856
rect 2922 133792 2931 133856
rect 2610 132768 2931 133792
rect 2610 132704 2618 132768
rect 2682 132704 2698 132768
rect 2762 132704 2778 132768
rect 2842 132704 2858 132768
rect 2922 132704 2931 132768
rect 2610 131680 2931 132704
rect 2610 131616 2618 131680
rect 2682 131616 2698 131680
rect 2762 131616 2778 131680
rect 2842 131616 2858 131680
rect 2922 131616 2931 131680
rect 2610 130592 2931 131616
rect 2610 130528 2618 130592
rect 2682 130528 2698 130592
rect 2762 130528 2778 130592
rect 2842 130528 2858 130592
rect 2922 130528 2931 130592
rect 2610 129504 2931 130528
rect 2610 129440 2618 129504
rect 2682 129440 2698 129504
rect 2762 129440 2778 129504
rect 2842 129440 2858 129504
rect 2922 129440 2931 129504
rect 2610 128416 2931 129440
rect 2610 128352 2618 128416
rect 2682 128352 2698 128416
rect 2762 128352 2778 128416
rect 2842 128352 2858 128416
rect 2922 128352 2931 128416
rect 2610 127328 2931 128352
rect 2610 127264 2618 127328
rect 2682 127264 2698 127328
rect 2762 127264 2778 127328
rect 2842 127264 2858 127328
rect 2922 127264 2931 127328
rect 2610 126240 2931 127264
rect 2610 126176 2618 126240
rect 2682 126176 2698 126240
rect 2762 126176 2778 126240
rect 2842 126176 2858 126240
rect 2922 126176 2931 126240
rect 2610 125152 2931 126176
rect 2610 125088 2618 125152
rect 2682 125088 2698 125152
rect 2762 125088 2778 125152
rect 2842 125088 2858 125152
rect 2922 125088 2931 125152
rect 2610 124064 2931 125088
rect 2610 124000 2618 124064
rect 2682 124000 2698 124064
rect 2762 124000 2778 124064
rect 2842 124000 2858 124064
rect 2922 124000 2931 124064
rect 2610 122976 2931 124000
rect 2610 122912 2618 122976
rect 2682 122912 2698 122976
rect 2762 122912 2778 122976
rect 2842 122912 2858 122976
rect 2922 122912 2931 122976
rect 2610 121888 2931 122912
rect 2610 121824 2618 121888
rect 2682 121824 2698 121888
rect 2762 121824 2778 121888
rect 2842 121824 2858 121888
rect 2922 121824 2931 121888
rect 2610 120800 2931 121824
rect 2610 120736 2618 120800
rect 2682 120736 2698 120800
rect 2762 120736 2778 120800
rect 2842 120736 2858 120800
rect 2922 120736 2931 120800
rect 2610 119712 2931 120736
rect 2610 119648 2618 119712
rect 2682 119648 2698 119712
rect 2762 119648 2778 119712
rect 2842 119648 2858 119712
rect 2922 119648 2931 119712
rect 2610 118624 2931 119648
rect 2610 118560 2618 118624
rect 2682 118560 2698 118624
rect 2762 118560 2778 118624
rect 2842 118560 2858 118624
rect 2922 118560 2931 118624
rect 2610 117536 2931 118560
rect 2610 117472 2618 117536
rect 2682 117472 2698 117536
rect 2762 117472 2778 117536
rect 2842 117472 2858 117536
rect 2922 117472 2931 117536
rect 2610 116448 2931 117472
rect 2610 116384 2618 116448
rect 2682 116384 2698 116448
rect 2762 116384 2778 116448
rect 2842 116384 2858 116448
rect 2922 116384 2931 116448
rect 2610 115360 2931 116384
rect 2610 115296 2618 115360
rect 2682 115296 2698 115360
rect 2762 115296 2778 115360
rect 2842 115296 2858 115360
rect 2922 115296 2931 115360
rect 2610 114272 2931 115296
rect 2610 114208 2618 114272
rect 2682 114208 2698 114272
rect 2762 114208 2778 114272
rect 2842 114208 2858 114272
rect 2922 114208 2931 114272
rect 2610 113184 2931 114208
rect 2610 113120 2618 113184
rect 2682 113120 2698 113184
rect 2762 113120 2778 113184
rect 2842 113120 2858 113184
rect 2922 113120 2931 113184
rect 2610 112096 2931 113120
rect 2610 112032 2618 112096
rect 2682 112032 2698 112096
rect 2762 112032 2778 112096
rect 2842 112032 2858 112096
rect 2922 112032 2931 112096
rect 2610 111008 2931 112032
rect 2610 110944 2618 111008
rect 2682 110944 2698 111008
rect 2762 110944 2778 111008
rect 2842 110944 2858 111008
rect 2922 110944 2931 111008
rect 2610 109920 2931 110944
rect 2610 109856 2618 109920
rect 2682 109856 2698 109920
rect 2762 109856 2778 109920
rect 2842 109856 2858 109920
rect 2922 109856 2931 109920
rect 2610 108832 2931 109856
rect 2610 108768 2618 108832
rect 2682 108768 2698 108832
rect 2762 108768 2778 108832
rect 2842 108768 2858 108832
rect 2922 108768 2931 108832
rect 2610 107744 2931 108768
rect 2610 107680 2618 107744
rect 2682 107680 2698 107744
rect 2762 107680 2778 107744
rect 2842 107680 2858 107744
rect 2922 107680 2931 107744
rect 2610 106656 2931 107680
rect 2610 106592 2618 106656
rect 2682 106592 2698 106656
rect 2762 106592 2778 106656
rect 2842 106592 2858 106656
rect 2922 106592 2931 106656
rect 2610 105568 2931 106592
rect 2610 105504 2618 105568
rect 2682 105504 2698 105568
rect 2762 105504 2778 105568
rect 2842 105504 2858 105568
rect 2922 105504 2931 105568
rect 2610 104480 2931 105504
rect 2610 104416 2618 104480
rect 2682 104416 2698 104480
rect 2762 104416 2778 104480
rect 2842 104416 2858 104480
rect 2922 104416 2931 104480
rect 2610 103392 2931 104416
rect 2610 103328 2618 103392
rect 2682 103328 2698 103392
rect 2762 103328 2778 103392
rect 2842 103328 2858 103392
rect 2922 103328 2931 103392
rect 2610 102304 2931 103328
rect 2610 102240 2618 102304
rect 2682 102240 2698 102304
rect 2762 102240 2778 102304
rect 2842 102240 2858 102304
rect 2922 102240 2931 102304
rect 2610 101216 2931 102240
rect 2610 101152 2618 101216
rect 2682 101152 2698 101216
rect 2762 101152 2778 101216
rect 2842 101152 2858 101216
rect 2922 101152 2931 101216
rect 2610 100128 2931 101152
rect 2610 100064 2618 100128
rect 2682 100064 2698 100128
rect 2762 100064 2778 100128
rect 2842 100064 2858 100128
rect 2922 100064 2931 100128
rect 2610 99040 2931 100064
rect 2610 98976 2618 99040
rect 2682 98976 2698 99040
rect 2762 98976 2778 99040
rect 2842 98976 2858 99040
rect 2922 98976 2931 99040
rect 2610 97952 2931 98976
rect 2610 97888 2618 97952
rect 2682 97888 2698 97952
rect 2762 97888 2778 97952
rect 2842 97888 2858 97952
rect 2922 97888 2931 97952
rect 2610 96864 2931 97888
rect 2610 96800 2618 96864
rect 2682 96800 2698 96864
rect 2762 96800 2778 96864
rect 2842 96800 2858 96864
rect 2922 96800 2931 96864
rect 2610 95776 2931 96800
rect 2610 95712 2618 95776
rect 2682 95712 2698 95776
rect 2762 95712 2778 95776
rect 2842 95712 2858 95776
rect 2922 95712 2931 95776
rect 2610 94688 2931 95712
rect 2610 94624 2618 94688
rect 2682 94624 2698 94688
rect 2762 94624 2778 94688
rect 2842 94624 2858 94688
rect 2922 94624 2931 94688
rect 2610 93600 2931 94624
rect 2610 93536 2618 93600
rect 2682 93536 2698 93600
rect 2762 93536 2778 93600
rect 2842 93536 2858 93600
rect 2922 93536 2931 93600
rect 2610 92512 2931 93536
rect 2610 92448 2618 92512
rect 2682 92448 2698 92512
rect 2762 92448 2778 92512
rect 2842 92448 2858 92512
rect 2922 92448 2931 92512
rect 2610 91424 2931 92448
rect 2610 91360 2618 91424
rect 2682 91360 2698 91424
rect 2762 91360 2778 91424
rect 2842 91360 2858 91424
rect 2922 91360 2931 91424
rect 2610 90336 2931 91360
rect 2610 90272 2618 90336
rect 2682 90272 2698 90336
rect 2762 90272 2778 90336
rect 2842 90272 2858 90336
rect 2922 90272 2931 90336
rect 2610 89248 2931 90272
rect 2610 89184 2618 89248
rect 2682 89184 2698 89248
rect 2762 89184 2778 89248
rect 2842 89184 2858 89248
rect 2922 89184 2931 89248
rect 2610 88160 2931 89184
rect 2610 88096 2618 88160
rect 2682 88096 2698 88160
rect 2762 88096 2778 88160
rect 2842 88096 2858 88160
rect 2922 88096 2931 88160
rect 2610 87072 2931 88096
rect 2610 87008 2618 87072
rect 2682 87008 2698 87072
rect 2762 87008 2778 87072
rect 2842 87008 2858 87072
rect 2922 87008 2931 87072
rect 2610 85984 2931 87008
rect 2610 85920 2618 85984
rect 2682 85920 2698 85984
rect 2762 85920 2778 85984
rect 2842 85920 2858 85984
rect 2922 85920 2931 85984
rect 2610 84896 2931 85920
rect 2610 84832 2618 84896
rect 2682 84832 2698 84896
rect 2762 84832 2778 84896
rect 2842 84832 2858 84896
rect 2922 84832 2931 84896
rect 2610 83808 2931 84832
rect 2610 83744 2618 83808
rect 2682 83744 2698 83808
rect 2762 83744 2778 83808
rect 2842 83744 2858 83808
rect 2922 83744 2931 83808
rect 2610 82720 2931 83744
rect 2610 82656 2618 82720
rect 2682 82656 2698 82720
rect 2762 82656 2778 82720
rect 2842 82656 2858 82720
rect 2922 82656 2931 82720
rect 2610 81632 2931 82656
rect 2610 81568 2618 81632
rect 2682 81568 2698 81632
rect 2762 81568 2778 81632
rect 2842 81568 2858 81632
rect 2922 81568 2931 81632
rect 2610 80544 2931 81568
rect 2610 80480 2618 80544
rect 2682 80480 2698 80544
rect 2762 80480 2778 80544
rect 2842 80480 2858 80544
rect 2922 80480 2931 80544
rect 2610 79456 2931 80480
rect 2610 79392 2618 79456
rect 2682 79392 2698 79456
rect 2762 79392 2778 79456
rect 2842 79392 2858 79456
rect 2922 79392 2931 79456
rect 2610 78368 2931 79392
rect 2610 78304 2618 78368
rect 2682 78304 2698 78368
rect 2762 78304 2778 78368
rect 2842 78304 2858 78368
rect 2922 78304 2931 78368
rect 2610 77280 2931 78304
rect 2610 77216 2618 77280
rect 2682 77216 2698 77280
rect 2762 77216 2778 77280
rect 2842 77216 2858 77280
rect 2922 77216 2931 77280
rect 2610 76192 2931 77216
rect 2610 76128 2618 76192
rect 2682 76128 2698 76192
rect 2762 76128 2778 76192
rect 2842 76128 2858 76192
rect 2922 76128 2931 76192
rect 2610 75104 2931 76128
rect 2610 75040 2618 75104
rect 2682 75040 2698 75104
rect 2762 75040 2778 75104
rect 2842 75040 2858 75104
rect 2922 75040 2931 75104
rect 2610 74016 2931 75040
rect 2610 73952 2618 74016
rect 2682 73952 2698 74016
rect 2762 73952 2778 74016
rect 2842 73952 2858 74016
rect 2922 73952 2931 74016
rect 2610 72928 2931 73952
rect 2610 72864 2618 72928
rect 2682 72864 2698 72928
rect 2762 72864 2778 72928
rect 2842 72864 2858 72928
rect 2922 72864 2931 72928
rect 2610 71840 2931 72864
rect 2610 71776 2618 71840
rect 2682 71776 2698 71840
rect 2762 71776 2778 71840
rect 2842 71776 2858 71840
rect 2922 71776 2931 71840
rect 2610 70752 2931 71776
rect 2610 70688 2618 70752
rect 2682 70688 2698 70752
rect 2762 70688 2778 70752
rect 2842 70688 2858 70752
rect 2922 70688 2931 70752
rect 2610 69664 2931 70688
rect 2610 69600 2618 69664
rect 2682 69600 2698 69664
rect 2762 69600 2778 69664
rect 2842 69600 2858 69664
rect 2922 69600 2931 69664
rect 2610 68576 2931 69600
rect 2610 68512 2618 68576
rect 2682 68512 2698 68576
rect 2762 68512 2778 68576
rect 2842 68512 2858 68576
rect 2922 68512 2931 68576
rect 2610 67488 2931 68512
rect 2610 67424 2618 67488
rect 2682 67424 2698 67488
rect 2762 67424 2778 67488
rect 2842 67424 2858 67488
rect 2922 67424 2931 67488
rect 2610 66400 2931 67424
rect 2610 66336 2618 66400
rect 2682 66336 2698 66400
rect 2762 66336 2778 66400
rect 2842 66336 2858 66400
rect 2922 66336 2931 66400
rect 2610 65312 2931 66336
rect 2610 65248 2618 65312
rect 2682 65248 2698 65312
rect 2762 65248 2778 65312
rect 2842 65248 2858 65312
rect 2922 65248 2931 65312
rect 2610 64224 2931 65248
rect 2610 64160 2618 64224
rect 2682 64160 2698 64224
rect 2762 64160 2778 64224
rect 2842 64160 2858 64224
rect 2922 64160 2931 64224
rect 2610 63136 2931 64160
rect 2610 63072 2618 63136
rect 2682 63072 2698 63136
rect 2762 63072 2778 63136
rect 2842 63072 2858 63136
rect 2922 63072 2931 63136
rect 2610 62048 2931 63072
rect 2610 61984 2618 62048
rect 2682 61984 2698 62048
rect 2762 61984 2778 62048
rect 2842 61984 2858 62048
rect 2922 61984 2931 62048
rect 2610 60960 2931 61984
rect 2610 60896 2618 60960
rect 2682 60896 2698 60960
rect 2762 60896 2778 60960
rect 2842 60896 2858 60960
rect 2922 60896 2931 60960
rect 2610 59872 2931 60896
rect 2610 59808 2618 59872
rect 2682 59808 2698 59872
rect 2762 59808 2778 59872
rect 2842 59808 2858 59872
rect 2922 59808 2931 59872
rect 2610 58784 2931 59808
rect 2610 58720 2618 58784
rect 2682 58720 2698 58784
rect 2762 58720 2778 58784
rect 2842 58720 2858 58784
rect 2922 58720 2931 58784
rect 2610 57696 2931 58720
rect 2610 57632 2618 57696
rect 2682 57632 2698 57696
rect 2762 57632 2778 57696
rect 2842 57632 2858 57696
rect 2922 57632 2931 57696
rect 2610 56608 2931 57632
rect 2610 56544 2618 56608
rect 2682 56544 2698 56608
rect 2762 56544 2778 56608
rect 2842 56544 2858 56608
rect 2922 56544 2931 56608
rect 2610 55520 2931 56544
rect 2610 55456 2618 55520
rect 2682 55456 2698 55520
rect 2762 55456 2778 55520
rect 2842 55456 2858 55520
rect 2922 55456 2931 55520
rect 2610 54432 2931 55456
rect 2610 54368 2618 54432
rect 2682 54368 2698 54432
rect 2762 54368 2778 54432
rect 2842 54368 2858 54432
rect 2922 54368 2931 54432
rect 2610 53344 2931 54368
rect 2610 53280 2618 53344
rect 2682 53280 2698 53344
rect 2762 53280 2778 53344
rect 2842 53280 2858 53344
rect 2922 53280 2931 53344
rect 2610 52256 2931 53280
rect 2610 52192 2618 52256
rect 2682 52192 2698 52256
rect 2762 52192 2778 52256
rect 2842 52192 2858 52256
rect 2922 52192 2931 52256
rect 2610 51168 2931 52192
rect 2610 51104 2618 51168
rect 2682 51104 2698 51168
rect 2762 51104 2778 51168
rect 2842 51104 2858 51168
rect 2922 51104 2931 51168
rect 2610 50080 2931 51104
rect 2610 50016 2618 50080
rect 2682 50016 2698 50080
rect 2762 50016 2778 50080
rect 2842 50016 2858 50080
rect 2922 50016 2931 50080
rect 2610 48992 2931 50016
rect 2610 48928 2618 48992
rect 2682 48928 2698 48992
rect 2762 48928 2778 48992
rect 2842 48928 2858 48992
rect 2922 48928 2931 48992
rect 2610 47904 2931 48928
rect 2610 47840 2618 47904
rect 2682 47840 2698 47904
rect 2762 47840 2778 47904
rect 2842 47840 2858 47904
rect 2922 47840 2931 47904
rect 2610 46816 2931 47840
rect 2610 46752 2618 46816
rect 2682 46752 2698 46816
rect 2762 46752 2778 46816
rect 2842 46752 2858 46816
rect 2922 46752 2931 46816
rect 2610 45728 2931 46752
rect 2610 45664 2618 45728
rect 2682 45664 2698 45728
rect 2762 45664 2778 45728
rect 2842 45664 2858 45728
rect 2922 45664 2931 45728
rect 2610 44640 2931 45664
rect 2610 44576 2618 44640
rect 2682 44576 2698 44640
rect 2762 44576 2778 44640
rect 2842 44576 2858 44640
rect 2922 44576 2931 44640
rect 2610 43552 2931 44576
rect 2610 43488 2618 43552
rect 2682 43488 2698 43552
rect 2762 43488 2778 43552
rect 2842 43488 2858 43552
rect 2922 43488 2931 43552
rect 2610 42464 2931 43488
rect 2610 42400 2618 42464
rect 2682 42400 2698 42464
rect 2762 42400 2778 42464
rect 2842 42400 2858 42464
rect 2922 42400 2931 42464
rect 2610 41376 2931 42400
rect 2610 41312 2618 41376
rect 2682 41312 2698 41376
rect 2762 41312 2778 41376
rect 2842 41312 2858 41376
rect 2922 41312 2931 41376
rect 2610 40288 2931 41312
rect 2610 40224 2618 40288
rect 2682 40224 2698 40288
rect 2762 40224 2778 40288
rect 2842 40224 2858 40288
rect 2922 40224 2931 40288
rect 2610 39200 2931 40224
rect 2610 39136 2618 39200
rect 2682 39136 2698 39200
rect 2762 39136 2778 39200
rect 2842 39136 2858 39200
rect 2922 39136 2931 39200
rect 2610 38112 2931 39136
rect 2610 38048 2618 38112
rect 2682 38048 2698 38112
rect 2762 38048 2778 38112
rect 2842 38048 2858 38112
rect 2922 38048 2931 38112
rect 2610 37024 2931 38048
rect 2610 36960 2618 37024
rect 2682 36960 2698 37024
rect 2762 36960 2778 37024
rect 2842 36960 2858 37024
rect 2922 36960 2931 37024
rect 2610 35936 2931 36960
rect 2610 35872 2618 35936
rect 2682 35872 2698 35936
rect 2762 35872 2778 35936
rect 2842 35872 2858 35936
rect 2922 35872 2931 35936
rect 2610 34848 2931 35872
rect 2610 34784 2618 34848
rect 2682 34784 2698 34848
rect 2762 34784 2778 34848
rect 2842 34784 2858 34848
rect 2922 34784 2931 34848
rect 2610 33760 2931 34784
rect 2610 33696 2618 33760
rect 2682 33696 2698 33760
rect 2762 33696 2778 33760
rect 2842 33696 2858 33760
rect 2922 33696 2931 33760
rect 2610 32672 2931 33696
rect 2610 32608 2618 32672
rect 2682 32608 2698 32672
rect 2762 32608 2778 32672
rect 2842 32608 2858 32672
rect 2922 32608 2931 32672
rect 2610 31584 2931 32608
rect 2610 31520 2618 31584
rect 2682 31520 2698 31584
rect 2762 31520 2778 31584
rect 2842 31520 2858 31584
rect 2922 31520 2931 31584
rect 2610 30496 2931 31520
rect 2610 30432 2618 30496
rect 2682 30432 2698 30496
rect 2762 30432 2778 30496
rect 2842 30432 2858 30496
rect 2922 30432 2931 30496
rect 2610 29408 2931 30432
rect 2610 29344 2618 29408
rect 2682 29344 2698 29408
rect 2762 29344 2778 29408
rect 2842 29344 2858 29408
rect 2922 29344 2931 29408
rect 2610 28320 2931 29344
rect 2610 28256 2618 28320
rect 2682 28256 2698 28320
rect 2762 28256 2778 28320
rect 2842 28256 2858 28320
rect 2922 28256 2931 28320
rect 2610 27232 2931 28256
rect 2610 27168 2618 27232
rect 2682 27168 2698 27232
rect 2762 27168 2778 27232
rect 2842 27168 2858 27232
rect 2922 27168 2931 27232
rect 2610 26144 2931 27168
rect 2610 26080 2618 26144
rect 2682 26080 2698 26144
rect 2762 26080 2778 26144
rect 2842 26080 2858 26144
rect 2922 26080 2931 26144
rect 2610 25056 2931 26080
rect 2610 24992 2618 25056
rect 2682 24992 2698 25056
rect 2762 24992 2778 25056
rect 2842 24992 2858 25056
rect 2922 24992 2931 25056
rect 2610 23968 2931 24992
rect 2610 23904 2618 23968
rect 2682 23904 2698 23968
rect 2762 23904 2778 23968
rect 2842 23904 2858 23968
rect 2922 23904 2931 23968
rect 2610 22880 2931 23904
rect 2610 22816 2618 22880
rect 2682 22816 2698 22880
rect 2762 22816 2778 22880
rect 2842 22816 2858 22880
rect 2922 22816 2931 22880
rect 2610 21792 2931 22816
rect 2610 21728 2618 21792
rect 2682 21728 2698 21792
rect 2762 21728 2778 21792
rect 2842 21728 2858 21792
rect 2922 21728 2931 21792
rect 2610 20704 2931 21728
rect 2610 20640 2618 20704
rect 2682 20640 2698 20704
rect 2762 20640 2778 20704
rect 2842 20640 2858 20704
rect 2922 20640 2931 20704
rect 2610 19616 2931 20640
rect 2610 19552 2618 19616
rect 2682 19552 2698 19616
rect 2762 19552 2778 19616
rect 2842 19552 2858 19616
rect 2922 19552 2931 19616
rect 2610 18528 2931 19552
rect 2610 18464 2618 18528
rect 2682 18464 2698 18528
rect 2762 18464 2778 18528
rect 2842 18464 2858 18528
rect 2922 18464 2931 18528
rect 2610 17440 2931 18464
rect 2610 17376 2618 17440
rect 2682 17376 2698 17440
rect 2762 17376 2778 17440
rect 2842 17376 2858 17440
rect 2922 17376 2931 17440
rect 2610 16352 2931 17376
rect 2610 16288 2618 16352
rect 2682 16288 2698 16352
rect 2762 16288 2778 16352
rect 2842 16288 2858 16352
rect 2922 16288 2931 16352
rect 2610 15264 2931 16288
rect 2610 15200 2618 15264
rect 2682 15200 2698 15264
rect 2762 15200 2778 15264
rect 2842 15200 2858 15264
rect 2922 15200 2931 15264
rect 2610 14176 2931 15200
rect 2610 14112 2618 14176
rect 2682 14112 2698 14176
rect 2762 14112 2778 14176
rect 2842 14112 2858 14176
rect 2922 14112 2931 14176
rect 2610 13088 2931 14112
rect 2610 13024 2618 13088
rect 2682 13024 2698 13088
rect 2762 13024 2778 13088
rect 2842 13024 2858 13088
rect 2922 13024 2931 13088
rect 2610 12000 2931 13024
rect 2610 11936 2618 12000
rect 2682 11936 2698 12000
rect 2762 11936 2778 12000
rect 2842 11936 2858 12000
rect 2922 11936 2931 12000
rect 2610 10912 2931 11936
rect 2610 10848 2618 10912
rect 2682 10848 2698 10912
rect 2762 10848 2778 10912
rect 2842 10848 2858 10912
rect 2922 10848 2931 10912
rect 2610 9824 2931 10848
rect 2610 9760 2618 9824
rect 2682 9760 2698 9824
rect 2762 9760 2778 9824
rect 2842 9760 2858 9824
rect 2922 9760 2931 9824
rect 2610 8736 2931 9760
rect 2610 8672 2618 8736
rect 2682 8672 2698 8736
rect 2762 8672 2778 8736
rect 2842 8672 2858 8736
rect 2922 8672 2931 8736
rect 2610 7648 2931 8672
rect 2610 7584 2618 7648
rect 2682 7584 2698 7648
rect 2762 7584 2778 7648
rect 2842 7584 2858 7648
rect 2922 7584 2931 7648
rect 2610 6560 2931 7584
rect 2610 6496 2618 6560
rect 2682 6496 2698 6560
rect 2762 6496 2778 6560
rect 2842 6496 2858 6560
rect 2922 6496 2931 6560
rect 2610 5472 2931 6496
rect 2610 5408 2618 5472
rect 2682 5408 2698 5472
rect 2762 5408 2778 5472
rect 2842 5408 2858 5472
rect 2922 5408 2931 5472
rect 2610 4384 2931 5408
rect 2610 4320 2618 4384
rect 2682 4320 2698 4384
rect 2762 4320 2778 4384
rect 2842 4320 2858 4384
rect 2922 4320 2931 4384
rect 2610 3296 2931 4320
rect 2610 3232 2618 3296
rect 2682 3232 2698 3296
rect 2762 3232 2778 3296
rect 2842 3232 2858 3296
rect 2922 3232 2931 3296
rect 2610 2208 2931 3232
rect 2610 2144 2618 2208
rect 2682 2144 2698 2208
rect 2762 2144 2778 2208
rect 2842 2144 2858 2208
rect 2922 2144 2931 2208
rect 2610 2128 2931 2144
rect 4277 330240 4597 330800
rect 4277 330176 4285 330240
rect 4349 330176 4365 330240
rect 4429 330176 4445 330240
rect 4509 330176 4525 330240
rect 4589 330176 4597 330240
rect 4277 329152 4597 330176
rect 4277 329088 4285 329152
rect 4349 329088 4365 329152
rect 4429 329088 4445 329152
rect 4509 329088 4525 329152
rect 4589 329088 4597 329152
rect 4277 328064 4597 329088
rect 4277 328000 4285 328064
rect 4349 328000 4365 328064
rect 4429 328000 4445 328064
rect 4509 328000 4525 328064
rect 4589 328000 4597 328064
rect 4277 326976 4597 328000
rect 4277 326912 4285 326976
rect 4349 326912 4365 326976
rect 4429 326912 4445 326976
rect 4509 326912 4525 326976
rect 4589 326912 4597 326976
rect 4277 325888 4597 326912
rect 4277 325824 4285 325888
rect 4349 325824 4365 325888
rect 4429 325824 4445 325888
rect 4509 325824 4525 325888
rect 4589 325824 4597 325888
rect 4277 324800 4597 325824
rect 4277 324736 4285 324800
rect 4349 324736 4365 324800
rect 4429 324736 4445 324800
rect 4509 324736 4525 324800
rect 4589 324736 4597 324800
rect 4277 323712 4597 324736
rect 4277 323648 4285 323712
rect 4349 323648 4365 323712
rect 4429 323648 4445 323712
rect 4509 323648 4525 323712
rect 4589 323648 4597 323712
rect 4277 322624 4597 323648
rect 4277 322560 4285 322624
rect 4349 322560 4365 322624
rect 4429 322560 4445 322624
rect 4509 322560 4525 322624
rect 4589 322560 4597 322624
rect 4277 321536 4597 322560
rect 4277 321472 4285 321536
rect 4349 321472 4365 321536
rect 4429 321472 4445 321536
rect 4509 321472 4525 321536
rect 4589 321472 4597 321536
rect 4277 320448 4597 321472
rect 4277 320384 4285 320448
rect 4349 320384 4365 320448
rect 4429 320384 4445 320448
rect 4509 320384 4525 320448
rect 4589 320384 4597 320448
rect 4277 319360 4597 320384
rect 4277 319296 4285 319360
rect 4349 319296 4365 319360
rect 4429 319296 4445 319360
rect 4509 319296 4525 319360
rect 4589 319296 4597 319360
rect 4277 318272 4597 319296
rect 4277 318208 4285 318272
rect 4349 318208 4365 318272
rect 4429 318208 4445 318272
rect 4509 318208 4525 318272
rect 4589 318208 4597 318272
rect 4277 317184 4597 318208
rect 4277 317120 4285 317184
rect 4349 317120 4365 317184
rect 4429 317120 4445 317184
rect 4509 317120 4525 317184
rect 4589 317120 4597 317184
rect 4277 316096 4597 317120
rect 4277 316032 4285 316096
rect 4349 316032 4365 316096
rect 4429 316032 4445 316096
rect 4509 316032 4525 316096
rect 4589 316032 4597 316096
rect 4277 315008 4597 316032
rect 4277 314944 4285 315008
rect 4349 314944 4365 315008
rect 4429 314944 4445 315008
rect 4509 314944 4525 315008
rect 4589 314944 4597 315008
rect 4277 313920 4597 314944
rect 4277 313856 4285 313920
rect 4349 313856 4365 313920
rect 4429 313856 4445 313920
rect 4509 313856 4525 313920
rect 4589 313856 4597 313920
rect 4277 312832 4597 313856
rect 4277 312768 4285 312832
rect 4349 312768 4365 312832
rect 4429 312768 4445 312832
rect 4509 312768 4525 312832
rect 4589 312768 4597 312832
rect 4277 311744 4597 312768
rect 4277 311680 4285 311744
rect 4349 311680 4365 311744
rect 4429 311680 4445 311744
rect 4509 311680 4525 311744
rect 4589 311680 4597 311744
rect 4277 310656 4597 311680
rect 4277 310592 4285 310656
rect 4349 310592 4365 310656
rect 4429 310592 4445 310656
rect 4509 310592 4525 310656
rect 4589 310592 4597 310656
rect 4277 309568 4597 310592
rect 4277 309504 4285 309568
rect 4349 309504 4365 309568
rect 4429 309504 4445 309568
rect 4509 309504 4525 309568
rect 4589 309504 4597 309568
rect 4277 308480 4597 309504
rect 4277 308416 4285 308480
rect 4349 308416 4365 308480
rect 4429 308416 4445 308480
rect 4509 308416 4525 308480
rect 4589 308416 4597 308480
rect 4277 307392 4597 308416
rect 4277 307328 4285 307392
rect 4349 307328 4365 307392
rect 4429 307328 4445 307392
rect 4509 307328 4525 307392
rect 4589 307328 4597 307392
rect 4277 306304 4597 307328
rect 4277 306240 4285 306304
rect 4349 306240 4365 306304
rect 4429 306240 4445 306304
rect 4509 306240 4525 306304
rect 4589 306240 4597 306304
rect 4277 305216 4597 306240
rect 4277 305152 4285 305216
rect 4349 305152 4365 305216
rect 4429 305152 4445 305216
rect 4509 305152 4525 305216
rect 4589 305152 4597 305216
rect 4277 304128 4597 305152
rect 4277 304064 4285 304128
rect 4349 304064 4365 304128
rect 4429 304064 4445 304128
rect 4509 304064 4525 304128
rect 4589 304064 4597 304128
rect 4277 303040 4597 304064
rect 4277 302976 4285 303040
rect 4349 302976 4365 303040
rect 4429 302976 4445 303040
rect 4509 302976 4525 303040
rect 4589 302976 4597 303040
rect 4277 301952 4597 302976
rect 4277 301888 4285 301952
rect 4349 301888 4365 301952
rect 4429 301888 4445 301952
rect 4509 301888 4525 301952
rect 4589 301888 4597 301952
rect 4277 300864 4597 301888
rect 4277 300800 4285 300864
rect 4349 300800 4365 300864
rect 4429 300800 4445 300864
rect 4509 300800 4525 300864
rect 4589 300800 4597 300864
rect 4277 299776 4597 300800
rect 4277 299712 4285 299776
rect 4349 299712 4365 299776
rect 4429 299712 4445 299776
rect 4509 299712 4525 299776
rect 4589 299712 4597 299776
rect 4277 298688 4597 299712
rect 4277 298624 4285 298688
rect 4349 298624 4365 298688
rect 4429 298624 4445 298688
rect 4509 298624 4525 298688
rect 4589 298624 4597 298688
rect 4277 297600 4597 298624
rect 4277 297536 4285 297600
rect 4349 297536 4365 297600
rect 4429 297536 4445 297600
rect 4509 297536 4525 297600
rect 4589 297536 4597 297600
rect 4277 296512 4597 297536
rect 4277 296448 4285 296512
rect 4349 296448 4365 296512
rect 4429 296448 4445 296512
rect 4509 296448 4525 296512
rect 4589 296448 4597 296512
rect 4277 295424 4597 296448
rect 4277 295360 4285 295424
rect 4349 295360 4365 295424
rect 4429 295360 4445 295424
rect 4509 295360 4525 295424
rect 4589 295360 4597 295424
rect 4277 294336 4597 295360
rect 4277 294272 4285 294336
rect 4349 294272 4365 294336
rect 4429 294272 4445 294336
rect 4509 294272 4525 294336
rect 4589 294272 4597 294336
rect 4277 293248 4597 294272
rect 4277 293184 4285 293248
rect 4349 293184 4365 293248
rect 4429 293184 4445 293248
rect 4509 293184 4525 293248
rect 4589 293184 4597 293248
rect 4277 292160 4597 293184
rect 4277 292096 4285 292160
rect 4349 292096 4365 292160
rect 4429 292096 4445 292160
rect 4509 292096 4525 292160
rect 4589 292096 4597 292160
rect 4277 291072 4597 292096
rect 4277 291008 4285 291072
rect 4349 291008 4365 291072
rect 4429 291008 4445 291072
rect 4509 291008 4525 291072
rect 4589 291008 4597 291072
rect 4277 289984 4597 291008
rect 4277 289920 4285 289984
rect 4349 289920 4365 289984
rect 4429 289920 4445 289984
rect 4509 289920 4525 289984
rect 4589 289920 4597 289984
rect 4277 288896 4597 289920
rect 4277 288832 4285 288896
rect 4349 288832 4365 288896
rect 4429 288832 4445 288896
rect 4509 288832 4525 288896
rect 4589 288832 4597 288896
rect 4277 287808 4597 288832
rect 4277 287744 4285 287808
rect 4349 287744 4365 287808
rect 4429 287744 4445 287808
rect 4509 287744 4525 287808
rect 4589 287744 4597 287808
rect 4277 286720 4597 287744
rect 4277 286656 4285 286720
rect 4349 286656 4365 286720
rect 4429 286656 4445 286720
rect 4509 286656 4525 286720
rect 4589 286656 4597 286720
rect 4277 285632 4597 286656
rect 4277 285568 4285 285632
rect 4349 285568 4365 285632
rect 4429 285568 4445 285632
rect 4509 285568 4525 285632
rect 4589 285568 4597 285632
rect 4277 284544 4597 285568
rect 4277 284480 4285 284544
rect 4349 284480 4365 284544
rect 4429 284480 4445 284544
rect 4509 284480 4525 284544
rect 4589 284480 4597 284544
rect 4277 283456 4597 284480
rect 4277 283392 4285 283456
rect 4349 283392 4365 283456
rect 4429 283392 4445 283456
rect 4509 283392 4525 283456
rect 4589 283392 4597 283456
rect 4277 282368 4597 283392
rect 4277 282304 4285 282368
rect 4349 282304 4365 282368
rect 4429 282304 4445 282368
rect 4509 282304 4525 282368
rect 4589 282304 4597 282368
rect 4277 281280 4597 282304
rect 4277 281216 4285 281280
rect 4349 281216 4365 281280
rect 4429 281216 4445 281280
rect 4509 281216 4525 281280
rect 4589 281216 4597 281280
rect 4277 280192 4597 281216
rect 4277 280128 4285 280192
rect 4349 280128 4365 280192
rect 4429 280128 4445 280192
rect 4509 280128 4525 280192
rect 4589 280128 4597 280192
rect 4277 279104 4597 280128
rect 4277 279040 4285 279104
rect 4349 279040 4365 279104
rect 4429 279040 4445 279104
rect 4509 279040 4525 279104
rect 4589 279040 4597 279104
rect 4277 278016 4597 279040
rect 4277 277952 4285 278016
rect 4349 277952 4365 278016
rect 4429 277952 4445 278016
rect 4509 277952 4525 278016
rect 4589 277952 4597 278016
rect 4277 276928 4597 277952
rect 4277 276864 4285 276928
rect 4349 276864 4365 276928
rect 4429 276864 4445 276928
rect 4509 276864 4525 276928
rect 4589 276864 4597 276928
rect 4277 275840 4597 276864
rect 4277 275776 4285 275840
rect 4349 275776 4365 275840
rect 4429 275776 4445 275840
rect 4509 275776 4525 275840
rect 4589 275776 4597 275840
rect 4277 274752 4597 275776
rect 4277 274688 4285 274752
rect 4349 274688 4365 274752
rect 4429 274688 4445 274752
rect 4509 274688 4525 274752
rect 4589 274688 4597 274752
rect 4277 273664 4597 274688
rect 4277 273600 4285 273664
rect 4349 273600 4365 273664
rect 4429 273600 4445 273664
rect 4509 273600 4525 273664
rect 4589 273600 4597 273664
rect 4277 272576 4597 273600
rect 4277 272512 4285 272576
rect 4349 272512 4365 272576
rect 4429 272512 4445 272576
rect 4509 272512 4525 272576
rect 4589 272512 4597 272576
rect 4277 271488 4597 272512
rect 4277 271424 4285 271488
rect 4349 271424 4365 271488
rect 4429 271424 4445 271488
rect 4509 271424 4525 271488
rect 4589 271424 4597 271488
rect 4277 270400 4597 271424
rect 4277 270336 4285 270400
rect 4349 270336 4365 270400
rect 4429 270336 4445 270400
rect 4509 270336 4525 270400
rect 4589 270336 4597 270400
rect 4277 269312 4597 270336
rect 4277 269248 4285 269312
rect 4349 269248 4365 269312
rect 4429 269248 4445 269312
rect 4509 269248 4525 269312
rect 4589 269248 4597 269312
rect 4277 268224 4597 269248
rect 4277 268160 4285 268224
rect 4349 268160 4365 268224
rect 4429 268160 4445 268224
rect 4509 268160 4525 268224
rect 4589 268160 4597 268224
rect 4277 267136 4597 268160
rect 4277 267072 4285 267136
rect 4349 267072 4365 267136
rect 4429 267072 4445 267136
rect 4509 267072 4525 267136
rect 4589 267072 4597 267136
rect 4277 266048 4597 267072
rect 4277 265984 4285 266048
rect 4349 265984 4365 266048
rect 4429 265984 4445 266048
rect 4509 265984 4525 266048
rect 4589 265984 4597 266048
rect 4277 264960 4597 265984
rect 4277 264896 4285 264960
rect 4349 264896 4365 264960
rect 4429 264896 4445 264960
rect 4509 264896 4525 264960
rect 4589 264896 4597 264960
rect 4277 263872 4597 264896
rect 4277 263808 4285 263872
rect 4349 263808 4365 263872
rect 4429 263808 4445 263872
rect 4509 263808 4525 263872
rect 4589 263808 4597 263872
rect 4277 262784 4597 263808
rect 4277 262720 4285 262784
rect 4349 262720 4365 262784
rect 4429 262720 4445 262784
rect 4509 262720 4525 262784
rect 4589 262720 4597 262784
rect 4277 261696 4597 262720
rect 4277 261632 4285 261696
rect 4349 261632 4365 261696
rect 4429 261632 4445 261696
rect 4509 261632 4525 261696
rect 4589 261632 4597 261696
rect 4277 260608 4597 261632
rect 4277 260544 4285 260608
rect 4349 260544 4365 260608
rect 4429 260544 4445 260608
rect 4509 260544 4525 260608
rect 4589 260544 4597 260608
rect 4277 259520 4597 260544
rect 4277 259456 4285 259520
rect 4349 259456 4365 259520
rect 4429 259456 4445 259520
rect 4509 259456 4525 259520
rect 4589 259456 4597 259520
rect 4277 258432 4597 259456
rect 4277 258368 4285 258432
rect 4349 258368 4365 258432
rect 4429 258368 4445 258432
rect 4509 258368 4525 258432
rect 4589 258368 4597 258432
rect 4277 257344 4597 258368
rect 4277 257280 4285 257344
rect 4349 257280 4365 257344
rect 4429 257280 4445 257344
rect 4509 257280 4525 257344
rect 4589 257280 4597 257344
rect 4277 256256 4597 257280
rect 4277 256192 4285 256256
rect 4349 256192 4365 256256
rect 4429 256192 4445 256256
rect 4509 256192 4525 256256
rect 4589 256192 4597 256256
rect 4277 255168 4597 256192
rect 4277 255104 4285 255168
rect 4349 255104 4365 255168
rect 4429 255104 4445 255168
rect 4509 255104 4525 255168
rect 4589 255104 4597 255168
rect 4277 254080 4597 255104
rect 4277 254016 4285 254080
rect 4349 254016 4365 254080
rect 4429 254016 4445 254080
rect 4509 254016 4525 254080
rect 4589 254016 4597 254080
rect 4277 252992 4597 254016
rect 4277 252928 4285 252992
rect 4349 252928 4365 252992
rect 4429 252928 4445 252992
rect 4509 252928 4525 252992
rect 4589 252928 4597 252992
rect 4277 251904 4597 252928
rect 4277 251840 4285 251904
rect 4349 251840 4365 251904
rect 4429 251840 4445 251904
rect 4509 251840 4525 251904
rect 4589 251840 4597 251904
rect 4277 250816 4597 251840
rect 4277 250752 4285 250816
rect 4349 250752 4365 250816
rect 4429 250752 4445 250816
rect 4509 250752 4525 250816
rect 4589 250752 4597 250816
rect 4277 249728 4597 250752
rect 4277 249664 4285 249728
rect 4349 249664 4365 249728
rect 4429 249664 4445 249728
rect 4509 249664 4525 249728
rect 4589 249664 4597 249728
rect 4277 248640 4597 249664
rect 4277 248576 4285 248640
rect 4349 248576 4365 248640
rect 4429 248576 4445 248640
rect 4509 248576 4525 248640
rect 4589 248576 4597 248640
rect 4277 247552 4597 248576
rect 4277 247488 4285 247552
rect 4349 247488 4365 247552
rect 4429 247488 4445 247552
rect 4509 247488 4525 247552
rect 4589 247488 4597 247552
rect 4277 246464 4597 247488
rect 4277 246400 4285 246464
rect 4349 246400 4365 246464
rect 4429 246400 4445 246464
rect 4509 246400 4525 246464
rect 4589 246400 4597 246464
rect 4277 245376 4597 246400
rect 4277 245312 4285 245376
rect 4349 245312 4365 245376
rect 4429 245312 4445 245376
rect 4509 245312 4525 245376
rect 4589 245312 4597 245376
rect 4277 244288 4597 245312
rect 4277 244224 4285 244288
rect 4349 244224 4365 244288
rect 4429 244224 4445 244288
rect 4509 244224 4525 244288
rect 4589 244224 4597 244288
rect 4277 243200 4597 244224
rect 4277 243136 4285 243200
rect 4349 243136 4365 243200
rect 4429 243136 4445 243200
rect 4509 243136 4525 243200
rect 4589 243136 4597 243200
rect 4277 242112 4597 243136
rect 4277 242048 4285 242112
rect 4349 242048 4365 242112
rect 4429 242048 4445 242112
rect 4509 242048 4525 242112
rect 4589 242048 4597 242112
rect 4277 241024 4597 242048
rect 4277 240960 4285 241024
rect 4349 240960 4365 241024
rect 4429 240960 4445 241024
rect 4509 240960 4525 241024
rect 4589 240960 4597 241024
rect 4277 239936 4597 240960
rect 4277 239872 4285 239936
rect 4349 239872 4365 239936
rect 4429 239872 4445 239936
rect 4509 239872 4525 239936
rect 4589 239872 4597 239936
rect 4277 238848 4597 239872
rect 4277 238784 4285 238848
rect 4349 238784 4365 238848
rect 4429 238784 4445 238848
rect 4509 238784 4525 238848
rect 4589 238784 4597 238848
rect 4277 237760 4597 238784
rect 4277 237696 4285 237760
rect 4349 237696 4365 237760
rect 4429 237696 4445 237760
rect 4509 237696 4525 237760
rect 4589 237696 4597 237760
rect 4277 236672 4597 237696
rect 4277 236608 4285 236672
rect 4349 236608 4365 236672
rect 4429 236608 4445 236672
rect 4509 236608 4525 236672
rect 4589 236608 4597 236672
rect 4277 235584 4597 236608
rect 4277 235520 4285 235584
rect 4349 235520 4365 235584
rect 4429 235520 4445 235584
rect 4509 235520 4525 235584
rect 4589 235520 4597 235584
rect 4277 234496 4597 235520
rect 4277 234432 4285 234496
rect 4349 234432 4365 234496
rect 4429 234432 4445 234496
rect 4509 234432 4525 234496
rect 4589 234432 4597 234496
rect 4277 233408 4597 234432
rect 4277 233344 4285 233408
rect 4349 233344 4365 233408
rect 4429 233344 4445 233408
rect 4509 233344 4525 233408
rect 4589 233344 4597 233408
rect 4277 232320 4597 233344
rect 4277 232256 4285 232320
rect 4349 232256 4365 232320
rect 4429 232256 4445 232320
rect 4509 232256 4525 232320
rect 4589 232256 4597 232320
rect 4277 231232 4597 232256
rect 4277 231168 4285 231232
rect 4349 231168 4365 231232
rect 4429 231168 4445 231232
rect 4509 231168 4525 231232
rect 4589 231168 4597 231232
rect 4277 230144 4597 231168
rect 4277 230080 4285 230144
rect 4349 230080 4365 230144
rect 4429 230080 4445 230144
rect 4509 230080 4525 230144
rect 4589 230080 4597 230144
rect 4277 229056 4597 230080
rect 4277 228992 4285 229056
rect 4349 228992 4365 229056
rect 4429 228992 4445 229056
rect 4509 228992 4525 229056
rect 4589 228992 4597 229056
rect 4277 227968 4597 228992
rect 4277 227904 4285 227968
rect 4349 227904 4365 227968
rect 4429 227904 4445 227968
rect 4509 227904 4525 227968
rect 4589 227904 4597 227968
rect 4277 226880 4597 227904
rect 4277 226816 4285 226880
rect 4349 226816 4365 226880
rect 4429 226816 4445 226880
rect 4509 226816 4525 226880
rect 4589 226816 4597 226880
rect 4277 225792 4597 226816
rect 4277 225728 4285 225792
rect 4349 225728 4365 225792
rect 4429 225728 4445 225792
rect 4509 225728 4525 225792
rect 4589 225728 4597 225792
rect 4277 224704 4597 225728
rect 4277 224640 4285 224704
rect 4349 224640 4365 224704
rect 4429 224640 4445 224704
rect 4509 224640 4525 224704
rect 4589 224640 4597 224704
rect 4277 223616 4597 224640
rect 4277 223552 4285 223616
rect 4349 223552 4365 223616
rect 4429 223552 4445 223616
rect 4509 223552 4525 223616
rect 4589 223552 4597 223616
rect 4277 222528 4597 223552
rect 4277 222464 4285 222528
rect 4349 222464 4365 222528
rect 4429 222464 4445 222528
rect 4509 222464 4525 222528
rect 4589 222464 4597 222528
rect 4277 221440 4597 222464
rect 4277 221376 4285 221440
rect 4349 221376 4365 221440
rect 4429 221376 4445 221440
rect 4509 221376 4525 221440
rect 4589 221376 4597 221440
rect 4277 220352 4597 221376
rect 4277 220288 4285 220352
rect 4349 220288 4365 220352
rect 4429 220288 4445 220352
rect 4509 220288 4525 220352
rect 4589 220288 4597 220352
rect 4277 219264 4597 220288
rect 4277 219200 4285 219264
rect 4349 219200 4365 219264
rect 4429 219200 4445 219264
rect 4509 219200 4525 219264
rect 4589 219200 4597 219264
rect 4277 218176 4597 219200
rect 4277 218112 4285 218176
rect 4349 218112 4365 218176
rect 4429 218112 4445 218176
rect 4509 218112 4525 218176
rect 4589 218112 4597 218176
rect 4277 217088 4597 218112
rect 4277 217024 4285 217088
rect 4349 217024 4365 217088
rect 4429 217024 4445 217088
rect 4509 217024 4525 217088
rect 4589 217024 4597 217088
rect 4277 216000 4597 217024
rect 4277 215936 4285 216000
rect 4349 215936 4365 216000
rect 4429 215936 4445 216000
rect 4509 215936 4525 216000
rect 4589 215936 4597 216000
rect 4277 214912 4597 215936
rect 4277 214848 4285 214912
rect 4349 214848 4365 214912
rect 4429 214848 4445 214912
rect 4509 214848 4525 214912
rect 4589 214848 4597 214912
rect 4277 213824 4597 214848
rect 4277 213760 4285 213824
rect 4349 213760 4365 213824
rect 4429 213760 4445 213824
rect 4509 213760 4525 213824
rect 4589 213760 4597 213824
rect 4277 212736 4597 213760
rect 4277 212672 4285 212736
rect 4349 212672 4365 212736
rect 4429 212672 4445 212736
rect 4509 212672 4525 212736
rect 4589 212672 4597 212736
rect 4277 211648 4597 212672
rect 4277 211584 4285 211648
rect 4349 211584 4365 211648
rect 4429 211584 4445 211648
rect 4509 211584 4525 211648
rect 4589 211584 4597 211648
rect 4277 210560 4597 211584
rect 4277 210496 4285 210560
rect 4349 210496 4365 210560
rect 4429 210496 4445 210560
rect 4509 210496 4525 210560
rect 4589 210496 4597 210560
rect 4277 209472 4597 210496
rect 4277 209408 4285 209472
rect 4349 209408 4365 209472
rect 4429 209408 4445 209472
rect 4509 209408 4525 209472
rect 4589 209408 4597 209472
rect 4277 208384 4597 209408
rect 4277 208320 4285 208384
rect 4349 208320 4365 208384
rect 4429 208320 4445 208384
rect 4509 208320 4525 208384
rect 4589 208320 4597 208384
rect 4277 207296 4597 208320
rect 4277 207232 4285 207296
rect 4349 207232 4365 207296
rect 4429 207232 4445 207296
rect 4509 207232 4525 207296
rect 4589 207232 4597 207296
rect 4277 206208 4597 207232
rect 4277 206144 4285 206208
rect 4349 206144 4365 206208
rect 4429 206144 4445 206208
rect 4509 206144 4525 206208
rect 4589 206144 4597 206208
rect 4277 205120 4597 206144
rect 4277 205056 4285 205120
rect 4349 205056 4365 205120
rect 4429 205056 4445 205120
rect 4509 205056 4525 205120
rect 4589 205056 4597 205120
rect 4277 204032 4597 205056
rect 4277 203968 4285 204032
rect 4349 203968 4365 204032
rect 4429 203968 4445 204032
rect 4509 203968 4525 204032
rect 4589 203968 4597 204032
rect 4277 202944 4597 203968
rect 4277 202880 4285 202944
rect 4349 202880 4365 202944
rect 4429 202880 4445 202944
rect 4509 202880 4525 202944
rect 4589 202880 4597 202944
rect 4277 201856 4597 202880
rect 4277 201792 4285 201856
rect 4349 201792 4365 201856
rect 4429 201792 4445 201856
rect 4509 201792 4525 201856
rect 4589 201792 4597 201856
rect 4277 200768 4597 201792
rect 4277 200704 4285 200768
rect 4349 200704 4365 200768
rect 4429 200704 4445 200768
rect 4509 200704 4525 200768
rect 4589 200704 4597 200768
rect 4277 199680 4597 200704
rect 4277 199616 4285 199680
rect 4349 199616 4365 199680
rect 4429 199616 4445 199680
rect 4509 199616 4525 199680
rect 4589 199616 4597 199680
rect 4277 198592 4597 199616
rect 4277 198528 4285 198592
rect 4349 198528 4365 198592
rect 4429 198528 4445 198592
rect 4509 198528 4525 198592
rect 4589 198528 4597 198592
rect 4277 197504 4597 198528
rect 4277 197440 4285 197504
rect 4349 197440 4365 197504
rect 4429 197440 4445 197504
rect 4509 197440 4525 197504
rect 4589 197440 4597 197504
rect 4277 196416 4597 197440
rect 4277 196352 4285 196416
rect 4349 196352 4365 196416
rect 4429 196352 4445 196416
rect 4509 196352 4525 196416
rect 4589 196352 4597 196416
rect 4277 195328 4597 196352
rect 4277 195264 4285 195328
rect 4349 195264 4365 195328
rect 4429 195264 4445 195328
rect 4509 195264 4525 195328
rect 4589 195264 4597 195328
rect 4277 194240 4597 195264
rect 4277 194176 4285 194240
rect 4349 194176 4365 194240
rect 4429 194176 4445 194240
rect 4509 194176 4525 194240
rect 4589 194176 4597 194240
rect 4277 193152 4597 194176
rect 4277 193088 4285 193152
rect 4349 193088 4365 193152
rect 4429 193088 4445 193152
rect 4509 193088 4525 193152
rect 4589 193088 4597 193152
rect 4277 192064 4597 193088
rect 4277 192000 4285 192064
rect 4349 192000 4365 192064
rect 4429 192000 4445 192064
rect 4509 192000 4525 192064
rect 4589 192000 4597 192064
rect 4277 190976 4597 192000
rect 4277 190912 4285 190976
rect 4349 190912 4365 190976
rect 4429 190912 4445 190976
rect 4509 190912 4525 190976
rect 4589 190912 4597 190976
rect 4277 189888 4597 190912
rect 4277 189824 4285 189888
rect 4349 189824 4365 189888
rect 4429 189824 4445 189888
rect 4509 189824 4525 189888
rect 4589 189824 4597 189888
rect 4277 188800 4597 189824
rect 4277 188736 4285 188800
rect 4349 188736 4365 188800
rect 4429 188736 4445 188800
rect 4509 188736 4525 188800
rect 4589 188736 4597 188800
rect 4277 187712 4597 188736
rect 4277 187648 4285 187712
rect 4349 187648 4365 187712
rect 4429 187648 4445 187712
rect 4509 187648 4525 187712
rect 4589 187648 4597 187712
rect 4277 186624 4597 187648
rect 4277 186560 4285 186624
rect 4349 186560 4365 186624
rect 4429 186560 4445 186624
rect 4509 186560 4525 186624
rect 4589 186560 4597 186624
rect 4277 185536 4597 186560
rect 4277 185472 4285 185536
rect 4349 185472 4365 185536
rect 4429 185472 4445 185536
rect 4509 185472 4525 185536
rect 4589 185472 4597 185536
rect 4277 184448 4597 185472
rect 4277 184384 4285 184448
rect 4349 184384 4365 184448
rect 4429 184384 4445 184448
rect 4509 184384 4525 184448
rect 4589 184384 4597 184448
rect 4277 183360 4597 184384
rect 4277 183296 4285 183360
rect 4349 183296 4365 183360
rect 4429 183296 4445 183360
rect 4509 183296 4525 183360
rect 4589 183296 4597 183360
rect 4277 182272 4597 183296
rect 4277 182208 4285 182272
rect 4349 182208 4365 182272
rect 4429 182208 4445 182272
rect 4509 182208 4525 182272
rect 4589 182208 4597 182272
rect 4277 181184 4597 182208
rect 4277 181120 4285 181184
rect 4349 181120 4365 181184
rect 4429 181120 4445 181184
rect 4509 181120 4525 181184
rect 4589 181120 4597 181184
rect 4277 180096 4597 181120
rect 4277 180032 4285 180096
rect 4349 180032 4365 180096
rect 4429 180032 4445 180096
rect 4509 180032 4525 180096
rect 4589 180032 4597 180096
rect 4277 179008 4597 180032
rect 4277 178944 4285 179008
rect 4349 178944 4365 179008
rect 4429 178944 4445 179008
rect 4509 178944 4525 179008
rect 4589 178944 4597 179008
rect 4277 177920 4597 178944
rect 4277 177856 4285 177920
rect 4349 177856 4365 177920
rect 4429 177856 4445 177920
rect 4509 177856 4525 177920
rect 4589 177856 4597 177920
rect 4277 176832 4597 177856
rect 4277 176768 4285 176832
rect 4349 176768 4365 176832
rect 4429 176768 4445 176832
rect 4509 176768 4525 176832
rect 4589 176768 4597 176832
rect 4277 175744 4597 176768
rect 4277 175680 4285 175744
rect 4349 175680 4365 175744
rect 4429 175680 4445 175744
rect 4509 175680 4525 175744
rect 4589 175680 4597 175744
rect 4277 174656 4597 175680
rect 4277 174592 4285 174656
rect 4349 174592 4365 174656
rect 4429 174592 4445 174656
rect 4509 174592 4525 174656
rect 4589 174592 4597 174656
rect 4277 173568 4597 174592
rect 4277 173504 4285 173568
rect 4349 173504 4365 173568
rect 4429 173504 4445 173568
rect 4509 173504 4525 173568
rect 4589 173504 4597 173568
rect 4277 172480 4597 173504
rect 4277 172416 4285 172480
rect 4349 172416 4365 172480
rect 4429 172416 4445 172480
rect 4509 172416 4525 172480
rect 4589 172416 4597 172480
rect 4277 171392 4597 172416
rect 4277 171328 4285 171392
rect 4349 171328 4365 171392
rect 4429 171328 4445 171392
rect 4509 171328 4525 171392
rect 4589 171328 4597 171392
rect 4277 170304 4597 171328
rect 4277 170240 4285 170304
rect 4349 170240 4365 170304
rect 4429 170240 4445 170304
rect 4509 170240 4525 170304
rect 4589 170240 4597 170304
rect 4277 169216 4597 170240
rect 4277 169152 4285 169216
rect 4349 169152 4365 169216
rect 4429 169152 4445 169216
rect 4509 169152 4525 169216
rect 4589 169152 4597 169216
rect 4277 168128 4597 169152
rect 4277 168064 4285 168128
rect 4349 168064 4365 168128
rect 4429 168064 4445 168128
rect 4509 168064 4525 168128
rect 4589 168064 4597 168128
rect 4277 167040 4597 168064
rect 4277 166976 4285 167040
rect 4349 166976 4365 167040
rect 4429 166976 4445 167040
rect 4509 166976 4525 167040
rect 4589 166976 4597 167040
rect 4277 165952 4597 166976
rect 4277 165888 4285 165952
rect 4349 165888 4365 165952
rect 4429 165888 4445 165952
rect 4509 165888 4525 165952
rect 4589 165888 4597 165952
rect 4277 164864 4597 165888
rect 4277 164800 4285 164864
rect 4349 164800 4365 164864
rect 4429 164800 4445 164864
rect 4509 164800 4525 164864
rect 4589 164800 4597 164864
rect 4277 163776 4597 164800
rect 4277 163712 4285 163776
rect 4349 163712 4365 163776
rect 4429 163712 4445 163776
rect 4509 163712 4525 163776
rect 4589 163712 4597 163776
rect 4277 162688 4597 163712
rect 4277 162624 4285 162688
rect 4349 162624 4365 162688
rect 4429 162624 4445 162688
rect 4509 162624 4525 162688
rect 4589 162624 4597 162688
rect 4277 161600 4597 162624
rect 4277 161536 4285 161600
rect 4349 161536 4365 161600
rect 4429 161536 4445 161600
rect 4509 161536 4525 161600
rect 4589 161536 4597 161600
rect 4277 160512 4597 161536
rect 4277 160448 4285 160512
rect 4349 160448 4365 160512
rect 4429 160448 4445 160512
rect 4509 160448 4525 160512
rect 4589 160448 4597 160512
rect 4277 159424 4597 160448
rect 4277 159360 4285 159424
rect 4349 159360 4365 159424
rect 4429 159360 4445 159424
rect 4509 159360 4525 159424
rect 4589 159360 4597 159424
rect 4277 158336 4597 159360
rect 4277 158272 4285 158336
rect 4349 158272 4365 158336
rect 4429 158272 4445 158336
rect 4509 158272 4525 158336
rect 4589 158272 4597 158336
rect 4277 157248 4597 158272
rect 4277 157184 4285 157248
rect 4349 157184 4365 157248
rect 4429 157184 4445 157248
rect 4509 157184 4525 157248
rect 4589 157184 4597 157248
rect 4277 156160 4597 157184
rect 4277 156096 4285 156160
rect 4349 156096 4365 156160
rect 4429 156096 4445 156160
rect 4509 156096 4525 156160
rect 4589 156096 4597 156160
rect 4277 155072 4597 156096
rect 4277 155008 4285 155072
rect 4349 155008 4365 155072
rect 4429 155008 4445 155072
rect 4509 155008 4525 155072
rect 4589 155008 4597 155072
rect 4277 153984 4597 155008
rect 4277 153920 4285 153984
rect 4349 153920 4365 153984
rect 4429 153920 4445 153984
rect 4509 153920 4525 153984
rect 4589 153920 4597 153984
rect 4277 152896 4597 153920
rect 4277 152832 4285 152896
rect 4349 152832 4365 152896
rect 4429 152832 4445 152896
rect 4509 152832 4525 152896
rect 4589 152832 4597 152896
rect 4277 151808 4597 152832
rect 4277 151744 4285 151808
rect 4349 151744 4365 151808
rect 4429 151744 4445 151808
rect 4509 151744 4525 151808
rect 4589 151744 4597 151808
rect 4277 150720 4597 151744
rect 4277 150656 4285 150720
rect 4349 150656 4365 150720
rect 4429 150656 4445 150720
rect 4509 150656 4525 150720
rect 4589 150656 4597 150720
rect 4277 149632 4597 150656
rect 4277 149568 4285 149632
rect 4349 149568 4365 149632
rect 4429 149568 4445 149632
rect 4509 149568 4525 149632
rect 4589 149568 4597 149632
rect 4277 148544 4597 149568
rect 4277 148480 4285 148544
rect 4349 148480 4365 148544
rect 4429 148480 4445 148544
rect 4509 148480 4525 148544
rect 4589 148480 4597 148544
rect 4277 147456 4597 148480
rect 4277 147392 4285 147456
rect 4349 147392 4365 147456
rect 4429 147392 4445 147456
rect 4509 147392 4525 147456
rect 4589 147392 4597 147456
rect 4277 146368 4597 147392
rect 4277 146304 4285 146368
rect 4349 146304 4365 146368
rect 4429 146304 4445 146368
rect 4509 146304 4525 146368
rect 4589 146304 4597 146368
rect 4277 145280 4597 146304
rect 4277 145216 4285 145280
rect 4349 145216 4365 145280
rect 4429 145216 4445 145280
rect 4509 145216 4525 145280
rect 4589 145216 4597 145280
rect 4277 144192 4597 145216
rect 4277 144128 4285 144192
rect 4349 144128 4365 144192
rect 4429 144128 4445 144192
rect 4509 144128 4525 144192
rect 4589 144128 4597 144192
rect 4277 143104 4597 144128
rect 4277 143040 4285 143104
rect 4349 143040 4365 143104
rect 4429 143040 4445 143104
rect 4509 143040 4525 143104
rect 4589 143040 4597 143104
rect 4277 142016 4597 143040
rect 4277 141952 4285 142016
rect 4349 141952 4365 142016
rect 4429 141952 4445 142016
rect 4509 141952 4525 142016
rect 4589 141952 4597 142016
rect 4277 140928 4597 141952
rect 4277 140864 4285 140928
rect 4349 140864 4365 140928
rect 4429 140864 4445 140928
rect 4509 140864 4525 140928
rect 4589 140864 4597 140928
rect 4277 139840 4597 140864
rect 4277 139776 4285 139840
rect 4349 139776 4365 139840
rect 4429 139776 4445 139840
rect 4509 139776 4525 139840
rect 4589 139776 4597 139840
rect 4277 138752 4597 139776
rect 4277 138688 4285 138752
rect 4349 138688 4365 138752
rect 4429 138688 4445 138752
rect 4509 138688 4525 138752
rect 4589 138688 4597 138752
rect 4277 137664 4597 138688
rect 4277 137600 4285 137664
rect 4349 137600 4365 137664
rect 4429 137600 4445 137664
rect 4509 137600 4525 137664
rect 4589 137600 4597 137664
rect 4277 136576 4597 137600
rect 4277 136512 4285 136576
rect 4349 136512 4365 136576
rect 4429 136512 4445 136576
rect 4509 136512 4525 136576
rect 4589 136512 4597 136576
rect 4277 135488 4597 136512
rect 4277 135424 4285 135488
rect 4349 135424 4365 135488
rect 4429 135424 4445 135488
rect 4509 135424 4525 135488
rect 4589 135424 4597 135488
rect 4277 134400 4597 135424
rect 4277 134336 4285 134400
rect 4349 134336 4365 134400
rect 4429 134336 4445 134400
rect 4509 134336 4525 134400
rect 4589 134336 4597 134400
rect 4277 133312 4597 134336
rect 4277 133248 4285 133312
rect 4349 133248 4365 133312
rect 4429 133248 4445 133312
rect 4509 133248 4525 133312
rect 4589 133248 4597 133312
rect 4277 132224 4597 133248
rect 4277 132160 4285 132224
rect 4349 132160 4365 132224
rect 4429 132160 4445 132224
rect 4509 132160 4525 132224
rect 4589 132160 4597 132224
rect 4277 131136 4597 132160
rect 4277 131072 4285 131136
rect 4349 131072 4365 131136
rect 4429 131072 4445 131136
rect 4509 131072 4525 131136
rect 4589 131072 4597 131136
rect 4277 130048 4597 131072
rect 4277 129984 4285 130048
rect 4349 129984 4365 130048
rect 4429 129984 4445 130048
rect 4509 129984 4525 130048
rect 4589 129984 4597 130048
rect 4277 128960 4597 129984
rect 4277 128896 4285 128960
rect 4349 128896 4365 128960
rect 4429 128896 4445 128960
rect 4509 128896 4525 128960
rect 4589 128896 4597 128960
rect 4277 127872 4597 128896
rect 4277 127808 4285 127872
rect 4349 127808 4365 127872
rect 4429 127808 4445 127872
rect 4509 127808 4525 127872
rect 4589 127808 4597 127872
rect 4277 126784 4597 127808
rect 4277 126720 4285 126784
rect 4349 126720 4365 126784
rect 4429 126720 4445 126784
rect 4509 126720 4525 126784
rect 4589 126720 4597 126784
rect 4277 125696 4597 126720
rect 4277 125632 4285 125696
rect 4349 125632 4365 125696
rect 4429 125632 4445 125696
rect 4509 125632 4525 125696
rect 4589 125632 4597 125696
rect 4277 124608 4597 125632
rect 4277 124544 4285 124608
rect 4349 124544 4365 124608
rect 4429 124544 4445 124608
rect 4509 124544 4525 124608
rect 4589 124544 4597 124608
rect 4277 123520 4597 124544
rect 4277 123456 4285 123520
rect 4349 123456 4365 123520
rect 4429 123456 4445 123520
rect 4509 123456 4525 123520
rect 4589 123456 4597 123520
rect 4277 122432 4597 123456
rect 4277 122368 4285 122432
rect 4349 122368 4365 122432
rect 4429 122368 4445 122432
rect 4509 122368 4525 122432
rect 4589 122368 4597 122432
rect 4277 121344 4597 122368
rect 4277 121280 4285 121344
rect 4349 121280 4365 121344
rect 4429 121280 4445 121344
rect 4509 121280 4525 121344
rect 4589 121280 4597 121344
rect 4277 120256 4597 121280
rect 4277 120192 4285 120256
rect 4349 120192 4365 120256
rect 4429 120192 4445 120256
rect 4509 120192 4525 120256
rect 4589 120192 4597 120256
rect 4277 119168 4597 120192
rect 4277 119104 4285 119168
rect 4349 119104 4365 119168
rect 4429 119104 4445 119168
rect 4509 119104 4525 119168
rect 4589 119104 4597 119168
rect 4277 118080 4597 119104
rect 4277 118016 4285 118080
rect 4349 118016 4365 118080
rect 4429 118016 4445 118080
rect 4509 118016 4525 118080
rect 4589 118016 4597 118080
rect 4277 116992 4597 118016
rect 4277 116928 4285 116992
rect 4349 116928 4365 116992
rect 4429 116928 4445 116992
rect 4509 116928 4525 116992
rect 4589 116928 4597 116992
rect 4277 115904 4597 116928
rect 4277 115840 4285 115904
rect 4349 115840 4365 115904
rect 4429 115840 4445 115904
rect 4509 115840 4525 115904
rect 4589 115840 4597 115904
rect 4277 114816 4597 115840
rect 4277 114752 4285 114816
rect 4349 114752 4365 114816
rect 4429 114752 4445 114816
rect 4509 114752 4525 114816
rect 4589 114752 4597 114816
rect 4277 113728 4597 114752
rect 4277 113664 4285 113728
rect 4349 113664 4365 113728
rect 4429 113664 4445 113728
rect 4509 113664 4525 113728
rect 4589 113664 4597 113728
rect 4277 112640 4597 113664
rect 4277 112576 4285 112640
rect 4349 112576 4365 112640
rect 4429 112576 4445 112640
rect 4509 112576 4525 112640
rect 4589 112576 4597 112640
rect 4277 111552 4597 112576
rect 4277 111488 4285 111552
rect 4349 111488 4365 111552
rect 4429 111488 4445 111552
rect 4509 111488 4525 111552
rect 4589 111488 4597 111552
rect 4277 110464 4597 111488
rect 4277 110400 4285 110464
rect 4349 110400 4365 110464
rect 4429 110400 4445 110464
rect 4509 110400 4525 110464
rect 4589 110400 4597 110464
rect 4277 109376 4597 110400
rect 4277 109312 4285 109376
rect 4349 109312 4365 109376
rect 4429 109312 4445 109376
rect 4509 109312 4525 109376
rect 4589 109312 4597 109376
rect 4277 108288 4597 109312
rect 4277 108224 4285 108288
rect 4349 108224 4365 108288
rect 4429 108224 4445 108288
rect 4509 108224 4525 108288
rect 4589 108224 4597 108288
rect 4277 107200 4597 108224
rect 4277 107136 4285 107200
rect 4349 107136 4365 107200
rect 4429 107136 4445 107200
rect 4509 107136 4525 107200
rect 4589 107136 4597 107200
rect 4277 106112 4597 107136
rect 4277 106048 4285 106112
rect 4349 106048 4365 106112
rect 4429 106048 4445 106112
rect 4509 106048 4525 106112
rect 4589 106048 4597 106112
rect 4277 105024 4597 106048
rect 4277 104960 4285 105024
rect 4349 104960 4365 105024
rect 4429 104960 4445 105024
rect 4509 104960 4525 105024
rect 4589 104960 4597 105024
rect 4277 103936 4597 104960
rect 4277 103872 4285 103936
rect 4349 103872 4365 103936
rect 4429 103872 4445 103936
rect 4509 103872 4525 103936
rect 4589 103872 4597 103936
rect 4277 102848 4597 103872
rect 4277 102784 4285 102848
rect 4349 102784 4365 102848
rect 4429 102784 4445 102848
rect 4509 102784 4525 102848
rect 4589 102784 4597 102848
rect 4277 101760 4597 102784
rect 4277 101696 4285 101760
rect 4349 101696 4365 101760
rect 4429 101696 4445 101760
rect 4509 101696 4525 101760
rect 4589 101696 4597 101760
rect 4277 100672 4597 101696
rect 4277 100608 4285 100672
rect 4349 100608 4365 100672
rect 4429 100608 4445 100672
rect 4509 100608 4525 100672
rect 4589 100608 4597 100672
rect 4277 99584 4597 100608
rect 4277 99520 4285 99584
rect 4349 99520 4365 99584
rect 4429 99520 4445 99584
rect 4509 99520 4525 99584
rect 4589 99520 4597 99584
rect 4277 98496 4597 99520
rect 4277 98432 4285 98496
rect 4349 98432 4365 98496
rect 4429 98432 4445 98496
rect 4509 98432 4525 98496
rect 4589 98432 4597 98496
rect 4277 97408 4597 98432
rect 4277 97344 4285 97408
rect 4349 97344 4365 97408
rect 4429 97344 4445 97408
rect 4509 97344 4525 97408
rect 4589 97344 4597 97408
rect 4277 96320 4597 97344
rect 4277 96256 4285 96320
rect 4349 96256 4365 96320
rect 4429 96256 4445 96320
rect 4509 96256 4525 96320
rect 4589 96256 4597 96320
rect 4277 95232 4597 96256
rect 4277 95168 4285 95232
rect 4349 95168 4365 95232
rect 4429 95168 4445 95232
rect 4509 95168 4525 95232
rect 4589 95168 4597 95232
rect 4277 94144 4597 95168
rect 4277 94080 4285 94144
rect 4349 94080 4365 94144
rect 4429 94080 4445 94144
rect 4509 94080 4525 94144
rect 4589 94080 4597 94144
rect 4277 93056 4597 94080
rect 4277 92992 4285 93056
rect 4349 92992 4365 93056
rect 4429 92992 4445 93056
rect 4509 92992 4525 93056
rect 4589 92992 4597 93056
rect 4277 91968 4597 92992
rect 4277 91904 4285 91968
rect 4349 91904 4365 91968
rect 4429 91904 4445 91968
rect 4509 91904 4525 91968
rect 4589 91904 4597 91968
rect 4277 90880 4597 91904
rect 4277 90816 4285 90880
rect 4349 90816 4365 90880
rect 4429 90816 4445 90880
rect 4509 90816 4525 90880
rect 4589 90816 4597 90880
rect 4277 89792 4597 90816
rect 4277 89728 4285 89792
rect 4349 89728 4365 89792
rect 4429 89728 4445 89792
rect 4509 89728 4525 89792
rect 4589 89728 4597 89792
rect 4277 88704 4597 89728
rect 4277 88640 4285 88704
rect 4349 88640 4365 88704
rect 4429 88640 4445 88704
rect 4509 88640 4525 88704
rect 4589 88640 4597 88704
rect 4277 87616 4597 88640
rect 4277 87552 4285 87616
rect 4349 87552 4365 87616
rect 4429 87552 4445 87616
rect 4509 87552 4525 87616
rect 4589 87552 4597 87616
rect 4277 86528 4597 87552
rect 4277 86464 4285 86528
rect 4349 86464 4365 86528
rect 4429 86464 4445 86528
rect 4509 86464 4525 86528
rect 4589 86464 4597 86528
rect 4277 85440 4597 86464
rect 4277 85376 4285 85440
rect 4349 85376 4365 85440
rect 4429 85376 4445 85440
rect 4509 85376 4525 85440
rect 4589 85376 4597 85440
rect 4277 84352 4597 85376
rect 4277 84288 4285 84352
rect 4349 84288 4365 84352
rect 4429 84288 4445 84352
rect 4509 84288 4525 84352
rect 4589 84288 4597 84352
rect 4277 83264 4597 84288
rect 4277 83200 4285 83264
rect 4349 83200 4365 83264
rect 4429 83200 4445 83264
rect 4509 83200 4525 83264
rect 4589 83200 4597 83264
rect 4277 82176 4597 83200
rect 4277 82112 4285 82176
rect 4349 82112 4365 82176
rect 4429 82112 4445 82176
rect 4509 82112 4525 82176
rect 4589 82112 4597 82176
rect 4277 81088 4597 82112
rect 4277 81024 4285 81088
rect 4349 81024 4365 81088
rect 4429 81024 4445 81088
rect 4509 81024 4525 81088
rect 4589 81024 4597 81088
rect 4277 80000 4597 81024
rect 4277 79936 4285 80000
rect 4349 79936 4365 80000
rect 4429 79936 4445 80000
rect 4509 79936 4525 80000
rect 4589 79936 4597 80000
rect 4277 78912 4597 79936
rect 4277 78848 4285 78912
rect 4349 78848 4365 78912
rect 4429 78848 4445 78912
rect 4509 78848 4525 78912
rect 4589 78848 4597 78912
rect 4277 77824 4597 78848
rect 4277 77760 4285 77824
rect 4349 77760 4365 77824
rect 4429 77760 4445 77824
rect 4509 77760 4525 77824
rect 4589 77760 4597 77824
rect 4277 76736 4597 77760
rect 4277 76672 4285 76736
rect 4349 76672 4365 76736
rect 4429 76672 4445 76736
rect 4509 76672 4525 76736
rect 4589 76672 4597 76736
rect 4277 75648 4597 76672
rect 4277 75584 4285 75648
rect 4349 75584 4365 75648
rect 4429 75584 4445 75648
rect 4509 75584 4525 75648
rect 4589 75584 4597 75648
rect 4277 74560 4597 75584
rect 4277 74496 4285 74560
rect 4349 74496 4365 74560
rect 4429 74496 4445 74560
rect 4509 74496 4525 74560
rect 4589 74496 4597 74560
rect 4277 73472 4597 74496
rect 4277 73408 4285 73472
rect 4349 73408 4365 73472
rect 4429 73408 4445 73472
rect 4509 73408 4525 73472
rect 4589 73408 4597 73472
rect 4277 72384 4597 73408
rect 4277 72320 4285 72384
rect 4349 72320 4365 72384
rect 4429 72320 4445 72384
rect 4509 72320 4525 72384
rect 4589 72320 4597 72384
rect 4277 71296 4597 72320
rect 4277 71232 4285 71296
rect 4349 71232 4365 71296
rect 4429 71232 4445 71296
rect 4509 71232 4525 71296
rect 4589 71232 4597 71296
rect 4277 70208 4597 71232
rect 4277 70144 4285 70208
rect 4349 70144 4365 70208
rect 4429 70144 4445 70208
rect 4509 70144 4525 70208
rect 4589 70144 4597 70208
rect 4277 69120 4597 70144
rect 4277 69056 4285 69120
rect 4349 69056 4365 69120
rect 4429 69056 4445 69120
rect 4509 69056 4525 69120
rect 4589 69056 4597 69120
rect 4277 68032 4597 69056
rect 4277 67968 4285 68032
rect 4349 67968 4365 68032
rect 4429 67968 4445 68032
rect 4509 67968 4525 68032
rect 4589 67968 4597 68032
rect 4277 66944 4597 67968
rect 4277 66880 4285 66944
rect 4349 66880 4365 66944
rect 4429 66880 4445 66944
rect 4509 66880 4525 66944
rect 4589 66880 4597 66944
rect 4277 65856 4597 66880
rect 4277 65792 4285 65856
rect 4349 65792 4365 65856
rect 4429 65792 4445 65856
rect 4509 65792 4525 65856
rect 4589 65792 4597 65856
rect 4277 64768 4597 65792
rect 4277 64704 4285 64768
rect 4349 64704 4365 64768
rect 4429 64704 4445 64768
rect 4509 64704 4525 64768
rect 4589 64704 4597 64768
rect 4277 63680 4597 64704
rect 4277 63616 4285 63680
rect 4349 63616 4365 63680
rect 4429 63616 4445 63680
rect 4509 63616 4525 63680
rect 4589 63616 4597 63680
rect 4277 62592 4597 63616
rect 4277 62528 4285 62592
rect 4349 62528 4365 62592
rect 4429 62528 4445 62592
rect 4509 62528 4525 62592
rect 4589 62528 4597 62592
rect 4277 61504 4597 62528
rect 4277 61440 4285 61504
rect 4349 61440 4365 61504
rect 4429 61440 4445 61504
rect 4509 61440 4525 61504
rect 4589 61440 4597 61504
rect 4277 60416 4597 61440
rect 4277 60352 4285 60416
rect 4349 60352 4365 60416
rect 4429 60352 4445 60416
rect 4509 60352 4525 60416
rect 4589 60352 4597 60416
rect 4277 59328 4597 60352
rect 4277 59264 4285 59328
rect 4349 59264 4365 59328
rect 4429 59264 4445 59328
rect 4509 59264 4525 59328
rect 4589 59264 4597 59328
rect 4277 58240 4597 59264
rect 4277 58176 4285 58240
rect 4349 58176 4365 58240
rect 4429 58176 4445 58240
rect 4509 58176 4525 58240
rect 4589 58176 4597 58240
rect 4277 57152 4597 58176
rect 4277 57088 4285 57152
rect 4349 57088 4365 57152
rect 4429 57088 4445 57152
rect 4509 57088 4525 57152
rect 4589 57088 4597 57152
rect 4277 56064 4597 57088
rect 4277 56000 4285 56064
rect 4349 56000 4365 56064
rect 4429 56000 4445 56064
rect 4509 56000 4525 56064
rect 4589 56000 4597 56064
rect 4277 54976 4597 56000
rect 4277 54912 4285 54976
rect 4349 54912 4365 54976
rect 4429 54912 4445 54976
rect 4509 54912 4525 54976
rect 4589 54912 4597 54976
rect 4277 53888 4597 54912
rect 4277 53824 4285 53888
rect 4349 53824 4365 53888
rect 4429 53824 4445 53888
rect 4509 53824 4525 53888
rect 4589 53824 4597 53888
rect 4277 52800 4597 53824
rect 4277 52736 4285 52800
rect 4349 52736 4365 52800
rect 4429 52736 4445 52800
rect 4509 52736 4525 52800
rect 4589 52736 4597 52800
rect 4277 51712 4597 52736
rect 4277 51648 4285 51712
rect 4349 51648 4365 51712
rect 4429 51648 4445 51712
rect 4509 51648 4525 51712
rect 4589 51648 4597 51712
rect 4277 50624 4597 51648
rect 4277 50560 4285 50624
rect 4349 50560 4365 50624
rect 4429 50560 4445 50624
rect 4509 50560 4525 50624
rect 4589 50560 4597 50624
rect 4277 49536 4597 50560
rect 4277 49472 4285 49536
rect 4349 49472 4365 49536
rect 4429 49472 4445 49536
rect 4509 49472 4525 49536
rect 4589 49472 4597 49536
rect 4277 48448 4597 49472
rect 4277 48384 4285 48448
rect 4349 48384 4365 48448
rect 4429 48384 4445 48448
rect 4509 48384 4525 48448
rect 4589 48384 4597 48448
rect 4277 47360 4597 48384
rect 4277 47296 4285 47360
rect 4349 47296 4365 47360
rect 4429 47296 4445 47360
rect 4509 47296 4525 47360
rect 4589 47296 4597 47360
rect 4277 46272 4597 47296
rect 4277 46208 4285 46272
rect 4349 46208 4365 46272
rect 4429 46208 4445 46272
rect 4509 46208 4525 46272
rect 4589 46208 4597 46272
rect 4277 45184 4597 46208
rect 4277 45120 4285 45184
rect 4349 45120 4365 45184
rect 4429 45120 4445 45184
rect 4509 45120 4525 45184
rect 4589 45120 4597 45184
rect 4277 44096 4597 45120
rect 4277 44032 4285 44096
rect 4349 44032 4365 44096
rect 4429 44032 4445 44096
rect 4509 44032 4525 44096
rect 4589 44032 4597 44096
rect 4277 43008 4597 44032
rect 4277 42944 4285 43008
rect 4349 42944 4365 43008
rect 4429 42944 4445 43008
rect 4509 42944 4525 43008
rect 4589 42944 4597 43008
rect 4277 41920 4597 42944
rect 4277 41856 4285 41920
rect 4349 41856 4365 41920
rect 4429 41856 4445 41920
rect 4509 41856 4525 41920
rect 4589 41856 4597 41920
rect 4277 40832 4597 41856
rect 4277 40768 4285 40832
rect 4349 40768 4365 40832
rect 4429 40768 4445 40832
rect 4509 40768 4525 40832
rect 4589 40768 4597 40832
rect 4277 39744 4597 40768
rect 4277 39680 4285 39744
rect 4349 39680 4365 39744
rect 4429 39680 4445 39744
rect 4509 39680 4525 39744
rect 4589 39680 4597 39744
rect 4277 38656 4597 39680
rect 4277 38592 4285 38656
rect 4349 38592 4365 38656
rect 4429 38592 4445 38656
rect 4509 38592 4525 38656
rect 4589 38592 4597 38656
rect 4277 37568 4597 38592
rect 4277 37504 4285 37568
rect 4349 37504 4365 37568
rect 4429 37504 4445 37568
rect 4509 37504 4525 37568
rect 4589 37504 4597 37568
rect 4277 36480 4597 37504
rect 4277 36416 4285 36480
rect 4349 36416 4365 36480
rect 4429 36416 4445 36480
rect 4509 36416 4525 36480
rect 4589 36416 4597 36480
rect 4277 35392 4597 36416
rect 4277 35328 4285 35392
rect 4349 35328 4365 35392
rect 4429 35328 4445 35392
rect 4509 35328 4525 35392
rect 4589 35328 4597 35392
rect 4277 34304 4597 35328
rect 4277 34240 4285 34304
rect 4349 34240 4365 34304
rect 4429 34240 4445 34304
rect 4509 34240 4525 34304
rect 4589 34240 4597 34304
rect 4277 33216 4597 34240
rect 4277 33152 4285 33216
rect 4349 33152 4365 33216
rect 4429 33152 4445 33216
rect 4509 33152 4525 33216
rect 4589 33152 4597 33216
rect 4277 32128 4597 33152
rect 4277 32064 4285 32128
rect 4349 32064 4365 32128
rect 4429 32064 4445 32128
rect 4509 32064 4525 32128
rect 4589 32064 4597 32128
rect 4277 31040 4597 32064
rect 4277 30976 4285 31040
rect 4349 30976 4365 31040
rect 4429 30976 4445 31040
rect 4509 30976 4525 31040
rect 4589 30976 4597 31040
rect 4277 29952 4597 30976
rect 4277 29888 4285 29952
rect 4349 29888 4365 29952
rect 4429 29888 4445 29952
rect 4509 29888 4525 29952
rect 4589 29888 4597 29952
rect 4277 28864 4597 29888
rect 4277 28800 4285 28864
rect 4349 28800 4365 28864
rect 4429 28800 4445 28864
rect 4509 28800 4525 28864
rect 4589 28800 4597 28864
rect 4277 27776 4597 28800
rect 4277 27712 4285 27776
rect 4349 27712 4365 27776
rect 4429 27712 4445 27776
rect 4509 27712 4525 27776
rect 4589 27712 4597 27776
rect 4277 26688 4597 27712
rect 4277 26624 4285 26688
rect 4349 26624 4365 26688
rect 4429 26624 4445 26688
rect 4509 26624 4525 26688
rect 4589 26624 4597 26688
rect 4277 25600 4597 26624
rect 4277 25536 4285 25600
rect 4349 25536 4365 25600
rect 4429 25536 4445 25600
rect 4509 25536 4525 25600
rect 4589 25536 4597 25600
rect 4277 24512 4597 25536
rect 4277 24448 4285 24512
rect 4349 24448 4365 24512
rect 4429 24448 4445 24512
rect 4509 24448 4525 24512
rect 4589 24448 4597 24512
rect 4277 23424 4597 24448
rect 4277 23360 4285 23424
rect 4349 23360 4365 23424
rect 4429 23360 4445 23424
rect 4509 23360 4525 23424
rect 4589 23360 4597 23424
rect 4277 22336 4597 23360
rect 4277 22272 4285 22336
rect 4349 22272 4365 22336
rect 4429 22272 4445 22336
rect 4509 22272 4525 22336
rect 4589 22272 4597 22336
rect 4277 21248 4597 22272
rect 4277 21184 4285 21248
rect 4349 21184 4365 21248
rect 4429 21184 4445 21248
rect 4509 21184 4525 21248
rect 4589 21184 4597 21248
rect 4277 20160 4597 21184
rect 4277 20096 4285 20160
rect 4349 20096 4365 20160
rect 4429 20096 4445 20160
rect 4509 20096 4525 20160
rect 4589 20096 4597 20160
rect 4277 19072 4597 20096
rect 4277 19008 4285 19072
rect 4349 19008 4365 19072
rect 4429 19008 4445 19072
rect 4509 19008 4525 19072
rect 4589 19008 4597 19072
rect 4277 17984 4597 19008
rect 4277 17920 4285 17984
rect 4349 17920 4365 17984
rect 4429 17920 4445 17984
rect 4509 17920 4525 17984
rect 4589 17920 4597 17984
rect 4277 16896 4597 17920
rect 4277 16832 4285 16896
rect 4349 16832 4365 16896
rect 4429 16832 4445 16896
rect 4509 16832 4525 16896
rect 4589 16832 4597 16896
rect 4277 15808 4597 16832
rect 4277 15744 4285 15808
rect 4349 15744 4365 15808
rect 4429 15744 4445 15808
rect 4509 15744 4525 15808
rect 4589 15744 4597 15808
rect 4277 14720 4597 15744
rect 4277 14656 4285 14720
rect 4349 14656 4365 14720
rect 4429 14656 4445 14720
rect 4509 14656 4525 14720
rect 4589 14656 4597 14720
rect 4277 13632 4597 14656
rect 4277 13568 4285 13632
rect 4349 13568 4365 13632
rect 4429 13568 4445 13632
rect 4509 13568 4525 13632
rect 4589 13568 4597 13632
rect 4277 12544 4597 13568
rect 4277 12480 4285 12544
rect 4349 12480 4365 12544
rect 4429 12480 4445 12544
rect 4509 12480 4525 12544
rect 4589 12480 4597 12544
rect 4277 11456 4597 12480
rect 4277 11392 4285 11456
rect 4349 11392 4365 11456
rect 4429 11392 4445 11456
rect 4509 11392 4525 11456
rect 4589 11392 4597 11456
rect 4277 10368 4597 11392
rect 4277 10304 4285 10368
rect 4349 10304 4365 10368
rect 4429 10304 4445 10368
rect 4509 10304 4525 10368
rect 4589 10304 4597 10368
rect 4277 9280 4597 10304
rect 4277 9216 4285 9280
rect 4349 9216 4365 9280
rect 4429 9216 4445 9280
rect 4509 9216 4525 9280
rect 4589 9216 4597 9280
rect 4277 8192 4597 9216
rect 4277 8128 4285 8192
rect 4349 8128 4365 8192
rect 4429 8128 4445 8192
rect 4509 8128 4525 8192
rect 4589 8128 4597 8192
rect 4277 7104 4597 8128
rect 4277 7040 4285 7104
rect 4349 7040 4365 7104
rect 4429 7040 4445 7104
rect 4509 7040 4525 7104
rect 4589 7040 4597 7104
rect 4277 6016 4597 7040
rect 4277 5952 4285 6016
rect 4349 5952 4365 6016
rect 4429 5952 4445 6016
rect 4509 5952 4525 6016
rect 4589 5952 4597 6016
rect 4277 4928 4597 5952
rect 4277 4864 4285 4928
rect 4349 4864 4365 4928
rect 4429 4864 4445 4928
rect 4509 4864 4525 4928
rect 4589 4864 4597 4928
rect 4277 3840 4597 4864
rect 4277 3776 4285 3840
rect 4349 3776 4365 3840
rect 4429 3776 4445 3840
rect 4509 3776 4525 3840
rect 4589 3776 4597 3840
rect 4277 2752 4597 3776
rect 4277 2688 4285 2752
rect 4349 2688 4365 2752
rect 4429 2688 4445 2752
rect 4509 2688 4525 2752
rect 4589 2688 4597 2752
rect 4277 2128 4597 2688
rect 5944 330784 6264 330800
rect 5944 330720 5952 330784
rect 6016 330720 6032 330784
rect 6096 330720 6112 330784
rect 6176 330720 6192 330784
rect 6256 330720 6264 330784
rect 5944 329696 6264 330720
rect 5944 329632 5952 329696
rect 6016 329632 6032 329696
rect 6096 329632 6112 329696
rect 6176 329632 6192 329696
rect 6256 329632 6264 329696
rect 5944 328608 6264 329632
rect 5944 328544 5952 328608
rect 6016 328544 6032 328608
rect 6096 328544 6112 328608
rect 6176 328544 6192 328608
rect 6256 328544 6264 328608
rect 5944 327520 6264 328544
rect 5944 327456 5952 327520
rect 6016 327456 6032 327520
rect 6096 327456 6112 327520
rect 6176 327456 6192 327520
rect 6256 327456 6264 327520
rect 5944 326432 6264 327456
rect 5944 326368 5952 326432
rect 6016 326368 6032 326432
rect 6096 326368 6112 326432
rect 6176 326368 6192 326432
rect 6256 326368 6264 326432
rect 5944 325344 6264 326368
rect 5944 325280 5952 325344
rect 6016 325280 6032 325344
rect 6096 325280 6112 325344
rect 6176 325280 6192 325344
rect 6256 325280 6264 325344
rect 5944 324256 6264 325280
rect 5944 324192 5952 324256
rect 6016 324192 6032 324256
rect 6096 324192 6112 324256
rect 6176 324192 6192 324256
rect 6256 324192 6264 324256
rect 5944 323168 6264 324192
rect 5944 323104 5952 323168
rect 6016 323104 6032 323168
rect 6096 323104 6112 323168
rect 6176 323104 6192 323168
rect 6256 323104 6264 323168
rect 5944 322080 6264 323104
rect 5944 322016 5952 322080
rect 6016 322016 6032 322080
rect 6096 322016 6112 322080
rect 6176 322016 6192 322080
rect 6256 322016 6264 322080
rect 5944 320992 6264 322016
rect 5944 320928 5952 320992
rect 6016 320928 6032 320992
rect 6096 320928 6112 320992
rect 6176 320928 6192 320992
rect 6256 320928 6264 320992
rect 5944 319904 6264 320928
rect 5944 319840 5952 319904
rect 6016 319840 6032 319904
rect 6096 319840 6112 319904
rect 6176 319840 6192 319904
rect 6256 319840 6264 319904
rect 5944 318816 6264 319840
rect 5944 318752 5952 318816
rect 6016 318752 6032 318816
rect 6096 318752 6112 318816
rect 6176 318752 6192 318816
rect 6256 318752 6264 318816
rect 5944 317728 6264 318752
rect 5944 317664 5952 317728
rect 6016 317664 6032 317728
rect 6096 317664 6112 317728
rect 6176 317664 6192 317728
rect 6256 317664 6264 317728
rect 5944 316640 6264 317664
rect 5944 316576 5952 316640
rect 6016 316576 6032 316640
rect 6096 316576 6112 316640
rect 6176 316576 6192 316640
rect 6256 316576 6264 316640
rect 5944 315552 6264 316576
rect 5944 315488 5952 315552
rect 6016 315488 6032 315552
rect 6096 315488 6112 315552
rect 6176 315488 6192 315552
rect 6256 315488 6264 315552
rect 5944 314464 6264 315488
rect 5944 314400 5952 314464
rect 6016 314400 6032 314464
rect 6096 314400 6112 314464
rect 6176 314400 6192 314464
rect 6256 314400 6264 314464
rect 5944 313376 6264 314400
rect 5944 313312 5952 313376
rect 6016 313312 6032 313376
rect 6096 313312 6112 313376
rect 6176 313312 6192 313376
rect 6256 313312 6264 313376
rect 5944 312288 6264 313312
rect 5944 312224 5952 312288
rect 6016 312224 6032 312288
rect 6096 312224 6112 312288
rect 6176 312224 6192 312288
rect 6256 312224 6264 312288
rect 5944 311200 6264 312224
rect 5944 311136 5952 311200
rect 6016 311136 6032 311200
rect 6096 311136 6112 311200
rect 6176 311136 6192 311200
rect 6256 311136 6264 311200
rect 5944 310112 6264 311136
rect 5944 310048 5952 310112
rect 6016 310048 6032 310112
rect 6096 310048 6112 310112
rect 6176 310048 6192 310112
rect 6256 310048 6264 310112
rect 5944 309024 6264 310048
rect 5944 308960 5952 309024
rect 6016 308960 6032 309024
rect 6096 308960 6112 309024
rect 6176 308960 6192 309024
rect 6256 308960 6264 309024
rect 5944 307936 6264 308960
rect 5944 307872 5952 307936
rect 6016 307872 6032 307936
rect 6096 307872 6112 307936
rect 6176 307872 6192 307936
rect 6256 307872 6264 307936
rect 5944 306848 6264 307872
rect 5944 306784 5952 306848
rect 6016 306784 6032 306848
rect 6096 306784 6112 306848
rect 6176 306784 6192 306848
rect 6256 306784 6264 306848
rect 5944 305760 6264 306784
rect 5944 305696 5952 305760
rect 6016 305696 6032 305760
rect 6096 305696 6112 305760
rect 6176 305696 6192 305760
rect 6256 305696 6264 305760
rect 5944 304672 6264 305696
rect 5944 304608 5952 304672
rect 6016 304608 6032 304672
rect 6096 304608 6112 304672
rect 6176 304608 6192 304672
rect 6256 304608 6264 304672
rect 5944 303584 6264 304608
rect 5944 303520 5952 303584
rect 6016 303520 6032 303584
rect 6096 303520 6112 303584
rect 6176 303520 6192 303584
rect 6256 303520 6264 303584
rect 5944 302496 6264 303520
rect 5944 302432 5952 302496
rect 6016 302432 6032 302496
rect 6096 302432 6112 302496
rect 6176 302432 6192 302496
rect 6256 302432 6264 302496
rect 5944 301408 6264 302432
rect 5944 301344 5952 301408
rect 6016 301344 6032 301408
rect 6096 301344 6112 301408
rect 6176 301344 6192 301408
rect 6256 301344 6264 301408
rect 5944 300320 6264 301344
rect 5944 300256 5952 300320
rect 6016 300256 6032 300320
rect 6096 300256 6112 300320
rect 6176 300256 6192 300320
rect 6256 300256 6264 300320
rect 5944 299232 6264 300256
rect 5944 299168 5952 299232
rect 6016 299168 6032 299232
rect 6096 299168 6112 299232
rect 6176 299168 6192 299232
rect 6256 299168 6264 299232
rect 5944 298144 6264 299168
rect 5944 298080 5952 298144
rect 6016 298080 6032 298144
rect 6096 298080 6112 298144
rect 6176 298080 6192 298144
rect 6256 298080 6264 298144
rect 5944 297056 6264 298080
rect 5944 296992 5952 297056
rect 6016 296992 6032 297056
rect 6096 296992 6112 297056
rect 6176 296992 6192 297056
rect 6256 296992 6264 297056
rect 5944 295968 6264 296992
rect 5944 295904 5952 295968
rect 6016 295904 6032 295968
rect 6096 295904 6112 295968
rect 6176 295904 6192 295968
rect 6256 295904 6264 295968
rect 5944 294880 6264 295904
rect 5944 294816 5952 294880
rect 6016 294816 6032 294880
rect 6096 294816 6112 294880
rect 6176 294816 6192 294880
rect 6256 294816 6264 294880
rect 5944 293792 6264 294816
rect 5944 293728 5952 293792
rect 6016 293728 6032 293792
rect 6096 293728 6112 293792
rect 6176 293728 6192 293792
rect 6256 293728 6264 293792
rect 5944 292704 6264 293728
rect 5944 292640 5952 292704
rect 6016 292640 6032 292704
rect 6096 292640 6112 292704
rect 6176 292640 6192 292704
rect 6256 292640 6264 292704
rect 5944 291616 6264 292640
rect 5944 291552 5952 291616
rect 6016 291552 6032 291616
rect 6096 291552 6112 291616
rect 6176 291552 6192 291616
rect 6256 291552 6264 291616
rect 5944 290528 6264 291552
rect 5944 290464 5952 290528
rect 6016 290464 6032 290528
rect 6096 290464 6112 290528
rect 6176 290464 6192 290528
rect 6256 290464 6264 290528
rect 5944 289440 6264 290464
rect 5944 289376 5952 289440
rect 6016 289376 6032 289440
rect 6096 289376 6112 289440
rect 6176 289376 6192 289440
rect 6256 289376 6264 289440
rect 5944 288352 6264 289376
rect 5944 288288 5952 288352
rect 6016 288288 6032 288352
rect 6096 288288 6112 288352
rect 6176 288288 6192 288352
rect 6256 288288 6264 288352
rect 5944 287264 6264 288288
rect 5944 287200 5952 287264
rect 6016 287200 6032 287264
rect 6096 287200 6112 287264
rect 6176 287200 6192 287264
rect 6256 287200 6264 287264
rect 5944 286176 6264 287200
rect 5944 286112 5952 286176
rect 6016 286112 6032 286176
rect 6096 286112 6112 286176
rect 6176 286112 6192 286176
rect 6256 286112 6264 286176
rect 5944 285088 6264 286112
rect 5944 285024 5952 285088
rect 6016 285024 6032 285088
rect 6096 285024 6112 285088
rect 6176 285024 6192 285088
rect 6256 285024 6264 285088
rect 5944 284000 6264 285024
rect 5944 283936 5952 284000
rect 6016 283936 6032 284000
rect 6096 283936 6112 284000
rect 6176 283936 6192 284000
rect 6256 283936 6264 284000
rect 5944 282912 6264 283936
rect 5944 282848 5952 282912
rect 6016 282848 6032 282912
rect 6096 282848 6112 282912
rect 6176 282848 6192 282912
rect 6256 282848 6264 282912
rect 5944 281824 6264 282848
rect 5944 281760 5952 281824
rect 6016 281760 6032 281824
rect 6096 281760 6112 281824
rect 6176 281760 6192 281824
rect 6256 281760 6264 281824
rect 5944 280736 6264 281760
rect 5944 280672 5952 280736
rect 6016 280672 6032 280736
rect 6096 280672 6112 280736
rect 6176 280672 6192 280736
rect 6256 280672 6264 280736
rect 5944 279648 6264 280672
rect 5944 279584 5952 279648
rect 6016 279584 6032 279648
rect 6096 279584 6112 279648
rect 6176 279584 6192 279648
rect 6256 279584 6264 279648
rect 5944 278560 6264 279584
rect 5944 278496 5952 278560
rect 6016 278496 6032 278560
rect 6096 278496 6112 278560
rect 6176 278496 6192 278560
rect 6256 278496 6264 278560
rect 5944 277472 6264 278496
rect 5944 277408 5952 277472
rect 6016 277408 6032 277472
rect 6096 277408 6112 277472
rect 6176 277408 6192 277472
rect 6256 277408 6264 277472
rect 5944 276384 6264 277408
rect 5944 276320 5952 276384
rect 6016 276320 6032 276384
rect 6096 276320 6112 276384
rect 6176 276320 6192 276384
rect 6256 276320 6264 276384
rect 5944 275296 6264 276320
rect 5944 275232 5952 275296
rect 6016 275232 6032 275296
rect 6096 275232 6112 275296
rect 6176 275232 6192 275296
rect 6256 275232 6264 275296
rect 5944 274208 6264 275232
rect 5944 274144 5952 274208
rect 6016 274144 6032 274208
rect 6096 274144 6112 274208
rect 6176 274144 6192 274208
rect 6256 274144 6264 274208
rect 5944 273120 6264 274144
rect 5944 273056 5952 273120
rect 6016 273056 6032 273120
rect 6096 273056 6112 273120
rect 6176 273056 6192 273120
rect 6256 273056 6264 273120
rect 5944 272032 6264 273056
rect 5944 271968 5952 272032
rect 6016 271968 6032 272032
rect 6096 271968 6112 272032
rect 6176 271968 6192 272032
rect 6256 271968 6264 272032
rect 5944 270944 6264 271968
rect 5944 270880 5952 270944
rect 6016 270880 6032 270944
rect 6096 270880 6112 270944
rect 6176 270880 6192 270944
rect 6256 270880 6264 270944
rect 5944 269856 6264 270880
rect 5944 269792 5952 269856
rect 6016 269792 6032 269856
rect 6096 269792 6112 269856
rect 6176 269792 6192 269856
rect 6256 269792 6264 269856
rect 5944 268768 6264 269792
rect 5944 268704 5952 268768
rect 6016 268704 6032 268768
rect 6096 268704 6112 268768
rect 6176 268704 6192 268768
rect 6256 268704 6264 268768
rect 5944 267680 6264 268704
rect 5944 267616 5952 267680
rect 6016 267616 6032 267680
rect 6096 267616 6112 267680
rect 6176 267616 6192 267680
rect 6256 267616 6264 267680
rect 5944 266592 6264 267616
rect 5944 266528 5952 266592
rect 6016 266528 6032 266592
rect 6096 266528 6112 266592
rect 6176 266528 6192 266592
rect 6256 266528 6264 266592
rect 5944 265504 6264 266528
rect 5944 265440 5952 265504
rect 6016 265440 6032 265504
rect 6096 265440 6112 265504
rect 6176 265440 6192 265504
rect 6256 265440 6264 265504
rect 5944 264416 6264 265440
rect 5944 264352 5952 264416
rect 6016 264352 6032 264416
rect 6096 264352 6112 264416
rect 6176 264352 6192 264416
rect 6256 264352 6264 264416
rect 5944 263328 6264 264352
rect 5944 263264 5952 263328
rect 6016 263264 6032 263328
rect 6096 263264 6112 263328
rect 6176 263264 6192 263328
rect 6256 263264 6264 263328
rect 5944 262240 6264 263264
rect 5944 262176 5952 262240
rect 6016 262176 6032 262240
rect 6096 262176 6112 262240
rect 6176 262176 6192 262240
rect 6256 262176 6264 262240
rect 5944 261152 6264 262176
rect 5944 261088 5952 261152
rect 6016 261088 6032 261152
rect 6096 261088 6112 261152
rect 6176 261088 6192 261152
rect 6256 261088 6264 261152
rect 5944 260064 6264 261088
rect 5944 260000 5952 260064
rect 6016 260000 6032 260064
rect 6096 260000 6112 260064
rect 6176 260000 6192 260064
rect 6256 260000 6264 260064
rect 5944 258976 6264 260000
rect 5944 258912 5952 258976
rect 6016 258912 6032 258976
rect 6096 258912 6112 258976
rect 6176 258912 6192 258976
rect 6256 258912 6264 258976
rect 5944 257888 6264 258912
rect 5944 257824 5952 257888
rect 6016 257824 6032 257888
rect 6096 257824 6112 257888
rect 6176 257824 6192 257888
rect 6256 257824 6264 257888
rect 5944 256800 6264 257824
rect 5944 256736 5952 256800
rect 6016 256736 6032 256800
rect 6096 256736 6112 256800
rect 6176 256736 6192 256800
rect 6256 256736 6264 256800
rect 5944 255712 6264 256736
rect 5944 255648 5952 255712
rect 6016 255648 6032 255712
rect 6096 255648 6112 255712
rect 6176 255648 6192 255712
rect 6256 255648 6264 255712
rect 5944 254624 6264 255648
rect 5944 254560 5952 254624
rect 6016 254560 6032 254624
rect 6096 254560 6112 254624
rect 6176 254560 6192 254624
rect 6256 254560 6264 254624
rect 5944 253536 6264 254560
rect 5944 253472 5952 253536
rect 6016 253472 6032 253536
rect 6096 253472 6112 253536
rect 6176 253472 6192 253536
rect 6256 253472 6264 253536
rect 5944 252448 6264 253472
rect 5944 252384 5952 252448
rect 6016 252384 6032 252448
rect 6096 252384 6112 252448
rect 6176 252384 6192 252448
rect 6256 252384 6264 252448
rect 5944 251360 6264 252384
rect 5944 251296 5952 251360
rect 6016 251296 6032 251360
rect 6096 251296 6112 251360
rect 6176 251296 6192 251360
rect 6256 251296 6264 251360
rect 5944 250272 6264 251296
rect 5944 250208 5952 250272
rect 6016 250208 6032 250272
rect 6096 250208 6112 250272
rect 6176 250208 6192 250272
rect 6256 250208 6264 250272
rect 5944 249184 6264 250208
rect 5944 249120 5952 249184
rect 6016 249120 6032 249184
rect 6096 249120 6112 249184
rect 6176 249120 6192 249184
rect 6256 249120 6264 249184
rect 5944 248096 6264 249120
rect 5944 248032 5952 248096
rect 6016 248032 6032 248096
rect 6096 248032 6112 248096
rect 6176 248032 6192 248096
rect 6256 248032 6264 248096
rect 5944 247008 6264 248032
rect 5944 246944 5952 247008
rect 6016 246944 6032 247008
rect 6096 246944 6112 247008
rect 6176 246944 6192 247008
rect 6256 246944 6264 247008
rect 5944 245920 6264 246944
rect 5944 245856 5952 245920
rect 6016 245856 6032 245920
rect 6096 245856 6112 245920
rect 6176 245856 6192 245920
rect 6256 245856 6264 245920
rect 5944 244832 6264 245856
rect 5944 244768 5952 244832
rect 6016 244768 6032 244832
rect 6096 244768 6112 244832
rect 6176 244768 6192 244832
rect 6256 244768 6264 244832
rect 5944 243744 6264 244768
rect 5944 243680 5952 243744
rect 6016 243680 6032 243744
rect 6096 243680 6112 243744
rect 6176 243680 6192 243744
rect 6256 243680 6264 243744
rect 5944 242656 6264 243680
rect 5944 242592 5952 242656
rect 6016 242592 6032 242656
rect 6096 242592 6112 242656
rect 6176 242592 6192 242656
rect 6256 242592 6264 242656
rect 5944 241568 6264 242592
rect 5944 241504 5952 241568
rect 6016 241504 6032 241568
rect 6096 241504 6112 241568
rect 6176 241504 6192 241568
rect 6256 241504 6264 241568
rect 5944 240480 6264 241504
rect 5944 240416 5952 240480
rect 6016 240416 6032 240480
rect 6096 240416 6112 240480
rect 6176 240416 6192 240480
rect 6256 240416 6264 240480
rect 5944 239392 6264 240416
rect 5944 239328 5952 239392
rect 6016 239328 6032 239392
rect 6096 239328 6112 239392
rect 6176 239328 6192 239392
rect 6256 239328 6264 239392
rect 5944 238304 6264 239328
rect 5944 238240 5952 238304
rect 6016 238240 6032 238304
rect 6096 238240 6112 238304
rect 6176 238240 6192 238304
rect 6256 238240 6264 238304
rect 5944 237216 6264 238240
rect 5944 237152 5952 237216
rect 6016 237152 6032 237216
rect 6096 237152 6112 237216
rect 6176 237152 6192 237216
rect 6256 237152 6264 237216
rect 5944 236128 6264 237152
rect 5944 236064 5952 236128
rect 6016 236064 6032 236128
rect 6096 236064 6112 236128
rect 6176 236064 6192 236128
rect 6256 236064 6264 236128
rect 5944 235040 6264 236064
rect 5944 234976 5952 235040
rect 6016 234976 6032 235040
rect 6096 234976 6112 235040
rect 6176 234976 6192 235040
rect 6256 234976 6264 235040
rect 5944 233952 6264 234976
rect 5944 233888 5952 233952
rect 6016 233888 6032 233952
rect 6096 233888 6112 233952
rect 6176 233888 6192 233952
rect 6256 233888 6264 233952
rect 5944 232864 6264 233888
rect 5944 232800 5952 232864
rect 6016 232800 6032 232864
rect 6096 232800 6112 232864
rect 6176 232800 6192 232864
rect 6256 232800 6264 232864
rect 5944 231776 6264 232800
rect 5944 231712 5952 231776
rect 6016 231712 6032 231776
rect 6096 231712 6112 231776
rect 6176 231712 6192 231776
rect 6256 231712 6264 231776
rect 5944 230688 6264 231712
rect 5944 230624 5952 230688
rect 6016 230624 6032 230688
rect 6096 230624 6112 230688
rect 6176 230624 6192 230688
rect 6256 230624 6264 230688
rect 5944 229600 6264 230624
rect 5944 229536 5952 229600
rect 6016 229536 6032 229600
rect 6096 229536 6112 229600
rect 6176 229536 6192 229600
rect 6256 229536 6264 229600
rect 5944 228512 6264 229536
rect 5944 228448 5952 228512
rect 6016 228448 6032 228512
rect 6096 228448 6112 228512
rect 6176 228448 6192 228512
rect 6256 228448 6264 228512
rect 5944 227424 6264 228448
rect 5944 227360 5952 227424
rect 6016 227360 6032 227424
rect 6096 227360 6112 227424
rect 6176 227360 6192 227424
rect 6256 227360 6264 227424
rect 5944 226336 6264 227360
rect 5944 226272 5952 226336
rect 6016 226272 6032 226336
rect 6096 226272 6112 226336
rect 6176 226272 6192 226336
rect 6256 226272 6264 226336
rect 5944 225248 6264 226272
rect 5944 225184 5952 225248
rect 6016 225184 6032 225248
rect 6096 225184 6112 225248
rect 6176 225184 6192 225248
rect 6256 225184 6264 225248
rect 5944 224160 6264 225184
rect 5944 224096 5952 224160
rect 6016 224096 6032 224160
rect 6096 224096 6112 224160
rect 6176 224096 6192 224160
rect 6256 224096 6264 224160
rect 5944 223072 6264 224096
rect 5944 223008 5952 223072
rect 6016 223008 6032 223072
rect 6096 223008 6112 223072
rect 6176 223008 6192 223072
rect 6256 223008 6264 223072
rect 5944 221984 6264 223008
rect 5944 221920 5952 221984
rect 6016 221920 6032 221984
rect 6096 221920 6112 221984
rect 6176 221920 6192 221984
rect 6256 221920 6264 221984
rect 5944 220896 6264 221920
rect 5944 220832 5952 220896
rect 6016 220832 6032 220896
rect 6096 220832 6112 220896
rect 6176 220832 6192 220896
rect 6256 220832 6264 220896
rect 5944 219808 6264 220832
rect 5944 219744 5952 219808
rect 6016 219744 6032 219808
rect 6096 219744 6112 219808
rect 6176 219744 6192 219808
rect 6256 219744 6264 219808
rect 5944 218720 6264 219744
rect 5944 218656 5952 218720
rect 6016 218656 6032 218720
rect 6096 218656 6112 218720
rect 6176 218656 6192 218720
rect 6256 218656 6264 218720
rect 5944 217632 6264 218656
rect 5944 217568 5952 217632
rect 6016 217568 6032 217632
rect 6096 217568 6112 217632
rect 6176 217568 6192 217632
rect 6256 217568 6264 217632
rect 5944 216544 6264 217568
rect 5944 216480 5952 216544
rect 6016 216480 6032 216544
rect 6096 216480 6112 216544
rect 6176 216480 6192 216544
rect 6256 216480 6264 216544
rect 5944 215456 6264 216480
rect 5944 215392 5952 215456
rect 6016 215392 6032 215456
rect 6096 215392 6112 215456
rect 6176 215392 6192 215456
rect 6256 215392 6264 215456
rect 5944 214368 6264 215392
rect 5944 214304 5952 214368
rect 6016 214304 6032 214368
rect 6096 214304 6112 214368
rect 6176 214304 6192 214368
rect 6256 214304 6264 214368
rect 5944 213280 6264 214304
rect 5944 213216 5952 213280
rect 6016 213216 6032 213280
rect 6096 213216 6112 213280
rect 6176 213216 6192 213280
rect 6256 213216 6264 213280
rect 5944 212192 6264 213216
rect 5944 212128 5952 212192
rect 6016 212128 6032 212192
rect 6096 212128 6112 212192
rect 6176 212128 6192 212192
rect 6256 212128 6264 212192
rect 5944 211104 6264 212128
rect 5944 211040 5952 211104
rect 6016 211040 6032 211104
rect 6096 211040 6112 211104
rect 6176 211040 6192 211104
rect 6256 211040 6264 211104
rect 5944 210016 6264 211040
rect 5944 209952 5952 210016
rect 6016 209952 6032 210016
rect 6096 209952 6112 210016
rect 6176 209952 6192 210016
rect 6256 209952 6264 210016
rect 5944 208928 6264 209952
rect 5944 208864 5952 208928
rect 6016 208864 6032 208928
rect 6096 208864 6112 208928
rect 6176 208864 6192 208928
rect 6256 208864 6264 208928
rect 5944 207840 6264 208864
rect 5944 207776 5952 207840
rect 6016 207776 6032 207840
rect 6096 207776 6112 207840
rect 6176 207776 6192 207840
rect 6256 207776 6264 207840
rect 5944 206752 6264 207776
rect 5944 206688 5952 206752
rect 6016 206688 6032 206752
rect 6096 206688 6112 206752
rect 6176 206688 6192 206752
rect 6256 206688 6264 206752
rect 5944 205664 6264 206688
rect 5944 205600 5952 205664
rect 6016 205600 6032 205664
rect 6096 205600 6112 205664
rect 6176 205600 6192 205664
rect 6256 205600 6264 205664
rect 5944 204576 6264 205600
rect 5944 204512 5952 204576
rect 6016 204512 6032 204576
rect 6096 204512 6112 204576
rect 6176 204512 6192 204576
rect 6256 204512 6264 204576
rect 5944 203488 6264 204512
rect 5944 203424 5952 203488
rect 6016 203424 6032 203488
rect 6096 203424 6112 203488
rect 6176 203424 6192 203488
rect 6256 203424 6264 203488
rect 5944 202400 6264 203424
rect 5944 202336 5952 202400
rect 6016 202336 6032 202400
rect 6096 202336 6112 202400
rect 6176 202336 6192 202400
rect 6256 202336 6264 202400
rect 5944 201312 6264 202336
rect 5944 201248 5952 201312
rect 6016 201248 6032 201312
rect 6096 201248 6112 201312
rect 6176 201248 6192 201312
rect 6256 201248 6264 201312
rect 5944 200224 6264 201248
rect 5944 200160 5952 200224
rect 6016 200160 6032 200224
rect 6096 200160 6112 200224
rect 6176 200160 6192 200224
rect 6256 200160 6264 200224
rect 5944 199136 6264 200160
rect 5944 199072 5952 199136
rect 6016 199072 6032 199136
rect 6096 199072 6112 199136
rect 6176 199072 6192 199136
rect 6256 199072 6264 199136
rect 5944 198048 6264 199072
rect 5944 197984 5952 198048
rect 6016 197984 6032 198048
rect 6096 197984 6112 198048
rect 6176 197984 6192 198048
rect 6256 197984 6264 198048
rect 5944 196960 6264 197984
rect 5944 196896 5952 196960
rect 6016 196896 6032 196960
rect 6096 196896 6112 196960
rect 6176 196896 6192 196960
rect 6256 196896 6264 196960
rect 5944 195872 6264 196896
rect 5944 195808 5952 195872
rect 6016 195808 6032 195872
rect 6096 195808 6112 195872
rect 6176 195808 6192 195872
rect 6256 195808 6264 195872
rect 5944 194784 6264 195808
rect 5944 194720 5952 194784
rect 6016 194720 6032 194784
rect 6096 194720 6112 194784
rect 6176 194720 6192 194784
rect 6256 194720 6264 194784
rect 5944 193696 6264 194720
rect 5944 193632 5952 193696
rect 6016 193632 6032 193696
rect 6096 193632 6112 193696
rect 6176 193632 6192 193696
rect 6256 193632 6264 193696
rect 5944 192608 6264 193632
rect 5944 192544 5952 192608
rect 6016 192544 6032 192608
rect 6096 192544 6112 192608
rect 6176 192544 6192 192608
rect 6256 192544 6264 192608
rect 5944 191520 6264 192544
rect 5944 191456 5952 191520
rect 6016 191456 6032 191520
rect 6096 191456 6112 191520
rect 6176 191456 6192 191520
rect 6256 191456 6264 191520
rect 5944 190432 6264 191456
rect 5944 190368 5952 190432
rect 6016 190368 6032 190432
rect 6096 190368 6112 190432
rect 6176 190368 6192 190432
rect 6256 190368 6264 190432
rect 5944 189344 6264 190368
rect 5944 189280 5952 189344
rect 6016 189280 6032 189344
rect 6096 189280 6112 189344
rect 6176 189280 6192 189344
rect 6256 189280 6264 189344
rect 5944 188256 6264 189280
rect 5944 188192 5952 188256
rect 6016 188192 6032 188256
rect 6096 188192 6112 188256
rect 6176 188192 6192 188256
rect 6256 188192 6264 188256
rect 5944 187168 6264 188192
rect 5944 187104 5952 187168
rect 6016 187104 6032 187168
rect 6096 187104 6112 187168
rect 6176 187104 6192 187168
rect 6256 187104 6264 187168
rect 5944 186080 6264 187104
rect 5944 186016 5952 186080
rect 6016 186016 6032 186080
rect 6096 186016 6112 186080
rect 6176 186016 6192 186080
rect 6256 186016 6264 186080
rect 5944 184992 6264 186016
rect 5944 184928 5952 184992
rect 6016 184928 6032 184992
rect 6096 184928 6112 184992
rect 6176 184928 6192 184992
rect 6256 184928 6264 184992
rect 5944 183904 6264 184928
rect 5944 183840 5952 183904
rect 6016 183840 6032 183904
rect 6096 183840 6112 183904
rect 6176 183840 6192 183904
rect 6256 183840 6264 183904
rect 5944 182816 6264 183840
rect 5944 182752 5952 182816
rect 6016 182752 6032 182816
rect 6096 182752 6112 182816
rect 6176 182752 6192 182816
rect 6256 182752 6264 182816
rect 5944 181728 6264 182752
rect 5944 181664 5952 181728
rect 6016 181664 6032 181728
rect 6096 181664 6112 181728
rect 6176 181664 6192 181728
rect 6256 181664 6264 181728
rect 5944 180640 6264 181664
rect 5944 180576 5952 180640
rect 6016 180576 6032 180640
rect 6096 180576 6112 180640
rect 6176 180576 6192 180640
rect 6256 180576 6264 180640
rect 5944 179552 6264 180576
rect 5944 179488 5952 179552
rect 6016 179488 6032 179552
rect 6096 179488 6112 179552
rect 6176 179488 6192 179552
rect 6256 179488 6264 179552
rect 5944 178464 6264 179488
rect 5944 178400 5952 178464
rect 6016 178400 6032 178464
rect 6096 178400 6112 178464
rect 6176 178400 6192 178464
rect 6256 178400 6264 178464
rect 5944 177376 6264 178400
rect 5944 177312 5952 177376
rect 6016 177312 6032 177376
rect 6096 177312 6112 177376
rect 6176 177312 6192 177376
rect 6256 177312 6264 177376
rect 5944 176288 6264 177312
rect 5944 176224 5952 176288
rect 6016 176224 6032 176288
rect 6096 176224 6112 176288
rect 6176 176224 6192 176288
rect 6256 176224 6264 176288
rect 5944 175200 6264 176224
rect 5944 175136 5952 175200
rect 6016 175136 6032 175200
rect 6096 175136 6112 175200
rect 6176 175136 6192 175200
rect 6256 175136 6264 175200
rect 5944 174112 6264 175136
rect 5944 174048 5952 174112
rect 6016 174048 6032 174112
rect 6096 174048 6112 174112
rect 6176 174048 6192 174112
rect 6256 174048 6264 174112
rect 5944 173024 6264 174048
rect 5944 172960 5952 173024
rect 6016 172960 6032 173024
rect 6096 172960 6112 173024
rect 6176 172960 6192 173024
rect 6256 172960 6264 173024
rect 5944 171936 6264 172960
rect 5944 171872 5952 171936
rect 6016 171872 6032 171936
rect 6096 171872 6112 171936
rect 6176 171872 6192 171936
rect 6256 171872 6264 171936
rect 5944 170848 6264 171872
rect 5944 170784 5952 170848
rect 6016 170784 6032 170848
rect 6096 170784 6112 170848
rect 6176 170784 6192 170848
rect 6256 170784 6264 170848
rect 5944 169760 6264 170784
rect 5944 169696 5952 169760
rect 6016 169696 6032 169760
rect 6096 169696 6112 169760
rect 6176 169696 6192 169760
rect 6256 169696 6264 169760
rect 5944 168672 6264 169696
rect 5944 168608 5952 168672
rect 6016 168608 6032 168672
rect 6096 168608 6112 168672
rect 6176 168608 6192 168672
rect 6256 168608 6264 168672
rect 5944 167584 6264 168608
rect 5944 167520 5952 167584
rect 6016 167520 6032 167584
rect 6096 167520 6112 167584
rect 6176 167520 6192 167584
rect 6256 167520 6264 167584
rect 5944 166496 6264 167520
rect 5944 166432 5952 166496
rect 6016 166432 6032 166496
rect 6096 166432 6112 166496
rect 6176 166432 6192 166496
rect 6256 166432 6264 166496
rect 5944 165408 6264 166432
rect 5944 165344 5952 165408
rect 6016 165344 6032 165408
rect 6096 165344 6112 165408
rect 6176 165344 6192 165408
rect 6256 165344 6264 165408
rect 5944 164320 6264 165344
rect 5944 164256 5952 164320
rect 6016 164256 6032 164320
rect 6096 164256 6112 164320
rect 6176 164256 6192 164320
rect 6256 164256 6264 164320
rect 5944 163232 6264 164256
rect 5944 163168 5952 163232
rect 6016 163168 6032 163232
rect 6096 163168 6112 163232
rect 6176 163168 6192 163232
rect 6256 163168 6264 163232
rect 5944 162144 6264 163168
rect 5944 162080 5952 162144
rect 6016 162080 6032 162144
rect 6096 162080 6112 162144
rect 6176 162080 6192 162144
rect 6256 162080 6264 162144
rect 5944 161056 6264 162080
rect 5944 160992 5952 161056
rect 6016 160992 6032 161056
rect 6096 160992 6112 161056
rect 6176 160992 6192 161056
rect 6256 160992 6264 161056
rect 5944 159968 6264 160992
rect 5944 159904 5952 159968
rect 6016 159904 6032 159968
rect 6096 159904 6112 159968
rect 6176 159904 6192 159968
rect 6256 159904 6264 159968
rect 5944 158880 6264 159904
rect 5944 158816 5952 158880
rect 6016 158816 6032 158880
rect 6096 158816 6112 158880
rect 6176 158816 6192 158880
rect 6256 158816 6264 158880
rect 5944 157792 6264 158816
rect 5944 157728 5952 157792
rect 6016 157728 6032 157792
rect 6096 157728 6112 157792
rect 6176 157728 6192 157792
rect 6256 157728 6264 157792
rect 5944 156704 6264 157728
rect 5944 156640 5952 156704
rect 6016 156640 6032 156704
rect 6096 156640 6112 156704
rect 6176 156640 6192 156704
rect 6256 156640 6264 156704
rect 5944 155616 6264 156640
rect 5944 155552 5952 155616
rect 6016 155552 6032 155616
rect 6096 155552 6112 155616
rect 6176 155552 6192 155616
rect 6256 155552 6264 155616
rect 5944 154528 6264 155552
rect 5944 154464 5952 154528
rect 6016 154464 6032 154528
rect 6096 154464 6112 154528
rect 6176 154464 6192 154528
rect 6256 154464 6264 154528
rect 5944 153440 6264 154464
rect 5944 153376 5952 153440
rect 6016 153376 6032 153440
rect 6096 153376 6112 153440
rect 6176 153376 6192 153440
rect 6256 153376 6264 153440
rect 5944 152352 6264 153376
rect 5944 152288 5952 152352
rect 6016 152288 6032 152352
rect 6096 152288 6112 152352
rect 6176 152288 6192 152352
rect 6256 152288 6264 152352
rect 5944 151264 6264 152288
rect 5944 151200 5952 151264
rect 6016 151200 6032 151264
rect 6096 151200 6112 151264
rect 6176 151200 6192 151264
rect 6256 151200 6264 151264
rect 5944 150176 6264 151200
rect 5944 150112 5952 150176
rect 6016 150112 6032 150176
rect 6096 150112 6112 150176
rect 6176 150112 6192 150176
rect 6256 150112 6264 150176
rect 5944 149088 6264 150112
rect 5944 149024 5952 149088
rect 6016 149024 6032 149088
rect 6096 149024 6112 149088
rect 6176 149024 6192 149088
rect 6256 149024 6264 149088
rect 5944 148000 6264 149024
rect 5944 147936 5952 148000
rect 6016 147936 6032 148000
rect 6096 147936 6112 148000
rect 6176 147936 6192 148000
rect 6256 147936 6264 148000
rect 5944 146912 6264 147936
rect 5944 146848 5952 146912
rect 6016 146848 6032 146912
rect 6096 146848 6112 146912
rect 6176 146848 6192 146912
rect 6256 146848 6264 146912
rect 5944 145824 6264 146848
rect 5944 145760 5952 145824
rect 6016 145760 6032 145824
rect 6096 145760 6112 145824
rect 6176 145760 6192 145824
rect 6256 145760 6264 145824
rect 5944 144736 6264 145760
rect 5944 144672 5952 144736
rect 6016 144672 6032 144736
rect 6096 144672 6112 144736
rect 6176 144672 6192 144736
rect 6256 144672 6264 144736
rect 5944 143648 6264 144672
rect 5944 143584 5952 143648
rect 6016 143584 6032 143648
rect 6096 143584 6112 143648
rect 6176 143584 6192 143648
rect 6256 143584 6264 143648
rect 5944 142560 6264 143584
rect 5944 142496 5952 142560
rect 6016 142496 6032 142560
rect 6096 142496 6112 142560
rect 6176 142496 6192 142560
rect 6256 142496 6264 142560
rect 5944 141472 6264 142496
rect 5944 141408 5952 141472
rect 6016 141408 6032 141472
rect 6096 141408 6112 141472
rect 6176 141408 6192 141472
rect 6256 141408 6264 141472
rect 5944 140384 6264 141408
rect 5944 140320 5952 140384
rect 6016 140320 6032 140384
rect 6096 140320 6112 140384
rect 6176 140320 6192 140384
rect 6256 140320 6264 140384
rect 5944 139296 6264 140320
rect 5944 139232 5952 139296
rect 6016 139232 6032 139296
rect 6096 139232 6112 139296
rect 6176 139232 6192 139296
rect 6256 139232 6264 139296
rect 5944 138208 6264 139232
rect 5944 138144 5952 138208
rect 6016 138144 6032 138208
rect 6096 138144 6112 138208
rect 6176 138144 6192 138208
rect 6256 138144 6264 138208
rect 5944 137120 6264 138144
rect 5944 137056 5952 137120
rect 6016 137056 6032 137120
rect 6096 137056 6112 137120
rect 6176 137056 6192 137120
rect 6256 137056 6264 137120
rect 5944 136032 6264 137056
rect 5944 135968 5952 136032
rect 6016 135968 6032 136032
rect 6096 135968 6112 136032
rect 6176 135968 6192 136032
rect 6256 135968 6264 136032
rect 5944 134944 6264 135968
rect 5944 134880 5952 134944
rect 6016 134880 6032 134944
rect 6096 134880 6112 134944
rect 6176 134880 6192 134944
rect 6256 134880 6264 134944
rect 5944 133856 6264 134880
rect 5944 133792 5952 133856
rect 6016 133792 6032 133856
rect 6096 133792 6112 133856
rect 6176 133792 6192 133856
rect 6256 133792 6264 133856
rect 5944 132768 6264 133792
rect 5944 132704 5952 132768
rect 6016 132704 6032 132768
rect 6096 132704 6112 132768
rect 6176 132704 6192 132768
rect 6256 132704 6264 132768
rect 5944 131680 6264 132704
rect 5944 131616 5952 131680
rect 6016 131616 6032 131680
rect 6096 131616 6112 131680
rect 6176 131616 6192 131680
rect 6256 131616 6264 131680
rect 5944 130592 6264 131616
rect 5944 130528 5952 130592
rect 6016 130528 6032 130592
rect 6096 130528 6112 130592
rect 6176 130528 6192 130592
rect 6256 130528 6264 130592
rect 5944 129504 6264 130528
rect 5944 129440 5952 129504
rect 6016 129440 6032 129504
rect 6096 129440 6112 129504
rect 6176 129440 6192 129504
rect 6256 129440 6264 129504
rect 5944 128416 6264 129440
rect 5944 128352 5952 128416
rect 6016 128352 6032 128416
rect 6096 128352 6112 128416
rect 6176 128352 6192 128416
rect 6256 128352 6264 128416
rect 5944 127328 6264 128352
rect 5944 127264 5952 127328
rect 6016 127264 6032 127328
rect 6096 127264 6112 127328
rect 6176 127264 6192 127328
rect 6256 127264 6264 127328
rect 5944 126240 6264 127264
rect 5944 126176 5952 126240
rect 6016 126176 6032 126240
rect 6096 126176 6112 126240
rect 6176 126176 6192 126240
rect 6256 126176 6264 126240
rect 5944 125152 6264 126176
rect 5944 125088 5952 125152
rect 6016 125088 6032 125152
rect 6096 125088 6112 125152
rect 6176 125088 6192 125152
rect 6256 125088 6264 125152
rect 5944 124064 6264 125088
rect 5944 124000 5952 124064
rect 6016 124000 6032 124064
rect 6096 124000 6112 124064
rect 6176 124000 6192 124064
rect 6256 124000 6264 124064
rect 5944 122976 6264 124000
rect 5944 122912 5952 122976
rect 6016 122912 6032 122976
rect 6096 122912 6112 122976
rect 6176 122912 6192 122976
rect 6256 122912 6264 122976
rect 5944 121888 6264 122912
rect 5944 121824 5952 121888
rect 6016 121824 6032 121888
rect 6096 121824 6112 121888
rect 6176 121824 6192 121888
rect 6256 121824 6264 121888
rect 5944 120800 6264 121824
rect 5944 120736 5952 120800
rect 6016 120736 6032 120800
rect 6096 120736 6112 120800
rect 6176 120736 6192 120800
rect 6256 120736 6264 120800
rect 5944 119712 6264 120736
rect 5944 119648 5952 119712
rect 6016 119648 6032 119712
rect 6096 119648 6112 119712
rect 6176 119648 6192 119712
rect 6256 119648 6264 119712
rect 5944 118624 6264 119648
rect 5944 118560 5952 118624
rect 6016 118560 6032 118624
rect 6096 118560 6112 118624
rect 6176 118560 6192 118624
rect 6256 118560 6264 118624
rect 5944 117536 6264 118560
rect 5944 117472 5952 117536
rect 6016 117472 6032 117536
rect 6096 117472 6112 117536
rect 6176 117472 6192 117536
rect 6256 117472 6264 117536
rect 5944 116448 6264 117472
rect 5944 116384 5952 116448
rect 6016 116384 6032 116448
rect 6096 116384 6112 116448
rect 6176 116384 6192 116448
rect 6256 116384 6264 116448
rect 5944 115360 6264 116384
rect 5944 115296 5952 115360
rect 6016 115296 6032 115360
rect 6096 115296 6112 115360
rect 6176 115296 6192 115360
rect 6256 115296 6264 115360
rect 5944 114272 6264 115296
rect 5944 114208 5952 114272
rect 6016 114208 6032 114272
rect 6096 114208 6112 114272
rect 6176 114208 6192 114272
rect 6256 114208 6264 114272
rect 5944 113184 6264 114208
rect 5944 113120 5952 113184
rect 6016 113120 6032 113184
rect 6096 113120 6112 113184
rect 6176 113120 6192 113184
rect 6256 113120 6264 113184
rect 5944 112096 6264 113120
rect 5944 112032 5952 112096
rect 6016 112032 6032 112096
rect 6096 112032 6112 112096
rect 6176 112032 6192 112096
rect 6256 112032 6264 112096
rect 5944 111008 6264 112032
rect 5944 110944 5952 111008
rect 6016 110944 6032 111008
rect 6096 110944 6112 111008
rect 6176 110944 6192 111008
rect 6256 110944 6264 111008
rect 5944 109920 6264 110944
rect 5944 109856 5952 109920
rect 6016 109856 6032 109920
rect 6096 109856 6112 109920
rect 6176 109856 6192 109920
rect 6256 109856 6264 109920
rect 5944 108832 6264 109856
rect 5944 108768 5952 108832
rect 6016 108768 6032 108832
rect 6096 108768 6112 108832
rect 6176 108768 6192 108832
rect 6256 108768 6264 108832
rect 5944 107744 6264 108768
rect 5944 107680 5952 107744
rect 6016 107680 6032 107744
rect 6096 107680 6112 107744
rect 6176 107680 6192 107744
rect 6256 107680 6264 107744
rect 5944 106656 6264 107680
rect 5944 106592 5952 106656
rect 6016 106592 6032 106656
rect 6096 106592 6112 106656
rect 6176 106592 6192 106656
rect 6256 106592 6264 106656
rect 5944 105568 6264 106592
rect 5944 105504 5952 105568
rect 6016 105504 6032 105568
rect 6096 105504 6112 105568
rect 6176 105504 6192 105568
rect 6256 105504 6264 105568
rect 5944 104480 6264 105504
rect 5944 104416 5952 104480
rect 6016 104416 6032 104480
rect 6096 104416 6112 104480
rect 6176 104416 6192 104480
rect 6256 104416 6264 104480
rect 5944 103392 6264 104416
rect 5944 103328 5952 103392
rect 6016 103328 6032 103392
rect 6096 103328 6112 103392
rect 6176 103328 6192 103392
rect 6256 103328 6264 103392
rect 5944 102304 6264 103328
rect 5944 102240 5952 102304
rect 6016 102240 6032 102304
rect 6096 102240 6112 102304
rect 6176 102240 6192 102304
rect 6256 102240 6264 102304
rect 5944 101216 6264 102240
rect 5944 101152 5952 101216
rect 6016 101152 6032 101216
rect 6096 101152 6112 101216
rect 6176 101152 6192 101216
rect 6256 101152 6264 101216
rect 5944 100128 6264 101152
rect 5944 100064 5952 100128
rect 6016 100064 6032 100128
rect 6096 100064 6112 100128
rect 6176 100064 6192 100128
rect 6256 100064 6264 100128
rect 5944 99040 6264 100064
rect 5944 98976 5952 99040
rect 6016 98976 6032 99040
rect 6096 98976 6112 99040
rect 6176 98976 6192 99040
rect 6256 98976 6264 99040
rect 5944 97952 6264 98976
rect 5944 97888 5952 97952
rect 6016 97888 6032 97952
rect 6096 97888 6112 97952
rect 6176 97888 6192 97952
rect 6256 97888 6264 97952
rect 5944 96864 6264 97888
rect 5944 96800 5952 96864
rect 6016 96800 6032 96864
rect 6096 96800 6112 96864
rect 6176 96800 6192 96864
rect 6256 96800 6264 96864
rect 5944 95776 6264 96800
rect 5944 95712 5952 95776
rect 6016 95712 6032 95776
rect 6096 95712 6112 95776
rect 6176 95712 6192 95776
rect 6256 95712 6264 95776
rect 5944 94688 6264 95712
rect 5944 94624 5952 94688
rect 6016 94624 6032 94688
rect 6096 94624 6112 94688
rect 6176 94624 6192 94688
rect 6256 94624 6264 94688
rect 5944 93600 6264 94624
rect 5944 93536 5952 93600
rect 6016 93536 6032 93600
rect 6096 93536 6112 93600
rect 6176 93536 6192 93600
rect 6256 93536 6264 93600
rect 5944 92512 6264 93536
rect 5944 92448 5952 92512
rect 6016 92448 6032 92512
rect 6096 92448 6112 92512
rect 6176 92448 6192 92512
rect 6256 92448 6264 92512
rect 5944 91424 6264 92448
rect 5944 91360 5952 91424
rect 6016 91360 6032 91424
rect 6096 91360 6112 91424
rect 6176 91360 6192 91424
rect 6256 91360 6264 91424
rect 5944 90336 6264 91360
rect 5944 90272 5952 90336
rect 6016 90272 6032 90336
rect 6096 90272 6112 90336
rect 6176 90272 6192 90336
rect 6256 90272 6264 90336
rect 5944 89248 6264 90272
rect 5944 89184 5952 89248
rect 6016 89184 6032 89248
rect 6096 89184 6112 89248
rect 6176 89184 6192 89248
rect 6256 89184 6264 89248
rect 5944 88160 6264 89184
rect 5944 88096 5952 88160
rect 6016 88096 6032 88160
rect 6096 88096 6112 88160
rect 6176 88096 6192 88160
rect 6256 88096 6264 88160
rect 5944 87072 6264 88096
rect 5944 87008 5952 87072
rect 6016 87008 6032 87072
rect 6096 87008 6112 87072
rect 6176 87008 6192 87072
rect 6256 87008 6264 87072
rect 5944 85984 6264 87008
rect 5944 85920 5952 85984
rect 6016 85920 6032 85984
rect 6096 85920 6112 85984
rect 6176 85920 6192 85984
rect 6256 85920 6264 85984
rect 5944 84896 6264 85920
rect 5944 84832 5952 84896
rect 6016 84832 6032 84896
rect 6096 84832 6112 84896
rect 6176 84832 6192 84896
rect 6256 84832 6264 84896
rect 5944 83808 6264 84832
rect 5944 83744 5952 83808
rect 6016 83744 6032 83808
rect 6096 83744 6112 83808
rect 6176 83744 6192 83808
rect 6256 83744 6264 83808
rect 5944 82720 6264 83744
rect 5944 82656 5952 82720
rect 6016 82656 6032 82720
rect 6096 82656 6112 82720
rect 6176 82656 6192 82720
rect 6256 82656 6264 82720
rect 5944 81632 6264 82656
rect 5944 81568 5952 81632
rect 6016 81568 6032 81632
rect 6096 81568 6112 81632
rect 6176 81568 6192 81632
rect 6256 81568 6264 81632
rect 5944 80544 6264 81568
rect 5944 80480 5952 80544
rect 6016 80480 6032 80544
rect 6096 80480 6112 80544
rect 6176 80480 6192 80544
rect 6256 80480 6264 80544
rect 5944 79456 6264 80480
rect 5944 79392 5952 79456
rect 6016 79392 6032 79456
rect 6096 79392 6112 79456
rect 6176 79392 6192 79456
rect 6256 79392 6264 79456
rect 5944 78368 6264 79392
rect 5944 78304 5952 78368
rect 6016 78304 6032 78368
rect 6096 78304 6112 78368
rect 6176 78304 6192 78368
rect 6256 78304 6264 78368
rect 5944 77280 6264 78304
rect 5944 77216 5952 77280
rect 6016 77216 6032 77280
rect 6096 77216 6112 77280
rect 6176 77216 6192 77280
rect 6256 77216 6264 77280
rect 5944 76192 6264 77216
rect 5944 76128 5952 76192
rect 6016 76128 6032 76192
rect 6096 76128 6112 76192
rect 6176 76128 6192 76192
rect 6256 76128 6264 76192
rect 5944 75104 6264 76128
rect 5944 75040 5952 75104
rect 6016 75040 6032 75104
rect 6096 75040 6112 75104
rect 6176 75040 6192 75104
rect 6256 75040 6264 75104
rect 5944 74016 6264 75040
rect 5944 73952 5952 74016
rect 6016 73952 6032 74016
rect 6096 73952 6112 74016
rect 6176 73952 6192 74016
rect 6256 73952 6264 74016
rect 5944 72928 6264 73952
rect 5944 72864 5952 72928
rect 6016 72864 6032 72928
rect 6096 72864 6112 72928
rect 6176 72864 6192 72928
rect 6256 72864 6264 72928
rect 5944 71840 6264 72864
rect 5944 71776 5952 71840
rect 6016 71776 6032 71840
rect 6096 71776 6112 71840
rect 6176 71776 6192 71840
rect 6256 71776 6264 71840
rect 5944 70752 6264 71776
rect 5944 70688 5952 70752
rect 6016 70688 6032 70752
rect 6096 70688 6112 70752
rect 6176 70688 6192 70752
rect 6256 70688 6264 70752
rect 5944 69664 6264 70688
rect 5944 69600 5952 69664
rect 6016 69600 6032 69664
rect 6096 69600 6112 69664
rect 6176 69600 6192 69664
rect 6256 69600 6264 69664
rect 5944 68576 6264 69600
rect 5944 68512 5952 68576
rect 6016 68512 6032 68576
rect 6096 68512 6112 68576
rect 6176 68512 6192 68576
rect 6256 68512 6264 68576
rect 5944 67488 6264 68512
rect 5944 67424 5952 67488
rect 6016 67424 6032 67488
rect 6096 67424 6112 67488
rect 6176 67424 6192 67488
rect 6256 67424 6264 67488
rect 5944 66400 6264 67424
rect 5944 66336 5952 66400
rect 6016 66336 6032 66400
rect 6096 66336 6112 66400
rect 6176 66336 6192 66400
rect 6256 66336 6264 66400
rect 5944 65312 6264 66336
rect 5944 65248 5952 65312
rect 6016 65248 6032 65312
rect 6096 65248 6112 65312
rect 6176 65248 6192 65312
rect 6256 65248 6264 65312
rect 5944 64224 6264 65248
rect 5944 64160 5952 64224
rect 6016 64160 6032 64224
rect 6096 64160 6112 64224
rect 6176 64160 6192 64224
rect 6256 64160 6264 64224
rect 5944 63136 6264 64160
rect 5944 63072 5952 63136
rect 6016 63072 6032 63136
rect 6096 63072 6112 63136
rect 6176 63072 6192 63136
rect 6256 63072 6264 63136
rect 5944 62048 6264 63072
rect 5944 61984 5952 62048
rect 6016 61984 6032 62048
rect 6096 61984 6112 62048
rect 6176 61984 6192 62048
rect 6256 61984 6264 62048
rect 5944 60960 6264 61984
rect 5944 60896 5952 60960
rect 6016 60896 6032 60960
rect 6096 60896 6112 60960
rect 6176 60896 6192 60960
rect 6256 60896 6264 60960
rect 5944 59872 6264 60896
rect 5944 59808 5952 59872
rect 6016 59808 6032 59872
rect 6096 59808 6112 59872
rect 6176 59808 6192 59872
rect 6256 59808 6264 59872
rect 5944 58784 6264 59808
rect 5944 58720 5952 58784
rect 6016 58720 6032 58784
rect 6096 58720 6112 58784
rect 6176 58720 6192 58784
rect 6256 58720 6264 58784
rect 5944 57696 6264 58720
rect 5944 57632 5952 57696
rect 6016 57632 6032 57696
rect 6096 57632 6112 57696
rect 6176 57632 6192 57696
rect 6256 57632 6264 57696
rect 5944 56608 6264 57632
rect 5944 56544 5952 56608
rect 6016 56544 6032 56608
rect 6096 56544 6112 56608
rect 6176 56544 6192 56608
rect 6256 56544 6264 56608
rect 5944 55520 6264 56544
rect 5944 55456 5952 55520
rect 6016 55456 6032 55520
rect 6096 55456 6112 55520
rect 6176 55456 6192 55520
rect 6256 55456 6264 55520
rect 5944 54432 6264 55456
rect 5944 54368 5952 54432
rect 6016 54368 6032 54432
rect 6096 54368 6112 54432
rect 6176 54368 6192 54432
rect 6256 54368 6264 54432
rect 5944 53344 6264 54368
rect 5944 53280 5952 53344
rect 6016 53280 6032 53344
rect 6096 53280 6112 53344
rect 6176 53280 6192 53344
rect 6256 53280 6264 53344
rect 5944 52256 6264 53280
rect 5944 52192 5952 52256
rect 6016 52192 6032 52256
rect 6096 52192 6112 52256
rect 6176 52192 6192 52256
rect 6256 52192 6264 52256
rect 5944 51168 6264 52192
rect 5944 51104 5952 51168
rect 6016 51104 6032 51168
rect 6096 51104 6112 51168
rect 6176 51104 6192 51168
rect 6256 51104 6264 51168
rect 5944 50080 6264 51104
rect 5944 50016 5952 50080
rect 6016 50016 6032 50080
rect 6096 50016 6112 50080
rect 6176 50016 6192 50080
rect 6256 50016 6264 50080
rect 5944 48992 6264 50016
rect 5944 48928 5952 48992
rect 6016 48928 6032 48992
rect 6096 48928 6112 48992
rect 6176 48928 6192 48992
rect 6256 48928 6264 48992
rect 5944 47904 6264 48928
rect 5944 47840 5952 47904
rect 6016 47840 6032 47904
rect 6096 47840 6112 47904
rect 6176 47840 6192 47904
rect 6256 47840 6264 47904
rect 5944 46816 6264 47840
rect 5944 46752 5952 46816
rect 6016 46752 6032 46816
rect 6096 46752 6112 46816
rect 6176 46752 6192 46816
rect 6256 46752 6264 46816
rect 5944 45728 6264 46752
rect 5944 45664 5952 45728
rect 6016 45664 6032 45728
rect 6096 45664 6112 45728
rect 6176 45664 6192 45728
rect 6256 45664 6264 45728
rect 5944 44640 6264 45664
rect 5944 44576 5952 44640
rect 6016 44576 6032 44640
rect 6096 44576 6112 44640
rect 6176 44576 6192 44640
rect 6256 44576 6264 44640
rect 5944 43552 6264 44576
rect 5944 43488 5952 43552
rect 6016 43488 6032 43552
rect 6096 43488 6112 43552
rect 6176 43488 6192 43552
rect 6256 43488 6264 43552
rect 5944 42464 6264 43488
rect 5944 42400 5952 42464
rect 6016 42400 6032 42464
rect 6096 42400 6112 42464
rect 6176 42400 6192 42464
rect 6256 42400 6264 42464
rect 5944 41376 6264 42400
rect 5944 41312 5952 41376
rect 6016 41312 6032 41376
rect 6096 41312 6112 41376
rect 6176 41312 6192 41376
rect 6256 41312 6264 41376
rect 5944 40288 6264 41312
rect 5944 40224 5952 40288
rect 6016 40224 6032 40288
rect 6096 40224 6112 40288
rect 6176 40224 6192 40288
rect 6256 40224 6264 40288
rect 5944 39200 6264 40224
rect 5944 39136 5952 39200
rect 6016 39136 6032 39200
rect 6096 39136 6112 39200
rect 6176 39136 6192 39200
rect 6256 39136 6264 39200
rect 5944 38112 6264 39136
rect 5944 38048 5952 38112
rect 6016 38048 6032 38112
rect 6096 38048 6112 38112
rect 6176 38048 6192 38112
rect 6256 38048 6264 38112
rect 5944 37024 6264 38048
rect 5944 36960 5952 37024
rect 6016 36960 6032 37024
rect 6096 36960 6112 37024
rect 6176 36960 6192 37024
rect 6256 36960 6264 37024
rect 5944 35936 6264 36960
rect 5944 35872 5952 35936
rect 6016 35872 6032 35936
rect 6096 35872 6112 35936
rect 6176 35872 6192 35936
rect 6256 35872 6264 35936
rect 5944 34848 6264 35872
rect 5944 34784 5952 34848
rect 6016 34784 6032 34848
rect 6096 34784 6112 34848
rect 6176 34784 6192 34848
rect 6256 34784 6264 34848
rect 5944 33760 6264 34784
rect 5944 33696 5952 33760
rect 6016 33696 6032 33760
rect 6096 33696 6112 33760
rect 6176 33696 6192 33760
rect 6256 33696 6264 33760
rect 5944 32672 6264 33696
rect 5944 32608 5952 32672
rect 6016 32608 6032 32672
rect 6096 32608 6112 32672
rect 6176 32608 6192 32672
rect 6256 32608 6264 32672
rect 5944 31584 6264 32608
rect 5944 31520 5952 31584
rect 6016 31520 6032 31584
rect 6096 31520 6112 31584
rect 6176 31520 6192 31584
rect 6256 31520 6264 31584
rect 5944 30496 6264 31520
rect 5944 30432 5952 30496
rect 6016 30432 6032 30496
rect 6096 30432 6112 30496
rect 6176 30432 6192 30496
rect 6256 30432 6264 30496
rect 5944 29408 6264 30432
rect 5944 29344 5952 29408
rect 6016 29344 6032 29408
rect 6096 29344 6112 29408
rect 6176 29344 6192 29408
rect 6256 29344 6264 29408
rect 5944 28320 6264 29344
rect 5944 28256 5952 28320
rect 6016 28256 6032 28320
rect 6096 28256 6112 28320
rect 6176 28256 6192 28320
rect 6256 28256 6264 28320
rect 5944 27232 6264 28256
rect 5944 27168 5952 27232
rect 6016 27168 6032 27232
rect 6096 27168 6112 27232
rect 6176 27168 6192 27232
rect 6256 27168 6264 27232
rect 5944 26144 6264 27168
rect 5944 26080 5952 26144
rect 6016 26080 6032 26144
rect 6096 26080 6112 26144
rect 6176 26080 6192 26144
rect 6256 26080 6264 26144
rect 5944 25056 6264 26080
rect 5944 24992 5952 25056
rect 6016 24992 6032 25056
rect 6096 24992 6112 25056
rect 6176 24992 6192 25056
rect 6256 24992 6264 25056
rect 5944 23968 6264 24992
rect 5944 23904 5952 23968
rect 6016 23904 6032 23968
rect 6096 23904 6112 23968
rect 6176 23904 6192 23968
rect 6256 23904 6264 23968
rect 5944 22880 6264 23904
rect 5944 22816 5952 22880
rect 6016 22816 6032 22880
rect 6096 22816 6112 22880
rect 6176 22816 6192 22880
rect 6256 22816 6264 22880
rect 5944 21792 6264 22816
rect 5944 21728 5952 21792
rect 6016 21728 6032 21792
rect 6096 21728 6112 21792
rect 6176 21728 6192 21792
rect 6256 21728 6264 21792
rect 5944 20704 6264 21728
rect 5944 20640 5952 20704
rect 6016 20640 6032 20704
rect 6096 20640 6112 20704
rect 6176 20640 6192 20704
rect 6256 20640 6264 20704
rect 5944 19616 6264 20640
rect 5944 19552 5952 19616
rect 6016 19552 6032 19616
rect 6096 19552 6112 19616
rect 6176 19552 6192 19616
rect 6256 19552 6264 19616
rect 5944 18528 6264 19552
rect 5944 18464 5952 18528
rect 6016 18464 6032 18528
rect 6096 18464 6112 18528
rect 6176 18464 6192 18528
rect 6256 18464 6264 18528
rect 5944 17440 6264 18464
rect 5944 17376 5952 17440
rect 6016 17376 6032 17440
rect 6096 17376 6112 17440
rect 6176 17376 6192 17440
rect 6256 17376 6264 17440
rect 5944 16352 6264 17376
rect 5944 16288 5952 16352
rect 6016 16288 6032 16352
rect 6096 16288 6112 16352
rect 6176 16288 6192 16352
rect 6256 16288 6264 16352
rect 5944 15264 6264 16288
rect 5944 15200 5952 15264
rect 6016 15200 6032 15264
rect 6096 15200 6112 15264
rect 6176 15200 6192 15264
rect 6256 15200 6264 15264
rect 5944 14176 6264 15200
rect 5944 14112 5952 14176
rect 6016 14112 6032 14176
rect 6096 14112 6112 14176
rect 6176 14112 6192 14176
rect 6256 14112 6264 14176
rect 5944 13088 6264 14112
rect 5944 13024 5952 13088
rect 6016 13024 6032 13088
rect 6096 13024 6112 13088
rect 6176 13024 6192 13088
rect 6256 13024 6264 13088
rect 5944 12000 6264 13024
rect 5944 11936 5952 12000
rect 6016 11936 6032 12000
rect 6096 11936 6112 12000
rect 6176 11936 6192 12000
rect 6256 11936 6264 12000
rect 5944 10912 6264 11936
rect 5944 10848 5952 10912
rect 6016 10848 6032 10912
rect 6096 10848 6112 10912
rect 6176 10848 6192 10912
rect 6256 10848 6264 10912
rect 5944 9824 6264 10848
rect 5944 9760 5952 9824
rect 6016 9760 6032 9824
rect 6096 9760 6112 9824
rect 6176 9760 6192 9824
rect 6256 9760 6264 9824
rect 5944 8736 6264 9760
rect 5944 8672 5952 8736
rect 6016 8672 6032 8736
rect 6096 8672 6112 8736
rect 6176 8672 6192 8736
rect 6256 8672 6264 8736
rect 5944 7648 6264 8672
rect 5944 7584 5952 7648
rect 6016 7584 6032 7648
rect 6096 7584 6112 7648
rect 6176 7584 6192 7648
rect 6256 7584 6264 7648
rect 5944 6560 6264 7584
rect 5944 6496 5952 6560
rect 6016 6496 6032 6560
rect 6096 6496 6112 6560
rect 6176 6496 6192 6560
rect 6256 6496 6264 6560
rect 5944 5472 6264 6496
rect 5944 5408 5952 5472
rect 6016 5408 6032 5472
rect 6096 5408 6112 5472
rect 6176 5408 6192 5472
rect 6256 5408 6264 5472
rect 5944 4384 6264 5408
rect 5944 4320 5952 4384
rect 6016 4320 6032 4384
rect 6096 4320 6112 4384
rect 6176 4320 6192 4384
rect 6256 4320 6264 4384
rect 5944 3296 6264 4320
rect 5944 3232 5952 3296
rect 6016 3232 6032 3296
rect 6096 3232 6112 3296
rect 6176 3232 6192 3296
rect 6256 3232 6264 3296
rect 5944 2208 6264 3232
rect 5944 2144 5952 2208
rect 6016 2144 6032 2208
rect 6096 2144 6112 2208
rect 6176 2144 6192 2208
rect 6256 2144 6264 2208
rect 5944 2128 6264 2144
rect 7610 330240 7930 330800
rect 7610 330176 7618 330240
rect 7682 330176 7698 330240
rect 7762 330176 7778 330240
rect 7842 330176 7858 330240
rect 7922 330176 7930 330240
rect 7610 329152 7930 330176
rect 7610 329088 7618 329152
rect 7682 329088 7698 329152
rect 7762 329088 7778 329152
rect 7842 329088 7858 329152
rect 7922 329088 7930 329152
rect 7610 328064 7930 329088
rect 7610 328000 7618 328064
rect 7682 328000 7698 328064
rect 7762 328000 7778 328064
rect 7842 328000 7858 328064
rect 7922 328000 7930 328064
rect 7610 326976 7930 328000
rect 7610 326912 7618 326976
rect 7682 326912 7698 326976
rect 7762 326912 7778 326976
rect 7842 326912 7858 326976
rect 7922 326912 7930 326976
rect 7610 325888 7930 326912
rect 7610 325824 7618 325888
rect 7682 325824 7698 325888
rect 7762 325824 7778 325888
rect 7842 325824 7858 325888
rect 7922 325824 7930 325888
rect 7610 324800 7930 325824
rect 7610 324736 7618 324800
rect 7682 324736 7698 324800
rect 7762 324736 7778 324800
rect 7842 324736 7858 324800
rect 7922 324736 7930 324800
rect 7610 323712 7930 324736
rect 7610 323648 7618 323712
rect 7682 323648 7698 323712
rect 7762 323648 7778 323712
rect 7842 323648 7858 323712
rect 7922 323648 7930 323712
rect 7610 322624 7930 323648
rect 7610 322560 7618 322624
rect 7682 322560 7698 322624
rect 7762 322560 7778 322624
rect 7842 322560 7858 322624
rect 7922 322560 7930 322624
rect 7610 321536 7930 322560
rect 7610 321472 7618 321536
rect 7682 321472 7698 321536
rect 7762 321472 7778 321536
rect 7842 321472 7858 321536
rect 7922 321472 7930 321536
rect 7610 320448 7930 321472
rect 7610 320384 7618 320448
rect 7682 320384 7698 320448
rect 7762 320384 7778 320448
rect 7842 320384 7858 320448
rect 7922 320384 7930 320448
rect 7610 319360 7930 320384
rect 7610 319296 7618 319360
rect 7682 319296 7698 319360
rect 7762 319296 7778 319360
rect 7842 319296 7858 319360
rect 7922 319296 7930 319360
rect 7610 318272 7930 319296
rect 7610 318208 7618 318272
rect 7682 318208 7698 318272
rect 7762 318208 7778 318272
rect 7842 318208 7858 318272
rect 7922 318208 7930 318272
rect 7610 317184 7930 318208
rect 7610 317120 7618 317184
rect 7682 317120 7698 317184
rect 7762 317120 7778 317184
rect 7842 317120 7858 317184
rect 7922 317120 7930 317184
rect 7610 316096 7930 317120
rect 7610 316032 7618 316096
rect 7682 316032 7698 316096
rect 7762 316032 7778 316096
rect 7842 316032 7858 316096
rect 7922 316032 7930 316096
rect 7610 315008 7930 316032
rect 7610 314944 7618 315008
rect 7682 314944 7698 315008
rect 7762 314944 7778 315008
rect 7842 314944 7858 315008
rect 7922 314944 7930 315008
rect 7610 313920 7930 314944
rect 7610 313856 7618 313920
rect 7682 313856 7698 313920
rect 7762 313856 7778 313920
rect 7842 313856 7858 313920
rect 7922 313856 7930 313920
rect 7610 312832 7930 313856
rect 7610 312768 7618 312832
rect 7682 312768 7698 312832
rect 7762 312768 7778 312832
rect 7842 312768 7858 312832
rect 7922 312768 7930 312832
rect 7610 311744 7930 312768
rect 7610 311680 7618 311744
rect 7682 311680 7698 311744
rect 7762 311680 7778 311744
rect 7842 311680 7858 311744
rect 7922 311680 7930 311744
rect 7610 310656 7930 311680
rect 7610 310592 7618 310656
rect 7682 310592 7698 310656
rect 7762 310592 7778 310656
rect 7842 310592 7858 310656
rect 7922 310592 7930 310656
rect 7610 309568 7930 310592
rect 7610 309504 7618 309568
rect 7682 309504 7698 309568
rect 7762 309504 7778 309568
rect 7842 309504 7858 309568
rect 7922 309504 7930 309568
rect 7610 308480 7930 309504
rect 7610 308416 7618 308480
rect 7682 308416 7698 308480
rect 7762 308416 7778 308480
rect 7842 308416 7858 308480
rect 7922 308416 7930 308480
rect 7610 307392 7930 308416
rect 7610 307328 7618 307392
rect 7682 307328 7698 307392
rect 7762 307328 7778 307392
rect 7842 307328 7858 307392
rect 7922 307328 7930 307392
rect 7610 306304 7930 307328
rect 7610 306240 7618 306304
rect 7682 306240 7698 306304
rect 7762 306240 7778 306304
rect 7842 306240 7858 306304
rect 7922 306240 7930 306304
rect 7610 305216 7930 306240
rect 7610 305152 7618 305216
rect 7682 305152 7698 305216
rect 7762 305152 7778 305216
rect 7842 305152 7858 305216
rect 7922 305152 7930 305216
rect 7610 304128 7930 305152
rect 7610 304064 7618 304128
rect 7682 304064 7698 304128
rect 7762 304064 7778 304128
rect 7842 304064 7858 304128
rect 7922 304064 7930 304128
rect 7610 303040 7930 304064
rect 7610 302976 7618 303040
rect 7682 302976 7698 303040
rect 7762 302976 7778 303040
rect 7842 302976 7858 303040
rect 7922 302976 7930 303040
rect 7610 301952 7930 302976
rect 7610 301888 7618 301952
rect 7682 301888 7698 301952
rect 7762 301888 7778 301952
rect 7842 301888 7858 301952
rect 7922 301888 7930 301952
rect 7610 300864 7930 301888
rect 7610 300800 7618 300864
rect 7682 300800 7698 300864
rect 7762 300800 7778 300864
rect 7842 300800 7858 300864
rect 7922 300800 7930 300864
rect 7610 299776 7930 300800
rect 7610 299712 7618 299776
rect 7682 299712 7698 299776
rect 7762 299712 7778 299776
rect 7842 299712 7858 299776
rect 7922 299712 7930 299776
rect 7610 298688 7930 299712
rect 7610 298624 7618 298688
rect 7682 298624 7698 298688
rect 7762 298624 7778 298688
rect 7842 298624 7858 298688
rect 7922 298624 7930 298688
rect 7610 297600 7930 298624
rect 7610 297536 7618 297600
rect 7682 297536 7698 297600
rect 7762 297536 7778 297600
rect 7842 297536 7858 297600
rect 7922 297536 7930 297600
rect 7610 296512 7930 297536
rect 7610 296448 7618 296512
rect 7682 296448 7698 296512
rect 7762 296448 7778 296512
rect 7842 296448 7858 296512
rect 7922 296448 7930 296512
rect 7610 295424 7930 296448
rect 7610 295360 7618 295424
rect 7682 295360 7698 295424
rect 7762 295360 7778 295424
rect 7842 295360 7858 295424
rect 7922 295360 7930 295424
rect 7610 294336 7930 295360
rect 7610 294272 7618 294336
rect 7682 294272 7698 294336
rect 7762 294272 7778 294336
rect 7842 294272 7858 294336
rect 7922 294272 7930 294336
rect 7610 293248 7930 294272
rect 7610 293184 7618 293248
rect 7682 293184 7698 293248
rect 7762 293184 7778 293248
rect 7842 293184 7858 293248
rect 7922 293184 7930 293248
rect 7610 292160 7930 293184
rect 7610 292096 7618 292160
rect 7682 292096 7698 292160
rect 7762 292096 7778 292160
rect 7842 292096 7858 292160
rect 7922 292096 7930 292160
rect 7610 291072 7930 292096
rect 7610 291008 7618 291072
rect 7682 291008 7698 291072
rect 7762 291008 7778 291072
rect 7842 291008 7858 291072
rect 7922 291008 7930 291072
rect 7610 289984 7930 291008
rect 7610 289920 7618 289984
rect 7682 289920 7698 289984
rect 7762 289920 7778 289984
rect 7842 289920 7858 289984
rect 7922 289920 7930 289984
rect 7610 288896 7930 289920
rect 7610 288832 7618 288896
rect 7682 288832 7698 288896
rect 7762 288832 7778 288896
rect 7842 288832 7858 288896
rect 7922 288832 7930 288896
rect 7610 287808 7930 288832
rect 7610 287744 7618 287808
rect 7682 287744 7698 287808
rect 7762 287744 7778 287808
rect 7842 287744 7858 287808
rect 7922 287744 7930 287808
rect 7610 286720 7930 287744
rect 7610 286656 7618 286720
rect 7682 286656 7698 286720
rect 7762 286656 7778 286720
rect 7842 286656 7858 286720
rect 7922 286656 7930 286720
rect 7610 285632 7930 286656
rect 7610 285568 7618 285632
rect 7682 285568 7698 285632
rect 7762 285568 7778 285632
rect 7842 285568 7858 285632
rect 7922 285568 7930 285632
rect 7610 284544 7930 285568
rect 7610 284480 7618 284544
rect 7682 284480 7698 284544
rect 7762 284480 7778 284544
rect 7842 284480 7858 284544
rect 7922 284480 7930 284544
rect 7610 283456 7930 284480
rect 7610 283392 7618 283456
rect 7682 283392 7698 283456
rect 7762 283392 7778 283456
rect 7842 283392 7858 283456
rect 7922 283392 7930 283456
rect 7610 282368 7930 283392
rect 7610 282304 7618 282368
rect 7682 282304 7698 282368
rect 7762 282304 7778 282368
rect 7842 282304 7858 282368
rect 7922 282304 7930 282368
rect 7610 281280 7930 282304
rect 7610 281216 7618 281280
rect 7682 281216 7698 281280
rect 7762 281216 7778 281280
rect 7842 281216 7858 281280
rect 7922 281216 7930 281280
rect 7610 280192 7930 281216
rect 7610 280128 7618 280192
rect 7682 280128 7698 280192
rect 7762 280128 7778 280192
rect 7842 280128 7858 280192
rect 7922 280128 7930 280192
rect 7610 279104 7930 280128
rect 7610 279040 7618 279104
rect 7682 279040 7698 279104
rect 7762 279040 7778 279104
rect 7842 279040 7858 279104
rect 7922 279040 7930 279104
rect 7610 278016 7930 279040
rect 7610 277952 7618 278016
rect 7682 277952 7698 278016
rect 7762 277952 7778 278016
rect 7842 277952 7858 278016
rect 7922 277952 7930 278016
rect 7610 276928 7930 277952
rect 7610 276864 7618 276928
rect 7682 276864 7698 276928
rect 7762 276864 7778 276928
rect 7842 276864 7858 276928
rect 7922 276864 7930 276928
rect 7610 275840 7930 276864
rect 7610 275776 7618 275840
rect 7682 275776 7698 275840
rect 7762 275776 7778 275840
rect 7842 275776 7858 275840
rect 7922 275776 7930 275840
rect 7610 274752 7930 275776
rect 7610 274688 7618 274752
rect 7682 274688 7698 274752
rect 7762 274688 7778 274752
rect 7842 274688 7858 274752
rect 7922 274688 7930 274752
rect 7610 273664 7930 274688
rect 7610 273600 7618 273664
rect 7682 273600 7698 273664
rect 7762 273600 7778 273664
rect 7842 273600 7858 273664
rect 7922 273600 7930 273664
rect 7610 272576 7930 273600
rect 7610 272512 7618 272576
rect 7682 272512 7698 272576
rect 7762 272512 7778 272576
rect 7842 272512 7858 272576
rect 7922 272512 7930 272576
rect 7610 271488 7930 272512
rect 7610 271424 7618 271488
rect 7682 271424 7698 271488
rect 7762 271424 7778 271488
rect 7842 271424 7858 271488
rect 7922 271424 7930 271488
rect 7610 270400 7930 271424
rect 7610 270336 7618 270400
rect 7682 270336 7698 270400
rect 7762 270336 7778 270400
rect 7842 270336 7858 270400
rect 7922 270336 7930 270400
rect 7610 269312 7930 270336
rect 7610 269248 7618 269312
rect 7682 269248 7698 269312
rect 7762 269248 7778 269312
rect 7842 269248 7858 269312
rect 7922 269248 7930 269312
rect 7610 268224 7930 269248
rect 7610 268160 7618 268224
rect 7682 268160 7698 268224
rect 7762 268160 7778 268224
rect 7842 268160 7858 268224
rect 7922 268160 7930 268224
rect 7610 267136 7930 268160
rect 7610 267072 7618 267136
rect 7682 267072 7698 267136
rect 7762 267072 7778 267136
rect 7842 267072 7858 267136
rect 7922 267072 7930 267136
rect 7610 266048 7930 267072
rect 7610 265984 7618 266048
rect 7682 265984 7698 266048
rect 7762 265984 7778 266048
rect 7842 265984 7858 266048
rect 7922 265984 7930 266048
rect 7610 264960 7930 265984
rect 7610 264896 7618 264960
rect 7682 264896 7698 264960
rect 7762 264896 7778 264960
rect 7842 264896 7858 264960
rect 7922 264896 7930 264960
rect 7610 263872 7930 264896
rect 7610 263808 7618 263872
rect 7682 263808 7698 263872
rect 7762 263808 7778 263872
rect 7842 263808 7858 263872
rect 7922 263808 7930 263872
rect 7610 262784 7930 263808
rect 7610 262720 7618 262784
rect 7682 262720 7698 262784
rect 7762 262720 7778 262784
rect 7842 262720 7858 262784
rect 7922 262720 7930 262784
rect 7610 261696 7930 262720
rect 7610 261632 7618 261696
rect 7682 261632 7698 261696
rect 7762 261632 7778 261696
rect 7842 261632 7858 261696
rect 7922 261632 7930 261696
rect 7610 260608 7930 261632
rect 7610 260544 7618 260608
rect 7682 260544 7698 260608
rect 7762 260544 7778 260608
rect 7842 260544 7858 260608
rect 7922 260544 7930 260608
rect 7610 259520 7930 260544
rect 7610 259456 7618 259520
rect 7682 259456 7698 259520
rect 7762 259456 7778 259520
rect 7842 259456 7858 259520
rect 7922 259456 7930 259520
rect 7610 258432 7930 259456
rect 7610 258368 7618 258432
rect 7682 258368 7698 258432
rect 7762 258368 7778 258432
rect 7842 258368 7858 258432
rect 7922 258368 7930 258432
rect 7610 257344 7930 258368
rect 7610 257280 7618 257344
rect 7682 257280 7698 257344
rect 7762 257280 7778 257344
rect 7842 257280 7858 257344
rect 7922 257280 7930 257344
rect 7610 256256 7930 257280
rect 7610 256192 7618 256256
rect 7682 256192 7698 256256
rect 7762 256192 7778 256256
rect 7842 256192 7858 256256
rect 7922 256192 7930 256256
rect 7610 255168 7930 256192
rect 7610 255104 7618 255168
rect 7682 255104 7698 255168
rect 7762 255104 7778 255168
rect 7842 255104 7858 255168
rect 7922 255104 7930 255168
rect 7610 254080 7930 255104
rect 7610 254016 7618 254080
rect 7682 254016 7698 254080
rect 7762 254016 7778 254080
rect 7842 254016 7858 254080
rect 7922 254016 7930 254080
rect 7610 252992 7930 254016
rect 7610 252928 7618 252992
rect 7682 252928 7698 252992
rect 7762 252928 7778 252992
rect 7842 252928 7858 252992
rect 7922 252928 7930 252992
rect 7610 251904 7930 252928
rect 7610 251840 7618 251904
rect 7682 251840 7698 251904
rect 7762 251840 7778 251904
rect 7842 251840 7858 251904
rect 7922 251840 7930 251904
rect 7610 250816 7930 251840
rect 7610 250752 7618 250816
rect 7682 250752 7698 250816
rect 7762 250752 7778 250816
rect 7842 250752 7858 250816
rect 7922 250752 7930 250816
rect 7610 249728 7930 250752
rect 7610 249664 7618 249728
rect 7682 249664 7698 249728
rect 7762 249664 7778 249728
rect 7842 249664 7858 249728
rect 7922 249664 7930 249728
rect 7610 248640 7930 249664
rect 7610 248576 7618 248640
rect 7682 248576 7698 248640
rect 7762 248576 7778 248640
rect 7842 248576 7858 248640
rect 7922 248576 7930 248640
rect 7610 247552 7930 248576
rect 7610 247488 7618 247552
rect 7682 247488 7698 247552
rect 7762 247488 7778 247552
rect 7842 247488 7858 247552
rect 7922 247488 7930 247552
rect 7610 246464 7930 247488
rect 7610 246400 7618 246464
rect 7682 246400 7698 246464
rect 7762 246400 7778 246464
rect 7842 246400 7858 246464
rect 7922 246400 7930 246464
rect 7610 245376 7930 246400
rect 7610 245312 7618 245376
rect 7682 245312 7698 245376
rect 7762 245312 7778 245376
rect 7842 245312 7858 245376
rect 7922 245312 7930 245376
rect 7610 244288 7930 245312
rect 7610 244224 7618 244288
rect 7682 244224 7698 244288
rect 7762 244224 7778 244288
rect 7842 244224 7858 244288
rect 7922 244224 7930 244288
rect 7610 243200 7930 244224
rect 7610 243136 7618 243200
rect 7682 243136 7698 243200
rect 7762 243136 7778 243200
rect 7842 243136 7858 243200
rect 7922 243136 7930 243200
rect 7610 242112 7930 243136
rect 7610 242048 7618 242112
rect 7682 242048 7698 242112
rect 7762 242048 7778 242112
rect 7842 242048 7858 242112
rect 7922 242048 7930 242112
rect 7610 241024 7930 242048
rect 7610 240960 7618 241024
rect 7682 240960 7698 241024
rect 7762 240960 7778 241024
rect 7842 240960 7858 241024
rect 7922 240960 7930 241024
rect 7610 239936 7930 240960
rect 7610 239872 7618 239936
rect 7682 239872 7698 239936
rect 7762 239872 7778 239936
rect 7842 239872 7858 239936
rect 7922 239872 7930 239936
rect 7610 238848 7930 239872
rect 7610 238784 7618 238848
rect 7682 238784 7698 238848
rect 7762 238784 7778 238848
rect 7842 238784 7858 238848
rect 7922 238784 7930 238848
rect 7610 237760 7930 238784
rect 7610 237696 7618 237760
rect 7682 237696 7698 237760
rect 7762 237696 7778 237760
rect 7842 237696 7858 237760
rect 7922 237696 7930 237760
rect 7610 236672 7930 237696
rect 7610 236608 7618 236672
rect 7682 236608 7698 236672
rect 7762 236608 7778 236672
rect 7842 236608 7858 236672
rect 7922 236608 7930 236672
rect 7610 235584 7930 236608
rect 7610 235520 7618 235584
rect 7682 235520 7698 235584
rect 7762 235520 7778 235584
rect 7842 235520 7858 235584
rect 7922 235520 7930 235584
rect 7610 234496 7930 235520
rect 7610 234432 7618 234496
rect 7682 234432 7698 234496
rect 7762 234432 7778 234496
rect 7842 234432 7858 234496
rect 7922 234432 7930 234496
rect 7610 233408 7930 234432
rect 7610 233344 7618 233408
rect 7682 233344 7698 233408
rect 7762 233344 7778 233408
rect 7842 233344 7858 233408
rect 7922 233344 7930 233408
rect 7610 232320 7930 233344
rect 7610 232256 7618 232320
rect 7682 232256 7698 232320
rect 7762 232256 7778 232320
rect 7842 232256 7858 232320
rect 7922 232256 7930 232320
rect 7610 231232 7930 232256
rect 7610 231168 7618 231232
rect 7682 231168 7698 231232
rect 7762 231168 7778 231232
rect 7842 231168 7858 231232
rect 7922 231168 7930 231232
rect 7610 230144 7930 231168
rect 7610 230080 7618 230144
rect 7682 230080 7698 230144
rect 7762 230080 7778 230144
rect 7842 230080 7858 230144
rect 7922 230080 7930 230144
rect 7610 229056 7930 230080
rect 7610 228992 7618 229056
rect 7682 228992 7698 229056
rect 7762 228992 7778 229056
rect 7842 228992 7858 229056
rect 7922 228992 7930 229056
rect 7610 227968 7930 228992
rect 7610 227904 7618 227968
rect 7682 227904 7698 227968
rect 7762 227904 7778 227968
rect 7842 227904 7858 227968
rect 7922 227904 7930 227968
rect 7610 226880 7930 227904
rect 7610 226816 7618 226880
rect 7682 226816 7698 226880
rect 7762 226816 7778 226880
rect 7842 226816 7858 226880
rect 7922 226816 7930 226880
rect 7610 225792 7930 226816
rect 7610 225728 7618 225792
rect 7682 225728 7698 225792
rect 7762 225728 7778 225792
rect 7842 225728 7858 225792
rect 7922 225728 7930 225792
rect 7610 224704 7930 225728
rect 7610 224640 7618 224704
rect 7682 224640 7698 224704
rect 7762 224640 7778 224704
rect 7842 224640 7858 224704
rect 7922 224640 7930 224704
rect 7610 223616 7930 224640
rect 7610 223552 7618 223616
rect 7682 223552 7698 223616
rect 7762 223552 7778 223616
rect 7842 223552 7858 223616
rect 7922 223552 7930 223616
rect 7610 222528 7930 223552
rect 7610 222464 7618 222528
rect 7682 222464 7698 222528
rect 7762 222464 7778 222528
rect 7842 222464 7858 222528
rect 7922 222464 7930 222528
rect 7610 221440 7930 222464
rect 7610 221376 7618 221440
rect 7682 221376 7698 221440
rect 7762 221376 7778 221440
rect 7842 221376 7858 221440
rect 7922 221376 7930 221440
rect 7610 220352 7930 221376
rect 7610 220288 7618 220352
rect 7682 220288 7698 220352
rect 7762 220288 7778 220352
rect 7842 220288 7858 220352
rect 7922 220288 7930 220352
rect 7610 219264 7930 220288
rect 7610 219200 7618 219264
rect 7682 219200 7698 219264
rect 7762 219200 7778 219264
rect 7842 219200 7858 219264
rect 7922 219200 7930 219264
rect 7610 218176 7930 219200
rect 7610 218112 7618 218176
rect 7682 218112 7698 218176
rect 7762 218112 7778 218176
rect 7842 218112 7858 218176
rect 7922 218112 7930 218176
rect 7610 217088 7930 218112
rect 7610 217024 7618 217088
rect 7682 217024 7698 217088
rect 7762 217024 7778 217088
rect 7842 217024 7858 217088
rect 7922 217024 7930 217088
rect 7610 216000 7930 217024
rect 7610 215936 7618 216000
rect 7682 215936 7698 216000
rect 7762 215936 7778 216000
rect 7842 215936 7858 216000
rect 7922 215936 7930 216000
rect 7610 214912 7930 215936
rect 7610 214848 7618 214912
rect 7682 214848 7698 214912
rect 7762 214848 7778 214912
rect 7842 214848 7858 214912
rect 7922 214848 7930 214912
rect 7610 213824 7930 214848
rect 7610 213760 7618 213824
rect 7682 213760 7698 213824
rect 7762 213760 7778 213824
rect 7842 213760 7858 213824
rect 7922 213760 7930 213824
rect 7610 212736 7930 213760
rect 7610 212672 7618 212736
rect 7682 212672 7698 212736
rect 7762 212672 7778 212736
rect 7842 212672 7858 212736
rect 7922 212672 7930 212736
rect 7610 211648 7930 212672
rect 7610 211584 7618 211648
rect 7682 211584 7698 211648
rect 7762 211584 7778 211648
rect 7842 211584 7858 211648
rect 7922 211584 7930 211648
rect 7610 210560 7930 211584
rect 7610 210496 7618 210560
rect 7682 210496 7698 210560
rect 7762 210496 7778 210560
rect 7842 210496 7858 210560
rect 7922 210496 7930 210560
rect 7610 209472 7930 210496
rect 7610 209408 7618 209472
rect 7682 209408 7698 209472
rect 7762 209408 7778 209472
rect 7842 209408 7858 209472
rect 7922 209408 7930 209472
rect 7610 208384 7930 209408
rect 7610 208320 7618 208384
rect 7682 208320 7698 208384
rect 7762 208320 7778 208384
rect 7842 208320 7858 208384
rect 7922 208320 7930 208384
rect 7610 207296 7930 208320
rect 7610 207232 7618 207296
rect 7682 207232 7698 207296
rect 7762 207232 7778 207296
rect 7842 207232 7858 207296
rect 7922 207232 7930 207296
rect 7610 206208 7930 207232
rect 7610 206144 7618 206208
rect 7682 206144 7698 206208
rect 7762 206144 7778 206208
rect 7842 206144 7858 206208
rect 7922 206144 7930 206208
rect 7610 205120 7930 206144
rect 7610 205056 7618 205120
rect 7682 205056 7698 205120
rect 7762 205056 7778 205120
rect 7842 205056 7858 205120
rect 7922 205056 7930 205120
rect 7610 204032 7930 205056
rect 7610 203968 7618 204032
rect 7682 203968 7698 204032
rect 7762 203968 7778 204032
rect 7842 203968 7858 204032
rect 7922 203968 7930 204032
rect 7610 202944 7930 203968
rect 7610 202880 7618 202944
rect 7682 202880 7698 202944
rect 7762 202880 7778 202944
rect 7842 202880 7858 202944
rect 7922 202880 7930 202944
rect 7610 201856 7930 202880
rect 7610 201792 7618 201856
rect 7682 201792 7698 201856
rect 7762 201792 7778 201856
rect 7842 201792 7858 201856
rect 7922 201792 7930 201856
rect 7610 200768 7930 201792
rect 7610 200704 7618 200768
rect 7682 200704 7698 200768
rect 7762 200704 7778 200768
rect 7842 200704 7858 200768
rect 7922 200704 7930 200768
rect 7610 199680 7930 200704
rect 7610 199616 7618 199680
rect 7682 199616 7698 199680
rect 7762 199616 7778 199680
rect 7842 199616 7858 199680
rect 7922 199616 7930 199680
rect 7610 198592 7930 199616
rect 7610 198528 7618 198592
rect 7682 198528 7698 198592
rect 7762 198528 7778 198592
rect 7842 198528 7858 198592
rect 7922 198528 7930 198592
rect 7610 197504 7930 198528
rect 7610 197440 7618 197504
rect 7682 197440 7698 197504
rect 7762 197440 7778 197504
rect 7842 197440 7858 197504
rect 7922 197440 7930 197504
rect 7610 196416 7930 197440
rect 7610 196352 7618 196416
rect 7682 196352 7698 196416
rect 7762 196352 7778 196416
rect 7842 196352 7858 196416
rect 7922 196352 7930 196416
rect 7610 195328 7930 196352
rect 7610 195264 7618 195328
rect 7682 195264 7698 195328
rect 7762 195264 7778 195328
rect 7842 195264 7858 195328
rect 7922 195264 7930 195328
rect 7610 194240 7930 195264
rect 7610 194176 7618 194240
rect 7682 194176 7698 194240
rect 7762 194176 7778 194240
rect 7842 194176 7858 194240
rect 7922 194176 7930 194240
rect 7610 193152 7930 194176
rect 7610 193088 7618 193152
rect 7682 193088 7698 193152
rect 7762 193088 7778 193152
rect 7842 193088 7858 193152
rect 7922 193088 7930 193152
rect 7610 192064 7930 193088
rect 7610 192000 7618 192064
rect 7682 192000 7698 192064
rect 7762 192000 7778 192064
rect 7842 192000 7858 192064
rect 7922 192000 7930 192064
rect 7610 190976 7930 192000
rect 7610 190912 7618 190976
rect 7682 190912 7698 190976
rect 7762 190912 7778 190976
rect 7842 190912 7858 190976
rect 7922 190912 7930 190976
rect 7610 189888 7930 190912
rect 7610 189824 7618 189888
rect 7682 189824 7698 189888
rect 7762 189824 7778 189888
rect 7842 189824 7858 189888
rect 7922 189824 7930 189888
rect 7610 188800 7930 189824
rect 7610 188736 7618 188800
rect 7682 188736 7698 188800
rect 7762 188736 7778 188800
rect 7842 188736 7858 188800
rect 7922 188736 7930 188800
rect 7610 187712 7930 188736
rect 7610 187648 7618 187712
rect 7682 187648 7698 187712
rect 7762 187648 7778 187712
rect 7842 187648 7858 187712
rect 7922 187648 7930 187712
rect 7610 186624 7930 187648
rect 7610 186560 7618 186624
rect 7682 186560 7698 186624
rect 7762 186560 7778 186624
rect 7842 186560 7858 186624
rect 7922 186560 7930 186624
rect 7610 185536 7930 186560
rect 7610 185472 7618 185536
rect 7682 185472 7698 185536
rect 7762 185472 7778 185536
rect 7842 185472 7858 185536
rect 7922 185472 7930 185536
rect 7610 184448 7930 185472
rect 7610 184384 7618 184448
rect 7682 184384 7698 184448
rect 7762 184384 7778 184448
rect 7842 184384 7858 184448
rect 7922 184384 7930 184448
rect 7610 183360 7930 184384
rect 7610 183296 7618 183360
rect 7682 183296 7698 183360
rect 7762 183296 7778 183360
rect 7842 183296 7858 183360
rect 7922 183296 7930 183360
rect 7610 182272 7930 183296
rect 7610 182208 7618 182272
rect 7682 182208 7698 182272
rect 7762 182208 7778 182272
rect 7842 182208 7858 182272
rect 7922 182208 7930 182272
rect 7610 181184 7930 182208
rect 7610 181120 7618 181184
rect 7682 181120 7698 181184
rect 7762 181120 7778 181184
rect 7842 181120 7858 181184
rect 7922 181120 7930 181184
rect 7610 180096 7930 181120
rect 7610 180032 7618 180096
rect 7682 180032 7698 180096
rect 7762 180032 7778 180096
rect 7842 180032 7858 180096
rect 7922 180032 7930 180096
rect 7610 179008 7930 180032
rect 7610 178944 7618 179008
rect 7682 178944 7698 179008
rect 7762 178944 7778 179008
rect 7842 178944 7858 179008
rect 7922 178944 7930 179008
rect 7610 177920 7930 178944
rect 7610 177856 7618 177920
rect 7682 177856 7698 177920
rect 7762 177856 7778 177920
rect 7842 177856 7858 177920
rect 7922 177856 7930 177920
rect 7610 176832 7930 177856
rect 7610 176768 7618 176832
rect 7682 176768 7698 176832
rect 7762 176768 7778 176832
rect 7842 176768 7858 176832
rect 7922 176768 7930 176832
rect 7610 175744 7930 176768
rect 7610 175680 7618 175744
rect 7682 175680 7698 175744
rect 7762 175680 7778 175744
rect 7842 175680 7858 175744
rect 7922 175680 7930 175744
rect 7610 174656 7930 175680
rect 7610 174592 7618 174656
rect 7682 174592 7698 174656
rect 7762 174592 7778 174656
rect 7842 174592 7858 174656
rect 7922 174592 7930 174656
rect 7610 173568 7930 174592
rect 7610 173504 7618 173568
rect 7682 173504 7698 173568
rect 7762 173504 7778 173568
rect 7842 173504 7858 173568
rect 7922 173504 7930 173568
rect 7610 172480 7930 173504
rect 7610 172416 7618 172480
rect 7682 172416 7698 172480
rect 7762 172416 7778 172480
rect 7842 172416 7858 172480
rect 7922 172416 7930 172480
rect 7610 171392 7930 172416
rect 7610 171328 7618 171392
rect 7682 171328 7698 171392
rect 7762 171328 7778 171392
rect 7842 171328 7858 171392
rect 7922 171328 7930 171392
rect 7610 170304 7930 171328
rect 7610 170240 7618 170304
rect 7682 170240 7698 170304
rect 7762 170240 7778 170304
rect 7842 170240 7858 170304
rect 7922 170240 7930 170304
rect 7610 169216 7930 170240
rect 7610 169152 7618 169216
rect 7682 169152 7698 169216
rect 7762 169152 7778 169216
rect 7842 169152 7858 169216
rect 7922 169152 7930 169216
rect 7610 168128 7930 169152
rect 7610 168064 7618 168128
rect 7682 168064 7698 168128
rect 7762 168064 7778 168128
rect 7842 168064 7858 168128
rect 7922 168064 7930 168128
rect 7610 167040 7930 168064
rect 7610 166976 7618 167040
rect 7682 166976 7698 167040
rect 7762 166976 7778 167040
rect 7842 166976 7858 167040
rect 7922 166976 7930 167040
rect 7610 165952 7930 166976
rect 7610 165888 7618 165952
rect 7682 165888 7698 165952
rect 7762 165888 7778 165952
rect 7842 165888 7858 165952
rect 7922 165888 7930 165952
rect 7610 164864 7930 165888
rect 7610 164800 7618 164864
rect 7682 164800 7698 164864
rect 7762 164800 7778 164864
rect 7842 164800 7858 164864
rect 7922 164800 7930 164864
rect 7610 163776 7930 164800
rect 7610 163712 7618 163776
rect 7682 163712 7698 163776
rect 7762 163712 7778 163776
rect 7842 163712 7858 163776
rect 7922 163712 7930 163776
rect 7610 162688 7930 163712
rect 7610 162624 7618 162688
rect 7682 162624 7698 162688
rect 7762 162624 7778 162688
rect 7842 162624 7858 162688
rect 7922 162624 7930 162688
rect 7610 161600 7930 162624
rect 7610 161536 7618 161600
rect 7682 161536 7698 161600
rect 7762 161536 7778 161600
rect 7842 161536 7858 161600
rect 7922 161536 7930 161600
rect 7610 160512 7930 161536
rect 7610 160448 7618 160512
rect 7682 160448 7698 160512
rect 7762 160448 7778 160512
rect 7842 160448 7858 160512
rect 7922 160448 7930 160512
rect 7610 159424 7930 160448
rect 7610 159360 7618 159424
rect 7682 159360 7698 159424
rect 7762 159360 7778 159424
rect 7842 159360 7858 159424
rect 7922 159360 7930 159424
rect 7610 158336 7930 159360
rect 7610 158272 7618 158336
rect 7682 158272 7698 158336
rect 7762 158272 7778 158336
rect 7842 158272 7858 158336
rect 7922 158272 7930 158336
rect 7610 157248 7930 158272
rect 7610 157184 7618 157248
rect 7682 157184 7698 157248
rect 7762 157184 7778 157248
rect 7842 157184 7858 157248
rect 7922 157184 7930 157248
rect 7610 156160 7930 157184
rect 7610 156096 7618 156160
rect 7682 156096 7698 156160
rect 7762 156096 7778 156160
rect 7842 156096 7858 156160
rect 7922 156096 7930 156160
rect 7610 155072 7930 156096
rect 7610 155008 7618 155072
rect 7682 155008 7698 155072
rect 7762 155008 7778 155072
rect 7842 155008 7858 155072
rect 7922 155008 7930 155072
rect 7610 153984 7930 155008
rect 7610 153920 7618 153984
rect 7682 153920 7698 153984
rect 7762 153920 7778 153984
rect 7842 153920 7858 153984
rect 7922 153920 7930 153984
rect 7610 152896 7930 153920
rect 7610 152832 7618 152896
rect 7682 152832 7698 152896
rect 7762 152832 7778 152896
rect 7842 152832 7858 152896
rect 7922 152832 7930 152896
rect 7610 151808 7930 152832
rect 7610 151744 7618 151808
rect 7682 151744 7698 151808
rect 7762 151744 7778 151808
rect 7842 151744 7858 151808
rect 7922 151744 7930 151808
rect 7610 150720 7930 151744
rect 7610 150656 7618 150720
rect 7682 150656 7698 150720
rect 7762 150656 7778 150720
rect 7842 150656 7858 150720
rect 7922 150656 7930 150720
rect 7610 149632 7930 150656
rect 7610 149568 7618 149632
rect 7682 149568 7698 149632
rect 7762 149568 7778 149632
rect 7842 149568 7858 149632
rect 7922 149568 7930 149632
rect 7610 148544 7930 149568
rect 7610 148480 7618 148544
rect 7682 148480 7698 148544
rect 7762 148480 7778 148544
rect 7842 148480 7858 148544
rect 7922 148480 7930 148544
rect 7610 147456 7930 148480
rect 7610 147392 7618 147456
rect 7682 147392 7698 147456
rect 7762 147392 7778 147456
rect 7842 147392 7858 147456
rect 7922 147392 7930 147456
rect 7610 146368 7930 147392
rect 7610 146304 7618 146368
rect 7682 146304 7698 146368
rect 7762 146304 7778 146368
rect 7842 146304 7858 146368
rect 7922 146304 7930 146368
rect 7610 145280 7930 146304
rect 7610 145216 7618 145280
rect 7682 145216 7698 145280
rect 7762 145216 7778 145280
rect 7842 145216 7858 145280
rect 7922 145216 7930 145280
rect 7610 144192 7930 145216
rect 7610 144128 7618 144192
rect 7682 144128 7698 144192
rect 7762 144128 7778 144192
rect 7842 144128 7858 144192
rect 7922 144128 7930 144192
rect 7610 143104 7930 144128
rect 7610 143040 7618 143104
rect 7682 143040 7698 143104
rect 7762 143040 7778 143104
rect 7842 143040 7858 143104
rect 7922 143040 7930 143104
rect 7610 142016 7930 143040
rect 7610 141952 7618 142016
rect 7682 141952 7698 142016
rect 7762 141952 7778 142016
rect 7842 141952 7858 142016
rect 7922 141952 7930 142016
rect 7610 140928 7930 141952
rect 7610 140864 7618 140928
rect 7682 140864 7698 140928
rect 7762 140864 7778 140928
rect 7842 140864 7858 140928
rect 7922 140864 7930 140928
rect 7610 139840 7930 140864
rect 7610 139776 7618 139840
rect 7682 139776 7698 139840
rect 7762 139776 7778 139840
rect 7842 139776 7858 139840
rect 7922 139776 7930 139840
rect 7610 138752 7930 139776
rect 7610 138688 7618 138752
rect 7682 138688 7698 138752
rect 7762 138688 7778 138752
rect 7842 138688 7858 138752
rect 7922 138688 7930 138752
rect 7610 137664 7930 138688
rect 7610 137600 7618 137664
rect 7682 137600 7698 137664
rect 7762 137600 7778 137664
rect 7842 137600 7858 137664
rect 7922 137600 7930 137664
rect 7610 136576 7930 137600
rect 7610 136512 7618 136576
rect 7682 136512 7698 136576
rect 7762 136512 7778 136576
rect 7842 136512 7858 136576
rect 7922 136512 7930 136576
rect 7610 135488 7930 136512
rect 7610 135424 7618 135488
rect 7682 135424 7698 135488
rect 7762 135424 7778 135488
rect 7842 135424 7858 135488
rect 7922 135424 7930 135488
rect 7610 134400 7930 135424
rect 7610 134336 7618 134400
rect 7682 134336 7698 134400
rect 7762 134336 7778 134400
rect 7842 134336 7858 134400
rect 7922 134336 7930 134400
rect 7610 133312 7930 134336
rect 7610 133248 7618 133312
rect 7682 133248 7698 133312
rect 7762 133248 7778 133312
rect 7842 133248 7858 133312
rect 7922 133248 7930 133312
rect 7610 132224 7930 133248
rect 7610 132160 7618 132224
rect 7682 132160 7698 132224
rect 7762 132160 7778 132224
rect 7842 132160 7858 132224
rect 7922 132160 7930 132224
rect 7610 131136 7930 132160
rect 7610 131072 7618 131136
rect 7682 131072 7698 131136
rect 7762 131072 7778 131136
rect 7842 131072 7858 131136
rect 7922 131072 7930 131136
rect 7610 130048 7930 131072
rect 7610 129984 7618 130048
rect 7682 129984 7698 130048
rect 7762 129984 7778 130048
rect 7842 129984 7858 130048
rect 7922 129984 7930 130048
rect 7610 128960 7930 129984
rect 7610 128896 7618 128960
rect 7682 128896 7698 128960
rect 7762 128896 7778 128960
rect 7842 128896 7858 128960
rect 7922 128896 7930 128960
rect 7610 127872 7930 128896
rect 7610 127808 7618 127872
rect 7682 127808 7698 127872
rect 7762 127808 7778 127872
rect 7842 127808 7858 127872
rect 7922 127808 7930 127872
rect 7610 126784 7930 127808
rect 7610 126720 7618 126784
rect 7682 126720 7698 126784
rect 7762 126720 7778 126784
rect 7842 126720 7858 126784
rect 7922 126720 7930 126784
rect 7610 125696 7930 126720
rect 7610 125632 7618 125696
rect 7682 125632 7698 125696
rect 7762 125632 7778 125696
rect 7842 125632 7858 125696
rect 7922 125632 7930 125696
rect 7610 124608 7930 125632
rect 7610 124544 7618 124608
rect 7682 124544 7698 124608
rect 7762 124544 7778 124608
rect 7842 124544 7858 124608
rect 7922 124544 7930 124608
rect 7610 123520 7930 124544
rect 7610 123456 7618 123520
rect 7682 123456 7698 123520
rect 7762 123456 7778 123520
rect 7842 123456 7858 123520
rect 7922 123456 7930 123520
rect 7610 122432 7930 123456
rect 7610 122368 7618 122432
rect 7682 122368 7698 122432
rect 7762 122368 7778 122432
rect 7842 122368 7858 122432
rect 7922 122368 7930 122432
rect 7610 121344 7930 122368
rect 7610 121280 7618 121344
rect 7682 121280 7698 121344
rect 7762 121280 7778 121344
rect 7842 121280 7858 121344
rect 7922 121280 7930 121344
rect 7610 120256 7930 121280
rect 7610 120192 7618 120256
rect 7682 120192 7698 120256
rect 7762 120192 7778 120256
rect 7842 120192 7858 120256
rect 7922 120192 7930 120256
rect 7610 119168 7930 120192
rect 7610 119104 7618 119168
rect 7682 119104 7698 119168
rect 7762 119104 7778 119168
rect 7842 119104 7858 119168
rect 7922 119104 7930 119168
rect 7610 118080 7930 119104
rect 7610 118016 7618 118080
rect 7682 118016 7698 118080
rect 7762 118016 7778 118080
rect 7842 118016 7858 118080
rect 7922 118016 7930 118080
rect 7610 116992 7930 118016
rect 7610 116928 7618 116992
rect 7682 116928 7698 116992
rect 7762 116928 7778 116992
rect 7842 116928 7858 116992
rect 7922 116928 7930 116992
rect 7610 115904 7930 116928
rect 7610 115840 7618 115904
rect 7682 115840 7698 115904
rect 7762 115840 7778 115904
rect 7842 115840 7858 115904
rect 7922 115840 7930 115904
rect 7610 114816 7930 115840
rect 7610 114752 7618 114816
rect 7682 114752 7698 114816
rect 7762 114752 7778 114816
rect 7842 114752 7858 114816
rect 7922 114752 7930 114816
rect 7610 113728 7930 114752
rect 7610 113664 7618 113728
rect 7682 113664 7698 113728
rect 7762 113664 7778 113728
rect 7842 113664 7858 113728
rect 7922 113664 7930 113728
rect 7610 112640 7930 113664
rect 7610 112576 7618 112640
rect 7682 112576 7698 112640
rect 7762 112576 7778 112640
rect 7842 112576 7858 112640
rect 7922 112576 7930 112640
rect 7610 111552 7930 112576
rect 7610 111488 7618 111552
rect 7682 111488 7698 111552
rect 7762 111488 7778 111552
rect 7842 111488 7858 111552
rect 7922 111488 7930 111552
rect 7610 110464 7930 111488
rect 7610 110400 7618 110464
rect 7682 110400 7698 110464
rect 7762 110400 7778 110464
rect 7842 110400 7858 110464
rect 7922 110400 7930 110464
rect 7610 109376 7930 110400
rect 7610 109312 7618 109376
rect 7682 109312 7698 109376
rect 7762 109312 7778 109376
rect 7842 109312 7858 109376
rect 7922 109312 7930 109376
rect 7610 108288 7930 109312
rect 7610 108224 7618 108288
rect 7682 108224 7698 108288
rect 7762 108224 7778 108288
rect 7842 108224 7858 108288
rect 7922 108224 7930 108288
rect 7610 107200 7930 108224
rect 7610 107136 7618 107200
rect 7682 107136 7698 107200
rect 7762 107136 7778 107200
rect 7842 107136 7858 107200
rect 7922 107136 7930 107200
rect 7610 106112 7930 107136
rect 7610 106048 7618 106112
rect 7682 106048 7698 106112
rect 7762 106048 7778 106112
rect 7842 106048 7858 106112
rect 7922 106048 7930 106112
rect 7610 105024 7930 106048
rect 7610 104960 7618 105024
rect 7682 104960 7698 105024
rect 7762 104960 7778 105024
rect 7842 104960 7858 105024
rect 7922 104960 7930 105024
rect 7610 103936 7930 104960
rect 7610 103872 7618 103936
rect 7682 103872 7698 103936
rect 7762 103872 7778 103936
rect 7842 103872 7858 103936
rect 7922 103872 7930 103936
rect 7610 102848 7930 103872
rect 7610 102784 7618 102848
rect 7682 102784 7698 102848
rect 7762 102784 7778 102848
rect 7842 102784 7858 102848
rect 7922 102784 7930 102848
rect 7610 101760 7930 102784
rect 7610 101696 7618 101760
rect 7682 101696 7698 101760
rect 7762 101696 7778 101760
rect 7842 101696 7858 101760
rect 7922 101696 7930 101760
rect 7610 100672 7930 101696
rect 7610 100608 7618 100672
rect 7682 100608 7698 100672
rect 7762 100608 7778 100672
rect 7842 100608 7858 100672
rect 7922 100608 7930 100672
rect 7610 99584 7930 100608
rect 7610 99520 7618 99584
rect 7682 99520 7698 99584
rect 7762 99520 7778 99584
rect 7842 99520 7858 99584
rect 7922 99520 7930 99584
rect 7610 98496 7930 99520
rect 7610 98432 7618 98496
rect 7682 98432 7698 98496
rect 7762 98432 7778 98496
rect 7842 98432 7858 98496
rect 7922 98432 7930 98496
rect 7610 97408 7930 98432
rect 7610 97344 7618 97408
rect 7682 97344 7698 97408
rect 7762 97344 7778 97408
rect 7842 97344 7858 97408
rect 7922 97344 7930 97408
rect 7610 96320 7930 97344
rect 7610 96256 7618 96320
rect 7682 96256 7698 96320
rect 7762 96256 7778 96320
rect 7842 96256 7858 96320
rect 7922 96256 7930 96320
rect 7610 95232 7930 96256
rect 7610 95168 7618 95232
rect 7682 95168 7698 95232
rect 7762 95168 7778 95232
rect 7842 95168 7858 95232
rect 7922 95168 7930 95232
rect 7610 94144 7930 95168
rect 7610 94080 7618 94144
rect 7682 94080 7698 94144
rect 7762 94080 7778 94144
rect 7842 94080 7858 94144
rect 7922 94080 7930 94144
rect 7610 93056 7930 94080
rect 7610 92992 7618 93056
rect 7682 92992 7698 93056
rect 7762 92992 7778 93056
rect 7842 92992 7858 93056
rect 7922 92992 7930 93056
rect 7610 91968 7930 92992
rect 7610 91904 7618 91968
rect 7682 91904 7698 91968
rect 7762 91904 7778 91968
rect 7842 91904 7858 91968
rect 7922 91904 7930 91968
rect 7610 90880 7930 91904
rect 7610 90816 7618 90880
rect 7682 90816 7698 90880
rect 7762 90816 7778 90880
rect 7842 90816 7858 90880
rect 7922 90816 7930 90880
rect 7610 89792 7930 90816
rect 7610 89728 7618 89792
rect 7682 89728 7698 89792
rect 7762 89728 7778 89792
rect 7842 89728 7858 89792
rect 7922 89728 7930 89792
rect 7610 88704 7930 89728
rect 7610 88640 7618 88704
rect 7682 88640 7698 88704
rect 7762 88640 7778 88704
rect 7842 88640 7858 88704
rect 7922 88640 7930 88704
rect 7610 87616 7930 88640
rect 7610 87552 7618 87616
rect 7682 87552 7698 87616
rect 7762 87552 7778 87616
rect 7842 87552 7858 87616
rect 7922 87552 7930 87616
rect 7610 86528 7930 87552
rect 7610 86464 7618 86528
rect 7682 86464 7698 86528
rect 7762 86464 7778 86528
rect 7842 86464 7858 86528
rect 7922 86464 7930 86528
rect 7610 85440 7930 86464
rect 7610 85376 7618 85440
rect 7682 85376 7698 85440
rect 7762 85376 7778 85440
rect 7842 85376 7858 85440
rect 7922 85376 7930 85440
rect 7610 84352 7930 85376
rect 7610 84288 7618 84352
rect 7682 84288 7698 84352
rect 7762 84288 7778 84352
rect 7842 84288 7858 84352
rect 7922 84288 7930 84352
rect 7610 83264 7930 84288
rect 7610 83200 7618 83264
rect 7682 83200 7698 83264
rect 7762 83200 7778 83264
rect 7842 83200 7858 83264
rect 7922 83200 7930 83264
rect 7610 82176 7930 83200
rect 7610 82112 7618 82176
rect 7682 82112 7698 82176
rect 7762 82112 7778 82176
rect 7842 82112 7858 82176
rect 7922 82112 7930 82176
rect 7610 81088 7930 82112
rect 7610 81024 7618 81088
rect 7682 81024 7698 81088
rect 7762 81024 7778 81088
rect 7842 81024 7858 81088
rect 7922 81024 7930 81088
rect 7610 80000 7930 81024
rect 7610 79936 7618 80000
rect 7682 79936 7698 80000
rect 7762 79936 7778 80000
rect 7842 79936 7858 80000
rect 7922 79936 7930 80000
rect 7610 78912 7930 79936
rect 7610 78848 7618 78912
rect 7682 78848 7698 78912
rect 7762 78848 7778 78912
rect 7842 78848 7858 78912
rect 7922 78848 7930 78912
rect 7610 77824 7930 78848
rect 7610 77760 7618 77824
rect 7682 77760 7698 77824
rect 7762 77760 7778 77824
rect 7842 77760 7858 77824
rect 7922 77760 7930 77824
rect 7610 76736 7930 77760
rect 7610 76672 7618 76736
rect 7682 76672 7698 76736
rect 7762 76672 7778 76736
rect 7842 76672 7858 76736
rect 7922 76672 7930 76736
rect 7610 75648 7930 76672
rect 7610 75584 7618 75648
rect 7682 75584 7698 75648
rect 7762 75584 7778 75648
rect 7842 75584 7858 75648
rect 7922 75584 7930 75648
rect 7610 74560 7930 75584
rect 7610 74496 7618 74560
rect 7682 74496 7698 74560
rect 7762 74496 7778 74560
rect 7842 74496 7858 74560
rect 7922 74496 7930 74560
rect 7610 73472 7930 74496
rect 7610 73408 7618 73472
rect 7682 73408 7698 73472
rect 7762 73408 7778 73472
rect 7842 73408 7858 73472
rect 7922 73408 7930 73472
rect 7610 72384 7930 73408
rect 7610 72320 7618 72384
rect 7682 72320 7698 72384
rect 7762 72320 7778 72384
rect 7842 72320 7858 72384
rect 7922 72320 7930 72384
rect 7610 71296 7930 72320
rect 7610 71232 7618 71296
rect 7682 71232 7698 71296
rect 7762 71232 7778 71296
rect 7842 71232 7858 71296
rect 7922 71232 7930 71296
rect 7610 70208 7930 71232
rect 7610 70144 7618 70208
rect 7682 70144 7698 70208
rect 7762 70144 7778 70208
rect 7842 70144 7858 70208
rect 7922 70144 7930 70208
rect 7610 69120 7930 70144
rect 7610 69056 7618 69120
rect 7682 69056 7698 69120
rect 7762 69056 7778 69120
rect 7842 69056 7858 69120
rect 7922 69056 7930 69120
rect 7610 68032 7930 69056
rect 7610 67968 7618 68032
rect 7682 67968 7698 68032
rect 7762 67968 7778 68032
rect 7842 67968 7858 68032
rect 7922 67968 7930 68032
rect 7610 66944 7930 67968
rect 7610 66880 7618 66944
rect 7682 66880 7698 66944
rect 7762 66880 7778 66944
rect 7842 66880 7858 66944
rect 7922 66880 7930 66944
rect 7610 65856 7930 66880
rect 7610 65792 7618 65856
rect 7682 65792 7698 65856
rect 7762 65792 7778 65856
rect 7842 65792 7858 65856
rect 7922 65792 7930 65856
rect 7610 64768 7930 65792
rect 7610 64704 7618 64768
rect 7682 64704 7698 64768
rect 7762 64704 7778 64768
rect 7842 64704 7858 64768
rect 7922 64704 7930 64768
rect 7610 63680 7930 64704
rect 7610 63616 7618 63680
rect 7682 63616 7698 63680
rect 7762 63616 7778 63680
rect 7842 63616 7858 63680
rect 7922 63616 7930 63680
rect 7610 62592 7930 63616
rect 7610 62528 7618 62592
rect 7682 62528 7698 62592
rect 7762 62528 7778 62592
rect 7842 62528 7858 62592
rect 7922 62528 7930 62592
rect 7610 61504 7930 62528
rect 7610 61440 7618 61504
rect 7682 61440 7698 61504
rect 7762 61440 7778 61504
rect 7842 61440 7858 61504
rect 7922 61440 7930 61504
rect 7610 60416 7930 61440
rect 7610 60352 7618 60416
rect 7682 60352 7698 60416
rect 7762 60352 7778 60416
rect 7842 60352 7858 60416
rect 7922 60352 7930 60416
rect 7610 59328 7930 60352
rect 7610 59264 7618 59328
rect 7682 59264 7698 59328
rect 7762 59264 7778 59328
rect 7842 59264 7858 59328
rect 7922 59264 7930 59328
rect 7610 58240 7930 59264
rect 7610 58176 7618 58240
rect 7682 58176 7698 58240
rect 7762 58176 7778 58240
rect 7842 58176 7858 58240
rect 7922 58176 7930 58240
rect 7610 57152 7930 58176
rect 7610 57088 7618 57152
rect 7682 57088 7698 57152
rect 7762 57088 7778 57152
rect 7842 57088 7858 57152
rect 7922 57088 7930 57152
rect 7610 56064 7930 57088
rect 7610 56000 7618 56064
rect 7682 56000 7698 56064
rect 7762 56000 7778 56064
rect 7842 56000 7858 56064
rect 7922 56000 7930 56064
rect 7610 54976 7930 56000
rect 7610 54912 7618 54976
rect 7682 54912 7698 54976
rect 7762 54912 7778 54976
rect 7842 54912 7858 54976
rect 7922 54912 7930 54976
rect 7610 53888 7930 54912
rect 7610 53824 7618 53888
rect 7682 53824 7698 53888
rect 7762 53824 7778 53888
rect 7842 53824 7858 53888
rect 7922 53824 7930 53888
rect 7610 52800 7930 53824
rect 7610 52736 7618 52800
rect 7682 52736 7698 52800
rect 7762 52736 7778 52800
rect 7842 52736 7858 52800
rect 7922 52736 7930 52800
rect 7610 51712 7930 52736
rect 7610 51648 7618 51712
rect 7682 51648 7698 51712
rect 7762 51648 7778 51712
rect 7842 51648 7858 51712
rect 7922 51648 7930 51712
rect 7610 50624 7930 51648
rect 7610 50560 7618 50624
rect 7682 50560 7698 50624
rect 7762 50560 7778 50624
rect 7842 50560 7858 50624
rect 7922 50560 7930 50624
rect 7610 49536 7930 50560
rect 7610 49472 7618 49536
rect 7682 49472 7698 49536
rect 7762 49472 7778 49536
rect 7842 49472 7858 49536
rect 7922 49472 7930 49536
rect 7610 48448 7930 49472
rect 7610 48384 7618 48448
rect 7682 48384 7698 48448
rect 7762 48384 7778 48448
rect 7842 48384 7858 48448
rect 7922 48384 7930 48448
rect 7610 47360 7930 48384
rect 7610 47296 7618 47360
rect 7682 47296 7698 47360
rect 7762 47296 7778 47360
rect 7842 47296 7858 47360
rect 7922 47296 7930 47360
rect 7610 46272 7930 47296
rect 7610 46208 7618 46272
rect 7682 46208 7698 46272
rect 7762 46208 7778 46272
rect 7842 46208 7858 46272
rect 7922 46208 7930 46272
rect 7610 45184 7930 46208
rect 7610 45120 7618 45184
rect 7682 45120 7698 45184
rect 7762 45120 7778 45184
rect 7842 45120 7858 45184
rect 7922 45120 7930 45184
rect 7610 44096 7930 45120
rect 7610 44032 7618 44096
rect 7682 44032 7698 44096
rect 7762 44032 7778 44096
rect 7842 44032 7858 44096
rect 7922 44032 7930 44096
rect 7610 43008 7930 44032
rect 7610 42944 7618 43008
rect 7682 42944 7698 43008
rect 7762 42944 7778 43008
rect 7842 42944 7858 43008
rect 7922 42944 7930 43008
rect 7610 41920 7930 42944
rect 7610 41856 7618 41920
rect 7682 41856 7698 41920
rect 7762 41856 7778 41920
rect 7842 41856 7858 41920
rect 7922 41856 7930 41920
rect 7610 40832 7930 41856
rect 7610 40768 7618 40832
rect 7682 40768 7698 40832
rect 7762 40768 7778 40832
rect 7842 40768 7858 40832
rect 7922 40768 7930 40832
rect 7610 39744 7930 40768
rect 7610 39680 7618 39744
rect 7682 39680 7698 39744
rect 7762 39680 7778 39744
rect 7842 39680 7858 39744
rect 7922 39680 7930 39744
rect 7610 38656 7930 39680
rect 7610 38592 7618 38656
rect 7682 38592 7698 38656
rect 7762 38592 7778 38656
rect 7842 38592 7858 38656
rect 7922 38592 7930 38656
rect 7610 37568 7930 38592
rect 7610 37504 7618 37568
rect 7682 37504 7698 37568
rect 7762 37504 7778 37568
rect 7842 37504 7858 37568
rect 7922 37504 7930 37568
rect 7610 36480 7930 37504
rect 7610 36416 7618 36480
rect 7682 36416 7698 36480
rect 7762 36416 7778 36480
rect 7842 36416 7858 36480
rect 7922 36416 7930 36480
rect 7610 35392 7930 36416
rect 7610 35328 7618 35392
rect 7682 35328 7698 35392
rect 7762 35328 7778 35392
rect 7842 35328 7858 35392
rect 7922 35328 7930 35392
rect 7610 34304 7930 35328
rect 7610 34240 7618 34304
rect 7682 34240 7698 34304
rect 7762 34240 7778 34304
rect 7842 34240 7858 34304
rect 7922 34240 7930 34304
rect 7610 33216 7930 34240
rect 7610 33152 7618 33216
rect 7682 33152 7698 33216
rect 7762 33152 7778 33216
rect 7842 33152 7858 33216
rect 7922 33152 7930 33216
rect 7610 32128 7930 33152
rect 7610 32064 7618 32128
rect 7682 32064 7698 32128
rect 7762 32064 7778 32128
rect 7842 32064 7858 32128
rect 7922 32064 7930 32128
rect 7610 31040 7930 32064
rect 7610 30976 7618 31040
rect 7682 30976 7698 31040
rect 7762 30976 7778 31040
rect 7842 30976 7858 31040
rect 7922 30976 7930 31040
rect 7610 29952 7930 30976
rect 7610 29888 7618 29952
rect 7682 29888 7698 29952
rect 7762 29888 7778 29952
rect 7842 29888 7858 29952
rect 7922 29888 7930 29952
rect 7610 28864 7930 29888
rect 7610 28800 7618 28864
rect 7682 28800 7698 28864
rect 7762 28800 7778 28864
rect 7842 28800 7858 28864
rect 7922 28800 7930 28864
rect 7610 27776 7930 28800
rect 7610 27712 7618 27776
rect 7682 27712 7698 27776
rect 7762 27712 7778 27776
rect 7842 27712 7858 27776
rect 7922 27712 7930 27776
rect 7610 26688 7930 27712
rect 7610 26624 7618 26688
rect 7682 26624 7698 26688
rect 7762 26624 7778 26688
rect 7842 26624 7858 26688
rect 7922 26624 7930 26688
rect 7610 25600 7930 26624
rect 7610 25536 7618 25600
rect 7682 25536 7698 25600
rect 7762 25536 7778 25600
rect 7842 25536 7858 25600
rect 7922 25536 7930 25600
rect 7610 24512 7930 25536
rect 7610 24448 7618 24512
rect 7682 24448 7698 24512
rect 7762 24448 7778 24512
rect 7842 24448 7858 24512
rect 7922 24448 7930 24512
rect 7610 23424 7930 24448
rect 7610 23360 7618 23424
rect 7682 23360 7698 23424
rect 7762 23360 7778 23424
rect 7842 23360 7858 23424
rect 7922 23360 7930 23424
rect 7610 22336 7930 23360
rect 7610 22272 7618 22336
rect 7682 22272 7698 22336
rect 7762 22272 7778 22336
rect 7842 22272 7858 22336
rect 7922 22272 7930 22336
rect 7610 21248 7930 22272
rect 7610 21184 7618 21248
rect 7682 21184 7698 21248
rect 7762 21184 7778 21248
rect 7842 21184 7858 21248
rect 7922 21184 7930 21248
rect 7610 20160 7930 21184
rect 7610 20096 7618 20160
rect 7682 20096 7698 20160
rect 7762 20096 7778 20160
rect 7842 20096 7858 20160
rect 7922 20096 7930 20160
rect 7610 19072 7930 20096
rect 7610 19008 7618 19072
rect 7682 19008 7698 19072
rect 7762 19008 7778 19072
rect 7842 19008 7858 19072
rect 7922 19008 7930 19072
rect 7610 17984 7930 19008
rect 7610 17920 7618 17984
rect 7682 17920 7698 17984
rect 7762 17920 7778 17984
rect 7842 17920 7858 17984
rect 7922 17920 7930 17984
rect 7610 16896 7930 17920
rect 7610 16832 7618 16896
rect 7682 16832 7698 16896
rect 7762 16832 7778 16896
rect 7842 16832 7858 16896
rect 7922 16832 7930 16896
rect 7610 15808 7930 16832
rect 7610 15744 7618 15808
rect 7682 15744 7698 15808
rect 7762 15744 7778 15808
rect 7842 15744 7858 15808
rect 7922 15744 7930 15808
rect 7610 14720 7930 15744
rect 7610 14656 7618 14720
rect 7682 14656 7698 14720
rect 7762 14656 7778 14720
rect 7842 14656 7858 14720
rect 7922 14656 7930 14720
rect 7610 13632 7930 14656
rect 7610 13568 7618 13632
rect 7682 13568 7698 13632
rect 7762 13568 7778 13632
rect 7842 13568 7858 13632
rect 7922 13568 7930 13632
rect 7610 12544 7930 13568
rect 7610 12480 7618 12544
rect 7682 12480 7698 12544
rect 7762 12480 7778 12544
rect 7842 12480 7858 12544
rect 7922 12480 7930 12544
rect 7610 11456 7930 12480
rect 7610 11392 7618 11456
rect 7682 11392 7698 11456
rect 7762 11392 7778 11456
rect 7842 11392 7858 11456
rect 7922 11392 7930 11456
rect 7610 10368 7930 11392
rect 7610 10304 7618 10368
rect 7682 10304 7698 10368
rect 7762 10304 7778 10368
rect 7842 10304 7858 10368
rect 7922 10304 7930 10368
rect 7610 9280 7930 10304
rect 7610 9216 7618 9280
rect 7682 9216 7698 9280
rect 7762 9216 7778 9280
rect 7842 9216 7858 9280
rect 7922 9216 7930 9280
rect 7610 8192 7930 9216
rect 7610 8128 7618 8192
rect 7682 8128 7698 8192
rect 7762 8128 7778 8192
rect 7842 8128 7858 8192
rect 7922 8128 7930 8192
rect 7610 7104 7930 8128
rect 7610 7040 7618 7104
rect 7682 7040 7698 7104
rect 7762 7040 7778 7104
rect 7842 7040 7858 7104
rect 7922 7040 7930 7104
rect 7610 6016 7930 7040
rect 7610 5952 7618 6016
rect 7682 5952 7698 6016
rect 7762 5952 7778 6016
rect 7842 5952 7858 6016
rect 7922 5952 7930 6016
rect 7610 4928 7930 5952
rect 7610 4864 7618 4928
rect 7682 4864 7698 4928
rect 7762 4864 7778 4928
rect 7842 4864 7858 4928
rect 7922 4864 7930 4928
rect 7610 3840 7930 4864
rect 7610 3776 7618 3840
rect 7682 3776 7698 3840
rect 7762 3776 7778 3840
rect 7842 3776 7858 3840
rect 7922 3776 7930 3840
rect 7610 2752 7930 3776
rect 7610 2688 7618 2752
rect 7682 2688 7698 2752
rect 7762 2688 7778 2752
rect 7842 2688 7858 2752
rect 7922 2688 7930 2752
rect 7610 2128 7930 2688
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1208 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_39
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_51 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1209
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_1210
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_59 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 8832 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 8832 0 1 2720
box -38 -48 314 592
use scs8hd_decap_6  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_6  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_1_80 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8464 0 1 2720
box -38 -48 130 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1211
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 8832 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_1  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1212
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 8832 0 1 3808
box -38 -48 314 592
use scs8hd_decap_6  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_3_80
timestamp 1586364061
transform 1 0 8464 0 1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1213
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 8832 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1214
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_59
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 8832 0 1 4896
box -38 -48 314 592
use scs8hd_decap_6  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_5_80
timestamp 1586364061
transform 1 0 8464 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1215
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1216
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 8832 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 8832 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_6  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_7_80
timestamp 1586364061
transform 1 0 8464 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1217
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 8832 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_80
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_39
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_51
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1218
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_59
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 8832 0 1 7072
box -38 -48 314 592
use scs8hd_decap_6  FILLER_9_74
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_9_80
timestamp 1586364061
transform 1 0 8464 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1219
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_56
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_68
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 8832 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_80
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_27
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_39
timestamp 1586364061
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_51
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1220
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_59
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 8832 0 1 8160
box -38 -48 314 592
use scs8hd_decap_6  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_11_80
timestamp 1586364061
transform 1 0 8464 0 1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1221
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 8832 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1223
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_39
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_51
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1222
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_59
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_68
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 8832 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 8832 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_6  FILLER_13_74
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_13_80
timestamp 1586364061
transform 1 0 8464 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1224
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_59
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 8832 0 1 10336
box -38 -48 314 592
use scs8hd_decap_6  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_15_80
timestamp 1586364061
transform 1 0 8464 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1225
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 8832 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_16_80
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1226
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 8832 0 1 11424
box -38 -48 314 592
use scs8hd_decap_6  FILLER_17_74
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_17_80
timestamp 1586364061
transform 1 0 8464 0 1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1227
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 8832 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_80
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1229
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_51
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1228
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_68
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 8832 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 8832 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_6  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_19_80
timestamp 1586364061
transform 1 0 8464 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_80
timestamp 1586364061
transform 1 0 8464 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_27
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_39
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_51
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1230
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_59
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 8832 0 1 13600
box -38 -48 314 592
use scs8hd_decap_6  FILLER_21_74
timestamp 1586364061
transform 1 0 7912 0 1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_21_80
timestamp 1586364061
transform 1 0 8464 0 1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1231
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_44
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_56
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_68
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 8832 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_1  FILLER_22_80
timestamp 1586364061
transform 1 0 8464 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_51
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1232
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_59
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 8832 0 1 14688
box -38 -48 314 592
use scs8hd_decap_6  FILLER_23_74
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_23_80
timestamp 1586364061
transform 1 0 8464 0 1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1233
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_44
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_56
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_68
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 8832 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_1  FILLER_24_80
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_39
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_51
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1234
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_59
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 8832 0 1 15776
box -38 -48 314 592
use scs8hd_decap_6  FILLER_25_74
timestamp 1586364061
transform 1 0 7912 0 1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_25_80
timestamp 1586364061
transform 1 0 8464 0 1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1235
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_27
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_44
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1236
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_56
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_59
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 8832 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 8832 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_26_80
timestamp 1586364061
transform 1 0 8464 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_27_80
timestamp 1586364061
transform 1 0 8464 0 1 16864
box -38 -48 130 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1237
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 8832 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_28_80
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_27
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_39
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_51
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1238
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 8832 0 1 17952
box -38 -48 314 592
use scs8hd_decap_6  FILLER_29_74
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_29_80
timestamp 1586364061
transform 1 0 8464 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1239
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 8832 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_1  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_39
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1240
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_59
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 8832 0 1 19040
box -38 -48 314 592
use scs8hd_decap_6  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_31_80
timestamp 1586364061
transform 1 0 8464 0 1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1241
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 8832 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1243
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_39
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_51
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1242
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 8832 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 8832 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_6  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_33_80
timestamp 1586364061
transform 1 0 8464 0 1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1244
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 8832 0 1 21216
box -38 -48 314 592
use scs8hd_decap_6  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_35_80
timestamp 1586364061
transform 1 0 8464 0 1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1245
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 8832 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_1  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_27
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_39
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_51
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1246
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 8832 0 1 22304
box -38 -48 314 592
use scs8hd_decap_6  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_37_80
timestamp 1586364061
transform 1 0 8464 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1247
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 8832 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_15
timestamp 1586364061
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1249
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_27
timestamp 1586364061
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_39
timestamp 1586364061
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_51
timestamp 1586364061
transform 1 0 5796 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1248
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 8832 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 8832 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_6  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_39_80
timestamp 1586364061
transform 1 0 8464 0 1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1250
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 8832 0 1 24480
box -38 -48 314 592
use scs8hd_decap_6  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 590 592
use scs8hd_fill_1  FILLER_41_80
timestamp 1586364061
transform 1 0 8464 0 1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1251
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_68
timestamp 1586364061
transform 1 0 7360 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 8832 0 -1 25568
box -38 -48 314 592
use scs8hd_fill_1  FILLER_42_80
timestamp 1586364061
transform 1 0 8464 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_3  PHY_86
timestamp 1586364061
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_43_3
timestamp 1586364061
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_15
timestamp 1586364061
transform 1 0 2484 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_27
timestamp 1586364061
transform 1 0 3588 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_39
timestamp 1586364061
transform 1 0 4692 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_43_51
timestamp 1586364061
transform 1 0 5796 0 1 25568
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1252
timestamp 1586364061
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_43_59
timestamp 1586364061
transform 1 0 6532 0 1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_43_62
timestamp 1586364061
transform 1 0 6808 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_87
timestamp 1586364061
transform -1 0 8832 0 1 25568
box -38 -48 314 592
use scs8hd_decap_6  FILLER_43_74
timestamp 1586364061
transform 1 0 7912 0 1 25568
box -38 -48 590 592
use scs8hd_fill_1  FILLER_43_80
timestamp 1586364061
transform 1 0 8464 0 1 25568
box -38 -48 130 592
use scs8hd_decap_3  PHY_88
timestamp 1586364061
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_44_3
timestamp 1586364061
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_15
timestamp 1586364061
transform 1 0 2484 0 -1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1253
timestamp 1586364061
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_4  FILLER_44_27
timestamp 1586364061
transform 1 0 3588 0 -1 26656
box -38 -48 406 592
use scs8hd_decap_12  FILLER_44_32
timestamp 1586364061
transform 1 0 4048 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_44
timestamp 1586364061
transform 1 0 5152 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_56
timestamp 1586364061
transform 1 0 6256 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_68
timestamp 1586364061
transform 1 0 7360 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_3  PHY_89
timestamp 1586364061
transform -1 0 8832 0 -1 26656
box -38 -48 314 592
use scs8hd_fill_1  FILLER_44_80
timestamp 1586364061
transform 1 0 8464 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_3  PHY_90
timestamp 1586364061
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_45_3
timestamp 1586364061
transform 1 0 1380 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_15
timestamp 1586364061
transform 1 0 2484 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_27
timestamp 1586364061
transform 1 0 3588 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_39
timestamp 1586364061
transform 1 0 4692 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_45_51
timestamp 1586364061
transform 1 0 5796 0 1 26656
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1254
timestamp 1586364061
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use scs8hd_fill_2  FILLER_45_59
timestamp 1586364061
transform 1 0 6532 0 1 26656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_45_62
timestamp 1586364061
transform 1 0 6808 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_3  PHY_91
timestamp 1586364061
transform -1 0 8832 0 1 26656
box -38 -48 314 592
use scs8hd_decap_6  FILLER_45_74
timestamp 1586364061
transform 1 0 7912 0 1 26656
box -38 -48 590 592
use scs8hd_fill_1  FILLER_45_80
timestamp 1586364061
transform 1 0 8464 0 1 26656
box -38 -48 130 592
use scs8hd_decap_3  PHY_92
timestamp 1586364061
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_94
timestamp 1586364061
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use scs8hd_decap_12  FILLER_46_3
timestamp 1586364061
transform 1 0 1380 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_15
timestamp 1586364061
transform 1 0 2484 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_3
timestamp 1586364061
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_15
timestamp 1586364061
transform 1 0 2484 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1255
timestamp 1586364061
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_46_27
timestamp 1586364061
transform 1 0 3588 0 -1 27744
box -38 -48 406 592
use scs8hd_decap_12  FILLER_46_32
timestamp 1586364061
transform 1 0 4048 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_27
timestamp 1586364061
transform 1 0 3588 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_44
timestamp 1586364061
transform 1 0 5152 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_39
timestamp 1586364061
transform 1 0 4692 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_47_51
timestamp 1586364061
transform 1 0 5796 0 1 27744
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1256
timestamp 1586364061
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_56
timestamp 1586364061
transform 1 0 6256 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_68
timestamp 1586364061
transform 1 0 7360 0 -1 27744
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_47_59
timestamp 1586364061
transform 1 0 6532 0 1 27744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_47_62
timestamp 1586364061
transform 1 0 6808 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_3  PHY_93
timestamp 1586364061
transform -1 0 8832 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_95
timestamp 1586364061
transform -1 0 8832 0 1 27744
box -38 -48 314 592
use scs8hd_fill_1  FILLER_46_80
timestamp 1586364061
transform 1 0 8464 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_6  FILLER_47_74
timestamp 1586364061
transform 1 0 7912 0 1 27744
box -38 -48 590 592
use scs8hd_fill_1  FILLER_47_80
timestamp 1586364061
transform 1 0 8464 0 1 27744
box -38 -48 130 592
use scs8hd_decap_3  PHY_96
timestamp 1586364061
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_48_3
timestamp 1586364061
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_15
timestamp 1586364061
transform 1 0 2484 0 -1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1257
timestamp 1586364061
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_4  FILLER_48_27
timestamp 1586364061
transform 1 0 3588 0 -1 28832
box -38 -48 406 592
use scs8hd_decap_12  FILLER_48_32
timestamp 1586364061
transform 1 0 4048 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_44
timestamp 1586364061
transform 1 0 5152 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_56
timestamp 1586364061
transform 1 0 6256 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_68
timestamp 1586364061
transform 1 0 7360 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_3  PHY_97
timestamp 1586364061
transform -1 0 8832 0 -1 28832
box -38 -48 314 592
use scs8hd_fill_1  FILLER_48_80
timestamp 1586364061
transform 1 0 8464 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_3  PHY_98
timestamp 1586364061
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_49_3
timestamp 1586364061
transform 1 0 1380 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_15
timestamp 1586364061
transform 1 0 2484 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_27
timestamp 1586364061
transform 1 0 3588 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_39
timestamp 1586364061
transform 1 0 4692 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_49_51
timestamp 1586364061
transform 1 0 5796 0 1 28832
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1258
timestamp 1586364061
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use scs8hd_fill_2  FILLER_49_59
timestamp 1586364061
transform 1 0 6532 0 1 28832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_49_62
timestamp 1586364061
transform 1 0 6808 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_3  PHY_99
timestamp 1586364061
transform -1 0 8832 0 1 28832
box -38 -48 314 592
use scs8hd_decap_6  FILLER_49_74
timestamp 1586364061
transform 1 0 7912 0 1 28832
box -38 -48 590 592
use scs8hd_fill_1  FILLER_49_80
timestamp 1586364061
transform 1 0 8464 0 1 28832
box -38 -48 130 592
use scs8hd_decap_3  PHY_100
timestamp 1586364061
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_50_3
timestamp 1586364061
transform 1 0 1380 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_15
timestamp 1586364061
transform 1 0 2484 0 -1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1259
timestamp 1586364061
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_4  FILLER_50_27
timestamp 1586364061
transform 1 0 3588 0 -1 29920
box -38 -48 406 592
use scs8hd_decap_12  FILLER_50_32
timestamp 1586364061
transform 1 0 4048 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_44
timestamp 1586364061
transform 1 0 5152 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_56
timestamp 1586364061
transform 1 0 6256 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_68
timestamp 1586364061
transform 1 0 7360 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_3  PHY_101
timestamp 1586364061
transform -1 0 8832 0 -1 29920
box -38 -48 314 592
use scs8hd_fill_1  FILLER_50_80
timestamp 1586364061
transform 1 0 8464 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_3  PHY_102
timestamp 1586364061
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_51_3
timestamp 1586364061
transform 1 0 1380 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_15
timestamp 1586364061
transform 1 0 2484 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_27
timestamp 1586364061
transform 1 0 3588 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_39
timestamp 1586364061
transform 1 0 4692 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_51_51
timestamp 1586364061
transform 1 0 5796 0 1 29920
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1260
timestamp 1586364061
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use scs8hd_fill_2  FILLER_51_59
timestamp 1586364061
transform 1 0 6532 0 1 29920
box -38 -48 222 592
use scs8hd_decap_12  FILLER_51_62
timestamp 1586364061
transform 1 0 6808 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_3  PHY_103
timestamp 1586364061
transform -1 0 8832 0 1 29920
box -38 -48 314 592
use scs8hd_decap_6  FILLER_51_74
timestamp 1586364061
transform 1 0 7912 0 1 29920
box -38 -48 590 592
use scs8hd_fill_1  FILLER_51_80
timestamp 1586364061
transform 1 0 8464 0 1 29920
box -38 -48 130 592
use scs8hd_decap_3  PHY_104
timestamp 1586364061
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_106
timestamp 1586364061
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use scs8hd_decap_12  FILLER_52_3
timestamp 1586364061
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_15
timestamp 1586364061
transform 1 0 2484 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_3
timestamp 1586364061
transform 1 0 1380 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_15
timestamp 1586364061
transform 1 0 2484 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1261
timestamp 1586364061
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_52_27
timestamp 1586364061
transform 1 0 3588 0 -1 31008
box -38 -48 406 592
use scs8hd_decap_12  FILLER_52_32
timestamp 1586364061
transform 1 0 4048 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_27
timestamp 1586364061
transform 1 0 3588 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_44
timestamp 1586364061
transform 1 0 5152 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_39
timestamp 1586364061
transform 1 0 4692 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_53_51
timestamp 1586364061
transform 1 0 5796 0 1 31008
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1262
timestamp 1586364061
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_56
timestamp 1586364061
transform 1 0 6256 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_68
timestamp 1586364061
transform 1 0 7360 0 -1 31008
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_53_59
timestamp 1586364061
transform 1 0 6532 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_53_62
timestamp 1586364061
transform 1 0 6808 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_3  PHY_105
timestamp 1586364061
transform -1 0 8832 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_107
timestamp 1586364061
transform -1 0 8832 0 1 31008
box -38 -48 314 592
use scs8hd_fill_1  FILLER_52_80
timestamp 1586364061
transform 1 0 8464 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_6  FILLER_53_74
timestamp 1586364061
transform 1 0 7912 0 1 31008
box -38 -48 590 592
use scs8hd_fill_1  FILLER_53_80
timestamp 1586364061
transform 1 0 8464 0 1 31008
box -38 -48 130 592
use scs8hd_decap_3  PHY_108
timestamp 1586364061
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_54_3
timestamp 1586364061
transform 1 0 1380 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_15
timestamp 1586364061
transform 1 0 2484 0 -1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1263
timestamp 1586364061
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_4  FILLER_54_27
timestamp 1586364061
transform 1 0 3588 0 -1 32096
box -38 -48 406 592
use scs8hd_decap_12  FILLER_54_32
timestamp 1586364061
transform 1 0 4048 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_44
timestamp 1586364061
transform 1 0 5152 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_56
timestamp 1586364061
transform 1 0 6256 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_68
timestamp 1586364061
transform 1 0 7360 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_3  PHY_109
timestamp 1586364061
transform -1 0 8832 0 -1 32096
box -38 -48 314 592
use scs8hd_fill_1  FILLER_54_80
timestamp 1586364061
transform 1 0 8464 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_3  PHY_110
timestamp 1586364061
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_55_3
timestamp 1586364061
transform 1 0 1380 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_15
timestamp 1586364061
transform 1 0 2484 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_27
timestamp 1586364061
transform 1 0 3588 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_39
timestamp 1586364061
transform 1 0 4692 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_55_51
timestamp 1586364061
transform 1 0 5796 0 1 32096
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1264
timestamp 1586364061
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use scs8hd_fill_2  FILLER_55_59
timestamp 1586364061
transform 1 0 6532 0 1 32096
box -38 -48 222 592
use scs8hd_decap_12  FILLER_55_62
timestamp 1586364061
transform 1 0 6808 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_3  PHY_111
timestamp 1586364061
transform -1 0 8832 0 1 32096
box -38 -48 314 592
use scs8hd_decap_6  FILLER_55_74
timestamp 1586364061
transform 1 0 7912 0 1 32096
box -38 -48 590 592
use scs8hd_fill_1  FILLER_55_80
timestamp 1586364061
transform 1 0 8464 0 1 32096
box -38 -48 130 592
use scs8hd_decap_3  PHY_112
timestamp 1586364061
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_56_3
timestamp 1586364061
transform 1 0 1380 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_15
timestamp 1586364061
transform 1 0 2484 0 -1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1265
timestamp 1586364061
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_4  FILLER_56_27
timestamp 1586364061
transform 1 0 3588 0 -1 33184
box -38 -48 406 592
use scs8hd_decap_12  FILLER_56_32
timestamp 1586364061
transform 1 0 4048 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_44
timestamp 1586364061
transform 1 0 5152 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_56
timestamp 1586364061
transform 1 0 6256 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_68
timestamp 1586364061
transform 1 0 7360 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_3  PHY_113
timestamp 1586364061
transform -1 0 8832 0 -1 33184
box -38 -48 314 592
use scs8hd_fill_1  FILLER_56_80
timestamp 1586364061
transform 1 0 8464 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_3  PHY_114
timestamp 1586364061
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_57_3
timestamp 1586364061
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_15
timestamp 1586364061
transform 1 0 2484 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_27
timestamp 1586364061
transform 1 0 3588 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_39
timestamp 1586364061
transform 1 0 4692 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_57_51
timestamp 1586364061
transform 1 0 5796 0 1 33184
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1266
timestamp 1586364061
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use scs8hd_fill_2  FILLER_57_59
timestamp 1586364061
transform 1 0 6532 0 1 33184
box -38 -48 222 592
use scs8hd_decap_12  FILLER_57_62
timestamp 1586364061
transform 1 0 6808 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_3  PHY_115
timestamp 1586364061
transform -1 0 8832 0 1 33184
box -38 -48 314 592
use scs8hd_decap_6  FILLER_57_74
timestamp 1586364061
transform 1 0 7912 0 1 33184
box -38 -48 590 592
use scs8hd_fill_1  FILLER_57_80
timestamp 1586364061
transform 1 0 8464 0 1 33184
box -38 -48 130 592
use scs8hd_decap_3  PHY_116
timestamp 1586364061
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_12  FILLER_58_3
timestamp 1586364061
transform 1 0 1380 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_15
timestamp 1586364061
transform 1 0 2484 0 -1 34272
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1267
timestamp 1586364061
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_4  FILLER_58_27
timestamp 1586364061
transform 1 0 3588 0 -1 34272
box -38 -48 406 592
use scs8hd_decap_12  FILLER_58_32
timestamp 1586364061
transform 1 0 4048 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_44
timestamp 1586364061
transform 1 0 5152 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_56
timestamp 1586364061
transform 1 0 6256 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_68
timestamp 1586364061
transform 1 0 7360 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_3  PHY_117
timestamp 1586364061
transform -1 0 8832 0 -1 34272
box -38 -48 314 592
use scs8hd_fill_1  FILLER_58_80
timestamp 1586364061
transform 1 0 8464 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_3  PHY_118
timestamp 1586364061
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_120
timestamp 1586364061
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_59_3
timestamp 1586364061
transform 1 0 1380 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_15
timestamp 1586364061
transform 1 0 2484 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_3
timestamp 1586364061
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_15
timestamp 1586364061
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1269
timestamp 1586364061
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_27
timestamp 1586364061
transform 1 0 3588 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_60_27
timestamp 1586364061
transform 1 0 3588 0 -1 35360
box -38 -48 406 592
use scs8hd_decap_12  FILLER_60_32
timestamp 1586364061
transform 1 0 4048 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_39
timestamp 1586364061
transform 1 0 4692 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_59_51
timestamp 1586364061
transform 1 0 5796 0 1 34272
box -38 -48 774 592
use scs8hd_decap_12  FILLER_60_44
timestamp 1586364061
transform 1 0 5152 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1268
timestamp 1586364061
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use scs8hd_fill_2  FILLER_59_59
timestamp 1586364061
transform 1 0 6532 0 1 34272
box -38 -48 222 592
use scs8hd_decap_12  FILLER_59_62
timestamp 1586364061
transform 1 0 6808 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_56
timestamp 1586364061
transform 1 0 6256 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_68
timestamp 1586364061
transform 1 0 7360 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_3  PHY_119
timestamp 1586364061
transform -1 0 8832 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_121
timestamp 1586364061
transform -1 0 8832 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_6  FILLER_59_74
timestamp 1586364061
transform 1 0 7912 0 1 34272
box -38 -48 590 592
use scs8hd_fill_1  FILLER_59_80
timestamp 1586364061
transform 1 0 8464 0 1 34272
box -38 -48 130 592
use scs8hd_fill_1  FILLER_60_80
timestamp 1586364061
transform 1 0 8464 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_3  PHY_122
timestamp 1586364061
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_61_3
timestamp 1586364061
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_15
timestamp 1586364061
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_27
timestamp 1586364061
transform 1 0 3588 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_39
timestamp 1586364061
transform 1 0 4692 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_61_51
timestamp 1586364061
transform 1 0 5796 0 1 35360
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1270
timestamp 1586364061
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use scs8hd_fill_2  FILLER_61_59
timestamp 1586364061
transform 1 0 6532 0 1 35360
box -38 -48 222 592
use scs8hd_decap_12  FILLER_61_62
timestamp 1586364061
transform 1 0 6808 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_3  PHY_123
timestamp 1586364061
transform -1 0 8832 0 1 35360
box -38 -48 314 592
use scs8hd_decap_6  FILLER_61_74
timestamp 1586364061
transform 1 0 7912 0 1 35360
box -38 -48 590 592
use scs8hd_fill_1  FILLER_61_80
timestamp 1586364061
transform 1 0 8464 0 1 35360
box -38 -48 130 592
use scs8hd_decap_3  PHY_124
timestamp 1586364061
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_62_3
timestamp 1586364061
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_15
timestamp 1586364061
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1271
timestamp 1586364061
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_4  FILLER_62_27
timestamp 1586364061
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use scs8hd_decap_12  FILLER_62_32
timestamp 1586364061
transform 1 0 4048 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_44
timestamp 1586364061
transform 1 0 5152 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_56
timestamp 1586364061
transform 1 0 6256 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_68
timestamp 1586364061
transform 1 0 7360 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_3  PHY_125
timestamp 1586364061
transform -1 0 8832 0 -1 36448
box -38 -48 314 592
use scs8hd_fill_1  FILLER_62_80
timestamp 1586364061
transform 1 0 8464 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_3  PHY_126
timestamp 1586364061
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_63_3
timestamp 1586364061
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_15
timestamp 1586364061
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_27
timestamp 1586364061
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_39
timestamp 1586364061
transform 1 0 4692 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_63_51
timestamp 1586364061
transform 1 0 5796 0 1 36448
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1272
timestamp 1586364061
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use scs8hd_fill_2  FILLER_63_59
timestamp 1586364061
transform 1 0 6532 0 1 36448
box -38 -48 222 592
use scs8hd_decap_12  FILLER_63_62
timestamp 1586364061
transform 1 0 6808 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_3  PHY_127
timestamp 1586364061
transform -1 0 8832 0 1 36448
box -38 -48 314 592
use scs8hd_decap_6  FILLER_63_74
timestamp 1586364061
transform 1 0 7912 0 1 36448
box -38 -48 590 592
use scs8hd_fill_1  FILLER_63_80
timestamp 1586364061
transform 1 0 8464 0 1 36448
box -38 -48 130 592
use scs8hd_decap_3  PHY_128
timestamp 1586364061
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use scs8hd_decap_12  FILLER_64_3
timestamp 1586364061
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_15
timestamp 1586364061
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1273
timestamp 1586364061
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_4  FILLER_64_27
timestamp 1586364061
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use scs8hd_decap_12  FILLER_64_32
timestamp 1586364061
transform 1 0 4048 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_44
timestamp 1586364061
transform 1 0 5152 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_56
timestamp 1586364061
transform 1 0 6256 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_68
timestamp 1586364061
transform 1 0 7360 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_3  PHY_129
timestamp 1586364061
transform -1 0 8832 0 -1 37536
box -38 -48 314 592
use scs8hd_fill_1  FILLER_64_80
timestamp 1586364061
transform 1 0 8464 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_3  PHY_130
timestamp 1586364061
transform 1 0 1104 0 1 37536
box -38 -48 314 592
use scs8hd_decap_12  FILLER_65_3
timestamp 1586364061
transform 1 0 1380 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_15
timestamp 1586364061
transform 1 0 2484 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_27
timestamp 1586364061
transform 1 0 3588 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_39
timestamp 1586364061
transform 1 0 4692 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_65_51
timestamp 1586364061
transform 1 0 5796 0 1 37536
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1274
timestamp 1586364061
transform 1 0 6716 0 1 37536
box -38 -48 130 592
use scs8hd_fill_2  FILLER_65_59
timestamp 1586364061
transform 1 0 6532 0 1 37536
box -38 -48 222 592
use scs8hd_decap_12  FILLER_65_62
timestamp 1586364061
transform 1 0 6808 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_3  PHY_131
timestamp 1586364061
transform -1 0 8832 0 1 37536
box -38 -48 314 592
use scs8hd_decap_6  FILLER_65_74
timestamp 1586364061
transform 1 0 7912 0 1 37536
box -38 -48 590 592
use scs8hd_fill_1  FILLER_65_80
timestamp 1586364061
transform 1 0 8464 0 1 37536
box -38 -48 130 592
use scs8hd_decap_3  PHY_132
timestamp 1586364061
transform 1 0 1104 0 -1 38624
box -38 -48 314 592
use scs8hd_decap_3  PHY_134
timestamp 1586364061
transform 1 0 1104 0 1 38624
box -38 -48 314 592
use scs8hd_decap_12  FILLER_66_3
timestamp 1586364061
transform 1 0 1380 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_15
timestamp 1586364061
transform 1 0 2484 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_3
timestamp 1586364061
transform 1 0 1380 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_15
timestamp 1586364061
transform 1 0 2484 0 1 38624
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1275
timestamp 1586364061
transform 1 0 3956 0 -1 38624
box -38 -48 130 592
use scs8hd_decap_4  FILLER_66_27
timestamp 1586364061
transform 1 0 3588 0 -1 38624
box -38 -48 406 592
use scs8hd_decap_12  FILLER_66_32
timestamp 1586364061
transform 1 0 4048 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_27
timestamp 1586364061
transform 1 0 3588 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_44
timestamp 1586364061
transform 1 0 5152 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_39
timestamp 1586364061
transform 1 0 4692 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_67_51
timestamp 1586364061
transform 1 0 5796 0 1 38624
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1276
timestamp 1586364061
transform 1 0 6716 0 1 38624
box -38 -48 130 592
use scs8hd_decap_12  FILLER_66_56
timestamp 1586364061
transform 1 0 6256 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_68
timestamp 1586364061
transform 1 0 7360 0 -1 38624
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_67_59
timestamp 1586364061
transform 1 0 6532 0 1 38624
box -38 -48 222 592
use scs8hd_decap_12  FILLER_67_62
timestamp 1586364061
transform 1 0 6808 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_3  PHY_133
timestamp 1586364061
transform -1 0 8832 0 -1 38624
box -38 -48 314 592
use scs8hd_decap_3  PHY_135
timestamp 1586364061
transform -1 0 8832 0 1 38624
box -38 -48 314 592
use scs8hd_fill_1  FILLER_66_80
timestamp 1586364061
transform 1 0 8464 0 -1 38624
box -38 -48 130 592
use scs8hd_decap_6  FILLER_67_74
timestamp 1586364061
transform 1 0 7912 0 1 38624
box -38 -48 590 592
use scs8hd_fill_1  FILLER_67_80
timestamp 1586364061
transform 1 0 8464 0 1 38624
box -38 -48 130 592
use scs8hd_decap_3  PHY_136
timestamp 1586364061
transform 1 0 1104 0 -1 39712
box -38 -48 314 592
use scs8hd_decap_12  FILLER_68_3
timestamp 1586364061
transform 1 0 1380 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_15
timestamp 1586364061
transform 1 0 2484 0 -1 39712
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1277
timestamp 1586364061
transform 1 0 3956 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_4  FILLER_68_27
timestamp 1586364061
transform 1 0 3588 0 -1 39712
box -38 -48 406 592
use scs8hd_decap_12  FILLER_68_32
timestamp 1586364061
transform 1 0 4048 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_44
timestamp 1586364061
transform 1 0 5152 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_56
timestamp 1586364061
transform 1 0 6256 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_68
timestamp 1586364061
transform 1 0 7360 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_3  PHY_137
timestamp 1586364061
transform -1 0 8832 0 -1 39712
box -38 -48 314 592
use scs8hd_fill_1  FILLER_68_80
timestamp 1586364061
transform 1 0 8464 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_3  PHY_138
timestamp 1586364061
transform 1 0 1104 0 1 39712
box -38 -48 314 592
use scs8hd_decap_12  FILLER_69_3
timestamp 1586364061
transform 1 0 1380 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_15
timestamp 1586364061
transform 1 0 2484 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_27
timestamp 1586364061
transform 1 0 3588 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_39
timestamp 1586364061
transform 1 0 4692 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_69_51
timestamp 1586364061
transform 1 0 5796 0 1 39712
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1278
timestamp 1586364061
transform 1 0 6716 0 1 39712
box -38 -48 130 592
use scs8hd_fill_2  FILLER_69_59
timestamp 1586364061
transform 1 0 6532 0 1 39712
box -38 -48 222 592
use scs8hd_decap_12  FILLER_69_62
timestamp 1586364061
transform 1 0 6808 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_3  PHY_139
timestamp 1586364061
transform -1 0 8832 0 1 39712
box -38 -48 314 592
use scs8hd_decap_6  FILLER_69_74
timestamp 1586364061
transform 1 0 7912 0 1 39712
box -38 -48 590 592
use scs8hd_fill_1  FILLER_69_80
timestamp 1586364061
transform 1 0 8464 0 1 39712
box -38 -48 130 592
use scs8hd_decap_3  PHY_140
timestamp 1586364061
transform 1 0 1104 0 -1 40800
box -38 -48 314 592
use scs8hd_decap_12  FILLER_70_3
timestamp 1586364061
transform 1 0 1380 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_15
timestamp 1586364061
transform 1 0 2484 0 -1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1279
timestamp 1586364061
transform 1 0 3956 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_4  FILLER_70_27
timestamp 1586364061
transform 1 0 3588 0 -1 40800
box -38 -48 406 592
use scs8hd_decap_12  FILLER_70_32
timestamp 1586364061
transform 1 0 4048 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_44
timestamp 1586364061
transform 1 0 5152 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_56
timestamp 1586364061
transform 1 0 6256 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_68
timestamp 1586364061
transform 1 0 7360 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_3  PHY_141
timestamp 1586364061
transform -1 0 8832 0 -1 40800
box -38 -48 314 592
use scs8hd_fill_1  FILLER_70_80
timestamp 1586364061
transform 1 0 8464 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_3  PHY_142
timestamp 1586364061
transform 1 0 1104 0 1 40800
box -38 -48 314 592
use scs8hd_decap_12  FILLER_71_3
timestamp 1586364061
transform 1 0 1380 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_15
timestamp 1586364061
transform 1 0 2484 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_27
timestamp 1586364061
transform 1 0 3588 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_39
timestamp 1586364061
transform 1 0 4692 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_71_51
timestamp 1586364061
transform 1 0 5796 0 1 40800
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1280
timestamp 1586364061
transform 1 0 6716 0 1 40800
box -38 -48 130 592
use scs8hd_fill_2  FILLER_71_59
timestamp 1586364061
transform 1 0 6532 0 1 40800
box -38 -48 222 592
use scs8hd_decap_12  FILLER_71_62
timestamp 1586364061
transform 1 0 6808 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_3  PHY_143
timestamp 1586364061
transform -1 0 8832 0 1 40800
box -38 -48 314 592
use scs8hd_decap_6  FILLER_71_74
timestamp 1586364061
transform 1 0 7912 0 1 40800
box -38 -48 590 592
use scs8hd_fill_1  FILLER_71_80
timestamp 1586364061
transform 1 0 8464 0 1 40800
box -38 -48 130 592
use scs8hd_decap_3  PHY_144
timestamp 1586364061
transform 1 0 1104 0 -1 41888
box -38 -48 314 592
use scs8hd_decap_3  PHY_146
timestamp 1586364061
transform 1 0 1104 0 1 41888
box -38 -48 314 592
use scs8hd_decap_12  FILLER_72_3
timestamp 1586364061
transform 1 0 1380 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_15
timestamp 1586364061
transform 1 0 2484 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_3
timestamp 1586364061
transform 1 0 1380 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_15
timestamp 1586364061
transform 1 0 2484 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1281
timestamp 1586364061
transform 1 0 3956 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_4  FILLER_72_27
timestamp 1586364061
transform 1 0 3588 0 -1 41888
box -38 -48 406 592
use scs8hd_decap_12  FILLER_72_32
timestamp 1586364061
transform 1 0 4048 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_27
timestamp 1586364061
transform 1 0 3588 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_44
timestamp 1586364061
transform 1 0 5152 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_39
timestamp 1586364061
transform 1 0 4692 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_73_51
timestamp 1586364061
transform 1 0 5796 0 1 41888
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1282
timestamp 1586364061
transform 1 0 6716 0 1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_56
timestamp 1586364061
transform 1 0 6256 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_68
timestamp 1586364061
transform 1 0 7360 0 -1 41888
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_73_59
timestamp 1586364061
transform 1 0 6532 0 1 41888
box -38 -48 222 592
use scs8hd_decap_12  FILLER_73_62
timestamp 1586364061
transform 1 0 6808 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_3  PHY_145
timestamp 1586364061
transform -1 0 8832 0 -1 41888
box -38 -48 314 592
use scs8hd_decap_3  PHY_147
timestamp 1586364061
transform -1 0 8832 0 1 41888
box -38 -48 314 592
use scs8hd_fill_1  FILLER_72_80
timestamp 1586364061
transform 1 0 8464 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_6  FILLER_73_74
timestamp 1586364061
transform 1 0 7912 0 1 41888
box -38 -48 590 592
use scs8hd_fill_1  FILLER_73_80
timestamp 1586364061
transform 1 0 8464 0 1 41888
box -38 -48 130 592
use scs8hd_decap_3  PHY_148
timestamp 1586364061
transform 1 0 1104 0 -1 42976
box -38 -48 314 592
use scs8hd_decap_12  FILLER_74_3
timestamp 1586364061
transform 1 0 1380 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_15
timestamp 1586364061
transform 1 0 2484 0 -1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1283
timestamp 1586364061
transform 1 0 3956 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_4  FILLER_74_27
timestamp 1586364061
transform 1 0 3588 0 -1 42976
box -38 -48 406 592
use scs8hd_decap_12  FILLER_74_32
timestamp 1586364061
transform 1 0 4048 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_44
timestamp 1586364061
transform 1 0 5152 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_56
timestamp 1586364061
transform 1 0 6256 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_68
timestamp 1586364061
transform 1 0 7360 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_3  PHY_149
timestamp 1586364061
transform -1 0 8832 0 -1 42976
box -38 -48 314 592
use scs8hd_fill_1  FILLER_74_80
timestamp 1586364061
transform 1 0 8464 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_3  PHY_150
timestamp 1586364061
transform 1 0 1104 0 1 42976
box -38 -48 314 592
use scs8hd_decap_12  FILLER_75_3
timestamp 1586364061
transform 1 0 1380 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_15
timestamp 1586364061
transform 1 0 2484 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_27
timestamp 1586364061
transform 1 0 3588 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_39
timestamp 1586364061
transform 1 0 4692 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_75_51
timestamp 1586364061
transform 1 0 5796 0 1 42976
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1284
timestamp 1586364061
transform 1 0 6716 0 1 42976
box -38 -48 130 592
use scs8hd_fill_2  FILLER_75_59
timestamp 1586364061
transform 1 0 6532 0 1 42976
box -38 -48 222 592
use scs8hd_decap_12  FILLER_75_62
timestamp 1586364061
transform 1 0 6808 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_3  PHY_151
timestamp 1586364061
transform -1 0 8832 0 1 42976
box -38 -48 314 592
use scs8hd_decap_6  FILLER_75_74
timestamp 1586364061
transform 1 0 7912 0 1 42976
box -38 -48 590 592
use scs8hd_fill_1  FILLER_75_80
timestamp 1586364061
transform 1 0 8464 0 1 42976
box -38 -48 130 592
use scs8hd_decap_3  PHY_152
timestamp 1586364061
transform 1 0 1104 0 -1 44064
box -38 -48 314 592
use scs8hd_decap_12  FILLER_76_3
timestamp 1586364061
transform 1 0 1380 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_15
timestamp 1586364061
transform 1 0 2484 0 -1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1285
timestamp 1586364061
transform 1 0 3956 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_4  FILLER_76_27
timestamp 1586364061
transform 1 0 3588 0 -1 44064
box -38 -48 406 592
use scs8hd_decap_12  FILLER_76_32
timestamp 1586364061
transform 1 0 4048 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_44
timestamp 1586364061
transform 1 0 5152 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_56
timestamp 1586364061
transform 1 0 6256 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_68
timestamp 1586364061
transform 1 0 7360 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_3  PHY_153
timestamp 1586364061
transform -1 0 8832 0 -1 44064
box -38 -48 314 592
use scs8hd_fill_1  FILLER_76_80
timestamp 1586364061
transform 1 0 8464 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_3  PHY_154
timestamp 1586364061
transform 1 0 1104 0 1 44064
box -38 -48 314 592
use scs8hd_decap_12  FILLER_77_3
timestamp 1586364061
transform 1 0 1380 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_15
timestamp 1586364061
transform 1 0 2484 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_27
timestamp 1586364061
transform 1 0 3588 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_39
timestamp 1586364061
transform 1 0 4692 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_77_51
timestamp 1586364061
transform 1 0 5796 0 1 44064
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1286
timestamp 1586364061
transform 1 0 6716 0 1 44064
box -38 -48 130 592
use scs8hd_fill_2  FILLER_77_59
timestamp 1586364061
transform 1 0 6532 0 1 44064
box -38 -48 222 592
use scs8hd_decap_12  FILLER_77_62
timestamp 1586364061
transform 1 0 6808 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_3  PHY_155
timestamp 1586364061
transform -1 0 8832 0 1 44064
box -38 -48 314 592
use scs8hd_decap_6  FILLER_77_74
timestamp 1586364061
transform 1 0 7912 0 1 44064
box -38 -48 590 592
use scs8hd_fill_1  FILLER_77_80
timestamp 1586364061
transform 1 0 8464 0 1 44064
box -38 -48 130 592
use scs8hd_decap_3  PHY_156
timestamp 1586364061
transform 1 0 1104 0 -1 45152
box -38 -48 314 592
use scs8hd_decap_12  FILLER_78_3
timestamp 1586364061
transform 1 0 1380 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_15
timestamp 1586364061
transform 1 0 2484 0 -1 45152
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1287
timestamp 1586364061
transform 1 0 3956 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_4  FILLER_78_27
timestamp 1586364061
transform 1 0 3588 0 -1 45152
box -38 -48 406 592
use scs8hd_decap_12  FILLER_78_32
timestamp 1586364061
transform 1 0 4048 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_44
timestamp 1586364061
transform 1 0 5152 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_56
timestamp 1586364061
transform 1 0 6256 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_68
timestamp 1586364061
transform 1 0 7360 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_3  PHY_157
timestamp 1586364061
transform -1 0 8832 0 -1 45152
box -38 -48 314 592
use scs8hd_fill_1  FILLER_78_80
timestamp 1586364061
transform 1 0 8464 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_3  PHY_158
timestamp 1586364061
transform 1 0 1104 0 1 45152
box -38 -48 314 592
use scs8hd_decap_3  PHY_160
timestamp 1586364061
transform 1 0 1104 0 -1 46240
box -38 -48 314 592
use scs8hd_decap_12  FILLER_79_3
timestamp 1586364061
transform 1 0 1380 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_15
timestamp 1586364061
transform 1 0 2484 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_3
timestamp 1586364061
transform 1 0 1380 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_15
timestamp 1586364061
transform 1 0 2484 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1289
timestamp 1586364061
transform 1 0 3956 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_27
timestamp 1586364061
transform 1 0 3588 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_80_27
timestamp 1586364061
transform 1 0 3588 0 -1 46240
box -38 -48 406 592
use scs8hd_decap_12  FILLER_80_32
timestamp 1586364061
transform 1 0 4048 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_39
timestamp 1586364061
transform 1 0 4692 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_79_51
timestamp 1586364061
transform 1 0 5796 0 1 45152
box -38 -48 774 592
use scs8hd_decap_12  FILLER_80_44
timestamp 1586364061
transform 1 0 5152 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1288
timestamp 1586364061
transform 1 0 6716 0 1 45152
box -38 -48 130 592
use scs8hd_fill_2  FILLER_79_59
timestamp 1586364061
transform 1 0 6532 0 1 45152
box -38 -48 222 592
use scs8hd_decap_12  FILLER_79_62
timestamp 1586364061
transform 1 0 6808 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_56
timestamp 1586364061
transform 1 0 6256 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_68
timestamp 1586364061
transform 1 0 7360 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_3  PHY_159
timestamp 1586364061
transform -1 0 8832 0 1 45152
box -38 -48 314 592
use scs8hd_decap_3  PHY_161
timestamp 1586364061
transform -1 0 8832 0 -1 46240
box -38 -48 314 592
use scs8hd_decap_6  FILLER_79_74
timestamp 1586364061
transform 1 0 7912 0 1 45152
box -38 -48 590 592
use scs8hd_fill_1  FILLER_79_80
timestamp 1586364061
transform 1 0 8464 0 1 45152
box -38 -48 130 592
use scs8hd_fill_1  FILLER_80_80
timestamp 1586364061
transform 1 0 8464 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_3  PHY_162
timestamp 1586364061
transform 1 0 1104 0 1 46240
box -38 -48 314 592
use scs8hd_decap_12  FILLER_81_3
timestamp 1586364061
transform 1 0 1380 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_15
timestamp 1586364061
transform 1 0 2484 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_27
timestamp 1586364061
transform 1 0 3588 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_39
timestamp 1586364061
transform 1 0 4692 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_81_51
timestamp 1586364061
transform 1 0 5796 0 1 46240
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1290
timestamp 1586364061
transform 1 0 6716 0 1 46240
box -38 -48 130 592
use scs8hd_fill_2  FILLER_81_59
timestamp 1586364061
transform 1 0 6532 0 1 46240
box -38 -48 222 592
use scs8hd_decap_12  FILLER_81_62
timestamp 1586364061
transform 1 0 6808 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_3  PHY_163
timestamp 1586364061
transform -1 0 8832 0 1 46240
box -38 -48 314 592
use scs8hd_decap_6  FILLER_81_74
timestamp 1586364061
transform 1 0 7912 0 1 46240
box -38 -48 590 592
use scs8hd_fill_1  FILLER_81_80
timestamp 1586364061
transform 1 0 8464 0 1 46240
box -38 -48 130 592
use scs8hd_decap_3  PHY_164
timestamp 1586364061
transform 1 0 1104 0 -1 47328
box -38 -48 314 592
use scs8hd_decap_12  FILLER_82_3
timestamp 1586364061
transform 1 0 1380 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_15
timestamp 1586364061
transform 1 0 2484 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1291
timestamp 1586364061
transform 1 0 3956 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_4  FILLER_82_27
timestamp 1586364061
transform 1 0 3588 0 -1 47328
box -38 -48 406 592
use scs8hd_decap_12  FILLER_82_32
timestamp 1586364061
transform 1 0 4048 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_44
timestamp 1586364061
transform 1 0 5152 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_56
timestamp 1586364061
transform 1 0 6256 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_68
timestamp 1586364061
transform 1 0 7360 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_3  PHY_165
timestamp 1586364061
transform -1 0 8832 0 -1 47328
box -38 -48 314 592
use scs8hd_fill_1  FILLER_82_80
timestamp 1586364061
transform 1 0 8464 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_3  PHY_166
timestamp 1586364061
transform 1 0 1104 0 1 47328
box -38 -48 314 592
use scs8hd_decap_12  FILLER_83_3
timestamp 1586364061
transform 1 0 1380 0 1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_83_15
timestamp 1586364061
transform 1 0 2484 0 1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_83_27
timestamp 1586364061
transform 1 0 3588 0 1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_83_39
timestamp 1586364061
transform 1 0 4692 0 1 47328
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_83_51
timestamp 1586364061
transform 1 0 5796 0 1 47328
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1292
timestamp 1586364061
transform 1 0 6716 0 1 47328
box -38 -48 130 592
use scs8hd_fill_2  FILLER_83_59
timestamp 1586364061
transform 1 0 6532 0 1 47328
box -38 -48 222 592
use scs8hd_decap_12  FILLER_83_62
timestamp 1586364061
transform 1 0 6808 0 1 47328
box -38 -48 1142 592
use scs8hd_decap_3  PHY_167
timestamp 1586364061
transform -1 0 8832 0 1 47328
box -38 -48 314 592
use scs8hd_decap_6  FILLER_83_74
timestamp 1586364061
transform 1 0 7912 0 1 47328
box -38 -48 590 592
use scs8hd_fill_1  FILLER_83_80
timestamp 1586364061
transform 1 0 8464 0 1 47328
box -38 -48 130 592
use scs8hd_decap_3  PHY_168
timestamp 1586364061
transform 1 0 1104 0 -1 48416
box -38 -48 314 592
use scs8hd_decap_12  FILLER_84_3
timestamp 1586364061
transform 1 0 1380 0 -1 48416
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_84_15
timestamp 1586364061
transform 1 0 2484 0 -1 48416
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1293
timestamp 1586364061
transform 1 0 3956 0 -1 48416
box -38 -48 130 592
use scs8hd_decap_4  FILLER_84_27
timestamp 1586364061
transform 1 0 3588 0 -1 48416
box -38 -48 406 592
use scs8hd_decap_12  FILLER_84_32
timestamp 1586364061
transform 1 0 4048 0 -1 48416
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_84_44
timestamp 1586364061
transform 1 0 5152 0 -1 48416
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_84_56
timestamp 1586364061
transform 1 0 6256 0 -1 48416
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_84_68
timestamp 1586364061
transform 1 0 7360 0 -1 48416
box -38 -48 1142 592
use scs8hd_decap_3  PHY_169
timestamp 1586364061
transform -1 0 8832 0 -1 48416
box -38 -48 314 592
use scs8hd_fill_1  FILLER_84_80
timestamp 1586364061
transform 1 0 8464 0 -1 48416
box -38 -48 130 592
use scs8hd_decap_3  PHY_170
timestamp 1586364061
transform 1 0 1104 0 1 48416
box -38 -48 314 592
use scs8hd_decap_3  PHY_172
timestamp 1586364061
transform 1 0 1104 0 -1 49504
box -38 -48 314 592
use scs8hd_decap_12  FILLER_85_3
timestamp 1586364061
transform 1 0 1380 0 1 48416
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_85_15
timestamp 1586364061
transform 1 0 2484 0 1 48416
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_86_3
timestamp 1586364061
transform 1 0 1380 0 -1 49504
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_86_15
timestamp 1586364061
transform 1 0 2484 0 -1 49504
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1295
timestamp 1586364061
transform 1 0 3956 0 -1 49504
box -38 -48 130 592
use scs8hd_decap_12  FILLER_85_27
timestamp 1586364061
transform 1 0 3588 0 1 48416
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_86_27
timestamp 1586364061
transform 1 0 3588 0 -1 49504
box -38 -48 406 592
use scs8hd_decap_12  FILLER_86_32
timestamp 1586364061
transform 1 0 4048 0 -1 49504
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_85_39
timestamp 1586364061
transform 1 0 4692 0 1 48416
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_85_51
timestamp 1586364061
transform 1 0 5796 0 1 48416
box -38 -48 774 592
use scs8hd_decap_12  FILLER_86_44
timestamp 1586364061
transform 1 0 5152 0 -1 49504
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1294
timestamp 1586364061
transform 1 0 6716 0 1 48416
box -38 -48 130 592
use scs8hd_fill_2  FILLER_85_59
timestamp 1586364061
transform 1 0 6532 0 1 48416
box -38 -48 222 592
use scs8hd_decap_12  FILLER_85_62
timestamp 1586364061
transform 1 0 6808 0 1 48416
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_86_56
timestamp 1586364061
transform 1 0 6256 0 -1 49504
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_86_68
timestamp 1586364061
transform 1 0 7360 0 -1 49504
box -38 -48 1142 592
use scs8hd_decap_3  PHY_171
timestamp 1586364061
transform -1 0 8832 0 1 48416
box -38 -48 314 592
use scs8hd_decap_3  PHY_173
timestamp 1586364061
transform -1 0 8832 0 -1 49504
box -38 -48 314 592
use scs8hd_decap_6  FILLER_85_74
timestamp 1586364061
transform 1 0 7912 0 1 48416
box -38 -48 590 592
use scs8hd_fill_1  FILLER_85_80
timestamp 1586364061
transform 1 0 8464 0 1 48416
box -38 -48 130 592
use scs8hd_fill_1  FILLER_86_80
timestamp 1586364061
transform 1 0 8464 0 -1 49504
box -38 -48 130 592
use scs8hd_decap_3  PHY_174
timestamp 1586364061
transform 1 0 1104 0 1 49504
box -38 -48 314 592
use scs8hd_decap_12  FILLER_87_3
timestamp 1586364061
transform 1 0 1380 0 1 49504
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_87_15
timestamp 1586364061
transform 1 0 2484 0 1 49504
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_87_27
timestamp 1586364061
transform 1 0 3588 0 1 49504
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_87_39
timestamp 1586364061
transform 1 0 4692 0 1 49504
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_87_51
timestamp 1586364061
transform 1 0 5796 0 1 49504
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1296
timestamp 1586364061
transform 1 0 6716 0 1 49504
box -38 -48 130 592
use scs8hd_fill_2  FILLER_87_59
timestamp 1586364061
transform 1 0 6532 0 1 49504
box -38 -48 222 592
use scs8hd_decap_12  FILLER_87_62
timestamp 1586364061
transform 1 0 6808 0 1 49504
box -38 -48 1142 592
use scs8hd_decap_3  PHY_175
timestamp 1586364061
transform -1 0 8832 0 1 49504
box -38 -48 314 592
use scs8hd_decap_6  FILLER_87_74
timestamp 1586364061
transform 1 0 7912 0 1 49504
box -38 -48 590 592
use scs8hd_fill_1  FILLER_87_80
timestamp 1586364061
transform 1 0 8464 0 1 49504
box -38 -48 130 592
use scs8hd_decap_3  PHY_176
timestamp 1586364061
transform 1 0 1104 0 -1 50592
box -38 -48 314 592
use scs8hd_decap_12  FILLER_88_3
timestamp 1586364061
transform 1 0 1380 0 -1 50592
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_88_15
timestamp 1586364061
transform 1 0 2484 0 -1 50592
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1297
timestamp 1586364061
transform 1 0 3956 0 -1 50592
box -38 -48 130 592
use scs8hd_decap_4  FILLER_88_27
timestamp 1586364061
transform 1 0 3588 0 -1 50592
box -38 -48 406 592
use scs8hd_decap_12  FILLER_88_32
timestamp 1586364061
transform 1 0 4048 0 -1 50592
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_88_44
timestamp 1586364061
transform 1 0 5152 0 -1 50592
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_88_56
timestamp 1586364061
transform 1 0 6256 0 -1 50592
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_88_68
timestamp 1586364061
transform 1 0 7360 0 -1 50592
box -38 -48 1142 592
use scs8hd_decap_3  PHY_177
timestamp 1586364061
transform -1 0 8832 0 -1 50592
box -38 -48 314 592
use scs8hd_fill_1  FILLER_88_80
timestamp 1586364061
transform 1 0 8464 0 -1 50592
box -38 -48 130 592
use scs8hd_decap_3  PHY_178
timestamp 1586364061
transform 1 0 1104 0 1 50592
box -38 -48 314 592
use scs8hd_decap_12  FILLER_89_3
timestamp 1586364061
transform 1 0 1380 0 1 50592
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_89_15
timestamp 1586364061
transform 1 0 2484 0 1 50592
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_89_27
timestamp 1586364061
transform 1 0 3588 0 1 50592
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_89_39
timestamp 1586364061
transform 1 0 4692 0 1 50592
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_89_51
timestamp 1586364061
transform 1 0 5796 0 1 50592
box -38 -48 774 592
use scs8hd_buf_2  _16_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6808 0 1 50592
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_1298
timestamp 1586364061
transform 1 0 6716 0 1 50592
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__16__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7360 0 1 50592
box -38 -48 222 592
use scs8hd_fill_2  FILLER_89_59
timestamp 1586364061
transform 1 0 6532 0 1 50592
box -38 -48 222 592
use scs8hd_fill_2  FILLER_89_66
timestamp 1586364061
transform 1 0 7176 0 1 50592
box -38 -48 222 592
use scs8hd_decap_8  FILLER_89_70
timestamp 1586364061
transform 1 0 7544 0 1 50592
box -38 -48 774 592
use scs8hd_decap_3  PHY_179
timestamp 1586364061
transform -1 0 8832 0 1 50592
box -38 -48 314 592
use scs8hd_decap_3  FILLER_89_78
timestamp 1586364061
transform 1 0 8280 0 1 50592
box -38 -48 314 592
use scs8hd_decap_3  PHY_180
timestamp 1586364061
transform 1 0 1104 0 -1 51680
box -38 -48 314 592
use scs8hd_decap_12  FILLER_90_3
timestamp 1586364061
transform 1 0 1380 0 -1 51680
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_90_15
timestamp 1586364061
transform 1 0 2484 0 -1 51680
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1299
timestamp 1586364061
transform 1 0 3956 0 -1 51680
box -38 -48 130 592
use scs8hd_decap_4  FILLER_90_27
timestamp 1586364061
transform 1 0 3588 0 -1 51680
box -38 -48 406 592
use scs8hd_decap_12  FILLER_90_32
timestamp 1586364061
transform 1 0 4048 0 -1 51680
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_90_44
timestamp 1586364061
transform 1 0 5152 0 -1 51680
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_90_56
timestamp 1586364061
transform 1 0 6256 0 -1 51680
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_90_68
timestamp 1586364061
transform 1 0 7360 0 -1 51680
box -38 -48 1142 592
use scs8hd_decap_3  PHY_181
timestamp 1586364061
transform -1 0 8832 0 -1 51680
box -38 -48 314 592
use scs8hd_fill_1  FILLER_90_80
timestamp 1586364061
transform 1 0 8464 0 -1 51680
box -38 -48 130 592
use scs8hd_decap_3  PHY_182
timestamp 1586364061
transform 1 0 1104 0 1 51680
box -38 -48 314 592
use scs8hd_decap_12  FILLER_91_3
timestamp 1586364061
transform 1 0 1380 0 1 51680
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_91_15
timestamp 1586364061
transform 1 0 2484 0 1 51680
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_91_27
timestamp 1586364061
transform 1 0 3588 0 1 51680
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_91_39
timestamp 1586364061
transform 1 0 4692 0 1 51680
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_91_51
timestamp 1586364061
transform 1 0 5796 0 1 51680
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1300
timestamp 1586364061
transform 1 0 6716 0 1 51680
box -38 -48 130 592
use scs8hd_fill_2  FILLER_91_59
timestamp 1586364061
transform 1 0 6532 0 1 51680
box -38 -48 222 592
use scs8hd_decap_12  FILLER_91_62
timestamp 1586364061
transform 1 0 6808 0 1 51680
box -38 -48 1142 592
use scs8hd_decap_3  PHY_183
timestamp 1586364061
transform -1 0 8832 0 1 51680
box -38 -48 314 592
use scs8hd_decap_6  FILLER_91_74
timestamp 1586364061
transform 1 0 7912 0 1 51680
box -38 -48 590 592
use scs8hd_fill_1  FILLER_91_80
timestamp 1586364061
transform 1 0 8464 0 1 51680
box -38 -48 130 592
use scs8hd_decap_3  PHY_184
timestamp 1586364061
transform 1 0 1104 0 -1 52768
box -38 -48 314 592
use scs8hd_decap_3  PHY_186
timestamp 1586364061
transform 1 0 1104 0 1 52768
box -38 -48 314 592
use scs8hd_decap_12  FILLER_92_3
timestamp 1586364061
transform 1 0 1380 0 -1 52768
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_92_15
timestamp 1586364061
transform 1 0 2484 0 -1 52768
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_93_3
timestamp 1586364061
transform 1 0 1380 0 1 52768
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_93_15
timestamp 1586364061
transform 1 0 2484 0 1 52768
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1301
timestamp 1586364061
transform 1 0 3956 0 -1 52768
box -38 -48 130 592
use scs8hd_decap_4  FILLER_92_27
timestamp 1586364061
transform 1 0 3588 0 -1 52768
box -38 -48 406 592
use scs8hd_decap_12  FILLER_92_32
timestamp 1586364061
transform 1 0 4048 0 -1 52768
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_93_27
timestamp 1586364061
transform 1 0 3588 0 1 52768
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_92_44
timestamp 1586364061
transform 1 0 5152 0 -1 52768
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_93_39
timestamp 1586364061
transform 1 0 4692 0 1 52768
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_93_51
timestamp 1586364061
transform 1 0 5796 0 1 52768
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1302
timestamp 1586364061
transform 1 0 6716 0 1 52768
box -38 -48 130 592
use scs8hd_decap_12  FILLER_92_56
timestamp 1586364061
transform 1 0 6256 0 -1 52768
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_92_68
timestamp 1586364061
transform 1 0 7360 0 -1 52768
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_93_59
timestamp 1586364061
transform 1 0 6532 0 1 52768
box -38 -48 222 592
use scs8hd_decap_12  FILLER_93_62
timestamp 1586364061
transform 1 0 6808 0 1 52768
box -38 -48 1142 592
use scs8hd_decap_3  PHY_185
timestamp 1586364061
transform -1 0 8832 0 -1 52768
box -38 -48 314 592
use scs8hd_decap_3  PHY_187
timestamp 1586364061
transform -1 0 8832 0 1 52768
box -38 -48 314 592
use scs8hd_fill_1  FILLER_92_80
timestamp 1586364061
transform 1 0 8464 0 -1 52768
box -38 -48 130 592
use scs8hd_decap_6  FILLER_93_74
timestamp 1586364061
transform 1 0 7912 0 1 52768
box -38 -48 590 592
use scs8hd_fill_1  FILLER_93_80
timestamp 1586364061
transform 1 0 8464 0 1 52768
box -38 -48 130 592
use scs8hd_decap_3  PHY_188
timestamp 1586364061
transform 1 0 1104 0 -1 53856
box -38 -48 314 592
use scs8hd_decap_12  FILLER_94_3
timestamp 1586364061
transform 1 0 1380 0 -1 53856
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_94_15
timestamp 1586364061
transform 1 0 2484 0 -1 53856
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1303
timestamp 1586364061
transform 1 0 3956 0 -1 53856
box -38 -48 130 592
use scs8hd_decap_4  FILLER_94_27
timestamp 1586364061
transform 1 0 3588 0 -1 53856
box -38 -48 406 592
use scs8hd_decap_12  FILLER_94_32
timestamp 1586364061
transform 1 0 4048 0 -1 53856
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_94_44
timestamp 1586364061
transform 1 0 5152 0 -1 53856
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_94_56
timestamp 1586364061
transform 1 0 6256 0 -1 53856
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_94_68
timestamp 1586364061
transform 1 0 7360 0 -1 53856
box -38 -48 1142 592
use scs8hd_decap_3  PHY_189
timestamp 1586364061
transform -1 0 8832 0 -1 53856
box -38 -48 314 592
use scs8hd_fill_1  FILLER_94_80
timestamp 1586364061
transform 1 0 8464 0 -1 53856
box -38 -48 130 592
use scs8hd_decap_3  PHY_190
timestamp 1586364061
transform 1 0 1104 0 1 53856
box -38 -48 314 592
use scs8hd_decap_12  FILLER_95_3
timestamp 1586364061
transform 1 0 1380 0 1 53856
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_95_15
timestamp 1586364061
transform 1 0 2484 0 1 53856
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_95_27
timestamp 1586364061
transform 1 0 3588 0 1 53856
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_95_39
timestamp 1586364061
transform 1 0 4692 0 1 53856
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_95_51
timestamp 1586364061
transform 1 0 5796 0 1 53856
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1304
timestamp 1586364061
transform 1 0 6716 0 1 53856
box -38 -48 130 592
use scs8hd_fill_2  FILLER_95_59
timestamp 1586364061
transform 1 0 6532 0 1 53856
box -38 -48 222 592
use scs8hd_decap_12  FILLER_95_62
timestamp 1586364061
transform 1 0 6808 0 1 53856
box -38 -48 1142 592
use scs8hd_decap_3  PHY_191
timestamp 1586364061
transform -1 0 8832 0 1 53856
box -38 -48 314 592
use scs8hd_decap_6  FILLER_95_74
timestamp 1586364061
transform 1 0 7912 0 1 53856
box -38 -48 590 592
use scs8hd_fill_1  FILLER_95_80
timestamp 1586364061
transform 1 0 8464 0 1 53856
box -38 -48 130 592
use scs8hd_decap_3  PHY_192
timestamp 1586364061
transform 1 0 1104 0 -1 54944
box -38 -48 314 592
use scs8hd_decap_12  FILLER_96_3
timestamp 1586364061
transform 1 0 1380 0 -1 54944
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_96_15
timestamp 1586364061
transform 1 0 2484 0 -1 54944
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1305
timestamp 1586364061
transform 1 0 3956 0 -1 54944
box -38 -48 130 592
use scs8hd_decap_4  FILLER_96_27
timestamp 1586364061
transform 1 0 3588 0 -1 54944
box -38 -48 406 592
use scs8hd_decap_12  FILLER_96_32
timestamp 1586364061
transform 1 0 4048 0 -1 54944
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_96_44
timestamp 1586364061
transform 1 0 5152 0 -1 54944
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_96_56
timestamp 1586364061
transform 1 0 6256 0 -1 54944
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_96_68
timestamp 1586364061
transform 1 0 7360 0 -1 54944
box -38 -48 1142 592
use scs8hd_decap_3  PHY_193
timestamp 1586364061
transform -1 0 8832 0 -1 54944
box -38 -48 314 592
use scs8hd_fill_1  FILLER_96_80
timestamp 1586364061
transform 1 0 8464 0 -1 54944
box -38 -48 130 592
use scs8hd_decap_3  PHY_194
timestamp 1586364061
transform 1 0 1104 0 1 54944
box -38 -48 314 592
use scs8hd_decap_12  FILLER_97_3
timestamp 1586364061
transform 1 0 1380 0 1 54944
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_97_15
timestamp 1586364061
transform 1 0 2484 0 1 54944
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_97_27
timestamp 1586364061
transform 1 0 3588 0 1 54944
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_97_39
timestamp 1586364061
transform 1 0 4692 0 1 54944
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_97_51
timestamp 1586364061
transform 1 0 5796 0 1 54944
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1306
timestamp 1586364061
transform 1 0 6716 0 1 54944
box -38 -48 130 592
use scs8hd_fill_2  FILLER_97_59
timestamp 1586364061
transform 1 0 6532 0 1 54944
box -38 -48 222 592
use scs8hd_decap_12  FILLER_97_62
timestamp 1586364061
transform 1 0 6808 0 1 54944
box -38 -48 1142 592
use scs8hd_decap_3  PHY_195
timestamp 1586364061
transform -1 0 8832 0 1 54944
box -38 -48 314 592
use scs8hd_decap_6  FILLER_97_74
timestamp 1586364061
transform 1 0 7912 0 1 54944
box -38 -48 590 592
use scs8hd_fill_1  FILLER_97_80
timestamp 1586364061
transform 1 0 8464 0 1 54944
box -38 -48 130 592
use scs8hd_decap_3  PHY_196
timestamp 1586364061
transform 1 0 1104 0 -1 56032
box -38 -48 314 592
use scs8hd_decap_12  FILLER_98_3
timestamp 1586364061
transform 1 0 1380 0 -1 56032
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_98_15
timestamp 1586364061
transform 1 0 2484 0 -1 56032
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1307
timestamp 1586364061
transform 1 0 3956 0 -1 56032
box -38 -48 130 592
use scs8hd_decap_4  FILLER_98_27
timestamp 1586364061
transform 1 0 3588 0 -1 56032
box -38 -48 406 592
use scs8hd_decap_12  FILLER_98_32
timestamp 1586364061
transform 1 0 4048 0 -1 56032
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_98_44
timestamp 1586364061
transform 1 0 5152 0 -1 56032
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_98_56
timestamp 1586364061
transform 1 0 6256 0 -1 56032
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_98_68
timestamp 1586364061
transform 1 0 7360 0 -1 56032
box -38 -48 1142 592
use scs8hd_decap_3  PHY_197
timestamp 1586364061
transform -1 0 8832 0 -1 56032
box -38 -48 314 592
use scs8hd_fill_1  FILLER_98_80
timestamp 1586364061
transform 1 0 8464 0 -1 56032
box -38 -48 130 592
use scs8hd_decap_3  PHY_198
timestamp 1586364061
transform 1 0 1104 0 1 56032
box -38 -48 314 592
use scs8hd_decap_3  PHY_200
timestamp 1586364061
transform 1 0 1104 0 -1 57120
box -38 -48 314 592
use scs8hd_decap_12  FILLER_99_3
timestamp 1586364061
transform 1 0 1380 0 1 56032
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_99_15
timestamp 1586364061
transform 1 0 2484 0 1 56032
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_100_3
timestamp 1586364061
transform 1 0 1380 0 -1 57120
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_100_15
timestamp 1586364061
transform 1 0 2484 0 -1 57120
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1309
timestamp 1586364061
transform 1 0 3956 0 -1 57120
box -38 -48 130 592
use scs8hd_decap_12  FILLER_99_27
timestamp 1586364061
transform 1 0 3588 0 1 56032
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_100_27
timestamp 1586364061
transform 1 0 3588 0 -1 57120
box -38 -48 406 592
use scs8hd_decap_12  FILLER_100_32
timestamp 1586364061
transform 1 0 4048 0 -1 57120
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_99_39
timestamp 1586364061
transform 1 0 4692 0 1 56032
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_99_51
timestamp 1586364061
transform 1 0 5796 0 1 56032
box -38 -48 774 592
use scs8hd_decap_12  FILLER_100_44
timestamp 1586364061
transform 1 0 5152 0 -1 57120
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1308
timestamp 1586364061
transform 1 0 6716 0 1 56032
box -38 -48 130 592
use scs8hd_fill_2  FILLER_99_59
timestamp 1586364061
transform 1 0 6532 0 1 56032
box -38 -48 222 592
use scs8hd_decap_12  FILLER_99_62
timestamp 1586364061
transform 1 0 6808 0 1 56032
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_100_56
timestamp 1586364061
transform 1 0 6256 0 -1 57120
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_100_68
timestamp 1586364061
transform 1 0 7360 0 -1 57120
box -38 -48 1142 592
use scs8hd_decap_3  PHY_199
timestamp 1586364061
transform -1 0 8832 0 1 56032
box -38 -48 314 592
use scs8hd_decap_3  PHY_201
timestamp 1586364061
transform -1 0 8832 0 -1 57120
box -38 -48 314 592
use scs8hd_decap_6  FILLER_99_74
timestamp 1586364061
transform 1 0 7912 0 1 56032
box -38 -48 590 592
use scs8hd_fill_1  FILLER_99_80
timestamp 1586364061
transform 1 0 8464 0 1 56032
box -38 -48 130 592
use scs8hd_fill_1  FILLER_100_80
timestamp 1586364061
transform 1 0 8464 0 -1 57120
box -38 -48 130 592
use scs8hd_decap_3  PHY_202
timestamp 1586364061
transform 1 0 1104 0 1 57120
box -38 -48 314 592
use scs8hd_decap_12  FILLER_101_3
timestamp 1586364061
transform 1 0 1380 0 1 57120
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_101_15
timestamp 1586364061
transform 1 0 2484 0 1 57120
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_101_27
timestamp 1586364061
transform 1 0 3588 0 1 57120
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_101_39
timestamp 1586364061
transform 1 0 4692 0 1 57120
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_101_51
timestamp 1586364061
transform 1 0 5796 0 1 57120
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1310
timestamp 1586364061
transform 1 0 6716 0 1 57120
box -38 -48 130 592
use scs8hd_fill_2  FILLER_101_59
timestamp 1586364061
transform 1 0 6532 0 1 57120
box -38 -48 222 592
use scs8hd_decap_12  FILLER_101_62
timestamp 1586364061
transform 1 0 6808 0 1 57120
box -38 -48 1142 592
use scs8hd_decap_3  PHY_203
timestamp 1586364061
transform -1 0 8832 0 1 57120
box -38 -48 314 592
use scs8hd_decap_6  FILLER_101_74
timestamp 1586364061
transform 1 0 7912 0 1 57120
box -38 -48 590 592
use scs8hd_fill_1  FILLER_101_80
timestamp 1586364061
transform 1 0 8464 0 1 57120
box -38 -48 130 592
use scs8hd_decap_3  PHY_204
timestamp 1586364061
transform 1 0 1104 0 -1 58208
box -38 -48 314 592
use scs8hd_decap_12  FILLER_102_3
timestamp 1586364061
transform 1 0 1380 0 -1 58208
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_102_15
timestamp 1586364061
transform 1 0 2484 0 -1 58208
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1311
timestamp 1586364061
transform 1 0 3956 0 -1 58208
box -38 -48 130 592
use scs8hd_decap_4  FILLER_102_27
timestamp 1586364061
transform 1 0 3588 0 -1 58208
box -38 -48 406 592
use scs8hd_decap_12  FILLER_102_32
timestamp 1586364061
transform 1 0 4048 0 -1 58208
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_102_44
timestamp 1586364061
transform 1 0 5152 0 -1 58208
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_102_56
timestamp 1586364061
transform 1 0 6256 0 -1 58208
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_102_68
timestamp 1586364061
transform 1 0 7360 0 -1 58208
box -38 -48 1142 592
use scs8hd_decap_3  PHY_205
timestamp 1586364061
transform -1 0 8832 0 -1 58208
box -38 -48 314 592
use scs8hd_fill_1  FILLER_102_80
timestamp 1586364061
transform 1 0 8464 0 -1 58208
box -38 -48 130 592
use scs8hd_decap_3  PHY_206
timestamp 1586364061
transform 1 0 1104 0 1 58208
box -38 -48 314 592
use scs8hd_decap_12  FILLER_103_3
timestamp 1586364061
transform 1 0 1380 0 1 58208
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_103_15
timestamp 1586364061
transform 1 0 2484 0 1 58208
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_103_27
timestamp 1586364061
transform 1 0 3588 0 1 58208
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_103_39
timestamp 1586364061
transform 1 0 4692 0 1 58208
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_103_51
timestamp 1586364061
transform 1 0 5796 0 1 58208
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1312
timestamp 1586364061
transform 1 0 6716 0 1 58208
box -38 -48 130 592
use scs8hd_fill_2  FILLER_103_59
timestamp 1586364061
transform 1 0 6532 0 1 58208
box -38 -48 222 592
use scs8hd_decap_12  FILLER_103_62
timestamp 1586364061
transform 1 0 6808 0 1 58208
box -38 -48 1142 592
use scs8hd_decap_3  PHY_207
timestamp 1586364061
transform -1 0 8832 0 1 58208
box -38 -48 314 592
use scs8hd_decap_6  FILLER_103_74
timestamp 1586364061
transform 1 0 7912 0 1 58208
box -38 -48 590 592
use scs8hd_fill_1  FILLER_103_80
timestamp 1586364061
transform 1 0 8464 0 1 58208
box -38 -48 130 592
use scs8hd_decap_3  PHY_208
timestamp 1586364061
transform 1 0 1104 0 -1 59296
box -38 -48 314 592
use scs8hd_decap_12  FILLER_104_3
timestamp 1586364061
transform 1 0 1380 0 -1 59296
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_104_15
timestamp 1586364061
transform 1 0 2484 0 -1 59296
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1313
timestamp 1586364061
transform 1 0 3956 0 -1 59296
box -38 -48 130 592
use scs8hd_decap_4  FILLER_104_27
timestamp 1586364061
transform 1 0 3588 0 -1 59296
box -38 -48 406 592
use scs8hd_decap_12  FILLER_104_32
timestamp 1586364061
transform 1 0 4048 0 -1 59296
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_104_44
timestamp 1586364061
transform 1 0 5152 0 -1 59296
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_104_56
timestamp 1586364061
transform 1 0 6256 0 -1 59296
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_104_68
timestamp 1586364061
transform 1 0 7360 0 -1 59296
box -38 -48 1142 592
use scs8hd_decap_3  PHY_209
timestamp 1586364061
transform -1 0 8832 0 -1 59296
box -38 -48 314 592
use scs8hd_fill_1  FILLER_104_80
timestamp 1586364061
transform 1 0 8464 0 -1 59296
box -38 -48 130 592
use scs8hd_decap_3  PHY_210
timestamp 1586364061
transform 1 0 1104 0 1 59296
box -38 -48 314 592
use scs8hd_decap_3  PHY_212
timestamp 1586364061
transform 1 0 1104 0 -1 60384
box -38 -48 314 592
use scs8hd_decap_12  FILLER_105_3
timestamp 1586364061
transform 1 0 1380 0 1 59296
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_105_15
timestamp 1586364061
transform 1 0 2484 0 1 59296
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_106_3
timestamp 1586364061
transform 1 0 1380 0 -1 60384
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_106_15
timestamp 1586364061
transform 1 0 2484 0 -1 60384
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1315
timestamp 1586364061
transform 1 0 3956 0 -1 60384
box -38 -48 130 592
use scs8hd_decap_12  FILLER_105_27
timestamp 1586364061
transform 1 0 3588 0 1 59296
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_106_27
timestamp 1586364061
transform 1 0 3588 0 -1 60384
box -38 -48 406 592
use scs8hd_decap_12  FILLER_106_32
timestamp 1586364061
transform 1 0 4048 0 -1 60384
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_105_39
timestamp 1586364061
transform 1 0 4692 0 1 59296
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_105_51
timestamp 1586364061
transform 1 0 5796 0 1 59296
box -38 -48 774 592
use scs8hd_decap_12  FILLER_106_44
timestamp 1586364061
transform 1 0 5152 0 -1 60384
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1314
timestamp 1586364061
transform 1 0 6716 0 1 59296
box -38 -48 130 592
use scs8hd_fill_2  FILLER_105_59
timestamp 1586364061
transform 1 0 6532 0 1 59296
box -38 -48 222 592
use scs8hd_decap_12  FILLER_105_62
timestamp 1586364061
transform 1 0 6808 0 1 59296
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_106_56
timestamp 1586364061
transform 1 0 6256 0 -1 60384
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_106_68
timestamp 1586364061
transform 1 0 7360 0 -1 60384
box -38 -48 1142 592
use scs8hd_decap_3  PHY_211
timestamp 1586364061
transform -1 0 8832 0 1 59296
box -38 -48 314 592
use scs8hd_decap_3  PHY_213
timestamp 1586364061
transform -1 0 8832 0 -1 60384
box -38 -48 314 592
use scs8hd_decap_6  FILLER_105_74
timestamp 1586364061
transform 1 0 7912 0 1 59296
box -38 -48 590 592
use scs8hd_fill_1  FILLER_105_80
timestamp 1586364061
transform 1 0 8464 0 1 59296
box -38 -48 130 592
use scs8hd_fill_1  FILLER_106_80
timestamp 1586364061
transform 1 0 8464 0 -1 60384
box -38 -48 130 592
use scs8hd_decap_3  PHY_214
timestamp 1586364061
transform 1 0 1104 0 1 60384
box -38 -48 314 592
use scs8hd_decap_12  FILLER_107_3
timestamp 1586364061
transform 1 0 1380 0 1 60384
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_107_15
timestamp 1586364061
transform 1 0 2484 0 1 60384
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_107_27
timestamp 1586364061
transform 1 0 3588 0 1 60384
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_107_39
timestamp 1586364061
transform 1 0 4692 0 1 60384
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_107_51
timestamp 1586364061
transform 1 0 5796 0 1 60384
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1316
timestamp 1586364061
transform 1 0 6716 0 1 60384
box -38 -48 130 592
use scs8hd_fill_2  FILLER_107_59
timestamp 1586364061
transform 1 0 6532 0 1 60384
box -38 -48 222 592
use scs8hd_decap_12  FILLER_107_62
timestamp 1586364061
transform 1 0 6808 0 1 60384
box -38 -48 1142 592
use scs8hd_decap_3  PHY_215
timestamp 1586364061
transform -1 0 8832 0 1 60384
box -38 -48 314 592
use scs8hd_decap_6  FILLER_107_74
timestamp 1586364061
transform 1 0 7912 0 1 60384
box -38 -48 590 592
use scs8hd_fill_1  FILLER_107_80
timestamp 1586364061
transform 1 0 8464 0 1 60384
box -38 -48 130 592
use scs8hd_decap_3  PHY_216
timestamp 1586364061
transform 1 0 1104 0 -1 61472
box -38 -48 314 592
use scs8hd_decap_12  FILLER_108_3
timestamp 1586364061
transform 1 0 1380 0 -1 61472
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_108_15
timestamp 1586364061
transform 1 0 2484 0 -1 61472
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1317
timestamp 1586364061
transform 1 0 3956 0 -1 61472
box -38 -48 130 592
use scs8hd_decap_4  FILLER_108_27
timestamp 1586364061
transform 1 0 3588 0 -1 61472
box -38 -48 406 592
use scs8hd_decap_12  FILLER_108_32
timestamp 1586364061
transform 1 0 4048 0 -1 61472
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_108_44
timestamp 1586364061
transform 1 0 5152 0 -1 61472
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_108_56
timestamp 1586364061
transform 1 0 6256 0 -1 61472
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_108_68
timestamp 1586364061
transform 1 0 7360 0 -1 61472
box -38 -48 1142 592
use scs8hd_decap_3  PHY_217
timestamp 1586364061
transform -1 0 8832 0 -1 61472
box -38 -48 314 592
use scs8hd_fill_1  FILLER_108_80
timestamp 1586364061
transform 1 0 8464 0 -1 61472
box -38 -48 130 592
use scs8hd_decap_3  PHY_218
timestamp 1586364061
transform 1 0 1104 0 1 61472
box -38 -48 314 592
use scs8hd_decap_12  FILLER_109_3
timestamp 1586364061
transform 1 0 1380 0 1 61472
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_109_15
timestamp 1586364061
transform 1 0 2484 0 1 61472
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_109_27
timestamp 1586364061
transform 1 0 3588 0 1 61472
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_109_39
timestamp 1586364061
transform 1 0 4692 0 1 61472
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_109_51
timestamp 1586364061
transform 1 0 5796 0 1 61472
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1318
timestamp 1586364061
transform 1 0 6716 0 1 61472
box -38 -48 130 592
use scs8hd_fill_2  FILLER_109_59
timestamp 1586364061
transform 1 0 6532 0 1 61472
box -38 -48 222 592
use scs8hd_decap_12  FILLER_109_62
timestamp 1586364061
transform 1 0 6808 0 1 61472
box -38 -48 1142 592
use scs8hd_decap_3  PHY_219
timestamp 1586364061
transform -1 0 8832 0 1 61472
box -38 -48 314 592
use scs8hd_decap_6  FILLER_109_74
timestamp 1586364061
transform 1 0 7912 0 1 61472
box -38 -48 590 592
use scs8hd_fill_1  FILLER_109_80
timestamp 1586364061
transform 1 0 8464 0 1 61472
box -38 -48 130 592
use scs8hd_decap_3  PHY_220
timestamp 1586364061
transform 1 0 1104 0 -1 62560
box -38 -48 314 592
use scs8hd_decap_12  FILLER_110_3
timestamp 1586364061
transform 1 0 1380 0 -1 62560
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_110_15
timestamp 1586364061
transform 1 0 2484 0 -1 62560
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1319
timestamp 1586364061
transform 1 0 3956 0 -1 62560
box -38 -48 130 592
use scs8hd_decap_4  FILLER_110_27
timestamp 1586364061
transform 1 0 3588 0 -1 62560
box -38 -48 406 592
use scs8hd_decap_12  FILLER_110_32
timestamp 1586364061
transform 1 0 4048 0 -1 62560
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_110_44
timestamp 1586364061
transform 1 0 5152 0 -1 62560
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_110_56
timestamp 1586364061
transform 1 0 6256 0 -1 62560
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_110_68
timestamp 1586364061
transform 1 0 7360 0 -1 62560
box -38 -48 1142 592
use scs8hd_decap_3  PHY_221
timestamp 1586364061
transform -1 0 8832 0 -1 62560
box -38 -48 314 592
use scs8hd_fill_1  FILLER_110_80
timestamp 1586364061
transform 1 0 8464 0 -1 62560
box -38 -48 130 592
use scs8hd_decap_3  PHY_222
timestamp 1586364061
transform 1 0 1104 0 1 62560
box -38 -48 314 592
use scs8hd_decap_12  FILLER_111_3
timestamp 1586364061
transform 1 0 1380 0 1 62560
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_111_15
timestamp 1586364061
transform 1 0 2484 0 1 62560
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_111_27
timestamp 1586364061
transform 1 0 3588 0 1 62560
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_111_39
timestamp 1586364061
transform 1 0 4692 0 1 62560
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_111_51
timestamp 1586364061
transform 1 0 5796 0 1 62560
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1320
timestamp 1586364061
transform 1 0 6716 0 1 62560
box -38 -48 130 592
use scs8hd_fill_2  FILLER_111_59
timestamp 1586364061
transform 1 0 6532 0 1 62560
box -38 -48 222 592
use scs8hd_decap_12  FILLER_111_62
timestamp 1586364061
transform 1 0 6808 0 1 62560
box -38 -48 1142 592
use scs8hd_decap_3  PHY_223
timestamp 1586364061
transform -1 0 8832 0 1 62560
box -38 -48 314 592
use scs8hd_decap_6  FILLER_111_74
timestamp 1586364061
transform 1 0 7912 0 1 62560
box -38 -48 590 592
use scs8hd_fill_1  FILLER_111_80
timestamp 1586364061
transform 1 0 8464 0 1 62560
box -38 -48 130 592
use scs8hd_decap_3  PHY_224
timestamp 1586364061
transform 1 0 1104 0 -1 63648
box -38 -48 314 592
use scs8hd_decap_3  PHY_226
timestamp 1586364061
transform 1 0 1104 0 1 63648
box -38 -48 314 592
use scs8hd_decap_12  FILLER_112_3
timestamp 1586364061
transform 1 0 1380 0 -1 63648
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_112_15
timestamp 1586364061
transform 1 0 2484 0 -1 63648
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_113_3
timestamp 1586364061
transform 1 0 1380 0 1 63648
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_113_15
timestamp 1586364061
transform 1 0 2484 0 1 63648
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1321
timestamp 1586364061
transform 1 0 3956 0 -1 63648
box -38 -48 130 592
use scs8hd_decap_4  FILLER_112_27
timestamp 1586364061
transform 1 0 3588 0 -1 63648
box -38 -48 406 592
use scs8hd_decap_12  FILLER_112_32
timestamp 1586364061
transform 1 0 4048 0 -1 63648
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_113_27
timestamp 1586364061
transform 1 0 3588 0 1 63648
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_112_44
timestamp 1586364061
transform 1 0 5152 0 -1 63648
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_113_39
timestamp 1586364061
transform 1 0 4692 0 1 63648
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_113_51
timestamp 1586364061
transform 1 0 5796 0 1 63648
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1322
timestamp 1586364061
transform 1 0 6716 0 1 63648
box -38 -48 130 592
use scs8hd_decap_12  FILLER_112_56
timestamp 1586364061
transform 1 0 6256 0 -1 63648
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_112_68
timestamp 1586364061
transform 1 0 7360 0 -1 63648
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_113_59
timestamp 1586364061
transform 1 0 6532 0 1 63648
box -38 -48 222 592
use scs8hd_decap_12  FILLER_113_62
timestamp 1586364061
transform 1 0 6808 0 1 63648
box -38 -48 1142 592
use scs8hd_decap_3  PHY_225
timestamp 1586364061
transform -1 0 8832 0 -1 63648
box -38 -48 314 592
use scs8hd_decap_3  PHY_227
timestamp 1586364061
transform -1 0 8832 0 1 63648
box -38 -48 314 592
use scs8hd_fill_1  FILLER_112_80
timestamp 1586364061
transform 1 0 8464 0 -1 63648
box -38 -48 130 592
use scs8hd_decap_6  FILLER_113_74
timestamp 1586364061
transform 1 0 7912 0 1 63648
box -38 -48 590 592
use scs8hd_fill_1  FILLER_113_80
timestamp 1586364061
transform 1 0 8464 0 1 63648
box -38 -48 130 592
use scs8hd_decap_3  PHY_228
timestamp 1586364061
transform 1 0 1104 0 -1 64736
box -38 -48 314 592
use scs8hd_decap_12  FILLER_114_3
timestamp 1586364061
transform 1 0 1380 0 -1 64736
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_114_15
timestamp 1586364061
transform 1 0 2484 0 -1 64736
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1323
timestamp 1586364061
transform 1 0 3956 0 -1 64736
box -38 -48 130 592
use scs8hd_decap_4  FILLER_114_27
timestamp 1586364061
transform 1 0 3588 0 -1 64736
box -38 -48 406 592
use scs8hd_decap_12  FILLER_114_32
timestamp 1586364061
transform 1 0 4048 0 -1 64736
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_114_44
timestamp 1586364061
transform 1 0 5152 0 -1 64736
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_114_56
timestamp 1586364061
transform 1 0 6256 0 -1 64736
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_114_68
timestamp 1586364061
transform 1 0 7360 0 -1 64736
box -38 -48 1142 592
use scs8hd_decap_3  PHY_229
timestamp 1586364061
transform -1 0 8832 0 -1 64736
box -38 -48 314 592
use scs8hd_fill_1  FILLER_114_80
timestamp 1586364061
transform 1 0 8464 0 -1 64736
box -38 -48 130 592
use scs8hd_decap_3  PHY_230
timestamp 1586364061
transform 1 0 1104 0 1 64736
box -38 -48 314 592
use scs8hd_decap_12  FILLER_115_3
timestamp 1586364061
transform 1 0 1380 0 1 64736
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_115_15
timestamp 1586364061
transform 1 0 2484 0 1 64736
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_115_27
timestamp 1586364061
transform 1 0 3588 0 1 64736
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_115_39
timestamp 1586364061
transform 1 0 4692 0 1 64736
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_115_51
timestamp 1586364061
transform 1 0 5796 0 1 64736
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1324
timestamp 1586364061
transform 1 0 6716 0 1 64736
box -38 -48 130 592
use scs8hd_fill_2  FILLER_115_59
timestamp 1586364061
transform 1 0 6532 0 1 64736
box -38 -48 222 592
use scs8hd_decap_12  FILLER_115_62
timestamp 1586364061
transform 1 0 6808 0 1 64736
box -38 -48 1142 592
use scs8hd_decap_3  PHY_231
timestamp 1586364061
transform -1 0 8832 0 1 64736
box -38 -48 314 592
use scs8hd_decap_6  FILLER_115_74
timestamp 1586364061
transform 1 0 7912 0 1 64736
box -38 -48 590 592
use scs8hd_fill_1  FILLER_115_80
timestamp 1586364061
transform 1 0 8464 0 1 64736
box -38 -48 130 592
use scs8hd_decap_3  PHY_232
timestamp 1586364061
transform 1 0 1104 0 -1 65824
box -38 -48 314 592
use scs8hd_decap_12  FILLER_116_3
timestamp 1586364061
transform 1 0 1380 0 -1 65824
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_116_15
timestamp 1586364061
transform 1 0 2484 0 -1 65824
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1325
timestamp 1586364061
transform 1 0 3956 0 -1 65824
box -38 -48 130 592
use scs8hd_decap_4  FILLER_116_27
timestamp 1586364061
transform 1 0 3588 0 -1 65824
box -38 -48 406 592
use scs8hd_decap_12  FILLER_116_32
timestamp 1586364061
transform 1 0 4048 0 -1 65824
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_116_44
timestamp 1586364061
transform 1 0 5152 0 -1 65824
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_116_56
timestamp 1586364061
transform 1 0 6256 0 -1 65824
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_116_68
timestamp 1586364061
transform 1 0 7360 0 -1 65824
box -38 -48 1142 592
use scs8hd_decap_3  PHY_233
timestamp 1586364061
transform -1 0 8832 0 -1 65824
box -38 -48 314 592
use scs8hd_fill_1  FILLER_116_80
timestamp 1586364061
transform 1 0 8464 0 -1 65824
box -38 -48 130 592
use scs8hd_decap_3  PHY_234
timestamp 1586364061
transform 1 0 1104 0 1 65824
box -38 -48 314 592
use scs8hd_decap_12  FILLER_117_3
timestamp 1586364061
transform 1 0 1380 0 1 65824
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_117_15
timestamp 1586364061
transform 1 0 2484 0 1 65824
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_117_27
timestamp 1586364061
transform 1 0 3588 0 1 65824
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_117_39
timestamp 1586364061
transform 1 0 4692 0 1 65824
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_117_51
timestamp 1586364061
transform 1 0 5796 0 1 65824
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1326
timestamp 1586364061
transform 1 0 6716 0 1 65824
box -38 -48 130 592
use scs8hd_fill_2  FILLER_117_59
timestamp 1586364061
transform 1 0 6532 0 1 65824
box -38 -48 222 592
use scs8hd_decap_12  FILLER_117_62
timestamp 1586364061
transform 1 0 6808 0 1 65824
box -38 -48 1142 592
use scs8hd_decap_3  PHY_235
timestamp 1586364061
transform -1 0 8832 0 1 65824
box -38 -48 314 592
use scs8hd_decap_6  FILLER_117_74
timestamp 1586364061
transform 1 0 7912 0 1 65824
box -38 -48 590 592
use scs8hd_fill_1  FILLER_117_80
timestamp 1586364061
transform 1 0 8464 0 1 65824
box -38 -48 130 592
use scs8hd_decap_3  PHY_236
timestamp 1586364061
transform 1 0 1104 0 -1 66912
box -38 -48 314 592
use scs8hd_decap_3  PHY_238
timestamp 1586364061
transform 1 0 1104 0 1 66912
box -38 -48 314 592
use scs8hd_decap_12  FILLER_118_3
timestamp 1586364061
transform 1 0 1380 0 -1 66912
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_118_15
timestamp 1586364061
transform 1 0 2484 0 -1 66912
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_119_3
timestamp 1586364061
transform 1 0 1380 0 1 66912
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_119_15
timestamp 1586364061
transform 1 0 2484 0 1 66912
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1327
timestamp 1586364061
transform 1 0 3956 0 -1 66912
box -38 -48 130 592
use scs8hd_decap_4  FILLER_118_27
timestamp 1586364061
transform 1 0 3588 0 -1 66912
box -38 -48 406 592
use scs8hd_decap_12  FILLER_118_32
timestamp 1586364061
transform 1 0 4048 0 -1 66912
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_119_27
timestamp 1586364061
transform 1 0 3588 0 1 66912
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_118_44
timestamp 1586364061
transform 1 0 5152 0 -1 66912
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_119_39
timestamp 1586364061
transform 1 0 4692 0 1 66912
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_119_51
timestamp 1586364061
transform 1 0 5796 0 1 66912
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1328
timestamp 1586364061
transform 1 0 6716 0 1 66912
box -38 -48 130 592
use scs8hd_decap_12  FILLER_118_56
timestamp 1586364061
transform 1 0 6256 0 -1 66912
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_118_68
timestamp 1586364061
transform 1 0 7360 0 -1 66912
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_119_59
timestamp 1586364061
transform 1 0 6532 0 1 66912
box -38 -48 222 592
use scs8hd_decap_12  FILLER_119_62
timestamp 1586364061
transform 1 0 6808 0 1 66912
box -38 -48 1142 592
use scs8hd_decap_3  PHY_237
timestamp 1586364061
transform -1 0 8832 0 -1 66912
box -38 -48 314 592
use scs8hd_decap_3  PHY_239
timestamp 1586364061
transform -1 0 8832 0 1 66912
box -38 -48 314 592
use scs8hd_fill_1  FILLER_118_80
timestamp 1586364061
transform 1 0 8464 0 -1 66912
box -38 -48 130 592
use scs8hd_decap_6  FILLER_119_74
timestamp 1586364061
transform 1 0 7912 0 1 66912
box -38 -48 590 592
use scs8hd_fill_1  FILLER_119_80
timestamp 1586364061
transform 1 0 8464 0 1 66912
box -38 -48 130 592
use scs8hd_decap_3  PHY_240
timestamp 1586364061
transform 1 0 1104 0 -1 68000
box -38 -48 314 592
use scs8hd_decap_12  FILLER_120_3
timestamp 1586364061
transform 1 0 1380 0 -1 68000
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_120_15
timestamp 1586364061
transform 1 0 2484 0 -1 68000
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1329
timestamp 1586364061
transform 1 0 3956 0 -1 68000
box -38 -48 130 592
use scs8hd_decap_4  FILLER_120_27
timestamp 1586364061
transform 1 0 3588 0 -1 68000
box -38 -48 406 592
use scs8hd_decap_12  FILLER_120_32
timestamp 1586364061
transform 1 0 4048 0 -1 68000
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_120_44
timestamp 1586364061
transform 1 0 5152 0 -1 68000
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_120_56
timestamp 1586364061
transform 1 0 6256 0 -1 68000
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_120_68
timestamp 1586364061
transform 1 0 7360 0 -1 68000
box -38 -48 1142 592
use scs8hd_decap_3  PHY_241
timestamp 1586364061
transform -1 0 8832 0 -1 68000
box -38 -48 314 592
use scs8hd_fill_1  FILLER_120_80
timestamp 1586364061
transform 1 0 8464 0 -1 68000
box -38 -48 130 592
use scs8hd_decap_3  PHY_242
timestamp 1586364061
transform 1 0 1104 0 1 68000
box -38 -48 314 592
use scs8hd_decap_12  FILLER_121_3
timestamp 1586364061
transform 1 0 1380 0 1 68000
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_121_15
timestamp 1586364061
transform 1 0 2484 0 1 68000
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_121_27
timestamp 1586364061
transform 1 0 3588 0 1 68000
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_121_39
timestamp 1586364061
transform 1 0 4692 0 1 68000
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_121_51
timestamp 1586364061
transform 1 0 5796 0 1 68000
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1330
timestamp 1586364061
transform 1 0 6716 0 1 68000
box -38 -48 130 592
use scs8hd_fill_2  FILLER_121_59
timestamp 1586364061
transform 1 0 6532 0 1 68000
box -38 -48 222 592
use scs8hd_decap_12  FILLER_121_62
timestamp 1586364061
transform 1 0 6808 0 1 68000
box -38 -48 1142 592
use scs8hd_decap_3  PHY_243
timestamp 1586364061
transform -1 0 8832 0 1 68000
box -38 -48 314 592
use scs8hd_decap_6  FILLER_121_74
timestamp 1586364061
transform 1 0 7912 0 1 68000
box -38 -48 590 592
use scs8hd_fill_1  FILLER_121_80
timestamp 1586364061
transform 1 0 8464 0 1 68000
box -38 -48 130 592
use scs8hd_decap_3  PHY_244
timestamp 1586364061
transform 1 0 1104 0 -1 69088
box -38 -48 314 592
use scs8hd_decap_12  FILLER_122_3
timestamp 1586364061
transform 1 0 1380 0 -1 69088
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_122_15
timestamp 1586364061
transform 1 0 2484 0 -1 69088
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1331
timestamp 1586364061
transform 1 0 3956 0 -1 69088
box -38 -48 130 592
use scs8hd_decap_4  FILLER_122_27
timestamp 1586364061
transform 1 0 3588 0 -1 69088
box -38 -48 406 592
use scs8hd_decap_12  FILLER_122_32
timestamp 1586364061
transform 1 0 4048 0 -1 69088
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_122_44
timestamp 1586364061
transform 1 0 5152 0 -1 69088
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_122_56
timestamp 1586364061
transform 1 0 6256 0 -1 69088
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_122_68
timestamp 1586364061
transform 1 0 7360 0 -1 69088
box -38 -48 1142 592
use scs8hd_decap_3  PHY_245
timestamp 1586364061
transform -1 0 8832 0 -1 69088
box -38 -48 314 592
use scs8hd_fill_1  FILLER_122_80
timestamp 1586364061
transform 1 0 8464 0 -1 69088
box -38 -48 130 592
use scs8hd_decap_3  PHY_246
timestamp 1586364061
transform 1 0 1104 0 1 69088
box -38 -48 314 592
use scs8hd_decap_12  FILLER_123_3
timestamp 1586364061
transform 1 0 1380 0 1 69088
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_123_15
timestamp 1586364061
transform 1 0 2484 0 1 69088
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_123_27
timestamp 1586364061
transform 1 0 3588 0 1 69088
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_123_39
timestamp 1586364061
transform 1 0 4692 0 1 69088
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_123_51
timestamp 1586364061
transform 1 0 5796 0 1 69088
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1332
timestamp 1586364061
transform 1 0 6716 0 1 69088
box -38 -48 130 592
use scs8hd_fill_2  FILLER_123_59
timestamp 1586364061
transform 1 0 6532 0 1 69088
box -38 -48 222 592
use scs8hd_decap_12  FILLER_123_62
timestamp 1586364061
transform 1 0 6808 0 1 69088
box -38 -48 1142 592
use scs8hd_decap_3  PHY_247
timestamp 1586364061
transform -1 0 8832 0 1 69088
box -38 -48 314 592
use scs8hd_decap_6  FILLER_123_74
timestamp 1586364061
transform 1 0 7912 0 1 69088
box -38 -48 590 592
use scs8hd_fill_1  FILLER_123_80
timestamp 1586364061
transform 1 0 8464 0 1 69088
box -38 -48 130 592
use scs8hd_decap_3  PHY_248
timestamp 1586364061
transform 1 0 1104 0 -1 70176
box -38 -48 314 592
use scs8hd_decap_12  FILLER_124_3
timestamp 1586364061
transform 1 0 1380 0 -1 70176
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_124_15
timestamp 1586364061
transform 1 0 2484 0 -1 70176
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1333
timestamp 1586364061
transform 1 0 3956 0 -1 70176
box -38 -48 130 592
use scs8hd_decap_4  FILLER_124_27
timestamp 1586364061
transform 1 0 3588 0 -1 70176
box -38 -48 406 592
use scs8hd_decap_12  FILLER_124_32
timestamp 1586364061
transform 1 0 4048 0 -1 70176
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_124_44
timestamp 1586364061
transform 1 0 5152 0 -1 70176
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_124_56
timestamp 1586364061
transform 1 0 6256 0 -1 70176
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_124_68
timestamp 1586364061
transform 1 0 7360 0 -1 70176
box -38 -48 1142 592
use scs8hd_decap_3  PHY_249
timestamp 1586364061
transform -1 0 8832 0 -1 70176
box -38 -48 314 592
use scs8hd_fill_1  FILLER_124_80
timestamp 1586364061
transform 1 0 8464 0 -1 70176
box -38 -48 130 592
use scs8hd_decap_3  PHY_250
timestamp 1586364061
transform 1 0 1104 0 1 70176
box -38 -48 314 592
use scs8hd_decap_3  PHY_252
timestamp 1586364061
transform 1 0 1104 0 -1 71264
box -38 -48 314 592
use scs8hd_decap_12  FILLER_125_3
timestamp 1586364061
transform 1 0 1380 0 1 70176
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_125_15
timestamp 1586364061
transform 1 0 2484 0 1 70176
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_126_3
timestamp 1586364061
transform 1 0 1380 0 -1 71264
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_126_15
timestamp 1586364061
transform 1 0 2484 0 -1 71264
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1335
timestamp 1586364061
transform 1 0 3956 0 -1 71264
box -38 -48 130 592
use scs8hd_decap_12  FILLER_125_27
timestamp 1586364061
transform 1 0 3588 0 1 70176
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_126_27
timestamp 1586364061
transform 1 0 3588 0 -1 71264
box -38 -48 406 592
use scs8hd_decap_12  FILLER_126_32
timestamp 1586364061
transform 1 0 4048 0 -1 71264
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_125_39
timestamp 1586364061
transform 1 0 4692 0 1 70176
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_125_51
timestamp 1586364061
transform 1 0 5796 0 1 70176
box -38 -48 774 592
use scs8hd_decap_12  FILLER_126_44
timestamp 1586364061
transform 1 0 5152 0 -1 71264
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1334
timestamp 1586364061
transform 1 0 6716 0 1 70176
box -38 -48 130 592
use scs8hd_fill_2  FILLER_125_59
timestamp 1586364061
transform 1 0 6532 0 1 70176
box -38 -48 222 592
use scs8hd_decap_12  FILLER_125_62
timestamp 1586364061
transform 1 0 6808 0 1 70176
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_126_56
timestamp 1586364061
transform 1 0 6256 0 -1 71264
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_126_68
timestamp 1586364061
transform 1 0 7360 0 -1 71264
box -38 -48 1142 592
use scs8hd_decap_3  PHY_251
timestamp 1586364061
transform -1 0 8832 0 1 70176
box -38 -48 314 592
use scs8hd_decap_3  PHY_253
timestamp 1586364061
transform -1 0 8832 0 -1 71264
box -38 -48 314 592
use scs8hd_decap_6  FILLER_125_74
timestamp 1586364061
transform 1 0 7912 0 1 70176
box -38 -48 590 592
use scs8hd_fill_1  FILLER_125_80
timestamp 1586364061
transform 1 0 8464 0 1 70176
box -38 -48 130 592
use scs8hd_fill_1  FILLER_126_80
timestamp 1586364061
transform 1 0 8464 0 -1 71264
box -38 -48 130 592
use scs8hd_decap_3  PHY_254
timestamp 1586364061
transform 1 0 1104 0 1 71264
box -38 -48 314 592
use scs8hd_decap_12  FILLER_127_3
timestamp 1586364061
transform 1 0 1380 0 1 71264
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_127_15
timestamp 1586364061
transform 1 0 2484 0 1 71264
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_127_27
timestamp 1586364061
transform 1 0 3588 0 1 71264
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_127_39
timestamp 1586364061
transform 1 0 4692 0 1 71264
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_127_51
timestamp 1586364061
transform 1 0 5796 0 1 71264
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1336
timestamp 1586364061
transform 1 0 6716 0 1 71264
box -38 -48 130 592
use scs8hd_fill_2  FILLER_127_59
timestamp 1586364061
transform 1 0 6532 0 1 71264
box -38 -48 222 592
use scs8hd_decap_12  FILLER_127_62
timestamp 1586364061
transform 1 0 6808 0 1 71264
box -38 -48 1142 592
use scs8hd_decap_3  PHY_255
timestamp 1586364061
transform -1 0 8832 0 1 71264
box -38 -48 314 592
use scs8hd_decap_6  FILLER_127_74
timestamp 1586364061
transform 1 0 7912 0 1 71264
box -38 -48 590 592
use scs8hd_fill_1  FILLER_127_80
timestamp 1586364061
transform 1 0 8464 0 1 71264
box -38 -48 130 592
use scs8hd_decap_3  PHY_256
timestamp 1586364061
transform 1 0 1104 0 -1 72352
box -38 -48 314 592
use scs8hd_decap_12  FILLER_128_3
timestamp 1586364061
transform 1 0 1380 0 -1 72352
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_128_15
timestamp 1586364061
transform 1 0 2484 0 -1 72352
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1337
timestamp 1586364061
transform 1 0 3956 0 -1 72352
box -38 -48 130 592
use scs8hd_decap_4  FILLER_128_27
timestamp 1586364061
transform 1 0 3588 0 -1 72352
box -38 -48 406 592
use scs8hd_decap_12  FILLER_128_32
timestamp 1586364061
transform 1 0 4048 0 -1 72352
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_128_44
timestamp 1586364061
transform 1 0 5152 0 -1 72352
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_128_56
timestamp 1586364061
transform 1 0 6256 0 -1 72352
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_128_68
timestamp 1586364061
transform 1 0 7360 0 -1 72352
box -38 -48 1142 592
use scs8hd_decap_3  PHY_257
timestamp 1586364061
transform -1 0 8832 0 -1 72352
box -38 -48 314 592
use scs8hd_fill_1  FILLER_128_80
timestamp 1586364061
transform 1 0 8464 0 -1 72352
box -38 -48 130 592
use scs8hd_decap_3  PHY_258
timestamp 1586364061
transform 1 0 1104 0 1 72352
box -38 -48 314 592
use scs8hd_decap_12  FILLER_129_3
timestamp 1586364061
transform 1 0 1380 0 1 72352
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_129_15
timestamp 1586364061
transform 1 0 2484 0 1 72352
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_129_27
timestamp 1586364061
transform 1 0 3588 0 1 72352
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_129_39
timestamp 1586364061
transform 1 0 4692 0 1 72352
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_129_51
timestamp 1586364061
transform 1 0 5796 0 1 72352
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1338
timestamp 1586364061
transform 1 0 6716 0 1 72352
box -38 -48 130 592
use scs8hd_fill_2  FILLER_129_59
timestamp 1586364061
transform 1 0 6532 0 1 72352
box -38 -48 222 592
use scs8hd_decap_12  FILLER_129_62
timestamp 1586364061
transform 1 0 6808 0 1 72352
box -38 -48 1142 592
use scs8hd_decap_3  PHY_259
timestamp 1586364061
transform -1 0 8832 0 1 72352
box -38 -48 314 592
use scs8hd_decap_6  FILLER_129_74
timestamp 1586364061
transform 1 0 7912 0 1 72352
box -38 -48 590 592
use scs8hd_fill_1  FILLER_129_80
timestamp 1586364061
transform 1 0 8464 0 1 72352
box -38 -48 130 592
use scs8hd_decap_3  PHY_260
timestamp 1586364061
transform 1 0 1104 0 -1 73440
box -38 -48 314 592
use scs8hd_decap_12  FILLER_130_3
timestamp 1586364061
transform 1 0 1380 0 -1 73440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_130_15
timestamp 1586364061
transform 1 0 2484 0 -1 73440
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1339
timestamp 1586364061
transform 1 0 3956 0 -1 73440
box -38 -48 130 592
use scs8hd_decap_4  FILLER_130_27
timestamp 1586364061
transform 1 0 3588 0 -1 73440
box -38 -48 406 592
use scs8hd_decap_12  FILLER_130_32
timestamp 1586364061
transform 1 0 4048 0 -1 73440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_130_44
timestamp 1586364061
transform 1 0 5152 0 -1 73440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_130_56
timestamp 1586364061
transform 1 0 6256 0 -1 73440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_130_68
timestamp 1586364061
transform 1 0 7360 0 -1 73440
box -38 -48 1142 592
use scs8hd_decap_3  PHY_261
timestamp 1586364061
transform -1 0 8832 0 -1 73440
box -38 -48 314 592
use scs8hd_fill_1  FILLER_130_80
timestamp 1586364061
transform 1 0 8464 0 -1 73440
box -38 -48 130 592
use scs8hd_decap_3  PHY_262
timestamp 1586364061
transform 1 0 1104 0 1 73440
box -38 -48 314 592
use scs8hd_decap_12  FILLER_131_3
timestamp 1586364061
transform 1 0 1380 0 1 73440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_131_15
timestamp 1586364061
transform 1 0 2484 0 1 73440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_131_27
timestamp 1586364061
transform 1 0 3588 0 1 73440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_131_39
timestamp 1586364061
transform 1 0 4692 0 1 73440
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_131_51
timestamp 1586364061
transform 1 0 5796 0 1 73440
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1340
timestamp 1586364061
transform 1 0 6716 0 1 73440
box -38 -48 130 592
use scs8hd_fill_2  FILLER_131_59
timestamp 1586364061
transform 1 0 6532 0 1 73440
box -38 -48 222 592
use scs8hd_decap_12  FILLER_131_62
timestamp 1586364061
transform 1 0 6808 0 1 73440
box -38 -48 1142 592
use scs8hd_decap_3  PHY_263
timestamp 1586364061
transform -1 0 8832 0 1 73440
box -38 -48 314 592
use scs8hd_decap_6  FILLER_131_74
timestamp 1586364061
transform 1 0 7912 0 1 73440
box -38 -48 590 592
use scs8hd_fill_1  FILLER_131_80
timestamp 1586364061
transform 1 0 8464 0 1 73440
box -38 -48 130 592
use scs8hd_decap_3  PHY_264
timestamp 1586364061
transform 1 0 1104 0 -1 74528
box -38 -48 314 592
use scs8hd_decap_3  PHY_266
timestamp 1586364061
transform 1 0 1104 0 1 74528
box -38 -48 314 592
use scs8hd_decap_12  FILLER_132_3
timestamp 1586364061
transform 1 0 1380 0 -1 74528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_132_15
timestamp 1586364061
transform 1 0 2484 0 -1 74528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_133_3
timestamp 1586364061
transform 1 0 1380 0 1 74528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_133_15
timestamp 1586364061
transform 1 0 2484 0 1 74528
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1341
timestamp 1586364061
transform 1 0 3956 0 -1 74528
box -38 -48 130 592
use scs8hd_decap_4  FILLER_132_27
timestamp 1586364061
transform 1 0 3588 0 -1 74528
box -38 -48 406 592
use scs8hd_decap_12  FILLER_132_32
timestamp 1586364061
transform 1 0 4048 0 -1 74528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_133_27
timestamp 1586364061
transform 1 0 3588 0 1 74528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_132_44
timestamp 1586364061
transform 1 0 5152 0 -1 74528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_133_39
timestamp 1586364061
transform 1 0 4692 0 1 74528
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_133_51
timestamp 1586364061
transform 1 0 5796 0 1 74528
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1342
timestamp 1586364061
transform 1 0 6716 0 1 74528
box -38 -48 130 592
use scs8hd_decap_12  FILLER_132_56
timestamp 1586364061
transform 1 0 6256 0 -1 74528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_132_68
timestamp 1586364061
transform 1 0 7360 0 -1 74528
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_133_59
timestamp 1586364061
transform 1 0 6532 0 1 74528
box -38 -48 222 592
use scs8hd_decap_12  FILLER_133_62
timestamp 1586364061
transform 1 0 6808 0 1 74528
box -38 -48 1142 592
use scs8hd_decap_3  PHY_265
timestamp 1586364061
transform -1 0 8832 0 -1 74528
box -38 -48 314 592
use scs8hd_decap_3  PHY_267
timestamp 1586364061
transform -1 0 8832 0 1 74528
box -38 -48 314 592
use scs8hd_fill_1  FILLER_132_80
timestamp 1586364061
transform 1 0 8464 0 -1 74528
box -38 -48 130 592
use scs8hd_decap_6  FILLER_133_74
timestamp 1586364061
transform 1 0 7912 0 1 74528
box -38 -48 590 592
use scs8hd_fill_1  FILLER_133_80
timestamp 1586364061
transform 1 0 8464 0 1 74528
box -38 -48 130 592
use scs8hd_decap_3  PHY_268
timestamp 1586364061
transform 1 0 1104 0 -1 75616
box -38 -48 314 592
use scs8hd_decap_12  FILLER_134_3
timestamp 1586364061
transform 1 0 1380 0 -1 75616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_134_15
timestamp 1586364061
transform 1 0 2484 0 -1 75616
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1343
timestamp 1586364061
transform 1 0 3956 0 -1 75616
box -38 -48 130 592
use scs8hd_decap_4  FILLER_134_27
timestamp 1586364061
transform 1 0 3588 0 -1 75616
box -38 -48 406 592
use scs8hd_decap_12  FILLER_134_32
timestamp 1586364061
transform 1 0 4048 0 -1 75616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_134_44
timestamp 1586364061
transform 1 0 5152 0 -1 75616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_134_56
timestamp 1586364061
transform 1 0 6256 0 -1 75616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_134_68
timestamp 1586364061
transform 1 0 7360 0 -1 75616
box -38 -48 1142 592
use scs8hd_decap_3  PHY_269
timestamp 1586364061
transform -1 0 8832 0 -1 75616
box -38 -48 314 592
use scs8hd_fill_1  FILLER_134_80
timestamp 1586364061
transform 1 0 8464 0 -1 75616
box -38 -48 130 592
use scs8hd_decap_3  PHY_270
timestamp 1586364061
transform 1 0 1104 0 1 75616
box -38 -48 314 592
use scs8hd_decap_12  FILLER_135_3
timestamp 1586364061
transform 1 0 1380 0 1 75616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_135_15
timestamp 1586364061
transform 1 0 2484 0 1 75616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_135_27
timestamp 1586364061
transform 1 0 3588 0 1 75616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_135_39
timestamp 1586364061
transform 1 0 4692 0 1 75616
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_135_51
timestamp 1586364061
transform 1 0 5796 0 1 75616
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1344
timestamp 1586364061
transform 1 0 6716 0 1 75616
box -38 -48 130 592
use scs8hd_fill_2  FILLER_135_59
timestamp 1586364061
transform 1 0 6532 0 1 75616
box -38 -48 222 592
use scs8hd_decap_12  FILLER_135_62
timestamp 1586364061
transform 1 0 6808 0 1 75616
box -38 -48 1142 592
use scs8hd_decap_3  PHY_271
timestamp 1586364061
transform -1 0 8832 0 1 75616
box -38 -48 314 592
use scs8hd_decap_6  FILLER_135_74
timestamp 1586364061
transform 1 0 7912 0 1 75616
box -38 -48 590 592
use scs8hd_fill_1  FILLER_135_80
timestamp 1586364061
transform 1 0 8464 0 1 75616
box -38 -48 130 592
use scs8hd_decap_3  PHY_272
timestamp 1586364061
transform 1 0 1104 0 -1 76704
box -38 -48 314 592
use scs8hd_decap_12  FILLER_136_3
timestamp 1586364061
transform 1 0 1380 0 -1 76704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_136_15
timestamp 1586364061
transform 1 0 2484 0 -1 76704
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1345
timestamp 1586364061
transform 1 0 3956 0 -1 76704
box -38 -48 130 592
use scs8hd_decap_4  FILLER_136_27
timestamp 1586364061
transform 1 0 3588 0 -1 76704
box -38 -48 406 592
use scs8hd_decap_12  FILLER_136_32
timestamp 1586364061
transform 1 0 4048 0 -1 76704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_136_44
timestamp 1586364061
transform 1 0 5152 0 -1 76704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_136_56
timestamp 1586364061
transform 1 0 6256 0 -1 76704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_136_68
timestamp 1586364061
transform 1 0 7360 0 -1 76704
box -38 -48 1142 592
use scs8hd_decap_3  PHY_273
timestamp 1586364061
transform -1 0 8832 0 -1 76704
box -38 -48 314 592
use scs8hd_fill_1  FILLER_136_80
timestamp 1586364061
transform 1 0 8464 0 -1 76704
box -38 -48 130 592
use scs8hd_decap_3  PHY_274
timestamp 1586364061
transform 1 0 1104 0 1 76704
box -38 -48 314 592
use scs8hd_decap_12  FILLER_137_3
timestamp 1586364061
transform 1 0 1380 0 1 76704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_137_15
timestamp 1586364061
transform 1 0 2484 0 1 76704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_137_27
timestamp 1586364061
transform 1 0 3588 0 1 76704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_137_39
timestamp 1586364061
transform 1 0 4692 0 1 76704
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_137_51
timestamp 1586364061
transform 1 0 5796 0 1 76704
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1346
timestamp 1586364061
transform 1 0 6716 0 1 76704
box -38 -48 130 592
use scs8hd_fill_2  FILLER_137_59
timestamp 1586364061
transform 1 0 6532 0 1 76704
box -38 -48 222 592
use scs8hd_decap_12  FILLER_137_62
timestamp 1586364061
transform 1 0 6808 0 1 76704
box -38 -48 1142 592
use scs8hd_decap_3  PHY_275
timestamp 1586364061
transform -1 0 8832 0 1 76704
box -38 -48 314 592
use scs8hd_decap_6  FILLER_137_74
timestamp 1586364061
transform 1 0 7912 0 1 76704
box -38 -48 590 592
use scs8hd_fill_1  FILLER_137_80
timestamp 1586364061
transform 1 0 8464 0 1 76704
box -38 -48 130 592
use scs8hd_decap_3  PHY_276
timestamp 1586364061
transform 1 0 1104 0 -1 77792
box -38 -48 314 592
use scs8hd_decap_3  PHY_278
timestamp 1586364061
transform 1 0 1104 0 1 77792
box -38 -48 314 592
use scs8hd_decap_12  FILLER_138_3
timestamp 1586364061
transform 1 0 1380 0 -1 77792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_138_15
timestamp 1586364061
transform 1 0 2484 0 -1 77792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_139_3
timestamp 1586364061
transform 1 0 1380 0 1 77792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_139_15
timestamp 1586364061
transform 1 0 2484 0 1 77792
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1347
timestamp 1586364061
transform 1 0 3956 0 -1 77792
box -38 -48 130 592
use scs8hd_decap_4  FILLER_138_27
timestamp 1586364061
transform 1 0 3588 0 -1 77792
box -38 -48 406 592
use scs8hd_decap_12  FILLER_138_32
timestamp 1586364061
transform 1 0 4048 0 -1 77792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_139_27
timestamp 1586364061
transform 1 0 3588 0 1 77792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_138_44
timestamp 1586364061
transform 1 0 5152 0 -1 77792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_139_39
timestamp 1586364061
transform 1 0 4692 0 1 77792
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_139_51
timestamp 1586364061
transform 1 0 5796 0 1 77792
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1348
timestamp 1586364061
transform 1 0 6716 0 1 77792
box -38 -48 130 592
use scs8hd_decap_12  FILLER_138_56
timestamp 1586364061
transform 1 0 6256 0 -1 77792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_138_68
timestamp 1586364061
transform 1 0 7360 0 -1 77792
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_139_59
timestamp 1586364061
transform 1 0 6532 0 1 77792
box -38 -48 222 592
use scs8hd_decap_12  FILLER_139_62
timestamp 1586364061
transform 1 0 6808 0 1 77792
box -38 -48 1142 592
use scs8hd_decap_3  PHY_277
timestamp 1586364061
transform -1 0 8832 0 -1 77792
box -38 -48 314 592
use scs8hd_decap_3  PHY_279
timestamp 1586364061
transform -1 0 8832 0 1 77792
box -38 -48 314 592
use scs8hd_fill_1  FILLER_138_80
timestamp 1586364061
transform 1 0 8464 0 -1 77792
box -38 -48 130 592
use scs8hd_decap_6  FILLER_139_74
timestamp 1586364061
transform 1 0 7912 0 1 77792
box -38 -48 590 592
use scs8hd_fill_1  FILLER_139_80
timestamp 1586364061
transform 1 0 8464 0 1 77792
box -38 -48 130 592
use scs8hd_decap_3  PHY_280
timestamp 1586364061
transform 1 0 1104 0 -1 78880
box -38 -48 314 592
use scs8hd_decap_12  FILLER_140_3
timestamp 1586364061
transform 1 0 1380 0 -1 78880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_140_15
timestamp 1586364061
transform 1 0 2484 0 -1 78880
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1349
timestamp 1586364061
transform 1 0 3956 0 -1 78880
box -38 -48 130 592
use scs8hd_decap_4  FILLER_140_27
timestamp 1586364061
transform 1 0 3588 0 -1 78880
box -38 -48 406 592
use scs8hd_decap_12  FILLER_140_32
timestamp 1586364061
transform 1 0 4048 0 -1 78880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_140_44
timestamp 1586364061
transform 1 0 5152 0 -1 78880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_140_56
timestamp 1586364061
transform 1 0 6256 0 -1 78880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_140_68
timestamp 1586364061
transform 1 0 7360 0 -1 78880
box -38 -48 1142 592
use scs8hd_decap_3  PHY_281
timestamp 1586364061
transform -1 0 8832 0 -1 78880
box -38 -48 314 592
use scs8hd_fill_1  FILLER_140_80
timestamp 1586364061
transform 1 0 8464 0 -1 78880
box -38 -48 130 592
use scs8hd_decap_3  PHY_282
timestamp 1586364061
transform 1 0 1104 0 1 78880
box -38 -48 314 592
use scs8hd_decap_12  FILLER_141_3
timestamp 1586364061
transform 1 0 1380 0 1 78880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_141_15
timestamp 1586364061
transform 1 0 2484 0 1 78880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_141_27
timestamp 1586364061
transform 1 0 3588 0 1 78880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_141_39
timestamp 1586364061
transform 1 0 4692 0 1 78880
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_141_51
timestamp 1586364061
transform 1 0 5796 0 1 78880
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1350
timestamp 1586364061
transform 1 0 6716 0 1 78880
box -38 -48 130 592
use scs8hd_fill_2  FILLER_141_59
timestamp 1586364061
transform 1 0 6532 0 1 78880
box -38 -48 222 592
use scs8hd_decap_12  FILLER_141_62
timestamp 1586364061
transform 1 0 6808 0 1 78880
box -38 -48 1142 592
use scs8hd_decap_3  PHY_283
timestamp 1586364061
transform -1 0 8832 0 1 78880
box -38 -48 314 592
use scs8hd_decap_6  FILLER_141_74
timestamp 1586364061
transform 1 0 7912 0 1 78880
box -38 -48 590 592
use scs8hd_fill_1  FILLER_141_80
timestamp 1586364061
transform 1 0 8464 0 1 78880
box -38 -48 130 592
use scs8hd_decap_3  PHY_284
timestamp 1586364061
transform 1 0 1104 0 -1 79968
box -38 -48 314 592
use scs8hd_decap_12  FILLER_142_3
timestamp 1586364061
transform 1 0 1380 0 -1 79968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_142_15
timestamp 1586364061
transform 1 0 2484 0 -1 79968
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1351
timestamp 1586364061
transform 1 0 3956 0 -1 79968
box -38 -48 130 592
use scs8hd_decap_4  FILLER_142_27
timestamp 1586364061
transform 1 0 3588 0 -1 79968
box -38 -48 406 592
use scs8hd_decap_12  FILLER_142_32
timestamp 1586364061
transform 1 0 4048 0 -1 79968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_142_44
timestamp 1586364061
transform 1 0 5152 0 -1 79968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_142_56
timestamp 1586364061
transform 1 0 6256 0 -1 79968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_142_68
timestamp 1586364061
transform 1 0 7360 0 -1 79968
box -38 -48 1142 592
use scs8hd_decap_3  PHY_285
timestamp 1586364061
transform -1 0 8832 0 -1 79968
box -38 -48 314 592
use scs8hd_fill_1  FILLER_142_80
timestamp 1586364061
transform 1 0 8464 0 -1 79968
box -38 -48 130 592
use scs8hd_decap_3  PHY_286
timestamp 1586364061
transform 1 0 1104 0 1 79968
box -38 -48 314 592
use scs8hd_decap_12  FILLER_143_3
timestamp 1586364061
transform 1 0 1380 0 1 79968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_143_15
timestamp 1586364061
transform 1 0 2484 0 1 79968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_143_27
timestamp 1586364061
transform 1 0 3588 0 1 79968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_143_39
timestamp 1586364061
transform 1 0 4692 0 1 79968
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_143_51
timestamp 1586364061
transform 1 0 5796 0 1 79968
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1352
timestamp 1586364061
transform 1 0 6716 0 1 79968
box -38 -48 130 592
use scs8hd_fill_2  FILLER_143_59
timestamp 1586364061
transform 1 0 6532 0 1 79968
box -38 -48 222 592
use scs8hd_decap_12  FILLER_143_62
timestamp 1586364061
transform 1 0 6808 0 1 79968
box -38 -48 1142 592
use scs8hd_decap_3  PHY_287
timestamp 1586364061
transform -1 0 8832 0 1 79968
box -38 -48 314 592
use scs8hd_decap_6  FILLER_143_74
timestamp 1586364061
transform 1 0 7912 0 1 79968
box -38 -48 590 592
use scs8hd_fill_1  FILLER_143_80
timestamp 1586364061
transform 1 0 8464 0 1 79968
box -38 -48 130 592
use scs8hd_decap_3  PHY_288
timestamp 1586364061
transform 1 0 1104 0 -1 81056
box -38 -48 314 592
use scs8hd_decap_12  FILLER_144_3
timestamp 1586364061
transform 1 0 1380 0 -1 81056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_144_15
timestamp 1586364061
transform 1 0 2484 0 -1 81056
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1353
timestamp 1586364061
transform 1 0 3956 0 -1 81056
box -38 -48 130 592
use scs8hd_decap_4  FILLER_144_27
timestamp 1586364061
transform 1 0 3588 0 -1 81056
box -38 -48 406 592
use scs8hd_decap_12  FILLER_144_32
timestamp 1586364061
transform 1 0 4048 0 -1 81056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_144_44
timestamp 1586364061
transform 1 0 5152 0 -1 81056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_144_56
timestamp 1586364061
transform 1 0 6256 0 -1 81056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_144_68
timestamp 1586364061
transform 1 0 7360 0 -1 81056
box -38 -48 1142 592
use scs8hd_decap_3  PHY_289
timestamp 1586364061
transform -1 0 8832 0 -1 81056
box -38 -48 314 592
use scs8hd_fill_1  FILLER_144_80
timestamp 1586364061
transform 1 0 8464 0 -1 81056
box -38 -48 130 592
use scs8hd_decap_3  PHY_290
timestamp 1586364061
transform 1 0 1104 0 1 81056
box -38 -48 314 592
use scs8hd_decap_3  PHY_292
timestamp 1586364061
transform 1 0 1104 0 -1 82144
box -38 -48 314 592
use scs8hd_decap_12  FILLER_145_3
timestamp 1586364061
transform 1 0 1380 0 1 81056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_145_15
timestamp 1586364061
transform 1 0 2484 0 1 81056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_146_3
timestamp 1586364061
transform 1 0 1380 0 -1 82144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_146_15
timestamp 1586364061
transform 1 0 2484 0 -1 82144
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1355
timestamp 1586364061
transform 1 0 3956 0 -1 82144
box -38 -48 130 592
use scs8hd_decap_12  FILLER_145_27
timestamp 1586364061
transform 1 0 3588 0 1 81056
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_146_27
timestamp 1586364061
transform 1 0 3588 0 -1 82144
box -38 -48 406 592
use scs8hd_decap_12  FILLER_146_32
timestamp 1586364061
transform 1 0 4048 0 -1 82144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_145_39
timestamp 1586364061
transform 1 0 4692 0 1 81056
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_145_51
timestamp 1586364061
transform 1 0 5796 0 1 81056
box -38 -48 774 592
use scs8hd_decap_12  FILLER_146_44
timestamp 1586364061
transform 1 0 5152 0 -1 82144
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1354
timestamp 1586364061
transform 1 0 6716 0 1 81056
box -38 -48 130 592
use scs8hd_fill_2  FILLER_145_59
timestamp 1586364061
transform 1 0 6532 0 1 81056
box -38 -48 222 592
use scs8hd_decap_12  FILLER_145_62
timestamp 1586364061
transform 1 0 6808 0 1 81056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_146_56
timestamp 1586364061
transform 1 0 6256 0 -1 82144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_146_68
timestamp 1586364061
transform 1 0 7360 0 -1 82144
box -38 -48 1142 592
use scs8hd_decap_3  PHY_291
timestamp 1586364061
transform -1 0 8832 0 1 81056
box -38 -48 314 592
use scs8hd_decap_3  PHY_293
timestamp 1586364061
transform -1 0 8832 0 -1 82144
box -38 -48 314 592
use scs8hd_decap_6  FILLER_145_74
timestamp 1586364061
transform 1 0 7912 0 1 81056
box -38 -48 590 592
use scs8hd_fill_1  FILLER_145_80
timestamp 1586364061
transform 1 0 8464 0 1 81056
box -38 -48 130 592
use scs8hd_fill_1  FILLER_146_80
timestamp 1586364061
transform 1 0 8464 0 -1 82144
box -38 -48 130 592
use scs8hd_decap_3  PHY_294
timestamp 1586364061
transform 1 0 1104 0 1 82144
box -38 -48 314 592
use scs8hd_decap_12  FILLER_147_3
timestamp 1586364061
transform 1 0 1380 0 1 82144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_147_15
timestamp 1586364061
transform 1 0 2484 0 1 82144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_147_27
timestamp 1586364061
transform 1 0 3588 0 1 82144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_147_39
timestamp 1586364061
transform 1 0 4692 0 1 82144
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_147_51
timestamp 1586364061
transform 1 0 5796 0 1 82144
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1356
timestamp 1586364061
transform 1 0 6716 0 1 82144
box -38 -48 130 592
use scs8hd_fill_2  FILLER_147_59
timestamp 1586364061
transform 1 0 6532 0 1 82144
box -38 -48 222 592
use scs8hd_decap_12  FILLER_147_62
timestamp 1586364061
transform 1 0 6808 0 1 82144
box -38 -48 1142 592
use scs8hd_decap_3  PHY_295
timestamp 1586364061
transform -1 0 8832 0 1 82144
box -38 -48 314 592
use scs8hd_decap_6  FILLER_147_74
timestamp 1586364061
transform 1 0 7912 0 1 82144
box -38 -48 590 592
use scs8hd_fill_1  FILLER_147_80
timestamp 1586364061
transform 1 0 8464 0 1 82144
box -38 -48 130 592
use scs8hd_decap_3  PHY_296
timestamp 1586364061
transform 1 0 1104 0 -1 83232
box -38 -48 314 592
use scs8hd_decap_12  FILLER_148_3
timestamp 1586364061
transform 1 0 1380 0 -1 83232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_148_15
timestamp 1586364061
transform 1 0 2484 0 -1 83232
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1357
timestamp 1586364061
transform 1 0 3956 0 -1 83232
box -38 -48 130 592
use scs8hd_decap_4  FILLER_148_27
timestamp 1586364061
transform 1 0 3588 0 -1 83232
box -38 -48 406 592
use scs8hd_decap_12  FILLER_148_32
timestamp 1586364061
transform 1 0 4048 0 -1 83232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_148_44
timestamp 1586364061
transform 1 0 5152 0 -1 83232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_148_56
timestamp 1586364061
transform 1 0 6256 0 -1 83232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_148_68
timestamp 1586364061
transform 1 0 7360 0 -1 83232
box -38 -48 1142 592
use scs8hd_decap_3  PHY_297
timestamp 1586364061
transform -1 0 8832 0 -1 83232
box -38 -48 314 592
use scs8hd_fill_1  FILLER_148_80
timestamp 1586364061
transform 1 0 8464 0 -1 83232
box -38 -48 130 592
use scs8hd_decap_3  PHY_298
timestamp 1586364061
transform 1 0 1104 0 1 83232
box -38 -48 314 592
use scs8hd_decap_12  FILLER_149_3
timestamp 1586364061
transform 1 0 1380 0 1 83232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_149_15
timestamp 1586364061
transform 1 0 2484 0 1 83232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_149_27
timestamp 1586364061
transform 1 0 3588 0 1 83232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_149_39
timestamp 1586364061
transform 1 0 4692 0 1 83232
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_149_51
timestamp 1586364061
transform 1 0 5796 0 1 83232
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1358
timestamp 1586364061
transform 1 0 6716 0 1 83232
box -38 -48 130 592
use scs8hd_fill_2  FILLER_149_59
timestamp 1586364061
transform 1 0 6532 0 1 83232
box -38 -48 222 592
use scs8hd_decap_12  FILLER_149_62
timestamp 1586364061
transform 1 0 6808 0 1 83232
box -38 -48 1142 592
use scs8hd_decap_3  PHY_299
timestamp 1586364061
transform -1 0 8832 0 1 83232
box -38 -48 314 592
use scs8hd_decap_6  FILLER_149_74
timestamp 1586364061
transform 1 0 7912 0 1 83232
box -38 -48 590 592
use scs8hd_fill_1  FILLER_149_80
timestamp 1586364061
transform 1 0 8464 0 1 83232
box -38 -48 130 592
use scs8hd_decap_3  PHY_300
timestamp 1586364061
transform 1 0 1104 0 -1 84320
box -38 -48 314 592
use scs8hd_decap_12  FILLER_150_3
timestamp 1586364061
transform 1 0 1380 0 -1 84320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_150_15
timestamp 1586364061
transform 1 0 2484 0 -1 84320
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1359
timestamp 1586364061
transform 1 0 3956 0 -1 84320
box -38 -48 130 592
use scs8hd_decap_4  FILLER_150_27
timestamp 1586364061
transform 1 0 3588 0 -1 84320
box -38 -48 406 592
use scs8hd_decap_12  FILLER_150_32
timestamp 1586364061
transform 1 0 4048 0 -1 84320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_150_44
timestamp 1586364061
transform 1 0 5152 0 -1 84320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_150_56
timestamp 1586364061
transform 1 0 6256 0 -1 84320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_150_68
timestamp 1586364061
transform 1 0 7360 0 -1 84320
box -38 -48 1142 592
use scs8hd_decap_3  PHY_301
timestamp 1586364061
transform -1 0 8832 0 -1 84320
box -38 -48 314 592
use scs8hd_fill_1  FILLER_150_80
timestamp 1586364061
transform 1 0 8464 0 -1 84320
box -38 -48 130 592
use scs8hd_decap_3  PHY_302
timestamp 1586364061
transform 1 0 1104 0 1 84320
box -38 -48 314 592
use scs8hd_decap_3  PHY_304
timestamp 1586364061
transform 1 0 1104 0 -1 85408
box -38 -48 314 592
use scs8hd_decap_12  FILLER_151_3
timestamp 1586364061
transform 1 0 1380 0 1 84320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_151_15
timestamp 1586364061
transform 1 0 2484 0 1 84320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_152_3
timestamp 1586364061
transform 1 0 1380 0 -1 85408
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_152_15
timestamp 1586364061
transform 1 0 2484 0 -1 85408
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1361
timestamp 1586364061
transform 1 0 3956 0 -1 85408
box -38 -48 130 592
use scs8hd_decap_12  FILLER_151_27
timestamp 1586364061
transform 1 0 3588 0 1 84320
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_152_27
timestamp 1586364061
transform 1 0 3588 0 -1 85408
box -38 -48 406 592
use scs8hd_decap_12  FILLER_152_32
timestamp 1586364061
transform 1 0 4048 0 -1 85408
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_151_39
timestamp 1586364061
transform 1 0 4692 0 1 84320
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_151_51
timestamp 1586364061
transform 1 0 5796 0 1 84320
box -38 -48 774 592
use scs8hd_decap_12  FILLER_152_44
timestamp 1586364061
transform 1 0 5152 0 -1 85408
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1360
timestamp 1586364061
transform 1 0 6716 0 1 84320
box -38 -48 130 592
use scs8hd_fill_2  FILLER_151_59
timestamp 1586364061
transform 1 0 6532 0 1 84320
box -38 -48 222 592
use scs8hd_decap_12  FILLER_151_62
timestamp 1586364061
transform 1 0 6808 0 1 84320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_152_56
timestamp 1586364061
transform 1 0 6256 0 -1 85408
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_152_68
timestamp 1586364061
transform 1 0 7360 0 -1 85408
box -38 -48 1142 592
use scs8hd_decap_3  PHY_303
timestamp 1586364061
transform -1 0 8832 0 1 84320
box -38 -48 314 592
use scs8hd_decap_3  PHY_305
timestamp 1586364061
transform -1 0 8832 0 -1 85408
box -38 -48 314 592
use scs8hd_decap_6  FILLER_151_74
timestamp 1586364061
transform 1 0 7912 0 1 84320
box -38 -48 590 592
use scs8hd_fill_1  FILLER_151_80
timestamp 1586364061
transform 1 0 8464 0 1 84320
box -38 -48 130 592
use scs8hd_fill_1  FILLER_152_80
timestamp 1586364061
transform 1 0 8464 0 -1 85408
box -38 -48 130 592
use scs8hd_decap_3  PHY_306
timestamp 1586364061
transform 1 0 1104 0 1 85408
box -38 -48 314 592
use scs8hd_decap_12  FILLER_153_3
timestamp 1586364061
transform 1 0 1380 0 1 85408
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_153_15
timestamp 1586364061
transform 1 0 2484 0 1 85408
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_153_27
timestamp 1586364061
transform 1 0 3588 0 1 85408
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_153_39
timestamp 1586364061
transform 1 0 4692 0 1 85408
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_153_51
timestamp 1586364061
transform 1 0 5796 0 1 85408
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1362
timestamp 1586364061
transform 1 0 6716 0 1 85408
box -38 -48 130 592
use scs8hd_fill_2  FILLER_153_59
timestamp 1586364061
transform 1 0 6532 0 1 85408
box -38 -48 222 592
use scs8hd_decap_12  FILLER_153_62
timestamp 1586364061
transform 1 0 6808 0 1 85408
box -38 -48 1142 592
use scs8hd_decap_3  PHY_307
timestamp 1586364061
transform -1 0 8832 0 1 85408
box -38 -48 314 592
use scs8hd_decap_6  FILLER_153_74
timestamp 1586364061
transform 1 0 7912 0 1 85408
box -38 -48 590 592
use scs8hd_fill_1  FILLER_153_80
timestamp 1586364061
transform 1 0 8464 0 1 85408
box -38 -48 130 592
use scs8hd_decap_3  PHY_308
timestamp 1586364061
transform 1 0 1104 0 -1 86496
box -38 -48 314 592
use scs8hd_decap_12  FILLER_154_3
timestamp 1586364061
transform 1 0 1380 0 -1 86496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_154_15
timestamp 1586364061
transform 1 0 2484 0 -1 86496
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1363
timestamp 1586364061
transform 1 0 3956 0 -1 86496
box -38 -48 130 592
use scs8hd_decap_4  FILLER_154_27
timestamp 1586364061
transform 1 0 3588 0 -1 86496
box -38 -48 406 592
use scs8hd_decap_12  FILLER_154_32
timestamp 1586364061
transform 1 0 4048 0 -1 86496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_154_44
timestamp 1586364061
transform 1 0 5152 0 -1 86496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_154_56
timestamp 1586364061
transform 1 0 6256 0 -1 86496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_154_68
timestamp 1586364061
transform 1 0 7360 0 -1 86496
box -38 -48 1142 592
use scs8hd_decap_3  PHY_309
timestamp 1586364061
transform -1 0 8832 0 -1 86496
box -38 -48 314 592
use scs8hd_fill_1  FILLER_154_80
timestamp 1586364061
transform 1 0 8464 0 -1 86496
box -38 -48 130 592
use scs8hd_decap_3  PHY_310
timestamp 1586364061
transform 1 0 1104 0 1 86496
box -38 -48 314 592
use scs8hd_decap_12  FILLER_155_3
timestamp 1586364061
transform 1 0 1380 0 1 86496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_155_15
timestamp 1586364061
transform 1 0 2484 0 1 86496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_155_27
timestamp 1586364061
transform 1 0 3588 0 1 86496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_155_39
timestamp 1586364061
transform 1 0 4692 0 1 86496
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_155_51
timestamp 1586364061
transform 1 0 5796 0 1 86496
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1364
timestamp 1586364061
transform 1 0 6716 0 1 86496
box -38 -48 130 592
use scs8hd_fill_2  FILLER_155_59
timestamp 1586364061
transform 1 0 6532 0 1 86496
box -38 -48 222 592
use scs8hd_decap_12  FILLER_155_62
timestamp 1586364061
transform 1 0 6808 0 1 86496
box -38 -48 1142 592
use scs8hd_decap_3  PHY_311
timestamp 1586364061
transform -1 0 8832 0 1 86496
box -38 -48 314 592
use scs8hd_decap_6  FILLER_155_74
timestamp 1586364061
transform 1 0 7912 0 1 86496
box -38 -48 590 592
use scs8hd_fill_1  FILLER_155_80
timestamp 1586364061
transform 1 0 8464 0 1 86496
box -38 -48 130 592
use scs8hd_decap_3  PHY_312
timestamp 1586364061
transform 1 0 1104 0 -1 87584
box -38 -48 314 592
use scs8hd_decap_12  FILLER_156_3
timestamp 1586364061
transform 1 0 1380 0 -1 87584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_156_15
timestamp 1586364061
transform 1 0 2484 0 -1 87584
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1365
timestamp 1586364061
transform 1 0 3956 0 -1 87584
box -38 -48 130 592
use scs8hd_decap_4  FILLER_156_27
timestamp 1586364061
transform 1 0 3588 0 -1 87584
box -38 -48 406 592
use scs8hd_decap_12  FILLER_156_32
timestamp 1586364061
transform 1 0 4048 0 -1 87584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_156_44
timestamp 1586364061
transform 1 0 5152 0 -1 87584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_156_56
timestamp 1586364061
transform 1 0 6256 0 -1 87584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_156_68
timestamp 1586364061
transform 1 0 7360 0 -1 87584
box -38 -48 1142 592
use scs8hd_decap_3  PHY_313
timestamp 1586364061
transform -1 0 8832 0 -1 87584
box -38 -48 314 592
use scs8hd_fill_1  FILLER_156_80
timestamp 1586364061
transform 1 0 8464 0 -1 87584
box -38 -48 130 592
use scs8hd_decap_3  PHY_314
timestamp 1586364061
transform 1 0 1104 0 1 87584
box -38 -48 314 592
use scs8hd_decap_12  FILLER_157_3
timestamp 1586364061
transform 1 0 1380 0 1 87584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_157_15
timestamp 1586364061
transform 1 0 2484 0 1 87584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_157_27
timestamp 1586364061
transform 1 0 3588 0 1 87584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_157_39
timestamp 1586364061
transform 1 0 4692 0 1 87584
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_157_51
timestamp 1586364061
transform 1 0 5796 0 1 87584
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1366
timestamp 1586364061
transform 1 0 6716 0 1 87584
box -38 -48 130 592
use scs8hd_fill_2  FILLER_157_59
timestamp 1586364061
transform 1 0 6532 0 1 87584
box -38 -48 222 592
use scs8hd_decap_12  FILLER_157_62
timestamp 1586364061
transform 1 0 6808 0 1 87584
box -38 -48 1142 592
use scs8hd_decap_3  PHY_315
timestamp 1586364061
transform -1 0 8832 0 1 87584
box -38 -48 314 592
use scs8hd_decap_6  FILLER_157_74
timestamp 1586364061
transform 1 0 7912 0 1 87584
box -38 -48 590 592
use scs8hd_fill_1  FILLER_157_80
timestamp 1586364061
transform 1 0 8464 0 1 87584
box -38 -48 130 592
use scs8hd_decap_3  PHY_316
timestamp 1586364061
transform 1 0 1104 0 -1 88672
box -38 -48 314 592
use scs8hd_decap_3  PHY_318
timestamp 1586364061
transform 1 0 1104 0 1 88672
box -38 -48 314 592
use scs8hd_decap_12  FILLER_158_3
timestamp 1586364061
transform 1 0 1380 0 -1 88672
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_158_15
timestamp 1586364061
transform 1 0 2484 0 -1 88672
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_159_3
timestamp 1586364061
transform 1 0 1380 0 1 88672
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_159_15
timestamp 1586364061
transform 1 0 2484 0 1 88672
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1367
timestamp 1586364061
transform 1 0 3956 0 -1 88672
box -38 -48 130 592
use scs8hd_decap_4  FILLER_158_27
timestamp 1586364061
transform 1 0 3588 0 -1 88672
box -38 -48 406 592
use scs8hd_decap_12  FILLER_158_32
timestamp 1586364061
transform 1 0 4048 0 -1 88672
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_159_27
timestamp 1586364061
transform 1 0 3588 0 1 88672
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_158_44
timestamp 1586364061
transform 1 0 5152 0 -1 88672
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_159_39
timestamp 1586364061
transform 1 0 4692 0 1 88672
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_159_51
timestamp 1586364061
transform 1 0 5796 0 1 88672
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1368
timestamp 1586364061
transform 1 0 6716 0 1 88672
box -38 -48 130 592
use scs8hd_decap_12  FILLER_158_56
timestamp 1586364061
transform 1 0 6256 0 -1 88672
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_158_68
timestamp 1586364061
transform 1 0 7360 0 -1 88672
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_159_59
timestamp 1586364061
transform 1 0 6532 0 1 88672
box -38 -48 222 592
use scs8hd_decap_12  FILLER_159_62
timestamp 1586364061
transform 1 0 6808 0 1 88672
box -38 -48 1142 592
use scs8hd_decap_3  PHY_317
timestamp 1586364061
transform -1 0 8832 0 -1 88672
box -38 -48 314 592
use scs8hd_decap_3  PHY_319
timestamp 1586364061
transform -1 0 8832 0 1 88672
box -38 -48 314 592
use scs8hd_fill_1  FILLER_158_80
timestamp 1586364061
transform 1 0 8464 0 -1 88672
box -38 -48 130 592
use scs8hd_decap_6  FILLER_159_74
timestamp 1586364061
transform 1 0 7912 0 1 88672
box -38 -48 590 592
use scs8hd_fill_1  FILLER_159_80
timestamp 1586364061
transform 1 0 8464 0 1 88672
box -38 -48 130 592
use scs8hd_decap_3  PHY_320
timestamp 1586364061
transform 1 0 1104 0 -1 89760
box -38 -48 314 592
use scs8hd_decap_12  FILLER_160_3
timestamp 1586364061
transform 1 0 1380 0 -1 89760
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_160_15
timestamp 1586364061
transform 1 0 2484 0 -1 89760
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1369
timestamp 1586364061
transform 1 0 3956 0 -1 89760
box -38 -48 130 592
use scs8hd_decap_4  FILLER_160_27
timestamp 1586364061
transform 1 0 3588 0 -1 89760
box -38 -48 406 592
use scs8hd_decap_12  FILLER_160_32
timestamp 1586364061
transform 1 0 4048 0 -1 89760
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_160_44
timestamp 1586364061
transform 1 0 5152 0 -1 89760
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_160_56
timestamp 1586364061
transform 1 0 6256 0 -1 89760
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_160_68
timestamp 1586364061
transform 1 0 7360 0 -1 89760
box -38 -48 1142 592
use scs8hd_decap_3  PHY_321
timestamp 1586364061
transform -1 0 8832 0 -1 89760
box -38 -48 314 592
use scs8hd_fill_1  FILLER_160_80
timestamp 1586364061
transform 1 0 8464 0 -1 89760
box -38 -48 130 592
use scs8hd_decap_3  PHY_322
timestamp 1586364061
transform 1 0 1104 0 1 89760
box -38 -48 314 592
use scs8hd_decap_12  FILLER_161_3
timestamp 1586364061
transform 1 0 1380 0 1 89760
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_161_15
timestamp 1586364061
transform 1 0 2484 0 1 89760
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_161_27
timestamp 1586364061
transform 1 0 3588 0 1 89760
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_161_39
timestamp 1586364061
transform 1 0 4692 0 1 89760
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_161_51
timestamp 1586364061
transform 1 0 5796 0 1 89760
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1370
timestamp 1586364061
transform 1 0 6716 0 1 89760
box -38 -48 130 592
use scs8hd_fill_2  FILLER_161_59
timestamp 1586364061
transform 1 0 6532 0 1 89760
box -38 -48 222 592
use scs8hd_decap_12  FILLER_161_62
timestamp 1586364061
transform 1 0 6808 0 1 89760
box -38 -48 1142 592
use scs8hd_decap_3  PHY_323
timestamp 1586364061
transform -1 0 8832 0 1 89760
box -38 -48 314 592
use scs8hd_decap_6  FILLER_161_74
timestamp 1586364061
transform 1 0 7912 0 1 89760
box -38 -48 590 592
use scs8hd_fill_1  FILLER_161_80
timestamp 1586364061
transform 1 0 8464 0 1 89760
box -38 -48 130 592
use scs8hd_decap_3  PHY_324
timestamp 1586364061
transform 1 0 1104 0 -1 90848
box -38 -48 314 592
use scs8hd_decap_12  FILLER_162_3
timestamp 1586364061
transform 1 0 1380 0 -1 90848
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_162_15
timestamp 1586364061
transform 1 0 2484 0 -1 90848
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1371
timestamp 1586364061
transform 1 0 3956 0 -1 90848
box -38 -48 130 592
use scs8hd_decap_4  FILLER_162_27
timestamp 1586364061
transform 1 0 3588 0 -1 90848
box -38 -48 406 592
use scs8hd_decap_12  FILLER_162_32
timestamp 1586364061
transform 1 0 4048 0 -1 90848
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_162_44
timestamp 1586364061
transform 1 0 5152 0 -1 90848
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_162_56
timestamp 1586364061
transform 1 0 6256 0 -1 90848
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_162_68
timestamp 1586364061
transform 1 0 7360 0 -1 90848
box -38 -48 1142 592
use scs8hd_decap_3  PHY_325
timestamp 1586364061
transform -1 0 8832 0 -1 90848
box -38 -48 314 592
use scs8hd_fill_1  FILLER_162_80
timestamp 1586364061
transform 1 0 8464 0 -1 90848
box -38 -48 130 592
use scs8hd_decap_3  PHY_326
timestamp 1586364061
transform 1 0 1104 0 1 90848
box -38 -48 314 592
use scs8hd_decap_12  FILLER_163_3
timestamp 1586364061
transform 1 0 1380 0 1 90848
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_163_15
timestamp 1586364061
transform 1 0 2484 0 1 90848
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_163_27
timestamp 1586364061
transform 1 0 3588 0 1 90848
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_163_39
timestamp 1586364061
transform 1 0 4692 0 1 90848
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_163_51
timestamp 1586364061
transform 1 0 5796 0 1 90848
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1372
timestamp 1586364061
transform 1 0 6716 0 1 90848
box -38 -48 130 592
use scs8hd_fill_2  FILLER_163_59
timestamp 1586364061
transform 1 0 6532 0 1 90848
box -38 -48 222 592
use scs8hd_decap_12  FILLER_163_62
timestamp 1586364061
transform 1 0 6808 0 1 90848
box -38 -48 1142 592
use scs8hd_decap_3  PHY_327
timestamp 1586364061
transform -1 0 8832 0 1 90848
box -38 -48 314 592
use scs8hd_decap_6  FILLER_163_74
timestamp 1586364061
transform 1 0 7912 0 1 90848
box -38 -48 590 592
use scs8hd_fill_1  FILLER_163_80
timestamp 1586364061
transform 1 0 8464 0 1 90848
box -38 -48 130 592
use scs8hd_decap_3  PHY_328
timestamp 1586364061
transform 1 0 1104 0 -1 91936
box -38 -48 314 592
use scs8hd_decap_12  FILLER_164_3
timestamp 1586364061
transform 1 0 1380 0 -1 91936
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_164_15
timestamp 1586364061
transform 1 0 2484 0 -1 91936
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1373
timestamp 1586364061
transform 1 0 3956 0 -1 91936
box -38 -48 130 592
use scs8hd_decap_4  FILLER_164_27
timestamp 1586364061
transform 1 0 3588 0 -1 91936
box -38 -48 406 592
use scs8hd_decap_12  FILLER_164_32
timestamp 1586364061
transform 1 0 4048 0 -1 91936
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_164_44
timestamp 1586364061
transform 1 0 5152 0 -1 91936
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_164_56
timestamp 1586364061
transform 1 0 6256 0 -1 91936
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_164_68
timestamp 1586364061
transform 1 0 7360 0 -1 91936
box -38 -48 1142 592
use scs8hd_decap_3  PHY_329
timestamp 1586364061
transform -1 0 8832 0 -1 91936
box -38 -48 314 592
use scs8hd_fill_1  FILLER_164_80
timestamp 1586364061
transform 1 0 8464 0 -1 91936
box -38 -48 130 592
use scs8hd_decap_3  PHY_330
timestamp 1586364061
transform 1 0 1104 0 1 91936
box -38 -48 314 592
use scs8hd_decap_3  PHY_332
timestamp 1586364061
transform 1 0 1104 0 -1 93024
box -38 -48 314 592
use scs8hd_decap_12  FILLER_165_3
timestamp 1586364061
transform 1 0 1380 0 1 91936
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_165_15
timestamp 1586364061
transform 1 0 2484 0 1 91936
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_166_3
timestamp 1586364061
transform 1 0 1380 0 -1 93024
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_166_15
timestamp 1586364061
transform 1 0 2484 0 -1 93024
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1375
timestamp 1586364061
transform 1 0 3956 0 -1 93024
box -38 -48 130 592
use scs8hd_decap_12  FILLER_165_27
timestamp 1586364061
transform 1 0 3588 0 1 91936
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_166_27
timestamp 1586364061
transform 1 0 3588 0 -1 93024
box -38 -48 406 592
use scs8hd_decap_12  FILLER_166_32
timestamp 1586364061
transform 1 0 4048 0 -1 93024
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_165_39
timestamp 1586364061
transform 1 0 4692 0 1 91936
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_165_51
timestamp 1586364061
transform 1 0 5796 0 1 91936
box -38 -48 774 592
use scs8hd_decap_12  FILLER_166_44
timestamp 1586364061
transform 1 0 5152 0 -1 93024
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1374
timestamp 1586364061
transform 1 0 6716 0 1 91936
box -38 -48 130 592
use scs8hd_fill_2  FILLER_165_59
timestamp 1586364061
transform 1 0 6532 0 1 91936
box -38 -48 222 592
use scs8hd_decap_12  FILLER_165_62
timestamp 1586364061
transform 1 0 6808 0 1 91936
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_166_56
timestamp 1586364061
transform 1 0 6256 0 -1 93024
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_166_68
timestamp 1586364061
transform 1 0 7360 0 -1 93024
box -38 -48 1142 592
use scs8hd_decap_3  PHY_331
timestamp 1586364061
transform -1 0 8832 0 1 91936
box -38 -48 314 592
use scs8hd_decap_3  PHY_333
timestamp 1586364061
transform -1 0 8832 0 -1 93024
box -38 -48 314 592
use scs8hd_decap_6  FILLER_165_74
timestamp 1586364061
transform 1 0 7912 0 1 91936
box -38 -48 590 592
use scs8hd_fill_1  FILLER_165_80
timestamp 1586364061
transform 1 0 8464 0 1 91936
box -38 -48 130 592
use scs8hd_fill_1  FILLER_166_80
timestamp 1586364061
transform 1 0 8464 0 -1 93024
box -38 -48 130 592
use scs8hd_decap_3  PHY_334
timestamp 1586364061
transform 1 0 1104 0 1 93024
box -38 -48 314 592
use scs8hd_decap_12  FILLER_167_3
timestamp 1586364061
transform 1 0 1380 0 1 93024
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_167_15
timestamp 1586364061
transform 1 0 2484 0 1 93024
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_167_27
timestamp 1586364061
transform 1 0 3588 0 1 93024
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_167_39
timestamp 1586364061
transform 1 0 4692 0 1 93024
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_167_51
timestamp 1586364061
transform 1 0 5796 0 1 93024
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1376
timestamp 1586364061
transform 1 0 6716 0 1 93024
box -38 -48 130 592
use scs8hd_fill_2  FILLER_167_59
timestamp 1586364061
transform 1 0 6532 0 1 93024
box -38 -48 222 592
use scs8hd_decap_12  FILLER_167_62
timestamp 1586364061
transform 1 0 6808 0 1 93024
box -38 -48 1142 592
use scs8hd_decap_3  PHY_335
timestamp 1586364061
transform -1 0 8832 0 1 93024
box -38 -48 314 592
use scs8hd_decap_6  FILLER_167_74
timestamp 1586364061
transform 1 0 7912 0 1 93024
box -38 -48 590 592
use scs8hd_fill_1  FILLER_167_80
timestamp 1586364061
transform 1 0 8464 0 1 93024
box -38 -48 130 592
use scs8hd_decap_3  PHY_336
timestamp 1586364061
transform 1 0 1104 0 -1 94112
box -38 -48 314 592
use scs8hd_decap_12  FILLER_168_3
timestamp 1586364061
transform 1 0 1380 0 -1 94112
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_168_15
timestamp 1586364061
transform 1 0 2484 0 -1 94112
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1377
timestamp 1586364061
transform 1 0 3956 0 -1 94112
box -38 -48 130 592
use scs8hd_decap_4  FILLER_168_27
timestamp 1586364061
transform 1 0 3588 0 -1 94112
box -38 -48 406 592
use scs8hd_decap_12  FILLER_168_32
timestamp 1586364061
transform 1 0 4048 0 -1 94112
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_168_44
timestamp 1586364061
transform 1 0 5152 0 -1 94112
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_168_56
timestamp 1586364061
transform 1 0 6256 0 -1 94112
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_168_68
timestamp 1586364061
transform 1 0 7360 0 -1 94112
box -38 -48 1142 592
use scs8hd_decap_3  PHY_337
timestamp 1586364061
transform -1 0 8832 0 -1 94112
box -38 -48 314 592
use scs8hd_fill_1  FILLER_168_80
timestamp 1586364061
transform 1 0 8464 0 -1 94112
box -38 -48 130 592
use scs8hd_decap_3  PHY_338
timestamp 1586364061
transform 1 0 1104 0 1 94112
box -38 -48 314 592
use scs8hd_decap_12  FILLER_169_3
timestamp 1586364061
transform 1 0 1380 0 1 94112
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_169_15
timestamp 1586364061
transform 1 0 2484 0 1 94112
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_169_27
timestamp 1586364061
transform 1 0 3588 0 1 94112
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_169_39
timestamp 1586364061
transform 1 0 4692 0 1 94112
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_169_51
timestamp 1586364061
transform 1 0 5796 0 1 94112
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1378
timestamp 1586364061
transform 1 0 6716 0 1 94112
box -38 -48 130 592
use scs8hd_fill_2  FILLER_169_59
timestamp 1586364061
transform 1 0 6532 0 1 94112
box -38 -48 222 592
use scs8hd_decap_12  FILLER_169_62
timestamp 1586364061
transform 1 0 6808 0 1 94112
box -38 -48 1142 592
use scs8hd_decap_3  PHY_339
timestamp 1586364061
transform -1 0 8832 0 1 94112
box -38 -48 314 592
use scs8hd_decap_6  FILLER_169_74
timestamp 1586364061
transform 1 0 7912 0 1 94112
box -38 -48 590 592
use scs8hd_fill_1  FILLER_169_80
timestamp 1586364061
transform 1 0 8464 0 1 94112
box -38 -48 130 592
use scs8hd_decap_3  PHY_340
timestamp 1586364061
transform 1 0 1104 0 -1 95200
box -38 -48 314 592
use scs8hd_decap_12  FILLER_170_3
timestamp 1586364061
transform 1 0 1380 0 -1 95200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_170_15
timestamp 1586364061
transform 1 0 2484 0 -1 95200
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1379
timestamp 1586364061
transform 1 0 3956 0 -1 95200
box -38 -48 130 592
use scs8hd_decap_4  FILLER_170_27
timestamp 1586364061
transform 1 0 3588 0 -1 95200
box -38 -48 406 592
use scs8hd_decap_12  FILLER_170_32
timestamp 1586364061
transform 1 0 4048 0 -1 95200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_170_44
timestamp 1586364061
transform 1 0 5152 0 -1 95200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_170_56
timestamp 1586364061
transform 1 0 6256 0 -1 95200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_170_68
timestamp 1586364061
transform 1 0 7360 0 -1 95200
box -38 -48 1142 592
use scs8hd_decap_3  PHY_341
timestamp 1586364061
transform -1 0 8832 0 -1 95200
box -38 -48 314 592
use scs8hd_fill_1  FILLER_170_80
timestamp 1586364061
transform 1 0 8464 0 -1 95200
box -38 -48 130 592
use scs8hd_decap_3  PHY_342
timestamp 1586364061
transform 1 0 1104 0 1 95200
box -38 -48 314 592
use scs8hd_decap_3  PHY_344
timestamp 1586364061
transform 1 0 1104 0 -1 96288
box -38 -48 314 592
use scs8hd_decap_12  FILLER_171_3
timestamp 1586364061
transform 1 0 1380 0 1 95200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_171_15
timestamp 1586364061
transform 1 0 2484 0 1 95200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_172_3
timestamp 1586364061
transform 1 0 1380 0 -1 96288
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_172_15
timestamp 1586364061
transform 1 0 2484 0 -1 96288
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1381
timestamp 1586364061
transform 1 0 3956 0 -1 96288
box -38 -48 130 592
use scs8hd_decap_12  FILLER_171_27
timestamp 1586364061
transform 1 0 3588 0 1 95200
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_172_27
timestamp 1586364061
transform 1 0 3588 0 -1 96288
box -38 -48 406 592
use scs8hd_decap_12  FILLER_172_32
timestamp 1586364061
transform 1 0 4048 0 -1 96288
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_171_39
timestamp 1586364061
transform 1 0 4692 0 1 95200
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_171_51
timestamp 1586364061
transform 1 0 5796 0 1 95200
box -38 -48 774 592
use scs8hd_decap_12  FILLER_172_44
timestamp 1586364061
transform 1 0 5152 0 -1 96288
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1380
timestamp 1586364061
transform 1 0 6716 0 1 95200
box -38 -48 130 592
use scs8hd_fill_2  FILLER_171_59
timestamp 1586364061
transform 1 0 6532 0 1 95200
box -38 -48 222 592
use scs8hd_decap_12  FILLER_171_62
timestamp 1586364061
transform 1 0 6808 0 1 95200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_172_56
timestamp 1586364061
transform 1 0 6256 0 -1 96288
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_172_68
timestamp 1586364061
transform 1 0 7360 0 -1 96288
box -38 -48 1142 592
use scs8hd_decap_3  PHY_343
timestamp 1586364061
transform -1 0 8832 0 1 95200
box -38 -48 314 592
use scs8hd_decap_3  PHY_345
timestamp 1586364061
transform -1 0 8832 0 -1 96288
box -38 -48 314 592
use scs8hd_decap_6  FILLER_171_74
timestamp 1586364061
transform 1 0 7912 0 1 95200
box -38 -48 590 592
use scs8hd_fill_1  FILLER_171_80
timestamp 1586364061
transform 1 0 8464 0 1 95200
box -38 -48 130 592
use scs8hd_fill_1  FILLER_172_80
timestamp 1586364061
transform 1 0 8464 0 -1 96288
box -38 -48 130 592
use scs8hd_decap_3  PHY_346
timestamp 1586364061
transform 1 0 1104 0 1 96288
box -38 -48 314 592
use scs8hd_decap_12  FILLER_173_3
timestamp 1586364061
transform 1 0 1380 0 1 96288
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_173_15
timestamp 1586364061
transform 1 0 2484 0 1 96288
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_173_27
timestamp 1586364061
transform 1 0 3588 0 1 96288
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_173_39
timestamp 1586364061
transform 1 0 4692 0 1 96288
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_173_51
timestamp 1586364061
transform 1 0 5796 0 1 96288
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1382
timestamp 1586364061
transform 1 0 6716 0 1 96288
box -38 -48 130 592
use scs8hd_fill_2  FILLER_173_59
timestamp 1586364061
transform 1 0 6532 0 1 96288
box -38 -48 222 592
use scs8hd_decap_12  FILLER_173_62
timestamp 1586364061
transform 1 0 6808 0 1 96288
box -38 -48 1142 592
use scs8hd_decap_3  PHY_347
timestamp 1586364061
transform -1 0 8832 0 1 96288
box -38 -48 314 592
use scs8hd_decap_6  FILLER_173_74
timestamp 1586364061
transform 1 0 7912 0 1 96288
box -38 -48 590 592
use scs8hd_fill_1  FILLER_173_80
timestamp 1586364061
transform 1 0 8464 0 1 96288
box -38 -48 130 592
use scs8hd_decap_3  PHY_348
timestamp 1586364061
transform 1 0 1104 0 -1 97376
box -38 -48 314 592
use scs8hd_decap_12  FILLER_174_3
timestamp 1586364061
transform 1 0 1380 0 -1 97376
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_174_15
timestamp 1586364061
transform 1 0 2484 0 -1 97376
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1383
timestamp 1586364061
transform 1 0 3956 0 -1 97376
box -38 -48 130 592
use scs8hd_decap_4  FILLER_174_27
timestamp 1586364061
transform 1 0 3588 0 -1 97376
box -38 -48 406 592
use scs8hd_decap_12  FILLER_174_32
timestamp 1586364061
transform 1 0 4048 0 -1 97376
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_174_44
timestamp 1586364061
transform 1 0 5152 0 -1 97376
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_174_56
timestamp 1586364061
transform 1 0 6256 0 -1 97376
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_174_68
timestamp 1586364061
transform 1 0 7360 0 -1 97376
box -38 -48 1142 592
use scs8hd_decap_3  PHY_349
timestamp 1586364061
transform -1 0 8832 0 -1 97376
box -38 -48 314 592
use scs8hd_fill_1  FILLER_174_80
timestamp 1586364061
transform 1 0 8464 0 -1 97376
box -38 -48 130 592
use scs8hd_decap_3  PHY_350
timestamp 1586364061
transform 1 0 1104 0 1 97376
box -38 -48 314 592
use scs8hd_decap_12  FILLER_175_3
timestamp 1586364061
transform 1 0 1380 0 1 97376
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_175_15
timestamp 1586364061
transform 1 0 2484 0 1 97376
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_175_27
timestamp 1586364061
transform 1 0 3588 0 1 97376
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_175_39
timestamp 1586364061
transform 1 0 4692 0 1 97376
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_175_51
timestamp 1586364061
transform 1 0 5796 0 1 97376
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1384
timestamp 1586364061
transform 1 0 6716 0 1 97376
box -38 -48 130 592
use scs8hd_fill_2  FILLER_175_59
timestamp 1586364061
transform 1 0 6532 0 1 97376
box -38 -48 222 592
use scs8hd_decap_12  FILLER_175_62
timestamp 1586364061
transform 1 0 6808 0 1 97376
box -38 -48 1142 592
use scs8hd_decap_3  PHY_351
timestamp 1586364061
transform -1 0 8832 0 1 97376
box -38 -48 314 592
use scs8hd_decap_6  FILLER_175_74
timestamp 1586364061
transform 1 0 7912 0 1 97376
box -38 -48 590 592
use scs8hd_fill_1  FILLER_175_80
timestamp 1586364061
transform 1 0 8464 0 1 97376
box -38 -48 130 592
use scs8hd_decap_3  PHY_352
timestamp 1586364061
transform 1 0 1104 0 -1 98464
box -38 -48 314 592
use scs8hd_decap_12  FILLER_176_3
timestamp 1586364061
transform 1 0 1380 0 -1 98464
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_176_15
timestamp 1586364061
transform 1 0 2484 0 -1 98464
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1385
timestamp 1586364061
transform 1 0 3956 0 -1 98464
box -38 -48 130 592
use scs8hd_decap_4  FILLER_176_27
timestamp 1586364061
transform 1 0 3588 0 -1 98464
box -38 -48 406 592
use scs8hd_decap_12  FILLER_176_32
timestamp 1586364061
transform 1 0 4048 0 -1 98464
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_176_44
timestamp 1586364061
transform 1 0 5152 0 -1 98464
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_176_56
timestamp 1586364061
transform 1 0 6256 0 -1 98464
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_176_68
timestamp 1586364061
transform 1 0 7360 0 -1 98464
box -38 -48 1142 592
use scs8hd_decap_3  PHY_353
timestamp 1586364061
transform -1 0 8832 0 -1 98464
box -38 -48 314 592
use scs8hd_fill_1  FILLER_176_80
timestamp 1586364061
transform 1 0 8464 0 -1 98464
box -38 -48 130 592
use scs8hd_decap_3  PHY_354
timestamp 1586364061
transform 1 0 1104 0 1 98464
box -38 -48 314 592
use scs8hd_decap_12  FILLER_177_3
timestamp 1586364061
transform 1 0 1380 0 1 98464
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_177_15
timestamp 1586364061
transform 1 0 2484 0 1 98464
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_177_27
timestamp 1586364061
transform 1 0 3588 0 1 98464
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_177_39
timestamp 1586364061
transform 1 0 4692 0 1 98464
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_177_51
timestamp 1586364061
transform 1 0 5796 0 1 98464
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1386
timestamp 1586364061
transform 1 0 6716 0 1 98464
box -38 -48 130 592
use scs8hd_fill_2  FILLER_177_59
timestamp 1586364061
transform 1 0 6532 0 1 98464
box -38 -48 222 592
use scs8hd_decap_12  FILLER_177_62
timestamp 1586364061
transform 1 0 6808 0 1 98464
box -38 -48 1142 592
use scs8hd_decap_3  PHY_355
timestamp 1586364061
transform -1 0 8832 0 1 98464
box -38 -48 314 592
use scs8hd_decap_6  FILLER_177_74
timestamp 1586364061
transform 1 0 7912 0 1 98464
box -38 -48 590 592
use scs8hd_fill_1  FILLER_177_80
timestamp 1586364061
transform 1 0 8464 0 1 98464
box -38 -48 130 592
use scs8hd_decap_3  PHY_356
timestamp 1586364061
transform 1 0 1104 0 -1 99552
box -38 -48 314 592
use scs8hd_decap_3  PHY_358
timestamp 1586364061
transform 1 0 1104 0 1 99552
box -38 -48 314 592
use scs8hd_decap_12  FILLER_178_3
timestamp 1586364061
transform 1 0 1380 0 -1 99552
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_178_15
timestamp 1586364061
transform 1 0 2484 0 -1 99552
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_179_3
timestamp 1586364061
transform 1 0 1380 0 1 99552
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_179_15
timestamp 1586364061
transform 1 0 2484 0 1 99552
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1387
timestamp 1586364061
transform 1 0 3956 0 -1 99552
box -38 -48 130 592
use scs8hd_decap_4  FILLER_178_27
timestamp 1586364061
transform 1 0 3588 0 -1 99552
box -38 -48 406 592
use scs8hd_decap_12  FILLER_178_32
timestamp 1586364061
transform 1 0 4048 0 -1 99552
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_179_27
timestamp 1586364061
transform 1 0 3588 0 1 99552
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_178_44
timestamp 1586364061
transform 1 0 5152 0 -1 99552
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_179_39
timestamp 1586364061
transform 1 0 4692 0 1 99552
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_179_51
timestamp 1586364061
transform 1 0 5796 0 1 99552
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1388
timestamp 1586364061
transform 1 0 6716 0 1 99552
box -38 -48 130 592
use scs8hd_decap_12  FILLER_178_56
timestamp 1586364061
transform 1 0 6256 0 -1 99552
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_178_68
timestamp 1586364061
transform 1 0 7360 0 -1 99552
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_179_59
timestamp 1586364061
transform 1 0 6532 0 1 99552
box -38 -48 222 592
use scs8hd_decap_12  FILLER_179_62
timestamp 1586364061
transform 1 0 6808 0 1 99552
box -38 -48 1142 592
use scs8hd_decap_3  PHY_357
timestamp 1586364061
transform -1 0 8832 0 -1 99552
box -38 -48 314 592
use scs8hd_decap_3  PHY_359
timestamp 1586364061
transform -1 0 8832 0 1 99552
box -38 -48 314 592
use scs8hd_fill_1  FILLER_178_80
timestamp 1586364061
transform 1 0 8464 0 -1 99552
box -38 -48 130 592
use scs8hd_decap_6  FILLER_179_74
timestamp 1586364061
transform 1 0 7912 0 1 99552
box -38 -48 590 592
use scs8hd_fill_1  FILLER_179_80
timestamp 1586364061
transform 1 0 8464 0 1 99552
box -38 -48 130 592
use scs8hd_decap_3  PHY_360
timestamp 1586364061
transform 1 0 1104 0 -1 100640
box -38 -48 314 592
use scs8hd_decap_12  FILLER_180_3
timestamp 1586364061
transform 1 0 1380 0 -1 100640
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_180_15
timestamp 1586364061
transform 1 0 2484 0 -1 100640
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1389
timestamp 1586364061
transform 1 0 3956 0 -1 100640
box -38 -48 130 592
use scs8hd_decap_4  FILLER_180_27
timestamp 1586364061
transform 1 0 3588 0 -1 100640
box -38 -48 406 592
use scs8hd_decap_12  FILLER_180_32
timestamp 1586364061
transform 1 0 4048 0 -1 100640
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_180_44
timestamp 1586364061
transform 1 0 5152 0 -1 100640
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_180_56
timestamp 1586364061
transform 1 0 6256 0 -1 100640
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_180_68
timestamp 1586364061
transform 1 0 7360 0 -1 100640
box -38 -48 1142 592
use scs8hd_decap_3  PHY_361
timestamp 1586364061
transform -1 0 8832 0 -1 100640
box -38 -48 314 592
use scs8hd_fill_1  FILLER_180_80
timestamp 1586364061
transform 1 0 8464 0 -1 100640
box -38 -48 130 592
use scs8hd_decap_3  PHY_362
timestamp 1586364061
transform 1 0 1104 0 1 100640
box -38 -48 314 592
use scs8hd_decap_12  FILLER_181_3
timestamp 1586364061
transform 1 0 1380 0 1 100640
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_181_15
timestamp 1586364061
transform 1 0 2484 0 1 100640
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_181_27
timestamp 1586364061
transform 1 0 3588 0 1 100640
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_181_39
timestamp 1586364061
transform 1 0 4692 0 1 100640
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_181_51
timestamp 1586364061
transform 1 0 5796 0 1 100640
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1390
timestamp 1586364061
transform 1 0 6716 0 1 100640
box -38 -48 130 592
use scs8hd_fill_2  FILLER_181_59
timestamp 1586364061
transform 1 0 6532 0 1 100640
box -38 -48 222 592
use scs8hd_decap_12  FILLER_181_62
timestamp 1586364061
transform 1 0 6808 0 1 100640
box -38 -48 1142 592
use scs8hd_decap_3  PHY_363
timestamp 1586364061
transform -1 0 8832 0 1 100640
box -38 -48 314 592
use scs8hd_decap_6  FILLER_181_74
timestamp 1586364061
transform 1 0 7912 0 1 100640
box -38 -48 590 592
use scs8hd_fill_1  FILLER_181_80
timestamp 1586364061
transform 1 0 8464 0 1 100640
box -38 -48 130 592
use scs8hd_decap_3  PHY_364
timestamp 1586364061
transform 1 0 1104 0 -1 101728
box -38 -48 314 592
use scs8hd_decap_12  FILLER_182_3
timestamp 1586364061
transform 1 0 1380 0 -1 101728
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_182_15
timestamp 1586364061
transform 1 0 2484 0 -1 101728
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1391
timestamp 1586364061
transform 1 0 3956 0 -1 101728
box -38 -48 130 592
use scs8hd_decap_4  FILLER_182_27
timestamp 1586364061
transform 1 0 3588 0 -1 101728
box -38 -48 406 592
use scs8hd_decap_12  FILLER_182_32
timestamp 1586364061
transform 1 0 4048 0 -1 101728
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_182_44
timestamp 1586364061
transform 1 0 5152 0 -1 101728
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_182_56
timestamp 1586364061
transform 1 0 6256 0 -1 101728
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_182_68
timestamp 1586364061
transform 1 0 7360 0 -1 101728
box -38 -48 1142 592
use scs8hd_decap_3  PHY_365
timestamp 1586364061
transform -1 0 8832 0 -1 101728
box -38 -48 314 592
use scs8hd_fill_1  FILLER_182_80
timestamp 1586364061
transform 1 0 8464 0 -1 101728
box -38 -48 130 592
use scs8hd_decap_3  PHY_366
timestamp 1586364061
transform 1 0 1104 0 1 101728
box -38 -48 314 592
use scs8hd_decap_12  FILLER_183_3
timestamp 1586364061
transform 1 0 1380 0 1 101728
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_183_15
timestamp 1586364061
transform 1 0 2484 0 1 101728
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_183_27
timestamp 1586364061
transform 1 0 3588 0 1 101728
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_183_39
timestamp 1586364061
transform 1 0 4692 0 1 101728
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_183_51
timestamp 1586364061
transform 1 0 5796 0 1 101728
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1392
timestamp 1586364061
transform 1 0 6716 0 1 101728
box -38 -48 130 592
use scs8hd_fill_2  FILLER_183_59
timestamp 1586364061
transform 1 0 6532 0 1 101728
box -38 -48 222 592
use scs8hd_decap_12  FILLER_183_62
timestamp 1586364061
transform 1 0 6808 0 1 101728
box -38 -48 1142 592
use scs8hd_decap_3  PHY_367
timestamp 1586364061
transform -1 0 8832 0 1 101728
box -38 -48 314 592
use scs8hd_decap_6  FILLER_183_74
timestamp 1586364061
transform 1 0 7912 0 1 101728
box -38 -48 590 592
use scs8hd_fill_1  FILLER_183_80
timestamp 1586364061
transform 1 0 8464 0 1 101728
box -38 -48 130 592
use scs8hd_decap_3  PHY_368
timestamp 1586364061
transform 1 0 1104 0 -1 102816
box -38 -48 314 592
use scs8hd_decap_12  FILLER_184_3
timestamp 1586364061
transform 1 0 1380 0 -1 102816
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_184_15
timestamp 1586364061
transform 1 0 2484 0 -1 102816
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1393
timestamp 1586364061
transform 1 0 3956 0 -1 102816
box -38 -48 130 592
use scs8hd_decap_4  FILLER_184_27
timestamp 1586364061
transform 1 0 3588 0 -1 102816
box -38 -48 406 592
use scs8hd_decap_12  FILLER_184_32
timestamp 1586364061
transform 1 0 4048 0 -1 102816
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_184_44
timestamp 1586364061
transform 1 0 5152 0 -1 102816
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_184_56
timestamp 1586364061
transform 1 0 6256 0 -1 102816
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_184_68
timestamp 1586364061
transform 1 0 7360 0 -1 102816
box -38 -48 1142 592
use scs8hd_decap_3  PHY_369
timestamp 1586364061
transform -1 0 8832 0 -1 102816
box -38 -48 314 592
use scs8hd_fill_1  FILLER_184_80
timestamp 1586364061
transform 1 0 8464 0 -1 102816
box -38 -48 130 592
use scs8hd_decap_3  PHY_370
timestamp 1586364061
transform 1 0 1104 0 1 102816
box -38 -48 314 592
use scs8hd_decap_3  PHY_372
timestamp 1586364061
transform 1 0 1104 0 -1 103904
box -38 -48 314 592
use scs8hd_decap_12  FILLER_185_3
timestamp 1586364061
transform 1 0 1380 0 1 102816
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_185_15
timestamp 1586364061
transform 1 0 2484 0 1 102816
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_186_3
timestamp 1586364061
transform 1 0 1380 0 -1 103904
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_186_15
timestamp 1586364061
transform 1 0 2484 0 -1 103904
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1395
timestamp 1586364061
transform 1 0 3956 0 -1 103904
box -38 -48 130 592
use scs8hd_decap_12  FILLER_185_27
timestamp 1586364061
transform 1 0 3588 0 1 102816
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_186_27
timestamp 1586364061
transform 1 0 3588 0 -1 103904
box -38 -48 406 592
use scs8hd_decap_12  FILLER_186_32
timestamp 1586364061
transform 1 0 4048 0 -1 103904
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_185_39
timestamp 1586364061
transform 1 0 4692 0 1 102816
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_185_51
timestamp 1586364061
transform 1 0 5796 0 1 102816
box -38 -48 774 592
use scs8hd_decap_12  FILLER_186_44
timestamp 1586364061
transform 1 0 5152 0 -1 103904
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1394
timestamp 1586364061
transform 1 0 6716 0 1 102816
box -38 -48 130 592
use scs8hd_fill_2  FILLER_185_59
timestamp 1586364061
transform 1 0 6532 0 1 102816
box -38 -48 222 592
use scs8hd_decap_12  FILLER_185_62
timestamp 1586364061
transform 1 0 6808 0 1 102816
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_186_56
timestamp 1586364061
transform 1 0 6256 0 -1 103904
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_186_68
timestamp 1586364061
transform 1 0 7360 0 -1 103904
box -38 -48 1142 592
use scs8hd_decap_3  PHY_371
timestamp 1586364061
transform -1 0 8832 0 1 102816
box -38 -48 314 592
use scs8hd_decap_3  PHY_373
timestamp 1586364061
transform -1 0 8832 0 -1 103904
box -38 -48 314 592
use scs8hd_decap_6  FILLER_185_74
timestamp 1586364061
transform 1 0 7912 0 1 102816
box -38 -48 590 592
use scs8hd_fill_1  FILLER_185_80
timestamp 1586364061
transform 1 0 8464 0 1 102816
box -38 -48 130 592
use scs8hd_fill_1  FILLER_186_80
timestamp 1586364061
transform 1 0 8464 0 -1 103904
box -38 -48 130 592
use scs8hd_decap_3  PHY_374
timestamp 1586364061
transform 1 0 1104 0 1 103904
box -38 -48 314 592
use scs8hd_decap_12  FILLER_187_3
timestamp 1586364061
transform 1 0 1380 0 1 103904
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_187_15
timestamp 1586364061
transform 1 0 2484 0 1 103904
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_187_27
timestamp 1586364061
transform 1 0 3588 0 1 103904
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_187_39
timestamp 1586364061
transform 1 0 4692 0 1 103904
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_187_51
timestamp 1586364061
transform 1 0 5796 0 1 103904
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1396
timestamp 1586364061
transform 1 0 6716 0 1 103904
box -38 -48 130 592
use scs8hd_fill_2  FILLER_187_59
timestamp 1586364061
transform 1 0 6532 0 1 103904
box -38 -48 222 592
use scs8hd_decap_12  FILLER_187_62
timestamp 1586364061
transform 1 0 6808 0 1 103904
box -38 -48 1142 592
use scs8hd_decap_3  PHY_375
timestamp 1586364061
transform -1 0 8832 0 1 103904
box -38 -48 314 592
use scs8hd_decap_6  FILLER_187_74
timestamp 1586364061
transform 1 0 7912 0 1 103904
box -38 -48 590 592
use scs8hd_fill_1  FILLER_187_80
timestamp 1586364061
transform 1 0 8464 0 1 103904
box -38 -48 130 592
use scs8hd_decap_3  PHY_376
timestamp 1586364061
transform 1 0 1104 0 -1 104992
box -38 -48 314 592
use scs8hd_decap_12  FILLER_188_3
timestamp 1586364061
transform 1 0 1380 0 -1 104992
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_188_15
timestamp 1586364061
transform 1 0 2484 0 -1 104992
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1397
timestamp 1586364061
transform 1 0 3956 0 -1 104992
box -38 -48 130 592
use scs8hd_decap_4  FILLER_188_27
timestamp 1586364061
transform 1 0 3588 0 -1 104992
box -38 -48 406 592
use scs8hd_decap_12  FILLER_188_32
timestamp 1586364061
transform 1 0 4048 0 -1 104992
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_188_44
timestamp 1586364061
transform 1 0 5152 0 -1 104992
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_188_56
timestamp 1586364061
transform 1 0 6256 0 -1 104992
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_188_68
timestamp 1586364061
transform 1 0 7360 0 -1 104992
box -38 -48 1142 592
use scs8hd_decap_3  PHY_377
timestamp 1586364061
transform -1 0 8832 0 -1 104992
box -38 -48 314 592
use scs8hd_fill_1  FILLER_188_80
timestamp 1586364061
transform 1 0 8464 0 -1 104992
box -38 -48 130 592
use scs8hd_decap_3  PHY_378
timestamp 1586364061
transform 1 0 1104 0 1 104992
box -38 -48 314 592
use scs8hd_decap_12  FILLER_189_3
timestamp 1586364061
transform 1 0 1380 0 1 104992
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_189_15
timestamp 1586364061
transform 1 0 2484 0 1 104992
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_189_27
timestamp 1586364061
transform 1 0 3588 0 1 104992
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_189_39
timestamp 1586364061
transform 1 0 4692 0 1 104992
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_189_51
timestamp 1586364061
transform 1 0 5796 0 1 104992
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1398
timestamp 1586364061
transform 1 0 6716 0 1 104992
box -38 -48 130 592
use scs8hd_fill_2  FILLER_189_59
timestamp 1586364061
transform 1 0 6532 0 1 104992
box -38 -48 222 592
use scs8hd_decap_12  FILLER_189_62
timestamp 1586364061
transform 1 0 6808 0 1 104992
box -38 -48 1142 592
use scs8hd_decap_3  PHY_379
timestamp 1586364061
transform -1 0 8832 0 1 104992
box -38 -48 314 592
use scs8hd_decap_6  FILLER_189_74
timestamp 1586364061
transform 1 0 7912 0 1 104992
box -38 -48 590 592
use scs8hd_fill_1  FILLER_189_80
timestamp 1586364061
transform 1 0 8464 0 1 104992
box -38 -48 130 592
use scs8hd_decap_3  PHY_380
timestamp 1586364061
transform 1 0 1104 0 -1 106080
box -38 -48 314 592
use scs8hd_decap_12  FILLER_190_3
timestamp 1586364061
transform 1 0 1380 0 -1 106080
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_190_15
timestamp 1586364061
transform 1 0 2484 0 -1 106080
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1399
timestamp 1586364061
transform 1 0 3956 0 -1 106080
box -38 -48 130 592
use scs8hd_decap_4  FILLER_190_27
timestamp 1586364061
transform 1 0 3588 0 -1 106080
box -38 -48 406 592
use scs8hd_decap_12  FILLER_190_32
timestamp 1586364061
transform 1 0 4048 0 -1 106080
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_190_44
timestamp 1586364061
transform 1 0 5152 0 -1 106080
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_190_56
timestamp 1586364061
transform 1 0 6256 0 -1 106080
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_190_68
timestamp 1586364061
transform 1 0 7360 0 -1 106080
box -38 -48 1142 592
use scs8hd_decap_3  PHY_381
timestamp 1586364061
transform -1 0 8832 0 -1 106080
box -38 -48 314 592
use scs8hd_fill_1  FILLER_190_80
timestamp 1586364061
transform 1 0 8464 0 -1 106080
box -38 -48 130 592
use scs8hd_decap_3  PHY_382
timestamp 1586364061
transform 1 0 1104 0 1 106080
box -38 -48 314 592
use scs8hd_decap_3  PHY_384
timestamp 1586364061
transform 1 0 1104 0 -1 107168
box -38 -48 314 592
use scs8hd_decap_12  FILLER_191_3
timestamp 1586364061
transform 1 0 1380 0 1 106080
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_191_15
timestamp 1586364061
transform 1 0 2484 0 1 106080
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_192_3
timestamp 1586364061
transform 1 0 1380 0 -1 107168
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_192_15
timestamp 1586364061
transform 1 0 2484 0 -1 107168
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1401
timestamp 1586364061
transform 1 0 3956 0 -1 107168
box -38 -48 130 592
use scs8hd_decap_12  FILLER_191_27
timestamp 1586364061
transform 1 0 3588 0 1 106080
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_192_27
timestamp 1586364061
transform 1 0 3588 0 -1 107168
box -38 -48 406 592
use scs8hd_decap_12  FILLER_192_32
timestamp 1586364061
transform 1 0 4048 0 -1 107168
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_191_39
timestamp 1586364061
transform 1 0 4692 0 1 106080
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_191_51
timestamp 1586364061
transform 1 0 5796 0 1 106080
box -38 -48 774 592
use scs8hd_decap_12  FILLER_192_44
timestamp 1586364061
transform 1 0 5152 0 -1 107168
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1400
timestamp 1586364061
transform 1 0 6716 0 1 106080
box -38 -48 130 592
use scs8hd_fill_2  FILLER_191_59
timestamp 1586364061
transform 1 0 6532 0 1 106080
box -38 -48 222 592
use scs8hd_decap_12  FILLER_191_62
timestamp 1586364061
transform 1 0 6808 0 1 106080
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_192_56
timestamp 1586364061
transform 1 0 6256 0 -1 107168
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_192_68
timestamp 1586364061
transform 1 0 7360 0 -1 107168
box -38 -48 1142 592
use scs8hd_decap_3  PHY_383
timestamp 1586364061
transform -1 0 8832 0 1 106080
box -38 -48 314 592
use scs8hd_decap_3  PHY_385
timestamp 1586364061
transform -1 0 8832 0 -1 107168
box -38 -48 314 592
use scs8hd_decap_6  FILLER_191_74
timestamp 1586364061
transform 1 0 7912 0 1 106080
box -38 -48 590 592
use scs8hd_fill_1  FILLER_191_80
timestamp 1586364061
transform 1 0 8464 0 1 106080
box -38 -48 130 592
use scs8hd_fill_1  FILLER_192_80
timestamp 1586364061
transform 1 0 8464 0 -1 107168
box -38 -48 130 592
use scs8hd_decap_3  PHY_386
timestamp 1586364061
transform 1 0 1104 0 1 107168
box -38 -48 314 592
use scs8hd_decap_12  FILLER_193_3
timestamp 1586364061
transform 1 0 1380 0 1 107168
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_193_15
timestamp 1586364061
transform 1 0 2484 0 1 107168
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_193_27
timestamp 1586364061
transform 1 0 3588 0 1 107168
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_193_39
timestamp 1586364061
transform 1 0 4692 0 1 107168
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_193_51
timestamp 1586364061
transform 1 0 5796 0 1 107168
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1402
timestamp 1586364061
transform 1 0 6716 0 1 107168
box -38 -48 130 592
use scs8hd_fill_2  FILLER_193_59
timestamp 1586364061
transform 1 0 6532 0 1 107168
box -38 -48 222 592
use scs8hd_decap_12  FILLER_193_62
timestamp 1586364061
transform 1 0 6808 0 1 107168
box -38 -48 1142 592
use scs8hd_decap_3  PHY_387
timestamp 1586364061
transform -1 0 8832 0 1 107168
box -38 -48 314 592
use scs8hd_decap_6  FILLER_193_74
timestamp 1586364061
transform 1 0 7912 0 1 107168
box -38 -48 590 592
use scs8hd_fill_1  FILLER_193_80
timestamp 1586364061
transform 1 0 8464 0 1 107168
box -38 -48 130 592
use scs8hd_decap_3  PHY_388
timestamp 1586364061
transform 1 0 1104 0 -1 108256
box -38 -48 314 592
use scs8hd_decap_12  FILLER_194_3
timestamp 1586364061
transform 1 0 1380 0 -1 108256
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_194_15
timestamp 1586364061
transform 1 0 2484 0 -1 108256
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1403
timestamp 1586364061
transform 1 0 3956 0 -1 108256
box -38 -48 130 592
use scs8hd_decap_4  FILLER_194_27
timestamp 1586364061
transform 1 0 3588 0 -1 108256
box -38 -48 406 592
use scs8hd_decap_12  FILLER_194_32
timestamp 1586364061
transform 1 0 4048 0 -1 108256
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_194_44
timestamp 1586364061
transform 1 0 5152 0 -1 108256
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_194_56
timestamp 1586364061
transform 1 0 6256 0 -1 108256
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_194_68
timestamp 1586364061
transform 1 0 7360 0 -1 108256
box -38 -48 1142 592
use scs8hd_decap_3  PHY_389
timestamp 1586364061
transform -1 0 8832 0 -1 108256
box -38 -48 314 592
use scs8hd_fill_1  FILLER_194_80
timestamp 1586364061
transform 1 0 8464 0 -1 108256
box -38 -48 130 592
use scs8hd_decap_3  PHY_390
timestamp 1586364061
transform 1 0 1104 0 1 108256
box -38 -48 314 592
use scs8hd_decap_12  FILLER_195_3
timestamp 1586364061
transform 1 0 1380 0 1 108256
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_195_15
timestamp 1586364061
transform 1 0 2484 0 1 108256
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_195_27
timestamp 1586364061
transform 1 0 3588 0 1 108256
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_195_39
timestamp 1586364061
transform 1 0 4692 0 1 108256
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_195_51
timestamp 1586364061
transform 1 0 5796 0 1 108256
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1404
timestamp 1586364061
transform 1 0 6716 0 1 108256
box -38 -48 130 592
use scs8hd_fill_2  FILLER_195_59
timestamp 1586364061
transform 1 0 6532 0 1 108256
box -38 -48 222 592
use scs8hd_decap_12  FILLER_195_62
timestamp 1586364061
transform 1 0 6808 0 1 108256
box -38 -48 1142 592
use scs8hd_decap_3  PHY_391
timestamp 1586364061
transform -1 0 8832 0 1 108256
box -38 -48 314 592
use scs8hd_decap_6  FILLER_195_74
timestamp 1586364061
transform 1 0 7912 0 1 108256
box -38 -48 590 592
use scs8hd_fill_1  FILLER_195_80
timestamp 1586364061
transform 1 0 8464 0 1 108256
box -38 -48 130 592
use scs8hd_decap_3  PHY_392
timestamp 1586364061
transform 1 0 1104 0 -1 109344
box -38 -48 314 592
use scs8hd_decap_12  FILLER_196_3
timestamp 1586364061
transform 1 0 1380 0 -1 109344
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_196_15
timestamp 1586364061
transform 1 0 2484 0 -1 109344
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1405
timestamp 1586364061
transform 1 0 3956 0 -1 109344
box -38 -48 130 592
use scs8hd_decap_4  FILLER_196_27
timestamp 1586364061
transform 1 0 3588 0 -1 109344
box -38 -48 406 592
use scs8hd_decap_12  FILLER_196_32
timestamp 1586364061
transform 1 0 4048 0 -1 109344
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_196_44
timestamp 1586364061
transform 1 0 5152 0 -1 109344
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_196_56
timestamp 1586364061
transform 1 0 6256 0 -1 109344
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_196_68
timestamp 1586364061
transform 1 0 7360 0 -1 109344
box -38 -48 1142 592
use scs8hd_decap_3  PHY_393
timestamp 1586364061
transform -1 0 8832 0 -1 109344
box -38 -48 314 592
use scs8hd_fill_1  FILLER_196_80
timestamp 1586364061
transform 1 0 8464 0 -1 109344
box -38 -48 130 592
use scs8hd_decap_3  PHY_394
timestamp 1586364061
transform 1 0 1104 0 1 109344
box -38 -48 314 592
use scs8hd_decap_12  FILLER_197_3
timestamp 1586364061
transform 1 0 1380 0 1 109344
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_197_15
timestamp 1586364061
transform 1 0 2484 0 1 109344
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_197_27
timestamp 1586364061
transform 1 0 3588 0 1 109344
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_197_39
timestamp 1586364061
transform 1 0 4692 0 1 109344
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_197_51
timestamp 1586364061
transform 1 0 5796 0 1 109344
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1406
timestamp 1586364061
transform 1 0 6716 0 1 109344
box -38 -48 130 592
use scs8hd_fill_2  FILLER_197_59
timestamp 1586364061
transform 1 0 6532 0 1 109344
box -38 -48 222 592
use scs8hd_decap_12  FILLER_197_62
timestamp 1586364061
transform 1 0 6808 0 1 109344
box -38 -48 1142 592
use scs8hd_decap_3  PHY_395
timestamp 1586364061
transform -1 0 8832 0 1 109344
box -38 -48 314 592
use scs8hd_decap_6  FILLER_197_74
timestamp 1586364061
transform 1 0 7912 0 1 109344
box -38 -48 590 592
use scs8hd_fill_1  FILLER_197_80
timestamp 1586364061
transform 1 0 8464 0 1 109344
box -38 -48 130 592
use scs8hd_decap_3  PHY_396
timestamp 1586364061
transform 1 0 1104 0 -1 110432
box -38 -48 314 592
use scs8hd_decap_3  PHY_398
timestamp 1586364061
transform 1 0 1104 0 1 110432
box -38 -48 314 592
use scs8hd_decap_12  FILLER_198_3
timestamp 1586364061
transform 1 0 1380 0 -1 110432
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_198_15
timestamp 1586364061
transform 1 0 2484 0 -1 110432
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_199_3
timestamp 1586364061
transform 1 0 1380 0 1 110432
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_199_15
timestamp 1586364061
transform 1 0 2484 0 1 110432
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1407
timestamp 1586364061
transform 1 0 3956 0 -1 110432
box -38 -48 130 592
use scs8hd_decap_4  FILLER_198_27
timestamp 1586364061
transform 1 0 3588 0 -1 110432
box -38 -48 406 592
use scs8hd_decap_12  FILLER_198_32
timestamp 1586364061
transform 1 0 4048 0 -1 110432
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_199_27
timestamp 1586364061
transform 1 0 3588 0 1 110432
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_198_44
timestamp 1586364061
transform 1 0 5152 0 -1 110432
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_199_39
timestamp 1586364061
transform 1 0 4692 0 1 110432
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_199_51
timestamp 1586364061
transform 1 0 5796 0 1 110432
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1408
timestamp 1586364061
transform 1 0 6716 0 1 110432
box -38 -48 130 592
use scs8hd_decap_12  FILLER_198_56
timestamp 1586364061
transform 1 0 6256 0 -1 110432
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_198_68
timestamp 1586364061
transform 1 0 7360 0 -1 110432
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_199_59
timestamp 1586364061
transform 1 0 6532 0 1 110432
box -38 -48 222 592
use scs8hd_decap_12  FILLER_199_62
timestamp 1586364061
transform 1 0 6808 0 1 110432
box -38 -48 1142 592
use scs8hd_decap_3  PHY_397
timestamp 1586364061
transform -1 0 8832 0 -1 110432
box -38 -48 314 592
use scs8hd_decap_3  PHY_399
timestamp 1586364061
transform -1 0 8832 0 1 110432
box -38 -48 314 592
use scs8hd_fill_1  FILLER_198_80
timestamp 1586364061
transform 1 0 8464 0 -1 110432
box -38 -48 130 592
use scs8hd_decap_6  FILLER_199_74
timestamp 1586364061
transform 1 0 7912 0 1 110432
box -38 -48 590 592
use scs8hd_fill_1  FILLER_199_80
timestamp 1586364061
transform 1 0 8464 0 1 110432
box -38 -48 130 592
use scs8hd_decap_3  PHY_400
timestamp 1586364061
transform 1 0 1104 0 -1 111520
box -38 -48 314 592
use scs8hd_decap_12  FILLER_200_3
timestamp 1586364061
transform 1 0 1380 0 -1 111520
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_200_15
timestamp 1586364061
transform 1 0 2484 0 -1 111520
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1409
timestamp 1586364061
transform 1 0 3956 0 -1 111520
box -38 -48 130 592
use scs8hd_decap_4  FILLER_200_27
timestamp 1586364061
transform 1 0 3588 0 -1 111520
box -38 -48 406 592
use scs8hd_decap_12  FILLER_200_32
timestamp 1586364061
transform 1 0 4048 0 -1 111520
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_200_44
timestamp 1586364061
transform 1 0 5152 0 -1 111520
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_200_56
timestamp 1586364061
transform 1 0 6256 0 -1 111520
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_200_68
timestamp 1586364061
transform 1 0 7360 0 -1 111520
box -38 -48 1142 592
use scs8hd_decap_3  PHY_401
timestamp 1586364061
transform -1 0 8832 0 -1 111520
box -38 -48 314 592
use scs8hd_fill_1  FILLER_200_80
timestamp 1586364061
transform 1 0 8464 0 -1 111520
box -38 -48 130 592
use scs8hd_decap_3  PHY_402
timestamp 1586364061
transform 1 0 1104 0 1 111520
box -38 -48 314 592
use scs8hd_decap_12  FILLER_201_3
timestamp 1586364061
transform 1 0 1380 0 1 111520
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_201_15
timestamp 1586364061
transform 1 0 2484 0 1 111520
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_201_27
timestamp 1586364061
transform 1 0 3588 0 1 111520
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_201_39
timestamp 1586364061
transform 1 0 4692 0 1 111520
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_201_51
timestamp 1586364061
transform 1 0 5796 0 1 111520
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1410
timestamp 1586364061
transform 1 0 6716 0 1 111520
box -38 -48 130 592
use scs8hd_fill_2  FILLER_201_59
timestamp 1586364061
transform 1 0 6532 0 1 111520
box -38 -48 222 592
use scs8hd_decap_12  FILLER_201_62
timestamp 1586364061
transform 1 0 6808 0 1 111520
box -38 -48 1142 592
use scs8hd_decap_3  PHY_403
timestamp 1586364061
transform -1 0 8832 0 1 111520
box -38 -48 314 592
use scs8hd_decap_6  FILLER_201_74
timestamp 1586364061
transform 1 0 7912 0 1 111520
box -38 -48 590 592
use scs8hd_fill_1  FILLER_201_80
timestamp 1586364061
transform 1 0 8464 0 1 111520
box -38 -48 130 592
use scs8hd_decap_3  PHY_404
timestamp 1586364061
transform 1 0 1104 0 -1 112608
box -38 -48 314 592
use scs8hd_decap_12  FILLER_202_3
timestamp 1586364061
transform 1 0 1380 0 -1 112608
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_202_15
timestamp 1586364061
transform 1 0 2484 0 -1 112608
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1411
timestamp 1586364061
transform 1 0 3956 0 -1 112608
box -38 -48 130 592
use scs8hd_decap_4  FILLER_202_27
timestamp 1586364061
transform 1 0 3588 0 -1 112608
box -38 -48 406 592
use scs8hd_decap_12  FILLER_202_32
timestamp 1586364061
transform 1 0 4048 0 -1 112608
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_202_44
timestamp 1586364061
transform 1 0 5152 0 -1 112608
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_202_56
timestamp 1586364061
transform 1 0 6256 0 -1 112608
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_202_68
timestamp 1586364061
transform 1 0 7360 0 -1 112608
box -38 -48 1142 592
use scs8hd_decap_3  PHY_405
timestamp 1586364061
transform -1 0 8832 0 -1 112608
box -38 -48 314 592
use scs8hd_fill_1  FILLER_202_80
timestamp 1586364061
transform 1 0 8464 0 -1 112608
box -38 -48 130 592
use scs8hd_decap_3  PHY_406
timestamp 1586364061
transform 1 0 1104 0 1 112608
box -38 -48 314 592
use scs8hd_decap_12  FILLER_203_3
timestamp 1586364061
transform 1 0 1380 0 1 112608
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_203_15
timestamp 1586364061
transform 1 0 2484 0 1 112608
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_203_27
timestamp 1586364061
transform 1 0 3588 0 1 112608
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_203_39
timestamp 1586364061
transform 1 0 4692 0 1 112608
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_203_51
timestamp 1586364061
transform 1 0 5796 0 1 112608
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1412
timestamp 1586364061
transform 1 0 6716 0 1 112608
box -38 -48 130 592
use scs8hd_fill_2  FILLER_203_59
timestamp 1586364061
transform 1 0 6532 0 1 112608
box -38 -48 222 592
use scs8hd_decap_12  FILLER_203_62
timestamp 1586364061
transform 1 0 6808 0 1 112608
box -38 -48 1142 592
use scs8hd_decap_3  PHY_407
timestamp 1586364061
transform -1 0 8832 0 1 112608
box -38 -48 314 592
use scs8hd_decap_6  FILLER_203_74
timestamp 1586364061
transform 1 0 7912 0 1 112608
box -38 -48 590 592
use scs8hd_fill_1  FILLER_203_80
timestamp 1586364061
transform 1 0 8464 0 1 112608
box -38 -48 130 592
use scs8hd_decap_3  PHY_408
timestamp 1586364061
transform 1 0 1104 0 -1 113696
box -38 -48 314 592
use scs8hd_decap_3  PHY_410
timestamp 1586364061
transform 1 0 1104 0 1 113696
box -38 -48 314 592
use scs8hd_decap_12  FILLER_204_3
timestamp 1586364061
transform 1 0 1380 0 -1 113696
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_204_15
timestamp 1586364061
transform 1 0 2484 0 -1 113696
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_205_3
timestamp 1586364061
transform 1 0 1380 0 1 113696
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_205_15
timestamp 1586364061
transform 1 0 2484 0 1 113696
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1413
timestamp 1586364061
transform 1 0 3956 0 -1 113696
box -38 -48 130 592
use scs8hd_decap_4  FILLER_204_27
timestamp 1586364061
transform 1 0 3588 0 -1 113696
box -38 -48 406 592
use scs8hd_decap_12  FILLER_204_32
timestamp 1586364061
transform 1 0 4048 0 -1 113696
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_205_27
timestamp 1586364061
transform 1 0 3588 0 1 113696
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_204_44
timestamp 1586364061
transform 1 0 5152 0 -1 113696
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_205_39
timestamp 1586364061
transform 1 0 4692 0 1 113696
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_205_51
timestamp 1586364061
transform 1 0 5796 0 1 113696
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1414
timestamp 1586364061
transform 1 0 6716 0 1 113696
box -38 -48 130 592
use scs8hd_decap_12  FILLER_204_56
timestamp 1586364061
transform 1 0 6256 0 -1 113696
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_204_68
timestamp 1586364061
transform 1 0 7360 0 -1 113696
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_205_59
timestamp 1586364061
transform 1 0 6532 0 1 113696
box -38 -48 222 592
use scs8hd_decap_12  FILLER_205_62
timestamp 1586364061
transform 1 0 6808 0 1 113696
box -38 -48 1142 592
use scs8hd_decap_3  PHY_409
timestamp 1586364061
transform -1 0 8832 0 -1 113696
box -38 -48 314 592
use scs8hd_decap_3  PHY_411
timestamp 1586364061
transform -1 0 8832 0 1 113696
box -38 -48 314 592
use scs8hd_fill_1  FILLER_204_80
timestamp 1586364061
transform 1 0 8464 0 -1 113696
box -38 -48 130 592
use scs8hd_decap_6  FILLER_205_74
timestamp 1586364061
transform 1 0 7912 0 1 113696
box -38 -48 590 592
use scs8hd_fill_1  FILLER_205_80
timestamp 1586364061
transform 1 0 8464 0 1 113696
box -38 -48 130 592
use scs8hd_decap_3  PHY_412
timestamp 1586364061
transform 1 0 1104 0 -1 114784
box -38 -48 314 592
use scs8hd_decap_12  FILLER_206_3
timestamp 1586364061
transform 1 0 1380 0 -1 114784
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_206_15
timestamp 1586364061
transform 1 0 2484 0 -1 114784
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1415
timestamp 1586364061
transform 1 0 3956 0 -1 114784
box -38 -48 130 592
use scs8hd_decap_4  FILLER_206_27
timestamp 1586364061
transform 1 0 3588 0 -1 114784
box -38 -48 406 592
use scs8hd_decap_12  FILLER_206_32
timestamp 1586364061
transform 1 0 4048 0 -1 114784
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_206_44
timestamp 1586364061
transform 1 0 5152 0 -1 114784
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_206_56
timestamp 1586364061
transform 1 0 6256 0 -1 114784
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_206_68
timestamp 1586364061
transform 1 0 7360 0 -1 114784
box -38 -48 1142 592
use scs8hd_decap_3  PHY_413
timestamp 1586364061
transform -1 0 8832 0 -1 114784
box -38 -48 314 592
use scs8hd_fill_1  FILLER_206_80
timestamp 1586364061
transform 1 0 8464 0 -1 114784
box -38 -48 130 592
use scs8hd_decap_3  PHY_414
timestamp 1586364061
transform 1 0 1104 0 1 114784
box -38 -48 314 592
use scs8hd_decap_12  FILLER_207_3
timestamp 1586364061
transform 1 0 1380 0 1 114784
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_207_15
timestamp 1586364061
transform 1 0 2484 0 1 114784
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_207_27
timestamp 1586364061
transform 1 0 3588 0 1 114784
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_207_39
timestamp 1586364061
transform 1 0 4692 0 1 114784
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_207_51
timestamp 1586364061
transform 1 0 5796 0 1 114784
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1416
timestamp 1586364061
transform 1 0 6716 0 1 114784
box -38 -48 130 592
use scs8hd_fill_2  FILLER_207_59
timestamp 1586364061
transform 1 0 6532 0 1 114784
box -38 -48 222 592
use scs8hd_decap_12  FILLER_207_62
timestamp 1586364061
transform 1 0 6808 0 1 114784
box -38 -48 1142 592
use scs8hd_decap_3  PHY_415
timestamp 1586364061
transform -1 0 8832 0 1 114784
box -38 -48 314 592
use scs8hd_decap_6  FILLER_207_74
timestamp 1586364061
transform 1 0 7912 0 1 114784
box -38 -48 590 592
use scs8hd_fill_1  FILLER_207_80
timestamp 1586364061
transform 1 0 8464 0 1 114784
box -38 -48 130 592
use scs8hd_decap_3  PHY_416
timestamp 1586364061
transform 1 0 1104 0 -1 115872
box -38 -48 314 592
use scs8hd_decap_12  FILLER_208_3
timestamp 1586364061
transform 1 0 1380 0 -1 115872
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_208_15
timestamp 1586364061
transform 1 0 2484 0 -1 115872
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1417
timestamp 1586364061
transform 1 0 3956 0 -1 115872
box -38 -48 130 592
use scs8hd_decap_4  FILLER_208_27
timestamp 1586364061
transform 1 0 3588 0 -1 115872
box -38 -48 406 592
use scs8hd_decap_12  FILLER_208_32
timestamp 1586364061
transform 1 0 4048 0 -1 115872
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_208_44
timestamp 1586364061
transform 1 0 5152 0 -1 115872
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_208_56
timestamp 1586364061
transform 1 0 6256 0 -1 115872
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_208_68
timestamp 1586364061
transform 1 0 7360 0 -1 115872
box -38 -48 1142 592
use scs8hd_decap_3  PHY_417
timestamp 1586364061
transform -1 0 8832 0 -1 115872
box -38 -48 314 592
use scs8hd_fill_1  FILLER_208_80
timestamp 1586364061
transform 1 0 8464 0 -1 115872
box -38 -48 130 592
use scs8hd_decap_3  PHY_418
timestamp 1586364061
transform 1 0 1104 0 1 115872
box -38 -48 314 592
use scs8hd_decap_12  FILLER_209_3
timestamp 1586364061
transform 1 0 1380 0 1 115872
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_209_15
timestamp 1586364061
transform 1 0 2484 0 1 115872
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_209_27
timestamp 1586364061
transform 1 0 3588 0 1 115872
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_209_39
timestamp 1586364061
transform 1 0 4692 0 1 115872
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_209_51
timestamp 1586364061
transform 1 0 5796 0 1 115872
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1418
timestamp 1586364061
transform 1 0 6716 0 1 115872
box -38 -48 130 592
use scs8hd_fill_2  FILLER_209_59
timestamp 1586364061
transform 1 0 6532 0 1 115872
box -38 -48 222 592
use scs8hd_decap_12  FILLER_209_62
timestamp 1586364061
transform 1 0 6808 0 1 115872
box -38 -48 1142 592
use scs8hd_decap_3  PHY_419
timestamp 1586364061
transform -1 0 8832 0 1 115872
box -38 -48 314 592
use scs8hd_decap_6  FILLER_209_74
timestamp 1586364061
transform 1 0 7912 0 1 115872
box -38 -48 590 592
use scs8hd_fill_1  FILLER_209_80
timestamp 1586364061
transform 1 0 8464 0 1 115872
box -38 -48 130 592
use scs8hd_decap_3  PHY_420
timestamp 1586364061
transform 1 0 1104 0 -1 116960
box -38 -48 314 592
use scs8hd_decap_12  FILLER_210_3
timestamp 1586364061
transform 1 0 1380 0 -1 116960
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_210_15
timestamp 1586364061
transform 1 0 2484 0 -1 116960
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1419
timestamp 1586364061
transform 1 0 3956 0 -1 116960
box -38 -48 130 592
use scs8hd_decap_4  FILLER_210_27
timestamp 1586364061
transform 1 0 3588 0 -1 116960
box -38 -48 406 592
use scs8hd_decap_12  FILLER_210_32
timestamp 1586364061
transform 1 0 4048 0 -1 116960
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_210_44
timestamp 1586364061
transform 1 0 5152 0 -1 116960
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_210_56
timestamp 1586364061
transform 1 0 6256 0 -1 116960
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_210_68
timestamp 1586364061
transform 1 0 7360 0 -1 116960
box -38 -48 1142 592
use scs8hd_decap_3  PHY_421
timestamp 1586364061
transform -1 0 8832 0 -1 116960
box -38 -48 314 592
use scs8hd_fill_1  FILLER_210_80
timestamp 1586364061
transform 1 0 8464 0 -1 116960
box -38 -48 130 592
use scs8hd_decap_3  PHY_422
timestamp 1586364061
transform 1 0 1104 0 1 116960
box -38 -48 314 592
use scs8hd_decap_3  PHY_424
timestamp 1586364061
transform 1 0 1104 0 -1 118048
box -38 -48 314 592
use scs8hd_decap_12  FILLER_211_3
timestamp 1586364061
transform 1 0 1380 0 1 116960
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_211_15
timestamp 1586364061
transform 1 0 2484 0 1 116960
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_212_3
timestamp 1586364061
transform 1 0 1380 0 -1 118048
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_212_15
timestamp 1586364061
transform 1 0 2484 0 -1 118048
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1421
timestamp 1586364061
transform 1 0 3956 0 -1 118048
box -38 -48 130 592
use scs8hd_decap_12  FILLER_211_27
timestamp 1586364061
transform 1 0 3588 0 1 116960
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_212_27
timestamp 1586364061
transform 1 0 3588 0 -1 118048
box -38 -48 406 592
use scs8hd_decap_12  FILLER_212_32
timestamp 1586364061
transform 1 0 4048 0 -1 118048
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_211_39
timestamp 1586364061
transform 1 0 4692 0 1 116960
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_211_51
timestamp 1586364061
transform 1 0 5796 0 1 116960
box -38 -48 774 592
use scs8hd_decap_12  FILLER_212_44
timestamp 1586364061
transform 1 0 5152 0 -1 118048
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1420
timestamp 1586364061
transform 1 0 6716 0 1 116960
box -38 -48 130 592
use scs8hd_fill_2  FILLER_211_59
timestamp 1586364061
transform 1 0 6532 0 1 116960
box -38 -48 222 592
use scs8hd_decap_12  FILLER_211_62
timestamp 1586364061
transform 1 0 6808 0 1 116960
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_212_56
timestamp 1586364061
transform 1 0 6256 0 -1 118048
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_212_68
timestamp 1586364061
transform 1 0 7360 0 -1 118048
box -38 -48 1142 592
use scs8hd_decap_3  PHY_423
timestamp 1586364061
transform -1 0 8832 0 1 116960
box -38 -48 314 592
use scs8hd_decap_3  PHY_425
timestamp 1586364061
transform -1 0 8832 0 -1 118048
box -38 -48 314 592
use scs8hd_decap_6  FILLER_211_74
timestamp 1586364061
transform 1 0 7912 0 1 116960
box -38 -48 590 592
use scs8hd_fill_1  FILLER_211_80
timestamp 1586364061
transform 1 0 8464 0 1 116960
box -38 -48 130 592
use scs8hd_fill_1  FILLER_212_80
timestamp 1586364061
transform 1 0 8464 0 -1 118048
box -38 -48 130 592
use scs8hd_decap_3  PHY_426
timestamp 1586364061
transform 1 0 1104 0 1 118048
box -38 -48 314 592
use scs8hd_decap_12  FILLER_213_3
timestamp 1586364061
transform 1 0 1380 0 1 118048
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_213_15
timestamp 1586364061
transform 1 0 2484 0 1 118048
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_213_27
timestamp 1586364061
transform 1 0 3588 0 1 118048
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_213_39
timestamp 1586364061
transform 1 0 4692 0 1 118048
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_213_51
timestamp 1586364061
transform 1 0 5796 0 1 118048
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1422
timestamp 1586364061
transform 1 0 6716 0 1 118048
box -38 -48 130 592
use scs8hd_fill_2  FILLER_213_59
timestamp 1586364061
transform 1 0 6532 0 1 118048
box -38 -48 222 592
use scs8hd_decap_12  FILLER_213_62
timestamp 1586364061
transform 1 0 6808 0 1 118048
box -38 -48 1142 592
use scs8hd_decap_3  PHY_427
timestamp 1586364061
transform -1 0 8832 0 1 118048
box -38 -48 314 592
use scs8hd_decap_6  FILLER_213_74
timestamp 1586364061
transform 1 0 7912 0 1 118048
box -38 -48 590 592
use scs8hd_fill_1  FILLER_213_80
timestamp 1586364061
transform 1 0 8464 0 1 118048
box -38 -48 130 592
use scs8hd_decap_3  PHY_428
timestamp 1586364061
transform 1 0 1104 0 -1 119136
box -38 -48 314 592
use scs8hd_decap_12  FILLER_214_3
timestamp 1586364061
transform 1 0 1380 0 -1 119136
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_214_15
timestamp 1586364061
transform 1 0 2484 0 -1 119136
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1423
timestamp 1586364061
transform 1 0 3956 0 -1 119136
box -38 -48 130 592
use scs8hd_decap_4  FILLER_214_27
timestamp 1586364061
transform 1 0 3588 0 -1 119136
box -38 -48 406 592
use scs8hd_decap_12  FILLER_214_32
timestamp 1586364061
transform 1 0 4048 0 -1 119136
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_214_44
timestamp 1586364061
transform 1 0 5152 0 -1 119136
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_214_56
timestamp 1586364061
transform 1 0 6256 0 -1 119136
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_214_68
timestamp 1586364061
transform 1 0 7360 0 -1 119136
box -38 -48 1142 592
use scs8hd_decap_3  PHY_429
timestamp 1586364061
transform -1 0 8832 0 -1 119136
box -38 -48 314 592
use scs8hd_fill_1  FILLER_214_80
timestamp 1586364061
transform 1 0 8464 0 -1 119136
box -38 -48 130 592
use scs8hd_decap_3  PHY_430
timestamp 1586364061
transform 1 0 1104 0 1 119136
box -38 -48 314 592
use scs8hd_decap_12  FILLER_215_3
timestamp 1586364061
transform 1 0 1380 0 1 119136
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_215_15
timestamp 1586364061
transform 1 0 2484 0 1 119136
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_215_27
timestamp 1586364061
transform 1 0 3588 0 1 119136
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_215_39
timestamp 1586364061
transform 1 0 4692 0 1 119136
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_215_51
timestamp 1586364061
transform 1 0 5796 0 1 119136
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1424
timestamp 1586364061
transform 1 0 6716 0 1 119136
box -38 -48 130 592
use scs8hd_fill_2  FILLER_215_59
timestamp 1586364061
transform 1 0 6532 0 1 119136
box -38 -48 222 592
use scs8hd_decap_12  FILLER_215_62
timestamp 1586364061
transform 1 0 6808 0 1 119136
box -38 -48 1142 592
use scs8hd_decap_3  PHY_431
timestamp 1586364061
transform -1 0 8832 0 1 119136
box -38 -48 314 592
use scs8hd_decap_6  FILLER_215_74
timestamp 1586364061
transform 1 0 7912 0 1 119136
box -38 -48 590 592
use scs8hd_fill_1  FILLER_215_80
timestamp 1586364061
transform 1 0 8464 0 1 119136
box -38 -48 130 592
use scs8hd_decap_3  PHY_432
timestamp 1586364061
transform 1 0 1104 0 -1 120224
box -38 -48 314 592
use scs8hd_decap_12  FILLER_216_3
timestamp 1586364061
transform 1 0 1380 0 -1 120224
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_216_15
timestamp 1586364061
transform 1 0 2484 0 -1 120224
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1425
timestamp 1586364061
transform 1 0 3956 0 -1 120224
box -38 -48 130 592
use scs8hd_decap_4  FILLER_216_27
timestamp 1586364061
transform 1 0 3588 0 -1 120224
box -38 -48 406 592
use scs8hd_decap_12  FILLER_216_32
timestamp 1586364061
transform 1 0 4048 0 -1 120224
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_216_44
timestamp 1586364061
transform 1 0 5152 0 -1 120224
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_216_56
timestamp 1586364061
transform 1 0 6256 0 -1 120224
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_216_68
timestamp 1586364061
transform 1 0 7360 0 -1 120224
box -38 -48 1142 592
use scs8hd_decap_3  PHY_433
timestamp 1586364061
transform -1 0 8832 0 -1 120224
box -38 -48 314 592
use scs8hd_fill_1  FILLER_216_80
timestamp 1586364061
transform 1 0 8464 0 -1 120224
box -38 -48 130 592
use scs8hd_decap_3  PHY_434
timestamp 1586364061
transform 1 0 1104 0 1 120224
box -38 -48 314 592
use scs8hd_decap_12  FILLER_217_3
timestamp 1586364061
transform 1 0 1380 0 1 120224
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_217_15
timestamp 1586364061
transform 1 0 2484 0 1 120224
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_217_27
timestamp 1586364061
transform 1 0 3588 0 1 120224
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_217_39
timestamp 1586364061
transform 1 0 4692 0 1 120224
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_217_51
timestamp 1586364061
transform 1 0 5796 0 1 120224
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1426
timestamp 1586364061
transform 1 0 6716 0 1 120224
box -38 -48 130 592
use scs8hd_fill_2  FILLER_217_59
timestamp 1586364061
transform 1 0 6532 0 1 120224
box -38 -48 222 592
use scs8hd_decap_12  FILLER_217_62
timestamp 1586364061
transform 1 0 6808 0 1 120224
box -38 -48 1142 592
use scs8hd_decap_3  PHY_435
timestamp 1586364061
transform -1 0 8832 0 1 120224
box -38 -48 314 592
use scs8hd_decap_6  FILLER_217_74
timestamp 1586364061
transform 1 0 7912 0 1 120224
box -38 -48 590 592
use scs8hd_fill_1  FILLER_217_80
timestamp 1586364061
transform 1 0 8464 0 1 120224
box -38 -48 130 592
use scs8hd_decap_3  PHY_436
timestamp 1586364061
transform 1 0 1104 0 -1 121312
box -38 -48 314 592
use scs8hd_decap_3  PHY_438
timestamp 1586364061
transform 1 0 1104 0 1 121312
box -38 -48 314 592
use scs8hd_decap_12  FILLER_218_3
timestamp 1586364061
transform 1 0 1380 0 -1 121312
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_218_15
timestamp 1586364061
transform 1 0 2484 0 -1 121312
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_219_3
timestamp 1586364061
transform 1 0 1380 0 1 121312
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_219_15
timestamp 1586364061
transform 1 0 2484 0 1 121312
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1427
timestamp 1586364061
transform 1 0 3956 0 -1 121312
box -38 -48 130 592
use scs8hd_decap_4  FILLER_218_27
timestamp 1586364061
transform 1 0 3588 0 -1 121312
box -38 -48 406 592
use scs8hd_decap_12  FILLER_218_32
timestamp 1586364061
transform 1 0 4048 0 -1 121312
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_219_27
timestamp 1586364061
transform 1 0 3588 0 1 121312
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_218_44
timestamp 1586364061
transform 1 0 5152 0 -1 121312
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_219_39
timestamp 1586364061
transform 1 0 4692 0 1 121312
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_219_51
timestamp 1586364061
transform 1 0 5796 0 1 121312
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1428
timestamp 1586364061
transform 1 0 6716 0 1 121312
box -38 -48 130 592
use scs8hd_decap_12  FILLER_218_56
timestamp 1586364061
transform 1 0 6256 0 -1 121312
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_218_68
timestamp 1586364061
transform 1 0 7360 0 -1 121312
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_219_59
timestamp 1586364061
transform 1 0 6532 0 1 121312
box -38 -48 222 592
use scs8hd_decap_12  FILLER_219_62
timestamp 1586364061
transform 1 0 6808 0 1 121312
box -38 -48 1142 592
use scs8hd_decap_3  PHY_437
timestamp 1586364061
transform -1 0 8832 0 -1 121312
box -38 -48 314 592
use scs8hd_decap_3  PHY_439
timestamp 1586364061
transform -1 0 8832 0 1 121312
box -38 -48 314 592
use scs8hd_fill_1  FILLER_218_80
timestamp 1586364061
transform 1 0 8464 0 -1 121312
box -38 -48 130 592
use scs8hd_decap_6  FILLER_219_74
timestamp 1586364061
transform 1 0 7912 0 1 121312
box -38 -48 590 592
use scs8hd_fill_1  FILLER_219_80
timestamp 1586364061
transform 1 0 8464 0 1 121312
box -38 -48 130 592
use scs8hd_decap_3  PHY_440
timestamp 1586364061
transform 1 0 1104 0 -1 122400
box -38 -48 314 592
use scs8hd_decap_12  FILLER_220_3
timestamp 1586364061
transform 1 0 1380 0 -1 122400
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_220_15
timestamp 1586364061
transform 1 0 2484 0 -1 122400
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1429
timestamp 1586364061
transform 1 0 3956 0 -1 122400
box -38 -48 130 592
use scs8hd_decap_4  FILLER_220_27
timestamp 1586364061
transform 1 0 3588 0 -1 122400
box -38 -48 406 592
use scs8hd_decap_12  FILLER_220_32
timestamp 1586364061
transform 1 0 4048 0 -1 122400
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_220_44
timestamp 1586364061
transform 1 0 5152 0 -1 122400
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_220_56
timestamp 1586364061
transform 1 0 6256 0 -1 122400
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_220_68
timestamp 1586364061
transform 1 0 7360 0 -1 122400
box -38 -48 1142 592
use scs8hd_decap_3  PHY_441
timestamp 1586364061
transform -1 0 8832 0 -1 122400
box -38 -48 314 592
use scs8hd_fill_1  FILLER_220_80
timestamp 1586364061
transform 1 0 8464 0 -1 122400
box -38 -48 130 592
use scs8hd_decap_3  PHY_442
timestamp 1586364061
transform 1 0 1104 0 1 122400
box -38 -48 314 592
use scs8hd_decap_12  FILLER_221_3
timestamp 1586364061
transform 1 0 1380 0 1 122400
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_221_15
timestamp 1586364061
transform 1 0 2484 0 1 122400
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_221_27
timestamp 1586364061
transform 1 0 3588 0 1 122400
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_221_39
timestamp 1586364061
transform 1 0 4692 0 1 122400
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_221_51
timestamp 1586364061
transform 1 0 5796 0 1 122400
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1430
timestamp 1586364061
transform 1 0 6716 0 1 122400
box -38 -48 130 592
use scs8hd_fill_2  FILLER_221_59
timestamp 1586364061
transform 1 0 6532 0 1 122400
box -38 -48 222 592
use scs8hd_decap_12  FILLER_221_62
timestamp 1586364061
transform 1 0 6808 0 1 122400
box -38 -48 1142 592
use scs8hd_decap_3  PHY_443
timestamp 1586364061
transform -1 0 8832 0 1 122400
box -38 -48 314 592
use scs8hd_decap_6  FILLER_221_74
timestamp 1586364061
transform 1 0 7912 0 1 122400
box -38 -48 590 592
use scs8hd_fill_1  FILLER_221_80
timestamp 1586364061
transform 1 0 8464 0 1 122400
box -38 -48 130 592
use scs8hd_decap_3  PHY_444
timestamp 1586364061
transform 1 0 1104 0 -1 123488
box -38 -48 314 592
use scs8hd_decap_12  FILLER_222_3
timestamp 1586364061
transform 1 0 1380 0 -1 123488
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_222_15
timestamp 1586364061
transform 1 0 2484 0 -1 123488
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1431
timestamp 1586364061
transform 1 0 3956 0 -1 123488
box -38 -48 130 592
use scs8hd_decap_4  FILLER_222_27
timestamp 1586364061
transform 1 0 3588 0 -1 123488
box -38 -48 406 592
use scs8hd_decap_12  FILLER_222_32
timestamp 1586364061
transform 1 0 4048 0 -1 123488
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_222_44
timestamp 1586364061
transform 1 0 5152 0 -1 123488
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_222_56
timestamp 1586364061
transform 1 0 6256 0 -1 123488
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_222_68
timestamp 1586364061
transform 1 0 7360 0 -1 123488
box -38 -48 1142 592
use scs8hd_decap_3  PHY_445
timestamp 1586364061
transform -1 0 8832 0 -1 123488
box -38 -48 314 592
use scs8hd_fill_1  FILLER_222_80
timestamp 1586364061
transform 1 0 8464 0 -1 123488
box -38 -48 130 592
use scs8hd_decap_3  PHY_446
timestamp 1586364061
transform 1 0 1104 0 1 123488
box -38 -48 314 592
use scs8hd_decap_12  FILLER_223_3
timestamp 1586364061
transform 1 0 1380 0 1 123488
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_223_15
timestamp 1586364061
transform 1 0 2484 0 1 123488
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_223_27
timestamp 1586364061
transform 1 0 3588 0 1 123488
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_223_39
timestamp 1586364061
transform 1 0 4692 0 1 123488
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_223_51
timestamp 1586364061
transform 1 0 5796 0 1 123488
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1432
timestamp 1586364061
transform 1 0 6716 0 1 123488
box -38 -48 130 592
use scs8hd_fill_2  FILLER_223_59
timestamp 1586364061
transform 1 0 6532 0 1 123488
box -38 -48 222 592
use scs8hd_decap_12  FILLER_223_62
timestamp 1586364061
transform 1 0 6808 0 1 123488
box -38 -48 1142 592
use scs8hd_decap_3  PHY_447
timestamp 1586364061
transform -1 0 8832 0 1 123488
box -38 -48 314 592
use scs8hd_decap_6  FILLER_223_74
timestamp 1586364061
transform 1 0 7912 0 1 123488
box -38 -48 590 592
use scs8hd_fill_1  FILLER_223_80
timestamp 1586364061
transform 1 0 8464 0 1 123488
box -38 -48 130 592
use scs8hd_decap_3  PHY_448
timestamp 1586364061
transform 1 0 1104 0 -1 124576
box -38 -48 314 592
use scs8hd_decap_3  PHY_450
timestamp 1586364061
transform 1 0 1104 0 1 124576
box -38 -48 314 592
use scs8hd_decap_12  FILLER_224_3
timestamp 1586364061
transform 1 0 1380 0 -1 124576
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_224_15
timestamp 1586364061
transform 1 0 2484 0 -1 124576
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_225_3
timestamp 1586364061
transform 1 0 1380 0 1 124576
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_225_15
timestamp 1586364061
transform 1 0 2484 0 1 124576
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1433
timestamp 1586364061
transform 1 0 3956 0 -1 124576
box -38 -48 130 592
use scs8hd_decap_4  FILLER_224_27
timestamp 1586364061
transform 1 0 3588 0 -1 124576
box -38 -48 406 592
use scs8hd_decap_12  FILLER_224_32
timestamp 1586364061
transform 1 0 4048 0 -1 124576
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_225_27
timestamp 1586364061
transform 1 0 3588 0 1 124576
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_224_44
timestamp 1586364061
transform 1 0 5152 0 -1 124576
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_225_39
timestamp 1586364061
transform 1 0 4692 0 1 124576
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_225_51
timestamp 1586364061
transform 1 0 5796 0 1 124576
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1434
timestamp 1586364061
transform 1 0 6716 0 1 124576
box -38 -48 130 592
use scs8hd_decap_12  FILLER_224_56
timestamp 1586364061
transform 1 0 6256 0 -1 124576
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_224_68
timestamp 1586364061
transform 1 0 7360 0 -1 124576
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_225_59
timestamp 1586364061
transform 1 0 6532 0 1 124576
box -38 -48 222 592
use scs8hd_decap_12  FILLER_225_62
timestamp 1586364061
transform 1 0 6808 0 1 124576
box -38 -48 1142 592
use scs8hd_decap_3  PHY_449
timestamp 1586364061
transform -1 0 8832 0 -1 124576
box -38 -48 314 592
use scs8hd_decap_3  PHY_451
timestamp 1586364061
transform -1 0 8832 0 1 124576
box -38 -48 314 592
use scs8hd_fill_1  FILLER_224_80
timestamp 1586364061
transform 1 0 8464 0 -1 124576
box -38 -48 130 592
use scs8hd_decap_6  FILLER_225_74
timestamp 1586364061
transform 1 0 7912 0 1 124576
box -38 -48 590 592
use scs8hd_fill_1  FILLER_225_80
timestamp 1586364061
transform 1 0 8464 0 1 124576
box -38 -48 130 592
use scs8hd_decap_3  PHY_452
timestamp 1586364061
transform 1 0 1104 0 -1 125664
box -38 -48 314 592
use scs8hd_decap_12  FILLER_226_3
timestamp 1586364061
transform 1 0 1380 0 -1 125664
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_226_15
timestamp 1586364061
transform 1 0 2484 0 -1 125664
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1435
timestamp 1586364061
transform 1 0 3956 0 -1 125664
box -38 -48 130 592
use scs8hd_decap_4  FILLER_226_27
timestamp 1586364061
transform 1 0 3588 0 -1 125664
box -38 -48 406 592
use scs8hd_decap_12  FILLER_226_32
timestamp 1586364061
transform 1 0 4048 0 -1 125664
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_226_44
timestamp 1586364061
transform 1 0 5152 0 -1 125664
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_226_56
timestamp 1586364061
transform 1 0 6256 0 -1 125664
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_226_68
timestamp 1586364061
transform 1 0 7360 0 -1 125664
box -38 -48 1142 592
use scs8hd_decap_3  PHY_453
timestamp 1586364061
transform -1 0 8832 0 -1 125664
box -38 -48 314 592
use scs8hd_fill_1  FILLER_226_80
timestamp 1586364061
transform 1 0 8464 0 -1 125664
box -38 -48 130 592
use scs8hd_decap_3  PHY_454
timestamp 1586364061
transform 1 0 1104 0 1 125664
box -38 -48 314 592
use scs8hd_decap_12  FILLER_227_3
timestamp 1586364061
transform 1 0 1380 0 1 125664
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_227_15
timestamp 1586364061
transform 1 0 2484 0 1 125664
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_227_27
timestamp 1586364061
transform 1 0 3588 0 1 125664
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_227_39
timestamp 1586364061
transform 1 0 4692 0 1 125664
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_227_51
timestamp 1586364061
transform 1 0 5796 0 1 125664
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1436
timestamp 1586364061
transform 1 0 6716 0 1 125664
box -38 -48 130 592
use scs8hd_fill_2  FILLER_227_59
timestamp 1586364061
transform 1 0 6532 0 1 125664
box -38 -48 222 592
use scs8hd_decap_12  FILLER_227_62
timestamp 1586364061
transform 1 0 6808 0 1 125664
box -38 -48 1142 592
use scs8hd_decap_3  PHY_455
timestamp 1586364061
transform -1 0 8832 0 1 125664
box -38 -48 314 592
use scs8hd_decap_6  FILLER_227_74
timestamp 1586364061
transform 1 0 7912 0 1 125664
box -38 -48 590 592
use scs8hd_fill_1  FILLER_227_80
timestamp 1586364061
transform 1 0 8464 0 1 125664
box -38 -48 130 592
use scs8hd_decap_3  PHY_456
timestamp 1586364061
transform 1 0 1104 0 -1 126752
box -38 -48 314 592
use scs8hd_decap_12  FILLER_228_3
timestamp 1586364061
transform 1 0 1380 0 -1 126752
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_228_15
timestamp 1586364061
transform 1 0 2484 0 -1 126752
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1437
timestamp 1586364061
transform 1 0 3956 0 -1 126752
box -38 -48 130 592
use scs8hd_decap_4  FILLER_228_27
timestamp 1586364061
transform 1 0 3588 0 -1 126752
box -38 -48 406 592
use scs8hd_decap_12  FILLER_228_32
timestamp 1586364061
transform 1 0 4048 0 -1 126752
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_228_44
timestamp 1586364061
transform 1 0 5152 0 -1 126752
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_228_56
timestamp 1586364061
transform 1 0 6256 0 -1 126752
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_228_68
timestamp 1586364061
transform 1 0 7360 0 -1 126752
box -38 -48 1142 592
use scs8hd_decap_3  PHY_457
timestamp 1586364061
transform -1 0 8832 0 -1 126752
box -38 -48 314 592
use scs8hd_fill_1  FILLER_228_80
timestamp 1586364061
transform 1 0 8464 0 -1 126752
box -38 -48 130 592
use scs8hd_decap_3  PHY_458
timestamp 1586364061
transform 1 0 1104 0 1 126752
box -38 -48 314 592
use scs8hd_decap_12  FILLER_229_3
timestamp 1586364061
transform 1 0 1380 0 1 126752
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_229_15
timestamp 1586364061
transform 1 0 2484 0 1 126752
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_229_27
timestamp 1586364061
transform 1 0 3588 0 1 126752
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_229_39
timestamp 1586364061
transform 1 0 4692 0 1 126752
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_229_51
timestamp 1586364061
transform 1 0 5796 0 1 126752
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1438
timestamp 1586364061
transform 1 0 6716 0 1 126752
box -38 -48 130 592
use scs8hd_fill_2  FILLER_229_59
timestamp 1586364061
transform 1 0 6532 0 1 126752
box -38 -48 222 592
use scs8hd_decap_12  FILLER_229_62
timestamp 1586364061
transform 1 0 6808 0 1 126752
box -38 -48 1142 592
use scs8hd_decap_3  PHY_459
timestamp 1586364061
transform -1 0 8832 0 1 126752
box -38 -48 314 592
use scs8hd_decap_6  FILLER_229_74
timestamp 1586364061
transform 1 0 7912 0 1 126752
box -38 -48 590 592
use scs8hd_fill_1  FILLER_229_80
timestamp 1586364061
transform 1 0 8464 0 1 126752
box -38 -48 130 592
use scs8hd_decap_3  PHY_460
timestamp 1586364061
transform 1 0 1104 0 -1 127840
box -38 -48 314 592
use scs8hd_decap_12  FILLER_230_3
timestamp 1586364061
transform 1 0 1380 0 -1 127840
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_230_15
timestamp 1586364061
transform 1 0 2484 0 -1 127840
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1439
timestamp 1586364061
transform 1 0 3956 0 -1 127840
box -38 -48 130 592
use scs8hd_decap_4  FILLER_230_27
timestamp 1586364061
transform 1 0 3588 0 -1 127840
box -38 -48 406 592
use scs8hd_decap_12  FILLER_230_32
timestamp 1586364061
transform 1 0 4048 0 -1 127840
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_230_44
timestamp 1586364061
transform 1 0 5152 0 -1 127840
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_230_56
timestamp 1586364061
transform 1 0 6256 0 -1 127840
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_230_68
timestamp 1586364061
transform 1 0 7360 0 -1 127840
box -38 -48 1142 592
use scs8hd_decap_3  PHY_461
timestamp 1586364061
transform -1 0 8832 0 -1 127840
box -38 -48 314 592
use scs8hd_fill_1  FILLER_230_80
timestamp 1586364061
transform 1 0 8464 0 -1 127840
box -38 -48 130 592
use scs8hd_decap_3  PHY_462
timestamp 1586364061
transform 1 0 1104 0 1 127840
box -38 -48 314 592
use scs8hd_decap_3  PHY_464
timestamp 1586364061
transform 1 0 1104 0 -1 128928
box -38 -48 314 592
use scs8hd_decap_12  FILLER_231_3
timestamp 1586364061
transform 1 0 1380 0 1 127840
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_231_15
timestamp 1586364061
transform 1 0 2484 0 1 127840
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_232_3
timestamp 1586364061
transform 1 0 1380 0 -1 128928
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_232_15
timestamp 1586364061
transform 1 0 2484 0 -1 128928
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1441
timestamp 1586364061
transform 1 0 3956 0 -1 128928
box -38 -48 130 592
use scs8hd_decap_12  FILLER_231_27
timestamp 1586364061
transform 1 0 3588 0 1 127840
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_232_27
timestamp 1586364061
transform 1 0 3588 0 -1 128928
box -38 -48 406 592
use scs8hd_decap_12  FILLER_232_32
timestamp 1586364061
transform 1 0 4048 0 -1 128928
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_231_39
timestamp 1586364061
transform 1 0 4692 0 1 127840
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_231_51
timestamp 1586364061
transform 1 0 5796 0 1 127840
box -38 -48 774 592
use scs8hd_decap_12  FILLER_232_44
timestamp 1586364061
transform 1 0 5152 0 -1 128928
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1440
timestamp 1586364061
transform 1 0 6716 0 1 127840
box -38 -48 130 592
use scs8hd_fill_2  FILLER_231_59
timestamp 1586364061
transform 1 0 6532 0 1 127840
box -38 -48 222 592
use scs8hd_decap_12  FILLER_231_62
timestamp 1586364061
transform 1 0 6808 0 1 127840
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_232_56
timestamp 1586364061
transform 1 0 6256 0 -1 128928
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_232_68
timestamp 1586364061
transform 1 0 7360 0 -1 128928
box -38 -48 1142 592
use scs8hd_decap_3  PHY_463
timestamp 1586364061
transform -1 0 8832 0 1 127840
box -38 -48 314 592
use scs8hd_decap_3  PHY_465
timestamp 1586364061
transform -1 0 8832 0 -1 128928
box -38 -48 314 592
use scs8hd_decap_6  FILLER_231_74
timestamp 1586364061
transform 1 0 7912 0 1 127840
box -38 -48 590 592
use scs8hd_fill_1  FILLER_231_80
timestamp 1586364061
transform 1 0 8464 0 1 127840
box -38 -48 130 592
use scs8hd_fill_1  FILLER_232_80
timestamp 1586364061
transform 1 0 8464 0 -1 128928
box -38 -48 130 592
use scs8hd_decap_3  PHY_466
timestamp 1586364061
transform 1 0 1104 0 1 128928
box -38 -48 314 592
use scs8hd_decap_12  FILLER_233_3
timestamp 1586364061
transform 1 0 1380 0 1 128928
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_233_15
timestamp 1586364061
transform 1 0 2484 0 1 128928
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_233_27
timestamp 1586364061
transform 1 0 3588 0 1 128928
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_233_39
timestamp 1586364061
transform 1 0 4692 0 1 128928
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_233_51
timestamp 1586364061
transform 1 0 5796 0 1 128928
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1442
timestamp 1586364061
transform 1 0 6716 0 1 128928
box -38 -48 130 592
use scs8hd_fill_2  FILLER_233_59
timestamp 1586364061
transform 1 0 6532 0 1 128928
box -38 -48 222 592
use scs8hd_decap_12  FILLER_233_62
timestamp 1586364061
transform 1 0 6808 0 1 128928
box -38 -48 1142 592
use scs8hd_decap_3  PHY_467
timestamp 1586364061
transform -1 0 8832 0 1 128928
box -38 -48 314 592
use scs8hd_decap_6  FILLER_233_74
timestamp 1586364061
transform 1 0 7912 0 1 128928
box -38 -48 590 592
use scs8hd_fill_1  FILLER_233_80
timestamp 1586364061
transform 1 0 8464 0 1 128928
box -38 -48 130 592
use scs8hd_decap_3  PHY_468
timestamp 1586364061
transform 1 0 1104 0 -1 130016
box -38 -48 314 592
use scs8hd_decap_12  FILLER_234_3
timestamp 1586364061
transform 1 0 1380 0 -1 130016
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_234_15
timestamp 1586364061
transform 1 0 2484 0 -1 130016
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1443
timestamp 1586364061
transform 1 0 3956 0 -1 130016
box -38 -48 130 592
use scs8hd_decap_4  FILLER_234_27
timestamp 1586364061
transform 1 0 3588 0 -1 130016
box -38 -48 406 592
use scs8hd_decap_12  FILLER_234_32
timestamp 1586364061
transform 1 0 4048 0 -1 130016
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_234_44
timestamp 1586364061
transform 1 0 5152 0 -1 130016
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_234_56
timestamp 1586364061
transform 1 0 6256 0 -1 130016
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_234_68
timestamp 1586364061
transform 1 0 7360 0 -1 130016
box -38 -48 1142 592
use scs8hd_decap_3  PHY_469
timestamp 1586364061
transform -1 0 8832 0 -1 130016
box -38 -48 314 592
use scs8hd_fill_1  FILLER_234_80
timestamp 1586364061
transform 1 0 8464 0 -1 130016
box -38 -48 130 592
use scs8hd_decap_3  PHY_470
timestamp 1586364061
transform 1 0 1104 0 1 130016
box -38 -48 314 592
use scs8hd_decap_12  FILLER_235_3
timestamp 1586364061
transform 1 0 1380 0 1 130016
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_235_15
timestamp 1586364061
transform 1 0 2484 0 1 130016
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_235_27
timestamp 1586364061
transform 1 0 3588 0 1 130016
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_235_39
timestamp 1586364061
transform 1 0 4692 0 1 130016
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_235_51
timestamp 1586364061
transform 1 0 5796 0 1 130016
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1444
timestamp 1586364061
transform 1 0 6716 0 1 130016
box -38 -48 130 592
use scs8hd_fill_2  FILLER_235_59
timestamp 1586364061
transform 1 0 6532 0 1 130016
box -38 -48 222 592
use scs8hd_decap_12  FILLER_235_62
timestamp 1586364061
transform 1 0 6808 0 1 130016
box -38 -48 1142 592
use scs8hd_decap_3  PHY_471
timestamp 1586364061
transform -1 0 8832 0 1 130016
box -38 -48 314 592
use scs8hd_decap_6  FILLER_235_74
timestamp 1586364061
transform 1 0 7912 0 1 130016
box -38 -48 590 592
use scs8hd_fill_1  FILLER_235_80
timestamp 1586364061
transform 1 0 8464 0 1 130016
box -38 -48 130 592
use scs8hd_decap_3  PHY_472
timestamp 1586364061
transform 1 0 1104 0 -1 131104
box -38 -48 314 592
use scs8hd_decap_12  FILLER_236_3
timestamp 1586364061
transform 1 0 1380 0 -1 131104
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_236_15
timestamp 1586364061
transform 1 0 2484 0 -1 131104
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1445
timestamp 1586364061
transform 1 0 3956 0 -1 131104
box -38 -48 130 592
use scs8hd_decap_4  FILLER_236_27
timestamp 1586364061
transform 1 0 3588 0 -1 131104
box -38 -48 406 592
use scs8hd_decap_12  FILLER_236_32
timestamp 1586364061
transform 1 0 4048 0 -1 131104
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_236_44
timestamp 1586364061
transform 1 0 5152 0 -1 131104
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_236_56
timestamp 1586364061
transform 1 0 6256 0 -1 131104
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_236_68
timestamp 1586364061
transform 1 0 7360 0 -1 131104
box -38 -48 1142 592
use scs8hd_decap_3  PHY_473
timestamp 1586364061
transform -1 0 8832 0 -1 131104
box -38 -48 314 592
use scs8hd_fill_1  FILLER_236_80
timestamp 1586364061
transform 1 0 8464 0 -1 131104
box -38 -48 130 592
use scs8hd_decap_3  PHY_474
timestamp 1586364061
transform 1 0 1104 0 1 131104
box -38 -48 314 592
use scs8hd_decap_3  PHY_476
timestamp 1586364061
transform 1 0 1104 0 -1 132192
box -38 -48 314 592
use scs8hd_decap_12  FILLER_237_3
timestamp 1586364061
transform 1 0 1380 0 1 131104
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_237_15
timestamp 1586364061
transform 1 0 2484 0 1 131104
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_238_3
timestamp 1586364061
transform 1 0 1380 0 -1 132192
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_238_15
timestamp 1586364061
transform 1 0 2484 0 -1 132192
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1447
timestamp 1586364061
transform 1 0 3956 0 -1 132192
box -38 -48 130 592
use scs8hd_decap_12  FILLER_237_27
timestamp 1586364061
transform 1 0 3588 0 1 131104
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_238_27
timestamp 1586364061
transform 1 0 3588 0 -1 132192
box -38 -48 406 592
use scs8hd_decap_12  FILLER_238_32
timestamp 1586364061
transform 1 0 4048 0 -1 132192
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_237_39
timestamp 1586364061
transform 1 0 4692 0 1 131104
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_237_51
timestamp 1586364061
transform 1 0 5796 0 1 131104
box -38 -48 774 592
use scs8hd_decap_12  FILLER_238_44
timestamp 1586364061
transform 1 0 5152 0 -1 132192
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1446
timestamp 1586364061
transform 1 0 6716 0 1 131104
box -38 -48 130 592
use scs8hd_fill_2  FILLER_237_59
timestamp 1586364061
transform 1 0 6532 0 1 131104
box -38 -48 222 592
use scs8hd_decap_12  FILLER_237_62
timestamp 1586364061
transform 1 0 6808 0 1 131104
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_238_56
timestamp 1586364061
transform 1 0 6256 0 -1 132192
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_238_68
timestamp 1586364061
transform 1 0 7360 0 -1 132192
box -38 -48 1142 592
use scs8hd_decap_3  PHY_475
timestamp 1586364061
transform -1 0 8832 0 1 131104
box -38 -48 314 592
use scs8hd_decap_3  PHY_477
timestamp 1586364061
transform -1 0 8832 0 -1 132192
box -38 -48 314 592
use scs8hd_decap_6  FILLER_237_74
timestamp 1586364061
transform 1 0 7912 0 1 131104
box -38 -48 590 592
use scs8hd_fill_1  FILLER_237_80
timestamp 1586364061
transform 1 0 8464 0 1 131104
box -38 -48 130 592
use scs8hd_fill_1  FILLER_238_80
timestamp 1586364061
transform 1 0 8464 0 -1 132192
box -38 -48 130 592
use scs8hd_decap_3  PHY_478
timestamp 1586364061
transform 1 0 1104 0 1 132192
box -38 -48 314 592
use scs8hd_decap_12  FILLER_239_3
timestamp 1586364061
transform 1 0 1380 0 1 132192
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_239_15
timestamp 1586364061
transform 1 0 2484 0 1 132192
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_239_27
timestamp 1586364061
transform 1 0 3588 0 1 132192
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_239_39
timestamp 1586364061
transform 1 0 4692 0 1 132192
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_239_51
timestamp 1586364061
transform 1 0 5796 0 1 132192
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1448
timestamp 1586364061
transform 1 0 6716 0 1 132192
box -38 -48 130 592
use scs8hd_fill_2  FILLER_239_59
timestamp 1586364061
transform 1 0 6532 0 1 132192
box -38 -48 222 592
use scs8hd_decap_12  FILLER_239_62
timestamp 1586364061
transform 1 0 6808 0 1 132192
box -38 -48 1142 592
use scs8hd_decap_3  PHY_479
timestamp 1586364061
transform -1 0 8832 0 1 132192
box -38 -48 314 592
use scs8hd_decap_6  FILLER_239_74
timestamp 1586364061
transform 1 0 7912 0 1 132192
box -38 -48 590 592
use scs8hd_fill_1  FILLER_239_80
timestamp 1586364061
transform 1 0 8464 0 1 132192
box -38 -48 130 592
use scs8hd_decap_3  PHY_480
timestamp 1586364061
transform 1 0 1104 0 -1 133280
box -38 -48 314 592
use scs8hd_decap_12  FILLER_240_3
timestamp 1586364061
transform 1 0 1380 0 -1 133280
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_240_15
timestamp 1586364061
transform 1 0 2484 0 -1 133280
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1449
timestamp 1586364061
transform 1 0 3956 0 -1 133280
box -38 -48 130 592
use scs8hd_decap_4  FILLER_240_27
timestamp 1586364061
transform 1 0 3588 0 -1 133280
box -38 -48 406 592
use scs8hd_decap_12  FILLER_240_32
timestamp 1586364061
transform 1 0 4048 0 -1 133280
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_240_44
timestamp 1586364061
transform 1 0 5152 0 -1 133280
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_240_56
timestamp 1586364061
transform 1 0 6256 0 -1 133280
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_240_68
timestamp 1586364061
transform 1 0 7360 0 -1 133280
box -38 -48 1142 592
use scs8hd_decap_3  PHY_481
timestamp 1586364061
transform -1 0 8832 0 -1 133280
box -38 -48 314 592
use scs8hd_fill_1  FILLER_240_80
timestamp 1586364061
transform 1 0 8464 0 -1 133280
box -38 -48 130 592
use scs8hd_decap_3  PHY_482
timestamp 1586364061
transform 1 0 1104 0 1 133280
box -38 -48 314 592
use scs8hd_decap_12  FILLER_241_3
timestamp 1586364061
transform 1 0 1380 0 1 133280
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_241_15
timestamp 1586364061
transform 1 0 2484 0 1 133280
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_241_27
timestamp 1586364061
transform 1 0 3588 0 1 133280
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_241_39
timestamp 1586364061
transform 1 0 4692 0 1 133280
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_241_51
timestamp 1586364061
transform 1 0 5796 0 1 133280
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1450
timestamp 1586364061
transform 1 0 6716 0 1 133280
box -38 -48 130 592
use scs8hd_fill_2  FILLER_241_59
timestamp 1586364061
transform 1 0 6532 0 1 133280
box -38 -48 222 592
use scs8hd_decap_12  FILLER_241_62
timestamp 1586364061
transform 1 0 6808 0 1 133280
box -38 -48 1142 592
use scs8hd_decap_3  PHY_483
timestamp 1586364061
transform -1 0 8832 0 1 133280
box -38 -48 314 592
use scs8hd_decap_6  FILLER_241_74
timestamp 1586364061
transform 1 0 7912 0 1 133280
box -38 -48 590 592
use scs8hd_fill_1  FILLER_241_80
timestamp 1586364061
transform 1 0 8464 0 1 133280
box -38 -48 130 592
use scs8hd_decap_3  PHY_484
timestamp 1586364061
transform 1 0 1104 0 -1 134368
box -38 -48 314 592
use scs8hd_decap_12  FILLER_242_3
timestamp 1586364061
transform 1 0 1380 0 -1 134368
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_242_15
timestamp 1586364061
transform 1 0 2484 0 -1 134368
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1451
timestamp 1586364061
transform 1 0 3956 0 -1 134368
box -38 -48 130 592
use scs8hd_decap_4  FILLER_242_27
timestamp 1586364061
transform 1 0 3588 0 -1 134368
box -38 -48 406 592
use scs8hd_decap_12  FILLER_242_32
timestamp 1586364061
transform 1 0 4048 0 -1 134368
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_242_44
timestamp 1586364061
transform 1 0 5152 0 -1 134368
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_242_56
timestamp 1586364061
transform 1 0 6256 0 -1 134368
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_242_68
timestamp 1586364061
transform 1 0 7360 0 -1 134368
box -38 -48 1142 592
use scs8hd_decap_3  PHY_485
timestamp 1586364061
transform -1 0 8832 0 -1 134368
box -38 -48 314 592
use scs8hd_fill_1  FILLER_242_80
timestamp 1586364061
transform 1 0 8464 0 -1 134368
box -38 -48 130 592
use scs8hd_decap_3  PHY_486
timestamp 1586364061
transform 1 0 1104 0 1 134368
box -38 -48 314 592
use scs8hd_decap_12  FILLER_243_3
timestamp 1586364061
transform 1 0 1380 0 1 134368
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_243_15
timestamp 1586364061
transform 1 0 2484 0 1 134368
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_243_27
timestamp 1586364061
transform 1 0 3588 0 1 134368
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_243_39
timestamp 1586364061
transform 1 0 4692 0 1 134368
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_243_51
timestamp 1586364061
transform 1 0 5796 0 1 134368
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1452
timestamp 1586364061
transform 1 0 6716 0 1 134368
box -38 -48 130 592
use scs8hd_fill_2  FILLER_243_59
timestamp 1586364061
transform 1 0 6532 0 1 134368
box -38 -48 222 592
use scs8hd_decap_12  FILLER_243_62
timestamp 1586364061
transform 1 0 6808 0 1 134368
box -38 -48 1142 592
use scs8hd_decap_3  PHY_487
timestamp 1586364061
transform -1 0 8832 0 1 134368
box -38 -48 314 592
use scs8hd_decap_6  FILLER_243_74
timestamp 1586364061
transform 1 0 7912 0 1 134368
box -38 -48 590 592
use scs8hd_fill_1  FILLER_243_80
timestamp 1586364061
transform 1 0 8464 0 1 134368
box -38 -48 130 592
use scs8hd_decap_3  PHY_488
timestamp 1586364061
transform 1 0 1104 0 -1 135456
box -38 -48 314 592
use scs8hd_decap_3  PHY_490
timestamp 1586364061
transform 1 0 1104 0 1 135456
box -38 -48 314 592
use scs8hd_decap_12  FILLER_244_3
timestamp 1586364061
transform 1 0 1380 0 -1 135456
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_244_15
timestamp 1586364061
transform 1 0 2484 0 -1 135456
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_245_3
timestamp 1586364061
transform 1 0 1380 0 1 135456
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_245_15
timestamp 1586364061
transform 1 0 2484 0 1 135456
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1453
timestamp 1586364061
transform 1 0 3956 0 -1 135456
box -38 -48 130 592
use scs8hd_decap_4  FILLER_244_27
timestamp 1586364061
transform 1 0 3588 0 -1 135456
box -38 -48 406 592
use scs8hd_decap_12  FILLER_244_32
timestamp 1586364061
transform 1 0 4048 0 -1 135456
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_245_27
timestamp 1586364061
transform 1 0 3588 0 1 135456
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_244_44
timestamp 1586364061
transform 1 0 5152 0 -1 135456
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_245_39
timestamp 1586364061
transform 1 0 4692 0 1 135456
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_245_51
timestamp 1586364061
transform 1 0 5796 0 1 135456
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1454
timestamp 1586364061
transform 1 0 6716 0 1 135456
box -38 -48 130 592
use scs8hd_decap_12  FILLER_244_56
timestamp 1586364061
transform 1 0 6256 0 -1 135456
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_244_68
timestamp 1586364061
transform 1 0 7360 0 -1 135456
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_245_59
timestamp 1586364061
transform 1 0 6532 0 1 135456
box -38 -48 222 592
use scs8hd_decap_12  FILLER_245_62
timestamp 1586364061
transform 1 0 6808 0 1 135456
box -38 -48 1142 592
use scs8hd_decap_3  PHY_489
timestamp 1586364061
transform -1 0 8832 0 -1 135456
box -38 -48 314 592
use scs8hd_decap_3  PHY_491
timestamp 1586364061
transform -1 0 8832 0 1 135456
box -38 -48 314 592
use scs8hd_fill_1  FILLER_244_80
timestamp 1586364061
transform 1 0 8464 0 -1 135456
box -38 -48 130 592
use scs8hd_decap_6  FILLER_245_74
timestamp 1586364061
transform 1 0 7912 0 1 135456
box -38 -48 590 592
use scs8hd_fill_1  FILLER_245_80
timestamp 1586364061
transform 1 0 8464 0 1 135456
box -38 -48 130 592
use scs8hd_decap_3  PHY_492
timestamp 1586364061
transform 1 0 1104 0 -1 136544
box -38 -48 314 592
use scs8hd_decap_12  FILLER_246_3
timestamp 1586364061
transform 1 0 1380 0 -1 136544
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_246_15
timestamp 1586364061
transform 1 0 2484 0 -1 136544
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1455
timestamp 1586364061
transform 1 0 3956 0 -1 136544
box -38 -48 130 592
use scs8hd_decap_4  FILLER_246_27
timestamp 1586364061
transform 1 0 3588 0 -1 136544
box -38 -48 406 592
use scs8hd_decap_12  FILLER_246_32
timestamp 1586364061
transform 1 0 4048 0 -1 136544
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_246_44
timestamp 1586364061
transform 1 0 5152 0 -1 136544
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_246_56
timestamp 1586364061
transform 1 0 6256 0 -1 136544
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_246_68
timestamp 1586364061
transform 1 0 7360 0 -1 136544
box -38 -48 1142 592
use scs8hd_decap_3  PHY_493
timestamp 1586364061
transform -1 0 8832 0 -1 136544
box -38 -48 314 592
use scs8hd_fill_1  FILLER_246_80
timestamp 1586364061
transform 1 0 8464 0 -1 136544
box -38 -48 130 592
use scs8hd_decap_3  PHY_494
timestamp 1586364061
transform 1 0 1104 0 1 136544
box -38 -48 314 592
use scs8hd_decap_12  FILLER_247_3
timestamp 1586364061
transform 1 0 1380 0 1 136544
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_247_15
timestamp 1586364061
transform 1 0 2484 0 1 136544
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_247_27
timestamp 1586364061
transform 1 0 3588 0 1 136544
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_247_39
timestamp 1586364061
transform 1 0 4692 0 1 136544
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_247_51
timestamp 1586364061
transform 1 0 5796 0 1 136544
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1456
timestamp 1586364061
transform 1 0 6716 0 1 136544
box -38 -48 130 592
use scs8hd_fill_2  FILLER_247_59
timestamp 1586364061
transform 1 0 6532 0 1 136544
box -38 -48 222 592
use scs8hd_decap_12  FILLER_247_62
timestamp 1586364061
transform 1 0 6808 0 1 136544
box -38 -48 1142 592
use scs8hd_decap_3  PHY_495
timestamp 1586364061
transform -1 0 8832 0 1 136544
box -38 -48 314 592
use scs8hd_decap_6  FILLER_247_74
timestamp 1586364061
transform 1 0 7912 0 1 136544
box -38 -48 590 592
use scs8hd_fill_1  FILLER_247_80
timestamp 1586364061
transform 1 0 8464 0 1 136544
box -38 -48 130 592
use scs8hd_decap_3  PHY_496
timestamp 1586364061
transform 1 0 1104 0 -1 137632
box -38 -48 314 592
use scs8hd_decap_12  FILLER_248_3
timestamp 1586364061
transform 1 0 1380 0 -1 137632
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_248_15
timestamp 1586364061
transform 1 0 2484 0 -1 137632
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1457
timestamp 1586364061
transform 1 0 3956 0 -1 137632
box -38 -48 130 592
use scs8hd_decap_4  FILLER_248_27
timestamp 1586364061
transform 1 0 3588 0 -1 137632
box -38 -48 406 592
use scs8hd_decap_12  FILLER_248_32
timestamp 1586364061
transform 1 0 4048 0 -1 137632
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_248_44
timestamp 1586364061
transform 1 0 5152 0 -1 137632
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_248_56
timestamp 1586364061
transform 1 0 6256 0 -1 137632
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_248_68
timestamp 1586364061
transform 1 0 7360 0 -1 137632
box -38 -48 1142 592
use scs8hd_decap_3  PHY_497
timestamp 1586364061
transform -1 0 8832 0 -1 137632
box -38 -48 314 592
use scs8hd_fill_1  FILLER_248_80
timestamp 1586364061
transform 1 0 8464 0 -1 137632
box -38 -48 130 592
use scs8hd_decap_3  PHY_498
timestamp 1586364061
transform 1 0 1104 0 1 137632
box -38 -48 314 592
use scs8hd_decap_12  FILLER_249_3
timestamp 1586364061
transform 1 0 1380 0 1 137632
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_249_15
timestamp 1586364061
transform 1 0 2484 0 1 137632
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_249_27
timestamp 1586364061
transform 1 0 3588 0 1 137632
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_249_39
timestamp 1586364061
transform 1 0 4692 0 1 137632
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_249_51
timestamp 1586364061
transform 1 0 5796 0 1 137632
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1458
timestamp 1586364061
transform 1 0 6716 0 1 137632
box -38 -48 130 592
use scs8hd_fill_2  FILLER_249_59
timestamp 1586364061
transform 1 0 6532 0 1 137632
box -38 -48 222 592
use scs8hd_decap_12  FILLER_249_62
timestamp 1586364061
transform 1 0 6808 0 1 137632
box -38 -48 1142 592
use scs8hd_decap_3  PHY_499
timestamp 1586364061
transform -1 0 8832 0 1 137632
box -38 -48 314 592
use scs8hd_decap_6  FILLER_249_74
timestamp 1586364061
transform 1 0 7912 0 1 137632
box -38 -48 590 592
use scs8hd_fill_1  FILLER_249_80
timestamp 1586364061
transform 1 0 8464 0 1 137632
box -38 -48 130 592
use scs8hd_decap_3  PHY_500
timestamp 1586364061
transform 1 0 1104 0 -1 138720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_250_3
timestamp 1586364061
transform 1 0 1380 0 -1 138720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_250_15
timestamp 1586364061
transform 1 0 2484 0 -1 138720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1459
timestamp 1586364061
transform 1 0 3956 0 -1 138720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_250_27
timestamp 1586364061
transform 1 0 3588 0 -1 138720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_250_32
timestamp 1586364061
transform 1 0 4048 0 -1 138720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_250_44
timestamp 1586364061
transform 1 0 5152 0 -1 138720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_250_56
timestamp 1586364061
transform 1 0 6256 0 -1 138720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_250_68
timestamp 1586364061
transform 1 0 7360 0 -1 138720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_501
timestamp 1586364061
transform -1 0 8832 0 -1 138720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_250_80
timestamp 1586364061
transform 1 0 8464 0 -1 138720
box -38 -48 130 592
use scs8hd_decap_3  PHY_502
timestamp 1586364061
transform 1 0 1104 0 1 138720
box -38 -48 314 592
use scs8hd_decap_3  PHY_504
timestamp 1586364061
transform 1 0 1104 0 -1 139808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_251_3
timestamp 1586364061
transform 1 0 1380 0 1 138720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_251_15
timestamp 1586364061
transform 1 0 2484 0 1 138720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_252_3
timestamp 1586364061
transform 1 0 1380 0 -1 139808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_252_15
timestamp 1586364061
transform 1 0 2484 0 -1 139808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1461
timestamp 1586364061
transform 1 0 3956 0 -1 139808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_251_27
timestamp 1586364061
transform 1 0 3588 0 1 138720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_252_27
timestamp 1586364061
transform 1 0 3588 0 -1 139808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_252_32
timestamp 1586364061
transform 1 0 4048 0 -1 139808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_251_39
timestamp 1586364061
transform 1 0 4692 0 1 138720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_251_51
timestamp 1586364061
transform 1 0 5796 0 1 138720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_252_44
timestamp 1586364061
transform 1 0 5152 0 -1 139808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1460
timestamp 1586364061
transform 1 0 6716 0 1 138720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_251_59
timestamp 1586364061
transform 1 0 6532 0 1 138720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_251_62
timestamp 1586364061
transform 1 0 6808 0 1 138720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_252_56
timestamp 1586364061
transform 1 0 6256 0 -1 139808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_252_68
timestamp 1586364061
transform 1 0 7360 0 -1 139808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_503
timestamp 1586364061
transform -1 0 8832 0 1 138720
box -38 -48 314 592
use scs8hd_decap_3  PHY_505
timestamp 1586364061
transform -1 0 8832 0 -1 139808
box -38 -48 314 592
use scs8hd_decap_6  FILLER_251_74
timestamp 1586364061
transform 1 0 7912 0 1 138720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_251_80
timestamp 1586364061
transform 1 0 8464 0 1 138720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_252_80
timestamp 1586364061
transform 1 0 8464 0 -1 139808
box -38 -48 130 592
use scs8hd_decap_3  PHY_506
timestamp 1586364061
transform 1 0 1104 0 1 139808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_253_3
timestamp 1586364061
transform 1 0 1380 0 1 139808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_253_15
timestamp 1586364061
transform 1 0 2484 0 1 139808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_253_27
timestamp 1586364061
transform 1 0 3588 0 1 139808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_253_39
timestamp 1586364061
transform 1 0 4692 0 1 139808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_253_51
timestamp 1586364061
transform 1 0 5796 0 1 139808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1462
timestamp 1586364061
transform 1 0 6716 0 1 139808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_253_59
timestamp 1586364061
transform 1 0 6532 0 1 139808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_253_62
timestamp 1586364061
transform 1 0 6808 0 1 139808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_507
timestamp 1586364061
transform -1 0 8832 0 1 139808
box -38 -48 314 592
use scs8hd_decap_6  FILLER_253_74
timestamp 1586364061
transform 1 0 7912 0 1 139808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_253_80
timestamp 1586364061
transform 1 0 8464 0 1 139808
box -38 -48 130 592
use scs8hd_decap_3  PHY_508
timestamp 1586364061
transform 1 0 1104 0 -1 140896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_254_3
timestamp 1586364061
transform 1 0 1380 0 -1 140896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_254_15
timestamp 1586364061
transform 1 0 2484 0 -1 140896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1463
timestamp 1586364061
transform 1 0 3956 0 -1 140896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_254_27
timestamp 1586364061
transform 1 0 3588 0 -1 140896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_254_32
timestamp 1586364061
transform 1 0 4048 0 -1 140896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_254_44
timestamp 1586364061
transform 1 0 5152 0 -1 140896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_254_56
timestamp 1586364061
transform 1 0 6256 0 -1 140896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_254_68
timestamp 1586364061
transform 1 0 7360 0 -1 140896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_509
timestamp 1586364061
transform -1 0 8832 0 -1 140896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_254_80
timestamp 1586364061
transform 1 0 8464 0 -1 140896
box -38 -48 130 592
use scs8hd_decap_3  PHY_510
timestamp 1586364061
transform 1 0 1104 0 1 140896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_255_3
timestamp 1586364061
transform 1 0 1380 0 1 140896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_255_15
timestamp 1586364061
transform 1 0 2484 0 1 140896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_255_27
timestamp 1586364061
transform 1 0 3588 0 1 140896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_255_39
timestamp 1586364061
transform 1 0 4692 0 1 140896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_255_51
timestamp 1586364061
transform 1 0 5796 0 1 140896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1464
timestamp 1586364061
transform 1 0 6716 0 1 140896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_255_59
timestamp 1586364061
transform 1 0 6532 0 1 140896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_255_62
timestamp 1586364061
transform 1 0 6808 0 1 140896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_511
timestamp 1586364061
transform -1 0 8832 0 1 140896
box -38 -48 314 592
use scs8hd_decap_6  FILLER_255_74
timestamp 1586364061
transform 1 0 7912 0 1 140896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_255_80
timestamp 1586364061
transform 1 0 8464 0 1 140896
box -38 -48 130 592
use scs8hd_decap_3  PHY_512
timestamp 1586364061
transform 1 0 1104 0 -1 141984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_256_3
timestamp 1586364061
transform 1 0 1380 0 -1 141984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_256_15
timestamp 1586364061
transform 1 0 2484 0 -1 141984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1465
timestamp 1586364061
transform 1 0 3956 0 -1 141984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_256_27
timestamp 1586364061
transform 1 0 3588 0 -1 141984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_256_32
timestamp 1586364061
transform 1 0 4048 0 -1 141984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_256_44
timestamp 1586364061
transform 1 0 5152 0 -1 141984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_256_56
timestamp 1586364061
transform 1 0 6256 0 -1 141984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_256_68
timestamp 1586364061
transform 1 0 7360 0 -1 141984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_513
timestamp 1586364061
transform -1 0 8832 0 -1 141984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_256_80
timestamp 1586364061
transform 1 0 8464 0 -1 141984
box -38 -48 130 592
use scs8hd_decap_3  PHY_514
timestamp 1586364061
transform 1 0 1104 0 1 141984
box -38 -48 314 592
use scs8hd_decap_3  PHY_516
timestamp 1586364061
transform 1 0 1104 0 -1 143072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_257_3
timestamp 1586364061
transform 1 0 1380 0 1 141984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_257_15
timestamp 1586364061
transform 1 0 2484 0 1 141984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_258_3
timestamp 1586364061
transform 1 0 1380 0 -1 143072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_258_15
timestamp 1586364061
transform 1 0 2484 0 -1 143072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1467
timestamp 1586364061
transform 1 0 3956 0 -1 143072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_257_27
timestamp 1586364061
transform 1 0 3588 0 1 141984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_258_27
timestamp 1586364061
transform 1 0 3588 0 -1 143072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_258_32
timestamp 1586364061
transform 1 0 4048 0 -1 143072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_257_39
timestamp 1586364061
transform 1 0 4692 0 1 141984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_257_51
timestamp 1586364061
transform 1 0 5796 0 1 141984
box -38 -48 774 592
use scs8hd_decap_12  FILLER_258_44
timestamp 1586364061
transform 1 0 5152 0 -1 143072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1466
timestamp 1586364061
transform 1 0 6716 0 1 141984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_257_59
timestamp 1586364061
transform 1 0 6532 0 1 141984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_257_62
timestamp 1586364061
transform 1 0 6808 0 1 141984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_258_56
timestamp 1586364061
transform 1 0 6256 0 -1 143072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_258_68
timestamp 1586364061
transform 1 0 7360 0 -1 143072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_515
timestamp 1586364061
transform -1 0 8832 0 1 141984
box -38 -48 314 592
use scs8hd_decap_3  PHY_517
timestamp 1586364061
transform -1 0 8832 0 -1 143072
box -38 -48 314 592
use scs8hd_decap_6  FILLER_257_74
timestamp 1586364061
transform 1 0 7912 0 1 141984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_257_80
timestamp 1586364061
transform 1 0 8464 0 1 141984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_258_80
timestamp 1586364061
transform 1 0 8464 0 -1 143072
box -38 -48 130 592
use scs8hd_decap_3  PHY_518
timestamp 1586364061
transform 1 0 1104 0 1 143072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_259_3
timestamp 1586364061
transform 1 0 1380 0 1 143072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_259_15
timestamp 1586364061
transform 1 0 2484 0 1 143072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_259_27
timestamp 1586364061
transform 1 0 3588 0 1 143072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_259_39
timestamp 1586364061
transform 1 0 4692 0 1 143072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_259_51
timestamp 1586364061
transform 1 0 5796 0 1 143072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1468
timestamp 1586364061
transform 1 0 6716 0 1 143072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_259_59
timestamp 1586364061
transform 1 0 6532 0 1 143072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_259_62
timestamp 1586364061
transform 1 0 6808 0 1 143072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_519
timestamp 1586364061
transform -1 0 8832 0 1 143072
box -38 -48 314 592
use scs8hd_decap_6  FILLER_259_74
timestamp 1586364061
transform 1 0 7912 0 1 143072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_259_80
timestamp 1586364061
transform 1 0 8464 0 1 143072
box -38 -48 130 592
use scs8hd_decap_3  PHY_520
timestamp 1586364061
transform 1 0 1104 0 -1 144160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_260_3
timestamp 1586364061
transform 1 0 1380 0 -1 144160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_260_15
timestamp 1586364061
transform 1 0 2484 0 -1 144160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1469
timestamp 1586364061
transform 1 0 3956 0 -1 144160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_260_27
timestamp 1586364061
transform 1 0 3588 0 -1 144160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_260_32
timestamp 1586364061
transform 1 0 4048 0 -1 144160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_260_44
timestamp 1586364061
transform 1 0 5152 0 -1 144160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_260_56
timestamp 1586364061
transform 1 0 6256 0 -1 144160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_260_68
timestamp 1586364061
transform 1 0 7360 0 -1 144160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_521
timestamp 1586364061
transform -1 0 8832 0 -1 144160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_260_80
timestamp 1586364061
transform 1 0 8464 0 -1 144160
box -38 -48 130 592
use scs8hd_decap_3  PHY_522
timestamp 1586364061
transform 1 0 1104 0 1 144160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_261_3
timestamp 1586364061
transform 1 0 1380 0 1 144160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_261_15
timestamp 1586364061
transform 1 0 2484 0 1 144160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_261_27
timestamp 1586364061
transform 1 0 3588 0 1 144160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_261_39
timestamp 1586364061
transform 1 0 4692 0 1 144160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_261_51
timestamp 1586364061
transform 1 0 5796 0 1 144160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1470
timestamp 1586364061
transform 1 0 6716 0 1 144160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_261_59
timestamp 1586364061
transform 1 0 6532 0 1 144160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_261_62
timestamp 1586364061
transform 1 0 6808 0 1 144160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_523
timestamp 1586364061
transform -1 0 8832 0 1 144160
box -38 -48 314 592
use scs8hd_decap_6  FILLER_261_74
timestamp 1586364061
transform 1 0 7912 0 1 144160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_261_80
timestamp 1586364061
transform 1 0 8464 0 1 144160
box -38 -48 130 592
use scs8hd_decap_3  PHY_524
timestamp 1586364061
transform 1 0 1104 0 -1 145248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_262_3
timestamp 1586364061
transform 1 0 1380 0 -1 145248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_262_15
timestamp 1586364061
transform 1 0 2484 0 -1 145248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1471
timestamp 1586364061
transform 1 0 3956 0 -1 145248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_262_27
timestamp 1586364061
transform 1 0 3588 0 -1 145248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_262_32
timestamp 1586364061
transform 1 0 4048 0 -1 145248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_262_44
timestamp 1586364061
transform 1 0 5152 0 -1 145248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_262_56
timestamp 1586364061
transform 1 0 6256 0 -1 145248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_262_68
timestamp 1586364061
transform 1 0 7360 0 -1 145248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_525
timestamp 1586364061
transform -1 0 8832 0 -1 145248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_262_80
timestamp 1586364061
transform 1 0 8464 0 -1 145248
box -38 -48 130 592
use scs8hd_decap_3  PHY_526
timestamp 1586364061
transform 1 0 1104 0 1 145248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_263_3
timestamp 1586364061
transform 1 0 1380 0 1 145248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_263_15
timestamp 1586364061
transform 1 0 2484 0 1 145248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_263_27
timestamp 1586364061
transform 1 0 3588 0 1 145248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_263_39
timestamp 1586364061
transform 1 0 4692 0 1 145248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_263_51
timestamp 1586364061
transform 1 0 5796 0 1 145248
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1472
timestamp 1586364061
transform 1 0 6716 0 1 145248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_263_59
timestamp 1586364061
transform 1 0 6532 0 1 145248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_263_62
timestamp 1586364061
transform 1 0 6808 0 1 145248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_527
timestamp 1586364061
transform -1 0 8832 0 1 145248
box -38 -48 314 592
use scs8hd_decap_6  FILLER_263_74
timestamp 1586364061
transform 1 0 7912 0 1 145248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_263_80
timestamp 1586364061
transform 1 0 8464 0 1 145248
box -38 -48 130 592
use scs8hd_decap_3  PHY_528
timestamp 1586364061
transform 1 0 1104 0 -1 146336
box -38 -48 314 592
use scs8hd_decap_3  PHY_530
timestamp 1586364061
transform 1 0 1104 0 1 146336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_264_3
timestamp 1586364061
transform 1 0 1380 0 -1 146336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_264_15
timestamp 1586364061
transform 1 0 2484 0 -1 146336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_265_3
timestamp 1586364061
transform 1 0 1380 0 1 146336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_265_15
timestamp 1586364061
transform 1 0 2484 0 1 146336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1473
timestamp 1586364061
transform 1 0 3956 0 -1 146336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_264_27
timestamp 1586364061
transform 1 0 3588 0 -1 146336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_264_32
timestamp 1586364061
transform 1 0 4048 0 -1 146336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_265_27
timestamp 1586364061
transform 1 0 3588 0 1 146336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_264_44
timestamp 1586364061
transform 1 0 5152 0 -1 146336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_265_39
timestamp 1586364061
transform 1 0 4692 0 1 146336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_265_51
timestamp 1586364061
transform 1 0 5796 0 1 146336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1474
timestamp 1586364061
transform 1 0 6716 0 1 146336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_264_56
timestamp 1586364061
transform 1 0 6256 0 -1 146336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_264_68
timestamp 1586364061
transform 1 0 7360 0 -1 146336
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_265_59
timestamp 1586364061
transform 1 0 6532 0 1 146336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_265_62
timestamp 1586364061
transform 1 0 6808 0 1 146336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_529
timestamp 1586364061
transform -1 0 8832 0 -1 146336
box -38 -48 314 592
use scs8hd_decap_3  PHY_531
timestamp 1586364061
transform -1 0 8832 0 1 146336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_264_80
timestamp 1586364061
transform 1 0 8464 0 -1 146336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_265_74
timestamp 1586364061
transform 1 0 7912 0 1 146336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_265_80
timestamp 1586364061
transform 1 0 8464 0 1 146336
box -38 -48 130 592
use scs8hd_decap_3  PHY_532
timestamp 1586364061
transform 1 0 1104 0 -1 147424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_266_3
timestamp 1586364061
transform 1 0 1380 0 -1 147424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_266_15
timestamp 1586364061
transform 1 0 2484 0 -1 147424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1475
timestamp 1586364061
transform 1 0 3956 0 -1 147424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_266_27
timestamp 1586364061
transform 1 0 3588 0 -1 147424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_266_32
timestamp 1586364061
transform 1 0 4048 0 -1 147424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_266_44
timestamp 1586364061
transform 1 0 5152 0 -1 147424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_266_56
timestamp 1586364061
transform 1 0 6256 0 -1 147424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_266_68
timestamp 1586364061
transform 1 0 7360 0 -1 147424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_533
timestamp 1586364061
transform -1 0 8832 0 -1 147424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_266_80
timestamp 1586364061
transform 1 0 8464 0 -1 147424
box -38 -48 130 592
use scs8hd_decap_3  PHY_534
timestamp 1586364061
transform 1 0 1104 0 1 147424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_267_3
timestamp 1586364061
transform 1 0 1380 0 1 147424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_267_15
timestamp 1586364061
transform 1 0 2484 0 1 147424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_267_27
timestamp 1586364061
transform 1 0 3588 0 1 147424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_267_39
timestamp 1586364061
transform 1 0 4692 0 1 147424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_267_51
timestamp 1586364061
transform 1 0 5796 0 1 147424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1476
timestamp 1586364061
transform 1 0 6716 0 1 147424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_267_59
timestamp 1586364061
transform 1 0 6532 0 1 147424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_267_62
timestamp 1586364061
transform 1 0 6808 0 1 147424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_535
timestamp 1586364061
transform -1 0 8832 0 1 147424
box -38 -48 314 592
use scs8hd_decap_6  FILLER_267_74
timestamp 1586364061
transform 1 0 7912 0 1 147424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_267_80
timestamp 1586364061
transform 1 0 8464 0 1 147424
box -38 -48 130 592
use scs8hd_decap_3  PHY_536
timestamp 1586364061
transform 1 0 1104 0 -1 148512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_268_3
timestamp 1586364061
transform 1 0 1380 0 -1 148512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_268_15
timestamp 1586364061
transform 1 0 2484 0 -1 148512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1477
timestamp 1586364061
transform 1 0 3956 0 -1 148512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_268_27
timestamp 1586364061
transform 1 0 3588 0 -1 148512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_268_32
timestamp 1586364061
transform 1 0 4048 0 -1 148512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_268_44
timestamp 1586364061
transform 1 0 5152 0 -1 148512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_268_56
timestamp 1586364061
transform 1 0 6256 0 -1 148512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_268_68
timestamp 1586364061
transform 1 0 7360 0 -1 148512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_537
timestamp 1586364061
transform -1 0 8832 0 -1 148512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_268_80
timestamp 1586364061
transform 1 0 8464 0 -1 148512
box -38 -48 130 592
use scs8hd_decap_3  PHY_538
timestamp 1586364061
transform 1 0 1104 0 1 148512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_269_3
timestamp 1586364061
transform 1 0 1380 0 1 148512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_269_15
timestamp 1586364061
transform 1 0 2484 0 1 148512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_269_27
timestamp 1586364061
transform 1 0 3588 0 1 148512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_269_39
timestamp 1586364061
transform 1 0 4692 0 1 148512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_269_51
timestamp 1586364061
transform 1 0 5796 0 1 148512
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1478
timestamp 1586364061
transform 1 0 6716 0 1 148512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_269_59
timestamp 1586364061
transform 1 0 6532 0 1 148512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_269_62
timestamp 1586364061
transform 1 0 6808 0 1 148512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_539
timestamp 1586364061
transform -1 0 8832 0 1 148512
box -38 -48 314 592
use scs8hd_decap_6  FILLER_269_74
timestamp 1586364061
transform 1 0 7912 0 1 148512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_269_80
timestamp 1586364061
transform 1 0 8464 0 1 148512
box -38 -48 130 592
use scs8hd_decap_3  PHY_540
timestamp 1586364061
transform 1 0 1104 0 -1 149600
box -38 -48 314 592
use scs8hd_decap_3  PHY_542
timestamp 1586364061
transform 1 0 1104 0 1 149600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_270_3
timestamp 1586364061
transform 1 0 1380 0 -1 149600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_270_15
timestamp 1586364061
transform 1 0 2484 0 -1 149600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_271_3
timestamp 1586364061
transform 1 0 1380 0 1 149600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_271_15
timestamp 1586364061
transform 1 0 2484 0 1 149600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1479
timestamp 1586364061
transform 1 0 3956 0 -1 149600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_270_27
timestamp 1586364061
transform 1 0 3588 0 -1 149600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_270_32
timestamp 1586364061
transform 1 0 4048 0 -1 149600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_271_27
timestamp 1586364061
transform 1 0 3588 0 1 149600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_270_44
timestamp 1586364061
transform 1 0 5152 0 -1 149600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_271_39
timestamp 1586364061
transform 1 0 4692 0 1 149600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_271_51
timestamp 1586364061
transform 1 0 5796 0 1 149600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1480
timestamp 1586364061
transform 1 0 6716 0 1 149600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_270_56
timestamp 1586364061
transform 1 0 6256 0 -1 149600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_270_68
timestamp 1586364061
transform 1 0 7360 0 -1 149600
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_271_59
timestamp 1586364061
transform 1 0 6532 0 1 149600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_271_62
timestamp 1586364061
transform 1 0 6808 0 1 149600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_541
timestamp 1586364061
transform -1 0 8832 0 -1 149600
box -38 -48 314 592
use scs8hd_decap_3  PHY_543
timestamp 1586364061
transform -1 0 8832 0 1 149600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_270_80
timestamp 1586364061
transform 1 0 8464 0 -1 149600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_271_74
timestamp 1586364061
transform 1 0 7912 0 1 149600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_271_80
timestamp 1586364061
transform 1 0 8464 0 1 149600
box -38 -48 130 592
use scs8hd_decap_3  PHY_544
timestamp 1586364061
transform 1 0 1104 0 -1 150688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_272_3
timestamp 1586364061
transform 1 0 1380 0 -1 150688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_272_15
timestamp 1586364061
transform 1 0 2484 0 -1 150688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1481
timestamp 1586364061
transform 1 0 3956 0 -1 150688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_272_27
timestamp 1586364061
transform 1 0 3588 0 -1 150688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_272_32
timestamp 1586364061
transform 1 0 4048 0 -1 150688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_272_44
timestamp 1586364061
transform 1 0 5152 0 -1 150688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_272_56
timestamp 1586364061
transform 1 0 6256 0 -1 150688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_272_68
timestamp 1586364061
transform 1 0 7360 0 -1 150688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_545
timestamp 1586364061
transform -1 0 8832 0 -1 150688
box -38 -48 314 592
use scs8hd_fill_1  FILLER_272_80
timestamp 1586364061
transform 1 0 8464 0 -1 150688
box -38 -48 130 592
use scs8hd_decap_3  PHY_546
timestamp 1586364061
transform 1 0 1104 0 1 150688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_273_3
timestamp 1586364061
transform 1 0 1380 0 1 150688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_273_15
timestamp 1586364061
transform 1 0 2484 0 1 150688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_273_27
timestamp 1586364061
transform 1 0 3588 0 1 150688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_273_39
timestamp 1586364061
transform 1 0 4692 0 1 150688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_273_51
timestamp 1586364061
transform 1 0 5796 0 1 150688
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1482
timestamp 1586364061
transform 1 0 6716 0 1 150688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_273_59
timestamp 1586364061
transform 1 0 6532 0 1 150688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_273_62
timestamp 1586364061
transform 1 0 6808 0 1 150688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_547
timestamp 1586364061
transform -1 0 8832 0 1 150688
box -38 -48 314 592
use scs8hd_decap_6  FILLER_273_74
timestamp 1586364061
transform 1 0 7912 0 1 150688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_273_80
timestamp 1586364061
transform 1 0 8464 0 1 150688
box -38 -48 130 592
use scs8hd_decap_3  PHY_548
timestamp 1586364061
transform 1 0 1104 0 -1 151776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_274_3
timestamp 1586364061
transform 1 0 1380 0 -1 151776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_274_15
timestamp 1586364061
transform 1 0 2484 0 -1 151776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1483
timestamp 1586364061
transform 1 0 3956 0 -1 151776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_274_27
timestamp 1586364061
transform 1 0 3588 0 -1 151776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_274_32
timestamp 1586364061
transform 1 0 4048 0 -1 151776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_274_44
timestamp 1586364061
transform 1 0 5152 0 -1 151776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_274_56
timestamp 1586364061
transform 1 0 6256 0 -1 151776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_274_68
timestamp 1586364061
transform 1 0 7360 0 -1 151776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_549
timestamp 1586364061
transform -1 0 8832 0 -1 151776
box -38 -48 314 592
use scs8hd_fill_1  FILLER_274_80
timestamp 1586364061
transform 1 0 8464 0 -1 151776
box -38 -48 130 592
use scs8hd_decap_3  PHY_550
timestamp 1586364061
transform 1 0 1104 0 1 151776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_275_3
timestamp 1586364061
transform 1 0 1380 0 1 151776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_275_15
timestamp 1586364061
transform 1 0 2484 0 1 151776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_275_27
timestamp 1586364061
transform 1 0 3588 0 1 151776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_275_39
timestamp 1586364061
transform 1 0 4692 0 1 151776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_275_51
timestamp 1586364061
transform 1 0 5796 0 1 151776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1484
timestamp 1586364061
transform 1 0 6716 0 1 151776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_275_59
timestamp 1586364061
transform 1 0 6532 0 1 151776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_275_62
timestamp 1586364061
transform 1 0 6808 0 1 151776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_551
timestamp 1586364061
transform -1 0 8832 0 1 151776
box -38 -48 314 592
use scs8hd_decap_6  FILLER_275_74
timestamp 1586364061
transform 1 0 7912 0 1 151776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_275_80
timestamp 1586364061
transform 1 0 8464 0 1 151776
box -38 -48 130 592
use scs8hd_decap_3  PHY_552
timestamp 1586364061
transform 1 0 1104 0 -1 152864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_276_3
timestamp 1586364061
transform 1 0 1380 0 -1 152864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_276_15
timestamp 1586364061
transform 1 0 2484 0 -1 152864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1485
timestamp 1586364061
transform 1 0 3956 0 -1 152864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_276_27
timestamp 1586364061
transform 1 0 3588 0 -1 152864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_276_32
timestamp 1586364061
transform 1 0 4048 0 -1 152864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_276_44
timestamp 1586364061
transform 1 0 5152 0 -1 152864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_276_56
timestamp 1586364061
transform 1 0 6256 0 -1 152864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_276_68
timestamp 1586364061
transform 1 0 7360 0 -1 152864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_553
timestamp 1586364061
transform -1 0 8832 0 -1 152864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_276_80
timestamp 1586364061
transform 1 0 8464 0 -1 152864
box -38 -48 130 592
use scs8hd_decap_3  PHY_554
timestamp 1586364061
transform 1 0 1104 0 1 152864
box -38 -48 314 592
use scs8hd_decap_3  PHY_556
timestamp 1586364061
transform 1 0 1104 0 -1 153952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_277_3
timestamp 1586364061
transform 1 0 1380 0 1 152864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_277_15
timestamp 1586364061
transform 1 0 2484 0 1 152864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_278_3
timestamp 1586364061
transform 1 0 1380 0 -1 153952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_278_15
timestamp 1586364061
transform 1 0 2484 0 -1 153952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1487
timestamp 1586364061
transform 1 0 3956 0 -1 153952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_277_27
timestamp 1586364061
transform 1 0 3588 0 1 152864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_278_27
timestamp 1586364061
transform 1 0 3588 0 -1 153952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_278_32
timestamp 1586364061
transform 1 0 4048 0 -1 153952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_277_39
timestamp 1586364061
transform 1 0 4692 0 1 152864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_277_51
timestamp 1586364061
transform 1 0 5796 0 1 152864
box -38 -48 774 592
use scs8hd_decap_12  FILLER_278_44
timestamp 1586364061
transform 1 0 5152 0 -1 153952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1486
timestamp 1586364061
transform 1 0 6716 0 1 152864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_277_59
timestamp 1586364061
transform 1 0 6532 0 1 152864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_277_62
timestamp 1586364061
transform 1 0 6808 0 1 152864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_278_56
timestamp 1586364061
transform 1 0 6256 0 -1 153952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_278_68
timestamp 1586364061
transform 1 0 7360 0 -1 153952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_555
timestamp 1586364061
transform -1 0 8832 0 1 152864
box -38 -48 314 592
use scs8hd_decap_3  PHY_557
timestamp 1586364061
transform -1 0 8832 0 -1 153952
box -38 -48 314 592
use scs8hd_decap_6  FILLER_277_74
timestamp 1586364061
transform 1 0 7912 0 1 152864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_277_80
timestamp 1586364061
transform 1 0 8464 0 1 152864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_278_80
timestamp 1586364061
transform 1 0 8464 0 -1 153952
box -38 -48 130 592
use scs8hd_decap_3  PHY_558
timestamp 1586364061
transform 1 0 1104 0 1 153952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_279_3
timestamp 1586364061
transform 1 0 1380 0 1 153952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_279_15
timestamp 1586364061
transform 1 0 2484 0 1 153952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_279_27
timestamp 1586364061
transform 1 0 3588 0 1 153952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_279_39
timestamp 1586364061
transform 1 0 4692 0 1 153952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_279_51
timestamp 1586364061
transform 1 0 5796 0 1 153952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1488
timestamp 1586364061
transform 1 0 6716 0 1 153952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_279_59
timestamp 1586364061
transform 1 0 6532 0 1 153952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_279_62
timestamp 1586364061
transform 1 0 6808 0 1 153952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_559
timestamp 1586364061
transform -1 0 8832 0 1 153952
box -38 -48 314 592
use scs8hd_decap_6  FILLER_279_74
timestamp 1586364061
transform 1 0 7912 0 1 153952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_279_80
timestamp 1586364061
transform 1 0 8464 0 1 153952
box -38 -48 130 592
use scs8hd_decap_3  PHY_560
timestamp 1586364061
transform 1 0 1104 0 -1 155040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_280_3
timestamp 1586364061
transform 1 0 1380 0 -1 155040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_280_15
timestamp 1586364061
transform 1 0 2484 0 -1 155040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1489
timestamp 1586364061
transform 1 0 3956 0 -1 155040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_280_27
timestamp 1586364061
transform 1 0 3588 0 -1 155040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_280_32
timestamp 1586364061
transform 1 0 4048 0 -1 155040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_280_44
timestamp 1586364061
transform 1 0 5152 0 -1 155040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_280_56
timestamp 1586364061
transform 1 0 6256 0 -1 155040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_280_68
timestamp 1586364061
transform 1 0 7360 0 -1 155040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_561
timestamp 1586364061
transform -1 0 8832 0 -1 155040
box -38 -48 314 592
use scs8hd_fill_1  FILLER_280_80
timestamp 1586364061
transform 1 0 8464 0 -1 155040
box -38 -48 130 592
use scs8hd_decap_3  PHY_562
timestamp 1586364061
transform 1 0 1104 0 1 155040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_281_3
timestamp 1586364061
transform 1 0 1380 0 1 155040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_281_15
timestamp 1586364061
transform 1 0 2484 0 1 155040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_281_27
timestamp 1586364061
transform 1 0 3588 0 1 155040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_281_39
timestamp 1586364061
transform 1 0 4692 0 1 155040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_281_51
timestamp 1586364061
transform 1 0 5796 0 1 155040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1490
timestamp 1586364061
transform 1 0 6716 0 1 155040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_281_59
timestamp 1586364061
transform 1 0 6532 0 1 155040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_281_62
timestamp 1586364061
transform 1 0 6808 0 1 155040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_563
timestamp 1586364061
transform -1 0 8832 0 1 155040
box -38 -48 314 592
use scs8hd_decap_6  FILLER_281_74
timestamp 1586364061
transform 1 0 7912 0 1 155040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_281_80
timestamp 1586364061
transform 1 0 8464 0 1 155040
box -38 -48 130 592
use scs8hd_decap_3  PHY_564
timestamp 1586364061
transform 1 0 1104 0 -1 156128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_282_3
timestamp 1586364061
transform 1 0 1380 0 -1 156128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_282_15
timestamp 1586364061
transform 1 0 2484 0 -1 156128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1491
timestamp 1586364061
transform 1 0 3956 0 -1 156128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_282_27
timestamp 1586364061
transform 1 0 3588 0 -1 156128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_282_32
timestamp 1586364061
transform 1 0 4048 0 -1 156128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_282_44
timestamp 1586364061
transform 1 0 5152 0 -1 156128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_282_56
timestamp 1586364061
transform 1 0 6256 0 -1 156128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_282_68
timestamp 1586364061
transform 1 0 7360 0 -1 156128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_565
timestamp 1586364061
transform -1 0 8832 0 -1 156128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_282_80
timestamp 1586364061
transform 1 0 8464 0 -1 156128
box -38 -48 130 592
use scs8hd_decap_3  PHY_566
timestamp 1586364061
transform 1 0 1104 0 1 156128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_283_3
timestamp 1586364061
transform 1 0 1380 0 1 156128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_283_15
timestamp 1586364061
transform 1 0 2484 0 1 156128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_283_27
timestamp 1586364061
transform 1 0 3588 0 1 156128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_283_39
timestamp 1586364061
transform 1 0 4692 0 1 156128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_283_51
timestamp 1586364061
transform 1 0 5796 0 1 156128
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1492
timestamp 1586364061
transform 1 0 6716 0 1 156128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_283_59
timestamp 1586364061
transform 1 0 6532 0 1 156128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_283_62
timestamp 1586364061
transform 1 0 6808 0 1 156128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_567
timestamp 1586364061
transform -1 0 8832 0 1 156128
box -38 -48 314 592
use scs8hd_decap_6  FILLER_283_74
timestamp 1586364061
transform 1 0 7912 0 1 156128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_283_80
timestamp 1586364061
transform 1 0 8464 0 1 156128
box -38 -48 130 592
use scs8hd_decap_3  PHY_568
timestamp 1586364061
transform 1 0 1104 0 -1 157216
box -38 -48 314 592
use scs8hd_decap_3  PHY_570
timestamp 1586364061
transform 1 0 1104 0 1 157216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_284_3
timestamp 1586364061
transform 1 0 1380 0 -1 157216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_284_15
timestamp 1586364061
transform 1 0 2484 0 -1 157216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_285_3
timestamp 1586364061
transform 1 0 1380 0 1 157216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_285_15
timestamp 1586364061
transform 1 0 2484 0 1 157216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1493
timestamp 1586364061
transform 1 0 3956 0 -1 157216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__23__A
timestamp 1586364061
transform 1 0 4048 0 1 157216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_284_27
timestamp 1586364061
transform 1 0 3588 0 -1 157216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_284_32
timestamp 1586364061
transform 1 0 4048 0 -1 157216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_285_27
timestamp 1586364061
transform 1 0 3588 0 1 157216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_285_31
timestamp 1586364061
transform 1 0 3956 0 1 157216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_285_34
timestamp 1586364061
transform 1 0 4232 0 1 157216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_284_44
timestamp 1586364061
transform 1 0 5152 0 -1 157216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_285_46
timestamp 1586364061
transform 1 0 5336 0 1 157216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1494
timestamp 1586364061
transform 1 0 6716 0 1 157216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_284_56
timestamp 1586364061
transform 1 0 6256 0 -1 157216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_284_68
timestamp 1586364061
transform 1 0 7360 0 -1 157216
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_285_58
timestamp 1586364061
transform 1 0 6440 0 1 157216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_285_62
timestamp 1586364061
transform 1 0 6808 0 1 157216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_569
timestamp 1586364061
transform -1 0 8832 0 -1 157216
box -38 -48 314 592
use scs8hd_decap_3  PHY_571
timestamp 1586364061
transform -1 0 8832 0 1 157216
box -38 -48 314 592
use scs8hd_fill_1  FILLER_284_80
timestamp 1586364061
transform 1 0 8464 0 -1 157216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_285_74
timestamp 1586364061
transform 1 0 7912 0 1 157216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_285_80
timestamp 1586364061
transform 1 0 8464 0 1 157216
box -38 -48 130 592
use scs8hd_decap_3  PHY_572
timestamp 1586364061
transform 1 0 1104 0 -1 158304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_286_3
timestamp 1586364061
transform 1 0 1380 0 -1 158304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_286_15
timestamp 1586364061
transform 1 0 2484 0 -1 158304
box -38 -48 1142 592
use scs8hd_buf_2  _23_
timestamp 1586364061
transform 1 0 4048 0 -1 158304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_1495
timestamp 1586364061
transform 1 0 3956 0 -1 158304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_286_27
timestamp 1586364061
transform 1 0 3588 0 -1 158304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_286_36
timestamp 1586364061
transform 1 0 4416 0 -1 158304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_286_48
timestamp 1586364061
transform 1 0 5520 0 -1 158304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_286_60
timestamp 1586364061
transform 1 0 6624 0 -1 158304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_573
timestamp 1586364061
transform -1 0 8832 0 -1 158304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_286_72
timestamp 1586364061
transform 1 0 7728 0 -1 158304
box -38 -48 774 592
use scs8hd_fill_1  FILLER_286_80
timestamp 1586364061
transform 1 0 8464 0 -1 158304
box -38 -48 130 592
use scs8hd_decap_3  PHY_574
timestamp 1586364061
transform 1 0 1104 0 1 158304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_287_3
timestamp 1586364061
transform 1 0 1380 0 1 158304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_287_15
timestamp 1586364061
transform 1 0 2484 0 1 158304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_287_27
timestamp 1586364061
transform 1 0 3588 0 1 158304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_287_39
timestamp 1586364061
transform 1 0 4692 0 1 158304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_287_51
timestamp 1586364061
transform 1 0 5796 0 1 158304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1496
timestamp 1586364061
transform 1 0 6716 0 1 158304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_287_59
timestamp 1586364061
transform 1 0 6532 0 1 158304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_287_62
timestamp 1586364061
transform 1 0 6808 0 1 158304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_575
timestamp 1586364061
transform -1 0 8832 0 1 158304
box -38 -48 314 592
use scs8hd_decap_6  FILLER_287_74
timestamp 1586364061
transform 1 0 7912 0 1 158304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_287_80
timestamp 1586364061
transform 1 0 8464 0 1 158304
box -38 -48 130 592
use scs8hd_decap_3  PHY_576
timestamp 1586364061
transform 1 0 1104 0 -1 159392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_288_3
timestamp 1586364061
transform 1 0 1380 0 -1 159392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_288_15
timestamp 1586364061
transform 1 0 2484 0 -1 159392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1497
timestamp 1586364061
transform 1 0 3956 0 -1 159392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_288_27
timestamp 1586364061
transform 1 0 3588 0 -1 159392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_288_32
timestamp 1586364061
transform 1 0 4048 0 -1 159392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_288_44
timestamp 1586364061
transform 1 0 5152 0 -1 159392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_288_56
timestamp 1586364061
transform 1 0 6256 0 -1 159392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_288_68
timestamp 1586364061
transform 1 0 7360 0 -1 159392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_577
timestamp 1586364061
transform -1 0 8832 0 -1 159392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_288_80
timestamp 1586364061
transform 1 0 8464 0 -1 159392
box -38 -48 130 592
use scs8hd_decap_3  PHY_578
timestamp 1586364061
transform 1 0 1104 0 1 159392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_289_3
timestamp 1586364061
transform 1 0 1380 0 1 159392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_289_15
timestamp 1586364061
transform 1 0 2484 0 1 159392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_289_27
timestamp 1586364061
transform 1 0 3588 0 1 159392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_289_39
timestamp 1586364061
transform 1 0 4692 0 1 159392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_289_51
timestamp 1586364061
transform 1 0 5796 0 1 159392
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1498
timestamp 1586364061
transform 1 0 6716 0 1 159392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_289_59
timestamp 1586364061
transform 1 0 6532 0 1 159392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_289_62
timestamp 1586364061
transform 1 0 6808 0 1 159392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_579
timestamp 1586364061
transform -1 0 8832 0 1 159392
box -38 -48 314 592
use scs8hd_decap_6  FILLER_289_74
timestamp 1586364061
transform 1 0 7912 0 1 159392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_289_80
timestamp 1586364061
transform 1 0 8464 0 1 159392
box -38 -48 130 592
use scs8hd_decap_3  PHY_580
timestamp 1586364061
transform 1 0 1104 0 -1 160480
box -38 -48 314 592
use scs8hd_decap_3  PHY_582
timestamp 1586364061
transform 1 0 1104 0 1 160480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_290_3
timestamp 1586364061
transform 1 0 1380 0 -1 160480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_290_15
timestamp 1586364061
transform 1 0 2484 0 -1 160480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_291_3
timestamp 1586364061
transform 1 0 1380 0 1 160480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_291_15
timestamp 1586364061
transform 1 0 2484 0 1 160480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1499
timestamp 1586364061
transform 1 0 3956 0 -1 160480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_290_27
timestamp 1586364061
transform 1 0 3588 0 -1 160480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_290_32
timestamp 1586364061
transform 1 0 4048 0 -1 160480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_291_27
timestamp 1586364061
transform 1 0 3588 0 1 160480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_290_44
timestamp 1586364061
transform 1 0 5152 0 -1 160480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_291_39
timestamp 1586364061
transform 1 0 4692 0 1 160480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_291_51
timestamp 1586364061
transform 1 0 5796 0 1 160480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1500
timestamp 1586364061
transform 1 0 6716 0 1 160480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_290_56
timestamp 1586364061
transform 1 0 6256 0 -1 160480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_290_68
timestamp 1586364061
transform 1 0 7360 0 -1 160480
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_291_59
timestamp 1586364061
transform 1 0 6532 0 1 160480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_291_62
timestamp 1586364061
transform 1 0 6808 0 1 160480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_581
timestamp 1586364061
transform -1 0 8832 0 -1 160480
box -38 -48 314 592
use scs8hd_decap_3  PHY_583
timestamp 1586364061
transform -1 0 8832 0 1 160480
box -38 -48 314 592
use scs8hd_fill_1  FILLER_290_80
timestamp 1586364061
transform 1 0 8464 0 -1 160480
box -38 -48 130 592
use scs8hd_decap_6  FILLER_291_74
timestamp 1586364061
transform 1 0 7912 0 1 160480
box -38 -48 590 592
use scs8hd_fill_1  FILLER_291_80
timestamp 1586364061
transform 1 0 8464 0 1 160480
box -38 -48 130 592
use scs8hd_decap_3  PHY_584
timestamp 1586364061
transform 1 0 1104 0 -1 161568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_292_3
timestamp 1586364061
transform 1 0 1380 0 -1 161568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_292_15
timestamp 1586364061
transform 1 0 2484 0 -1 161568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1501
timestamp 1586364061
transform 1 0 3956 0 -1 161568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_292_27
timestamp 1586364061
transform 1 0 3588 0 -1 161568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_292_32
timestamp 1586364061
transform 1 0 4048 0 -1 161568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_292_44
timestamp 1586364061
transform 1 0 5152 0 -1 161568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_292_56
timestamp 1586364061
transform 1 0 6256 0 -1 161568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_292_68
timestamp 1586364061
transform 1 0 7360 0 -1 161568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_585
timestamp 1586364061
transform -1 0 8832 0 -1 161568
box -38 -48 314 592
use scs8hd_fill_1  FILLER_292_80
timestamp 1586364061
transform 1 0 8464 0 -1 161568
box -38 -48 130 592
use scs8hd_decap_3  PHY_586
timestamp 1586364061
transform 1 0 1104 0 1 161568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_293_3
timestamp 1586364061
transform 1 0 1380 0 1 161568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_293_15
timestamp 1586364061
transform 1 0 2484 0 1 161568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_293_27
timestamp 1586364061
transform 1 0 3588 0 1 161568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_293_39
timestamp 1586364061
transform 1 0 4692 0 1 161568
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_293_51
timestamp 1586364061
transform 1 0 5796 0 1 161568
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1502
timestamp 1586364061
transform 1 0 6716 0 1 161568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_293_59
timestamp 1586364061
transform 1 0 6532 0 1 161568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_293_62
timestamp 1586364061
transform 1 0 6808 0 1 161568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_587
timestamp 1586364061
transform -1 0 8832 0 1 161568
box -38 -48 314 592
use scs8hd_decap_6  FILLER_293_74
timestamp 1586364061
transform 1 0 7912 0 1 161568
box -38 -48 590 592
use scs8hd_fill_1  FILLER_293_80
timestamp 1586364061
transform 1 0 8464 0 1 161568
box -38 -48 130 592
use scs8hd_decap_3  PHY_588
timestamp 1586364061
transform 1 0 1104 0 -1 162656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_294_3
timestamp 1586364061
transform 1 0 1380 0 -1 162656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_294_15
timestamp 1586364061
transform 1 0 2484 0 -1 162656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1503
timestamp 1586364061
transform 1 0 3956 0 -1 162656
box -38 -48 130 592
use scs8hd_decap_4  FILLER_294_27
timestamp 1586364061
transform 1 0 3588 0 -1 162656
box -38 -48 406 592
use scs8hd_decap_12  FILLER_294_32
timestamp 1586364061
transform 1 0 4048 0 -1 162656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_294_44
timestamp 1586364061
transform 1 0 5152 0 -1 162656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_294_56
timestamp 1586364061
transform 1 0 6256 0 -1 162656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_294_68
timestamp 1586364061
transform 1 0 7360 0 -1 162656
box -38 -48 1142 592
use scs8hd_decap_3  PHY_589
timestamp 1586364061
transform -1 0 8832 0 -1 162656
box -38 -48 314 592
use scs8hd_fill_1  FILLER_294_80
timestamp 1586364061
transform 1 0 8464 0 -1 162656
box -38 -48 130 592
use scs8hd_decap_3  PHY_590
timestamp 1586364061
transform 1 0 1104 0 1 162656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_295_3
timestamp 1586364061
transform 1 0 1380 0 1 162656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_295_15
timestamp 1586364061
transform 1 0 2484 0 1 162656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_295_27
timestamp 1586364061
transform 1 0 3588 0 1 162656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_295_39
timestamp 1586364061
transform 1 0 4692 0 1 162656
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_295_51
timestamp 1586364061
transform 1 0 5796 0 1 162656
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1504
timestamp 1586364061
transform 1 0 6716 0 1 162656
box -38 -48 130 592
use scs8hd_fill_2  FILLER_295_59
timestamp 1586364061
transform 1 0 6532 0 1 162656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_295_62
timestamp 1586364061
transform 1 0 6808 0 1 162656
box -38 -48 1142 592
use scs8hd_decap_3  PHY_591
timestamp 1586364061
transform -1 0 8832 0 1 162656
box -38 -48 314 592
use scs8hd_decap_6  FILLER_295_74
timestamp 1586364061
transform 1 0 7912 0 1 162656
box -38 -48 590 592
use scs8hd_fill_1  FILLER_295_80
timestamp 1586364061
transform 1 0 8464 0 1 162656
box -38 -48 130 592
use scs8hd_decap_3  PHY_592
timestamp 1586364061
transform 1 0 1104 0 -1 163744
box -38 -48 314 592
use scs8hd_decap_12  FILLER_296_3
timestamp 1586364061
transform 1 0 1380 0 -1 163744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_296_15
timestamp 1586364061
transform 1 0 2484 0 -1 163744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1505
timestamp 1586364061
transform 1 0 3956 0 -1 163744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_296_27
timestamp 1586364061
transform 1 0 3588 0 -1 163744
box -38 -48 406 592
use scs8hd_decap_12  FILLER_296_32
timestamp 1586364061
transform 1 0 4048 0 -1 163744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_296_44
timestamp 1586364061
transform 1 0 5152 0 -1 163744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_296_56
timestamp 1586364061
transform 1 0 6256 0 -1 163744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_296_68
timestamp 1586364061
transform 1 0 7360 0 -1 163744
box -38 -48 1142 592
use scs8hd_decap_3  PHY_593
timestamp 1586364061
transform -1 0 8832 0 -1 163744
box -38 -48 314 592
use scs8hd_fill_1  FILLER_296_80
timestamp 1586364061
transform 1 0 8464 0 -1 163744
box -38 -48 130 592
use scs8hd_decap_3  PHY_594
timestamp 1586364061
transform 1 0 1104 0 1 163744
box -38 -48 314 592
use scs8hd_decap_3  PHY_596
timestamp 1586364061
transform 1 0 1104 0 -1 164832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_297_3
timestamp 1586364061
transform 1 0 1380 0 1 163744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_297_15
timestamp 1586364061
transform 1 0 2484 0 1 163744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_298_3
timestamp 1586364061
transform 1 0 1380 0 -1 164832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_298_15
timestamp 1586364061
transform 1 0 2484 0 -1 164832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1507
timestamp 1586364061
transform 1 0 3956 0 -1 164832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_297_27
timestamp 1586364061
transform 1 0 3588 0 1 163744
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_298_27
timestamp 1586364061
transform 1 0 3588 0 -1 164832
box -38 -48 406 592
use scs8hd_decap_12  FILLER_298_32
timestamp 1586364061
transform 1 0 4048 0 -1 164832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_297_39
timestamp 1586364061
transform 1 0 4692 0 1 163744
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_297_51
timestamp 1586364061
transform 1 0 5796 0 1 163744
box -38 -48 774 592
use scs8hd_decap_12  FILLER_298_44
timestamp 1586364061
transform 1 0 5152 0 -1 164832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1506
timestamp 1586364061
transform 1 0 6716 0 1 163744
box -38 -48 130 592
use scs8hd_fill_2  FILLER_297_59
timestamp 1586364061
transform 1 0 6532 0 1 163744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_297_62
timestamp 1586364061
transform 1 0 6808 0 1 163744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_298_56
timestamp 1586364061
transform 1 0 6256 0 -1 164832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_298_68
timestamp 1586364061
transform 1 0 7360 0 -1 164832
box -38 -48 1142 592
use scs8hd_decap_3  PHY_595
timestamp 1586364061
transform -1 0 8832 0 1 163744
box -38 -48 314 592
use scs8hd_decap_3  PHY_597
timestamp 1586364061
transform -1 0 8832 0 -1 164832
box -38 -48 314 592
use scs8hd_decap_6  FILLER_297_74
timestamp 1586364061
transform 1 0 7912 0 1 163744
box -38 -48 590 592
use scs8hd_fill_1  FILLER_297_80
timestamp 1586364061
transform 1 0 8464 0 1 163744
box -38 -48 130 592
use scs8hd_fill_1  FILLER_298_80
timestamp 1586364061
transform 1 0 8464 0 -1 164832
box -38 -48 130 592
use scs8hd_decap_3  PHY_598
timestamp 1586364061
transform 1 0 1104 0 1 164832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_299_3
timestamp 1586364061
transform 1 0 1380 0 1 164832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_299_15
timestamp 1586364061
transform 1 0 2484 0 1 164832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_299_27
timestamp 1586364061
transform 1 0 3588 0 1 164832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_299_39
timestamp 1586364061
transform 1 0 4692 0 1 164832
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_299_51
timestamp 1586364061
transform 1 0 5796 0 1 164832
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1508
timestamp 1586364061
transform 1 0 6716 0 1 164832
box -38 -48 130 592
use scs8hd_fill_2  FILLER_299_59
timestamp 1586364061
transform 1 0 6532 0 1 164832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_299_62
timestamp 1586364061
transform 1 0 6808 0 1 164832
box -38 -48 1142 592
use scs8hd_decap_3  PHY_599
timestamp 1586364061
transform -1 0 8832 0 1 164832
box -38 -48 314 592
use scs8hd_decap_6  FILLER_299_74
timestamp 1586364061
transform 1 0 7912 0 1 164832
box -38 -48 590 592
use scs8hd_fill_1  FILLER_299_80
timestamp 1586364061
transform 1 0 8464 0 1 164832
box -38 -48 130 592
use scs8hd_decap_3  PHY_600
timestamp 1586364061
transform 1 0 1104 0 -1 165920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_300_3
timestamp 1586364061
transform 1 0 1380 0 -1 165920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_300_15
timestamp 1586364061
transform 1 0 2484 0 -1 165920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1509
timestamp 1586364061
transform 1 0 3956 0 -1 165920
box -38 -48 130 592
use scs8hd_decap_4  FILLER_300_27
timestamp 1586364061
transform 1 0 3588 0 -1 165920
box -38 -48 406 592
use scs8hd_decap_12  FILLER_300_32
timestamp 1586364061
transform 1 0 4048 0 -1 165920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_300_44
timestamp 1586364061
transform 1 0 5152 0 -1 165920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_300_56
timestamp 1586364061
transform 1 0 6256 0 -1 165920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_300_68
timestamp 1586364061
transform 1 0 7360 0 -1 165920
box -38 -48 1142 592
use scs8hd_decap_3  PHY_601
timestamp 1586364061
transform -1 0 8832 0 -1 165920
box -38 -48 314 592
use scs8hd_fill_1  FILLER_300_80
timestamp 1586364061
transform 1 0 8464 0 -1 165920
box -38 -48 130 592
use scs8hd_decap_3  PHY_602
timestamp 1586364061
transform 1 0 1104 0 1 165920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_301_3
timestamp 1586364061
transform 1 0 1380 0 1 165920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_301_15
timestamp 1586364061
transform 1 0 2484 0 1 165920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_301_27
timestamp 1586364061
transform 1 0 3588 0 1 165920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_301_39
timestamp 1586364061
transform 1 0 4692 0 1 165920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_301_51
timestamp 1586364061
transform 1 0 5796 0 1 165920
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1510
timestamp 1586364061
transform 1 0 6716 0 1 165920
box -38 -48 130 592
use scs8hd_fill_2  FILLER_301_59
timestamp 1586364061
transform 1 0 6532 0 1 165920
box -38 -48 222 592
use scs8hd_decap_12  FILLER_301_62
timestamp 1586364061
transform 1 0 6808 0 1 165920
box -38 -48 1142 592
use scs8hd_decap_3  PHY_603
timestamp 1586364061
transform -1 0 8832 0 1 165920
box -38 -48 314 592
use scs8hd_decap_6  FILLER_301_74
timestamp 1586364061
transform 1 0 7912 0 1 165920
box -38 -48 590 592
use scs8hd_fill_1  FILLER_301_80
timestamp 1586364061
transform 1 0 8464 0 1 165920
box -38 -48 130 592
use scs8hd_decap_3  PHY_604
timestamp 1586364061
transform 1 0 1104 0 -1 167008
box -38 -48 314 592
use scs8hd_decap_12  FILLER_302_3
timestamp 1586364061
transform 1 0 1380 0 -1 167008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_302_15
timestamp 1586364061
transform 1 0 2484 0 -1 167008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1511
timestamp 1586364061
transform 1 0 3956 0 -1 167008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_302_27
timestamp 1586364061
transform 1 0 3588 0 -1 167008
box -38 -48 406 592
use scs8hd_decap_12  FILLER_302_32
timestamp 1586364061
transform 1 0 4048 0 -1 167008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_302_44
timestamp 1586364061
transform 1 0 5152 0 -1 167008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_302_56
timestamp 1586364061
transform 1 0 6256 0 -1 167008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_302_68
timestamp 1586364061
transform 1 0 7360 0 -1 167008
box -38 -48 1142 592
use scs8hd_decap_3  PHY_605
timestamp 1586364061
transform -1 0 8832 0 -1 167008
box -38 -48 314 592
use scs8hd_fill_1  FILLER_302_80
timestamp 1586364061
transform 1 0 8464 0 -1 167008
box -38 -48 130 592
use scs8hd_decap_3  PHY_606
timestamp 1586364061
transform 1 0 1104 0 1 167008
box -38 -48 314 592
use scs8hd_decap_3  PHY_608
timestamp 1586364061
transform 1 0 1104 0 -1 168096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_303_3
timestamp 1586364061
transform 1 0 1380 0 1 167008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_303_15
timestamp 1586364061
transform 1 0 2484 0 1 167008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_304_3
timestamp 1586364061
transform 1 0 1380 0 -1 168096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_304_15
timestamp 1586364061
transform 1 0 2484 0 -1 168096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1513
timestamp 1586364061
transform 1 0 3956 0 -1 168096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_303_27
timestamp 1586364061
transform 1 0 3588 0 1 167008
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_304_27
timestamp 1586364061
transform 1 0 3588 0 -1 168096
box -38 -48 406 592
use scs8hd_decap_12  FILLER_304_32
timestamp 1586364061
transform 1 0 4048 0 -1 168096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_303_39
timestamp 1586364061
transform 1 0 4692 0 1 167008
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_303_51
timestamp 1586364061
transform 1 0 5796 0 1 167008
box -38 -48 774 592
use scs8hd_decap_12  FILLER_304_44
timestamp 1586364061
transform 1 0 5152 0 -1 168096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1512
timestamp 1586364061
transform 1 0 6716 0 1 167008
box -38 -48 130 592
use scs8hd_fill_2  FILLER_303_59
timestamp 1586364061
transform 1 0 6532 0 1 167008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_303_62
timestamp 1586364061
transform 1 0 6808 0 1 167008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_304_56
timestamp 1586364061
transform 1 0 6256 0 -1 168096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_304_68
timestamp 1586364061
transform 1 0 7360 0 -1 168096
box -38 -48 1142 592
use scs8hd_decap_3  PHY_607
timestamp 1586364061
transform -1 0 8832 0 1 167008
box -38 -48 314 592
use scs8hd_decap_3  PHY_609
timestamp 1586364061
transform -1 0 8832 0 -1 168096
box -38 -48 314 592
use scs8hd_decap_6  FILLER_303_74
timestamp 1586364061
transform 1 0 7912 0 1 167008
box -38 -48 590 592
use scs8hd_fill_1  FILLER_303_80
timestamp 1586364061
transform 1 0 8464 0 1 167008
box -38 -48 130 592
use scs8hd_fill_1  FILLER_304_80
timestamp 1586364061
transform 1 0 8464 0 -1 168096
box -38 -48 130 592
use scs8hd_decap_3  PHY_610
timestamp 1586364061
transform 1 0 1104 0 1 168096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_305_3
timestamp 1586364061
transform 1 0 1380 0 1 168096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_305_15
timestamp 1586364061
transform 1 0 2484 0 1 168096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_305_27
timestamp 1586364061
transform 1 0 3588 0 1 168096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_305_39
timestamp 1586364061
transform 1 0 4692 0 1 168096
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_305_51
timestamp 1586364061
transform 1 0 5796 0 1 168096
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1514
timestamp 1586364061
transform 1 0 6716 0 1 168096
box -38 -48 130 592
use scs8hd_fill_2  FILLER_305_59
timestamp 1586364061
transform 1 0 6532 0 1 168096
box -38 -48 222 592
use scs8hd_decap_12  FILLER_305_62
timestamp 1586364061
transform 1 0 6808 0 1 168096
box -38 -48 1142 592
use scs8hd_decap_3  PHY_611
timestamp 1586364061
transform -1 0 8832 0 1 168096
box -38 -48 314 592
use scs8hd_decap_6  FILLER_305_74
timestamp 1586364061
transform 1 0 7912 0 1 168096
box -38 -48 590 592
use scs8hd_fill_1  FILLER_305_80
timestamp 1586364061
transform 1 0 8464 0 1 168096
box -38 -48 130 592
use scs8hd_decap_3  PHY_612
timestamp 1586364061
transform 1 0 1104 0 -1 169184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_306_3
timestamp 1586364061
transform 1 0 1380 0 -1 169184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_306_15
timestamp 1586364061
transform 1 0 2484 0 -1 169184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1515
timestamp 1586364061
transform 1 0 3956 0 -1 169184
box -38 -48 130 592
use scs8hd_decap_4  FILLER_306_27
timestamp 1586364061
transform 1 0 3588 0 -1 169184
box -38 -48 406 592
use scs8hd_decap_12  FILLER_306_32
timestamp 1586364061
transform 1 0 4048 0 -1 169184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_306_44
timestamp 1586364061
transform 1 0 5152 0 -1 169184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_306_56
timestamp 1586364061
transform 1 0 6256 0 -1 169184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_306_68
timestamp 1586364061
transform 1 0 7360 0 -1 169184
box -38 -48 1142 592
use scs8hd_decap_3  PHY_613
timestamp 1586364061
transform -1 0 8832 0 -1 169184
box -38 -48 314 592
use scs8hd_fill_1  FILLER_306_80
timestamp 1586364061
transform 1 0 8464 0 -1 169184
box -38 -48 130 592
use scs8hd_decap_3  PHY_614
timestamp 1586364061
transform 1 0 1104 0 1 169184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_307_3
timestamp 1586364061
transform 1 0 1380 0 1 169184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_307_15
timestamp 1586364061
transform 1 0 2484 0 1 169184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_307_27
timestamp 1586364061
transform 1 0 3588 0 1 169184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_307_39
timestamp 1586364061
transform 1 0 4692 0 1 169184
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_307_51
timestamp 1586364061
transform 1 0 5796 0 1 169184
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1516
timestamp 1586364061
transform 1 0 6716 0 1 169184
box -38 -48 130 592
use scs8hd_fill_2  FILLER_307_59
timestamp 1586364061
transform 1 0 6532 0 1 169184
box -38 -48 222 592
use scs8hd_decap_12  FILLER_307_62
timestamp 1586364061
transform 1 0 6808 0 1 169184
box -38 -48 1142 592
use scs8hd_decap_3  PHY_615
timestamp 1586364061
transform -1 0 8832 0 1 169184
box -38 -48 314 592
use scs8hd_decap_6  FILLER_307_74
timestamp 1586364061
transform 1 0 7912 0 1 169184
box -38 -48 590 592
use scs8hd_fill_1  FILLER_307_80
timestamp 1586364061
transform 1 0 8464 0 1 169184
box -38 -48 130 592
use scs8hd_decap_3  PHY_616
timestamp 1586364061
transform 1 0 1104 0 -1 170272
box -38 -48 314 592
use scs8hd_decap_12  FILLER_308_3
timestamp 1586364061
transform 1 0 1380 0 -1 170272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_308_15
timestamp 1586364061
transform 1 0 2484 0 -1 170272
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1517
timestamp 1586364061
transform 1 0 3956 0 -1 170272
box -38 -48 130 592
use scs8hd_decap_4  FILLER_308_27
timestamp 1586364061
transform 1 0 3588 0 -1 170272
box -38 -48 406 592
use scs8hd_decap_12  FILLER_308_32
timestamp 1586364061
transform 1 0 4048 0 -1 170272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_308_44
timestamp 1586364061
transform 1 0 5152 0 -1 170272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_308_56
timestamp 1586364061
transform 1 0 6256 0 -1 170272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_308_68
timestamp 1586364061
transform 1 0 7360 0 -1 170272
box -38 -48 1142 592
use scs8hd_decap_3  PHY_617
timestamp 1586364061
transform -1 0 8832 0 -1 170272
box -38 -48 314 592
use scs8hd_fill_1  FILLER_308_80
timestamp 1586364061
transform 1 0 8464 0 -1 170272
box -38 -48 130 592
use scs8hd_decap_3  PHY_618
timestamp 1586364061
transform 1 0 1104 0 1 170272
box -38 -48 314 592
use scs8hd_decap_12  FILLER_309_3
timestamp 1586364061
transform 1 0 1380 0 1 170272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_309_15
timestamp 1586364061
transform 1 0 2484 0 1 170272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_309_27
timestamp 1586364061
transform 1 0 3588 0 1 170272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_309_39
timestamp 1586364061
transform 1 0 4692 0 1 170272
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_309_51
timestamp 1586364061
transform 1 0 5796 0 1 170272
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1518
timestamp 1586364061
transform 1 0 6716 0 1 170272
box -38 -48 130 592
use scs8hd_fill_2  FILLER_309_59
timestamp 1586364061
transform 1 0 6532 0 1 170272
box -38 -48 222 592
use scs8hd_decap_12  FILLER_309_62
timestamp 1586364061
transform 1 0 6808 0 1 170272
box -38 -48 1142 592
use scs8hd_decap_3  PHY_619
timestamp 1586364061
transform -1 0 8832 0 1 170272
box -38 -48 314 592
use scs8hd_decap_6  FILLER_309_74
timestamp 1586364061
transform 1 0 7912 0 1 170272
box -38 -48 590 592
use scs8hd_fill_1  FILLER_309_80
timestamp 1586364061
transform 1 0 8464 0 1 170272
box -38 -48 130 592
use scs8hd_decap_3  PHY_620
timestamp 1586364061
transform 1 0 1104 0 -1 171360
box -38 -48 314 592
use scs8hd_decap_3  PHY_622
timestamp 1586364061
transform 1 0 1104 0 1 171360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_310_3
timestamp 1586364061
transform 1 0 1380 0 -1 171360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_310_15
timestamp 1586364061
transform 1 0 2484 0 -1 171360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_311_3
timestamp 1586364061
transform 1 0 1380 0 1 171360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_311_15
timestamp 1586364061
transform 1 0 2484 0 1 171360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1519
timestamp 1586364061
transform 1 0 3956 0 -1 171360
box -38 -48 130 592
use scs8hd_decap_4  FILLER_310_27
timestamp 1586364061
transform 1 0 3588 0 -1 171360
box -38 -48 406 592
use scs8hd_decap_12  FILLER_310_32
timestamp 1586364061
transform 1 0 4048 0 -1 171360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_311_27
timestamp 1586364061
transform 1 0 3588 0 1 171360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_310_44
timestamp 1586364061
transform 1 0 5152 0 -1 171360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_311_39
timestamp 1586364061
transform 1 0 4692 0 1 171360
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_311_51
timestamp 1586364061
transform 1 0 5796 0 1 171360
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1520
timestamp 1586364061
transform 1 0 6716 0 1 171360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__19__A
timestamp 1586364061
transform 1 0 7452 0 1 171360
box -38 -48 222 592
use scs8hd_decap_12  FILLER_310_56
timestamp 1586364061
transform 1 0 6256 0 -1 171360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_310_68
timestamp 1586364061
transform 1 0 7360 0 -1 171360
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_311_59
timestamp 1586364061
transform 1 0 6532 0 1 171360
box -38 -48 222 592
use scs8hd_decap_6  FILLER_311_62
timestamp 1586364061
transform 1 0 6808 0 1 171360
box -38 -48 590 592
use scs8hd_fill_1  FILLER_311_68
timestamp 1586364061
transform 1 0 7360 0 1 171360
box -38 -48 130 592
use scs8hd_decap_8  FILLER_311_71
timestamp 1586364061
transform 1 0 7636 0 1 171360
box -38 -48 774 592
use scs8hd_decap_3  PHY_621
timestamp 1586364061
transform -1 0 8832 0 -1 171360
box -38 -48 314 592
use scs8hd_decap_3  PHY_623
timestamp 1586364061
transform -1 0 8832 0 1 171360
box -38 -48 314 592
use scs8hd_fill_1  FILLER_310_80
timestamp 1586364061
transform 1 0 8464 0 -1 171360
box -38 -48 130 592
use scs8hd_fill_2  FILLER_311_79
timestamp 1586364061
transform 1 0 8372 0 1 171360
box -38 -48 222 592
use scs8hd_decap_3  PHY_624
timestamp 1586364061
transform 1 0 1104 0 -1 172448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_312_3
timestamp 1586364061
transform 1 0 1380 0 -1 172448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_312_15
timestamp 1586364061
transform 1 0 2484 0 -1 172448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1521
timestamp 1586364061
transform 1 0 3956 0 -1 172448
box -38 -48 130 592
use scs8hd_decap_4  FILLER_312_27
timestamp 1586364061
transform 1 0 3588 0 -1 172448
box -38 -48 406 592
use scs8hd_decap_12  FILLER_312_32
timestamp 1586364061
transform 1 0 4048 0 -1 172448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_312_44
timestamp 1586364061
transform 1 0 5152 0 -1 172448
box -38 -48 1142 592
use scs8hd_buf_2  _19_
timestamp 1586364061
transform 1 0 7452 0 -1 172448
box -38 -48 406 592
use scs8hd_decap_12  FILLER_312_56
timestamp 1586364061
transform 1 0 6256 0 -1 172448
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_312_68
timestamp 1586364061
transform 1 0 7360 0 -1 172448
box -38 -48 130 592
use scs8hd_decap_3  PHY_625
timestamp 1586364061
transform -1 0 8832 0 -1 172448
box -38 -48 314 592
use scs8hd_decap_8  FILLER_312_73
timestamp 1586364061
transform 1 0 7820 0 -1 172448
box -38 -48 774 592
use scs8hd_decap_3  PHY_626
timestamp 1586364061
transform 1 0 1104 0 1 172448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_313_3
timestamp 1586364061
transform 1 0 1380 0 1 172448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_313_15
timestamp 1586364061
transform 1 0 2484 0 1 172448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_313_27
timestamp 1586364061
transform 1 0 3588 0 1 172448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_313_39
timestamp 1586364061
transform 1 0 4692 0 1 172448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_313_51
timestamp 1586364061
transform 1 0 5796 0 1 172448
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1522
timestamp 1586364061
transform 1 0 6716 0 1 172448
box -38 -48 130 592
use scs8hd_fill_2  FILLER_313_59
timestamp 1586364061
transform 1 0 6532 0 1 172448
box -38 -48 222 592
use scs8hd_decap_12  FILLER_313_62
timestamp 1586364061
transform 1 0 6808 0 1 172448
box -38 -48 1142 592
use scs8hd_decap_3  PHY_627
timestamp 1586364061
transform -1 0 8832 0 1 172448
box -38 -48 314 592
use scs8hd_decap_6  FILLER_313_74
timestamp 1586364061
transform 1 0 7912 0 1 172448
box -38 -48 590 592
use scs8hd_fill_1  FILLER_313_80
timestamp 1586364061
transform 1 0 8464 0 1 172448
box -38 -48 130 592
use scs8hd_decap_3  PHY_628
timestamp 1586364061
transform 1 0 1104 0 -1 173536
box -38 -48 314 592
use scs8hd_decap_12  FILLER_314_3
timestamp 1586364061
transform 1 0 1380 0 -1 173536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_314_15
timestamp 1586364061
transform 1 0 2484 0 -1 173536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1523
timestamp 1586364061
transform 1 0 3956 0 -1 173536
box -38 -48 130 592
use scs8hd_decap_4  FILLER_314_27
timestamp 1586364061
transform 1 0 3588 0 -1 173536
box -38 -48 406 592
use scs8hd_decap_12  FILLER_314_32
timestamp 1586364061
transform 1 0 4048 0 -1 173536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_314_44
timestamp 1586364061
transform 1 0 5152 0 -1 173536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_314_56
timestamp 1586364061
transform 1 0 6256 0 -1 173536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_314_68
timestamp 1586364061
transform 1 0 7360 0 -1 173536
box -38 -48 1142 592
use scs8hd_decap_3  PHY_629
timestamp 1586364061
transform -1 0 8832 0 -1 173536
box -38 -48 314 592
use scs8hd_fill_1  FILLER_314_80
timestamp 1586364061
transform 1 0 8464 0 -1 173536
box -38 -48 130 592
use scs8hd_decap_3  PHY_630
timestamp 1586364061
transform 1 0 1104 0 1 173536
box -38 -48 314 592
use scs8hd_decap_12  FILLER_315_3
timestamp 1586364061
transform 1 0 1380 0 1 173536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_315_15
timestamp 1586364061
transform 1 0 2484 0 1 173536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_315_27
timestamp 1586364061
transform 1 0 3588 0 1 173536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_315_39
timestamp 1586364061
transform 1 0 4692 0 1 173536
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_315_51
timestamp 1586364061
transform 1 0 5796 0 1 173536
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1524
timestamp 1586364061
transform 1 0 6716 0 1 173536
box -38 -48 130 592
use scs8hd_fill_2  FILLER_315_59
timestamp 1586364061
transform 1 0 6532 0 1 173536
box -38 -48 222 592
use scs8hd_decap_12  FILLER_315_62
timestamp 1586364061
transform 1 0 6808 0 1 173536
box -38 -48 1142 592
use scs8hd_decap_3  PHY_631
timestamp 1586364061
transform -1 0 8832 0 1 173536
box -38 -48 314 592
use scs8hd_decap_6  FILLER_315_74
timestamp 1586364061
transform 1 0 7912 0 1 173536
box -38 -48 590 592
use scs8hd_fill_1  FILLER_315_80
timestamp 1586364061
transform 1 0 8464 0 1 173536
box -38 -48 130 592
use scs8hd_decap_3  PHY_632
timestamp 1586364061
transform 1 0 1104 0 -1 174624
box -38 -48 314 592
use scs8hd_decap_12  FILLER_316_3
timestamp 1586364061
transform 1 0 1380 0 -1 174624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_316_15
timestamp 1586364061
transform 1 0 2484 0 -1 174624
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1525
timestamp 1586364061
transform 1 0 3956 0 -1 174624
box -38 -48 130 592
use scs8hd_decap_4  FILLER_316_27
timestamp 1586364061
transform 1 0 3588 0 -1 174624
box -38 -48 406 592
use scs8hd_decap_12  FILLER_316_32
timestamp 1586364061
transform 1 0 4048 0 -1 174624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_316_44
timestamp 1586364061
transform 1 0 5152 0 -1 174624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_316_56
timestamp 1586364061
transform 1 0 6256 0 -1 174624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_316_68
timestamp 1586364061
transform 1 0 7360 0 -1 174624
box -38 -48 1142 592
use scs8hd_decap_3  PHY_633
timestamp 1586364061
transform -1 0 8832 0 -1 174624
box -38 -48 314 592
use scs8hd_fill_1  FILLER_316_80
timestamp 1586364061
transform 1 0 8464 0 -1 174624
box -38 -48 130 592
use scs8hd_decap_3  PHY_634
timestamp 1586364061
transform 1 0 1104 0 1 174624
box -38 -48 314 592
use scs8hd_decap_3  PHY_636
timestamp 1586364061
transform 1 0 1104 0 -1 175712
box -38 -48 314 592
use scs8hd_decap_12  FILLER_317_3
timestamp 1586364061
transform 1 0 1380 0 1 174624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_317_15
timestamp 1586364061
transform 1 0 2484 0 1 174624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_318_3
timestamp 1586364061
transform 1 0 1380 0 -1 175712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_318_15
timestamp 1586364061
transform 1 0 2484 0 -1 175712
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1527
timestamp 1586364061
transform 1 0 3956 0 -1 175712
box -38 -48 130 592
use scs8hd_decap_12  FILLER_317_27
timestamp 1586364061
transform 1 0 3588 0 1 174624
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_318_27
timestamp 1586364061
transform 1 0 3588 0 -1 175712
box -38 -48 406 592
use scs8hd_decap_12  FILLER_318_32
timestamp 1586364061
transform 1 0 4048 0 -1 175712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_317_39
timestamp 1586364061
transform 1 0 4692 0 1 174624
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_317_51
timestamp 1586364061
transform 1 0 5796 0 1 174624
box -38 -48 774 592
use scs8hd_decap_12  FILLER_318_44
timestamp 1586364061
transform 1 0 5152 0 -1 175712
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1526
timestamp 1586364061
transform 1 0 6716 0 1 174624
box -38 -48 130 592
use scs8hd_fill_2  FILLER_317_59
timestamp 1586364061
transform 1 0 6532 0 1 174624
box -38 -48 222 592
use scs8hd_decap_12  FILLER_317_62
timestamp 1586364061
transform 1 0 6808 0 1 174624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_318_56
timestamp 1586364061
transform 1 0 6256 0 -1 175712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_318_68
timestamp 1586364061
transform 1 0 7360 0 -1 175712
box -38 -48 1142 592
use scs8hd_decap_3  PHY_635
timestamp 1586364061
transform -1 0 8832 0 1 174624
box -38 -48 314 592
use scs8hd_decap_3  PHY_637
timestamp 1586364061
transform -1 0 8832 0 -1 175712
box -38 -48 314 592
use scs8hd_decap_6  FILLER_317_74
timestamp 1586364061
transform 1 0 7912 0 1 174624
box -38 -48 590 592
use scs8hd_fill_1  FILLER_317_80
timestamp 1586364061
transform 1 0 8464 0 1 174624
box -38 -48 130 592
use scs8hd_fill_1  FILLER_318_80
timestamp 1586364061
transform 1 0 8464 0 -1 175712
box -38 -48 130 592
use scs8hd_decap_3  PHY_638
timestamp 1586364061
transform 1 0 1104 0 1 175712
box -38 -48 314 592
use scs8hd_decap_12  FILLER_319_3
timestamp 1586364061
transform 1 0 1380 0 1 175712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_319_15
timestamp 1586364061
transform 1 0 2484 0 1 175712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_319_27
timestamp 1586364061
transform 1 0 3588 0 1 175712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_319_39
timestamp 1586364061
transform 1 0 4692 0 1 175712
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_319_51
timestamp 1586364061
transform 1 0 5796 0 1 175712
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1528
timestamp 1586364061
transform 1 0 6716 0 1 175712
box -38 -48 130 592
use scs8hd_fill_2  FILLER_319_59
timestamp 1586364061
transform 1 0 6532 0 1 175712
box -38 -48 222 592
use scs8hd_decap_12  FILLER_319_62
timestamp 1586364061
transform 1 0 6808 0 1 175712
box -38 -48 1142 592
use scs8hd_decap_3  PHY_639
timestamp 1586364061
transform -1 0 8832 0 1 175712
box -38 -48 314 592
use scs8hd_decap_6  FILLER_319_74
timestamp 1586364061
transform 1 0 7912 0 1 175712
box -38 -48 590 592
use scs8hd_fill_1  FILLER_319_80
timestamp 1586364061
transform 1 0 8464 0 1 175712
box -38 -48 130 592
use scs8hd_decap_3  PHY_640
timestamp 1586364061
transform 1 0 1104 0 -1 176800
box -38 -48 314 592
use scs8hd_decap_12  FILLER_320_3
timestamp 1586364061
transform 1 0 1380 0 -1 176800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_320_15
timestamp 1586364061
transform 1 0 2484 0 -1 176800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1529
timestamp 1586364061
transform 1 0 3956 0 -1 176800
box -38 -48 130 592
use scs8hd_decap_4  FILLER_320_27
timestamp 1586364061
transform 1 0 3588 0 -1 176800
box -38 -48 406 592
use scs8hd_decap_12  FILLER_320_32
timestamp 1586364061
transform 1 0 4048 0 -1 176800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_320_44
timestamp 1586364061
transform 1 0 5152 0 -1 176800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_320_56
timestamp 1586364061
transform 1 0 6256 0 -1 176800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_320_68
timestamp 1586364061
transform 1 0 7360 0 -1 176800
box -38 -48 1142 592
use scs8hd_decap_3  PHY_641
timestamp 1586364061
transform -1 0 8832 0 -1 176800
box -38 -48 314 592
use scs8hd_fill_1  FILLER_320_80
timestamp 1586364061
transform 1 0 8464 0 -1 176800
box -38 -48 130 592
use scs8hd_decap_3  PHY_642
timestamp 1586364061
transform 1 0 1104 0 1 176800
box -38 -48 314 592
use scs8hd_decap_12  FILLER_321_3
timestamp 1586364061
transform 1 0 1380 0 1 176800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_321_15
timestamp 1586364061
transform 1 0 2484 0 1 176800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_321_27
timestamp 1586364061
transform 1 0 3588 0 1 176800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_321_39
timestamp 1586364061
transform 1 0 4692 0 1 176800
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_321_51
timestamp 1586364061
transform 1 0 5796 0 1 176800
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1530
timestamp 1586364061
transform 1 0 6716 0 1 176800
box -38 -48 130 592
use scs8hd_fill_2  FILLER_321_59
timestamp 1586364061
transform 1 0 6532 0 1 176800
box -38 -48 222 592
use scs8hd_decap_12  FILLER_321_62
timestamp 1586364061
transform 1 0 6808 0 1 176800
box -38 -48 1142 592
use scs8hd_decap_3  PHY_643
timestamp 1586364061
transform -1 0 8832 0 1 176800
box -38 -48 314 592
use scs8hd_decap_6  FILLER_321_74
timestamp 1586364061
transform 1 0 7912 0 1 176800
box -38 -48 590 592
use scs8hd_fill_1  FILLER_321_80
timestamp 1586364061
transform 1 0 8464 0 1 176800
box -38 -48 130 592
use scs8hd_decap_3  PHY_644
timestamp 1586364061
transform 1 0 1104 0 -1 177888
box -38 -48 314 592
use scs8hd_decap_12  FILLER_322_3
timestamp 1586364061
transform 1 0 1380 0 -1 177888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_322_15
timestamp 1586364061
transform 1 0 2484 0 -1 177888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1531
timestamp 1586364061
transform 1 0 3956 0 -1 177888
box -38 -48 130 592
use scs8hd_decap_4  FILLER_322_27
timestamp 1586364061
transform 1 0 3588 0 -1 177888
box -38 -48 406 592
use scs8hd_decap_12  FILLER_322_32
timestamp 1586364061
transform 1 0 4048 0 -1 177888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_322_44
timestamp 1586364061
transform 1 0 5152 0 -1 177888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_322_56
timestamp 1586364061
transform 1 0 6256 0 -1 177888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_322_68
timestamp 1586364061
transform 1 0 7360 0 -1 177888
box -38 -48 1142 592
use scs8hd_decap_3  PHY_645
timestamp 1586364061
transform -1 0 8832 0 -1 177888
box -38 -48 314 592
use scs8hd_fill_1  FILLER_322_80
timestamp 1586364061
transform 1 0 8464 0 -1 177888
box -38 -48 130 592
use scs8hd_decap_3  PHY_646
timestamp 1586364061
transform 1 0 1104 0 1 177888
box -38 -48 314 592
use scs8hd_decap_3  PHY_648
timestamp 1586364061
transform 1 0 1104 0 -1 178976
box -38 -48 314 592
use scs8hd_decap_12  FILLER_323_3
timestamp 1586364061
transform 1 0 1380 0 1 177888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_323_15
timestamp 1586364061
transform 1 0 2484 0 1 177888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_324_3
timestamp 1586364061
transform 1 0 1380 0 -1 178976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_324_15
timestamp 1586364061
transform 1 0 2484 0 -1 178976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1533
timestamp 1586364061
transform 1 0 3956 0 -1 178976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_323_27
timestamp 1586364061
transform 1 0 3588 0 1 177888
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_324_27
timestamp 1586364061
transform 1 0 3588 0 -1 178976
box -38 -48 406 592
use scs8hd_decap_12  FILLER_324_32
timestamp 1586364061
transform 1 0 4048 0 -1 178976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_323_39
timestamp 1586364061
transform 1 0 4692 0 1 177888
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_323_51
timestamp 1586364061
transform 1 0 5796 0 1 177888
box -38 -48 774 592
use scs8hd_decap_12  FILLER_324_44
timestamp 1586364061
transform 1 0 5152 0 -1 178976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1532
timestamp 1586364061
transform 1 0 6716 0 1 177888
box -38 -48 130 592
use scs8hd_fill_2  FILLER_323_59
timestamp 1586364061
transform 1 0 6532 0 1 177888
box -38 -48 222 592
use scs8hd_decap_12  FILLER_323_62
timestamp 1586364061
transform 1 0 6808 0 1 177888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_324_56
timestamp 1586364061
transform 1 0 6256 0 -1 178976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_324_68
timestamp 1586364061
transform 1 0 7360 0 -1 178976
box -38 -48 1142 592
use scs8hd_decap_3  PHY_647
timestamp 1586364061
transform -1 0 8832 0 1 177888
box -38 -48 314 592
use scs8hd_decap_3  PHY_649
timestamp 1586364061
transform -1 0 8832 0 -1 178976
box -38 -48 314 592
use scs8hd_decap_6  FILLER_323_74
timestamp 1586364061
transform 1 0 7912 0 1 177888
box -38 -48 590 592
use scs8hd_fill_1  FILLER_323_80
timestamp 1586364061
transform 1 0 8464 0 1 177888
box -38 -48 130 592
use scs8hd_fill_1  FILLER_324_80
timestamp 1586364061
transform 1 0 8464 0 -1 178976
box -38 -48 130 592
use scs8hd_decap_3  PHY_650
timestamp 1586364061
transform 1 0 1104 0 1 178976
box -38 -48 314 592
use scs8hd_decap_12  FILLER_325_3
timestamp 1586364061
transform 1 0 1380 0 1 178976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_325_15
timestamp 1586364061
transform 1 0 2484 0 1 178976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_325_27
timestamp 1586364061
transform 1 0 3588 0 1 178976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_325_39
timestamp 1586364061
transform 1 0 4692 0 1 178976
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_325_51
timestamp 1586364061
transform 1 0 5796 0 1 178976
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1534
timestamp 1586364061
transform 1 0 6716 0 1 178976
box -38 -48 130 592
use scs8hd_fill_2  FILLER_325_59
timestamp 1586364061
transform 1 0 6532 0 1 178976
box -38 -48 222 592
use scs8hd_decap_12  FILLER_325_62
timestamp 1586364061
transform 1 0 6808 0 1 178976
box -38 -48 1142 592
use scs8hd_decap_3  PHY_651
timestamp 1586364061
transform -1 0 8832 0 1 178976
box -38 -48 314 592
use scs8hd_decap_6  FILLER_325_74
timestamp 1586364061
transform 1 0 7912 0 1 178976
box -38 -48 590 592
use scs8hd_fill_1  FILLER_325_80
timestamp 1586364061
transform 1 0 8464 0 1 178976
box -38 -48 130 592
use scs8hd_decap_3  PHY_652
timestamp 1586364061
transform 1 0 1104 0 -1 180064
box -38 -48 314 592
use scs8hd_decap_12  FILLER_326_3
timestamp 1586364061
transform 1 0 1380 0 -1 180064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_326_15
timestamp 1586364061
transform 1 0 2484 0 -1 180064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1535
timestamp 1586364061
transform 1 0 3956 0 -1 180064
box -38 -48 130 592
use scs8hd_decap_4  FILLER_326_27
timestamp 1586364061
transform 1 0 3588 0 -1 180064
box -38 -48 406 592
use scs8hd_decap_12  FILLER_326_32
timestamp 1586364061
transform 1 0 4048 0 -1 180064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_326_44
timestamp 1586364061
transform 1 0 5152 0 -1 180064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_326_56
timestamp 1586364061
transform 1 0 6256 0 -1 180064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_326_68
timestamp 1586364061
transform 1 0 7360 0 -1 180064
box -38 -48 1142 592
use scs8hd_decap_3  PHY_653
timestamp 1586364061
transform -1 0 8832 0 -1 180064
box -38 -48 314 592
use scs8hd_fill_1  FILLER_326_80
timestamp 1586364061
transform 1 0 8464 0 -1 180064
box -38 -48 130 592
use scs8hd_decap_3  PHY_654
timestamp 1586364061
transform 1 0 1104 0 1 180064
box -38 -48 314 592
use scs8hd_decap_12  FILLER_327_3
timestamp 1586364061
transform 1 0 1380 0 1 180064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_327_15
timestamp 1586364061
transform 1 0 2484 0 1 180064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_327_27
timestamp 1586364061
transform 1 0 3588 0 1 180064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_327_39
timestamp 1586364061
transform 1 0 4692 0 1 180064
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_327_51
timestamp 1586364061
transform 1 0 5796 0 1 180064
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1536
timestamp 1586364061
transform 1 0 6716 0 1 180064
box -38 -48 130 592
use scs8hd_fill_2  FILLER_327_59
timestamp 1586364061
transform 1 0 6532 0 1 180064
box -38 -48 222 592
use scs8hd_decap_12  FILLER_327_62
timestamp 1586364061
transform 1 0 6808 0 1 180064
box -38 -48 1142 592
use scs8hd_decap_3  PHY_655
timestamp 1586364061
transform -1 0 8832 0 1 180064
box -38 -48 314 592
use scs8hd_decap_6  FILLER_327_74
timestamp 1586364061
transform 1 0 7912 0 1 180064
box -38 -48 590 592
use scs8hd_fill_1  FILLER_327_80
timestamp 1586364061
transform 1 0 8464 0 1 180064
box -38 -48 130 592
use scs8hd_decap_3  PHY_656
timestamp 1586364061
transform 1 0 1104 0 -1 181152
box -38 -48 314 592
use scs8hd_decap_12  FILLER_328_3
timestamp 1586364061
transform 1 0 1380 0 -1 181152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_328_15
timestamp 1586364061
transform 1 0 2484 0 -1 181152
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1537
timestamp 1586364061
transform 1 0 3956 0 -1 181152
box -38 -48 130 592
use scs8hd_decap_4  FILLER_328_27
timestamp 1586364061
transform 1 0 3588 0 -1 181152
box -38 -48 406 592
use scs8hd_decap_12  FILLER_328_32
timestamp 1586364061
transform 1 0 4048 0 -1 181152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_328_44
timestamp 1586364061
transform 1 0 5152 0 -1 181152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_328_56
timestamp 1586364061
transform 1 0 6256 0 -1 181152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_328_68
timestamp 1586364061
transform 1 0 7360 0 -1 181152
box -38 -48 1142 592
use scs8hd_decap_3  PHY_657
timestamp 1586364061
transform -1 0 8832 0 -1 181152
box -38 -48 314 592
use scs8hd_fill_1  FILLER_328_80
timestamp 1586364061
transform 1 0 8464 0 -1 181152
box -38 -48 130 592
use scs8hd_decap_3  PHY_658
timestamp 1586364061
transform 1 0 1104 0 1 181152
box -38 -48 314 592
use scs8hd_decap_12  FILLER_329_3
timestamp 1586364061
transform 1 0 1380 0 1 181152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_329_15
timestamp 1586364061
transform 1 0 2484 0 1 181152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_329_27
timestamp 1586364061
transform 1 0 3588 0 1 181152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_329_39
timestamp 1586364061
transform 1 0 4692 0 1 181152
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_329_51
timestamp 1586364061
transform 1 0 5796 0 1 181152
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1538
timestamp 1586364061
transform 1 0 6716 0 1 181152
box -38 -48 130 592
use scs8hd_fill_2  FILLER_329_59
timestamp 1586364061
transform 1 0 6532 0 1 181152
box -38 -48 222 592
use scs8hd_decap_12  FILLER_329_62
timestamp 1586364061
transform 1 0 6808 0 1 181152
box -38 -48 1142 592
use scs8hd_decap_3  PHY_659
timestamp 1586364061
transform -1 0 8832 0 1 181152
box -38 -48 314 592
use scs8hd_decap_6  FILLER_329_74
timestamp 1586364061
transform 1 0 7912 0 1 181152
box -38 -48 590 592
use scs8hd_fill_1  FILLER_329_80
timestamp 1586364061
transform 1 0 8464 0 1 181152
box -38 -48 130 592
use scs8hd_decap_3  PHY_660
timestamp 1586364061
transform 1 0 1104 0 -1 182240
box -38 -48 314 592
use scs8hd_decap_3  PHY_662
timestamp 1586364061
transform 1 0 1104 0 1 182240
box -38 -48 314 592
use scs8hd_decap_12  FILLER_330_3
timestamp 1586364061
transform 1 0 1380 0 -1 182240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_330_15
timestamp 1586364061
transform 1 0 2484 0 -1 182240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_331_3
timestamp 1586364061
transform 1 0 1380 0 1 182240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_331_15
timestamp 1586364061
transform 1 0 2484 0 1 182240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1539
timestamp 1586364061
transform 1 0 3956 0 -1 182240
box -38 -48 130 592
use scs8hd_decap_4  FILLER_330_27
timestamp 1586364061
transform 1 0 3588 0 -1 182240
box -38 -48 406 592
use scs8hd_decap_12  FILLER_330_32
timestamp 1586364061
transform 1 0 4048 0 -1 182240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_331_27
timestamp 1586364061
transform 1 0 3588 0 1 182240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_330_44
timestamp 1586364061
transform 1 0 5152 0 -1 182240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_331_39
timestamp 1586364061
transform 1 0 4692 0 1 182240
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_331_51
timestamp 1586364061
transform 1 0 5796 0 1 182240
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1540
timestamp 1586364061
transform 1 0 6716 0 1 182240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_330_56
timestamp 1586364061
transform 1 0 6256 0 -1 182240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_330_68
timestamp 1586364061
transform 1 0 7360 0 -1 182240
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_331_59
timestamp 1586364061
transform 1 0 6532 0 1 182240
box -38 -48 222 592
use scs8hd_decap_12  FILLER_331_62
timestamp 1586364061
transform 1 0 6808 0 1 182240
box -38 -48 1142 592
use scs8hd_decap_3  PHY_661
timestamp 1586364061
transform -1 0 8832 0 -1 182240
box -38 -48 314 592
use scs8hd_decap_3  PHY_663
timestamp 1586364061
transform -1 0 8832 0 1 182240
box -38 -48 314 592
use scs8hd_fill_1  FILLER_330_80
timestamp 1586364061
transform 1 0 8464 0 -1 182240
box -38 -48 130 592
use scs8hd_decap_6  FILLER_331_74
timestamp 1586364061
transform 1 0 7912 0 1 182240
box -38 -48 590 592
use scs8hd_fill_1  FILLER_331_80
timestamp 1586364061
transform 1 0 8464 0 1 182240
box -38 -48 130 592
use scs8hd_decap_3  PHY_664
timestamp 1586364061
transform 1 0 1104 0 -1 183328
box -38 -48 314 592
use scs8hd_decap_12  FILLER_332_3
timestamp 1586364061
transform 1 0 1380 0 -1 183328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_332_15
timestamp 1586364061
transform 1 0 2484 0 -1 183328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1541
timestamp 1586364061
transform 1 0 3956 0 -1 183328
box -38 -48 130 592
use scs8hd_decap_4  FILLER_332_27
timestamp 1586364061
transform 1 0 3588 0 -1 183328
box -38 -48 406 592
use scs8hd_decap_12  FILLER_332_32
timestamp 1586364061
transform 1 0 4048 0 -1 183328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_332_44
timestamp 1586364061
transform 1 0 5152 0 -1 183328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_332_56
timestamp 1586364061
transform 1 0 6256 0 -1 183328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_332_68
timestamp 1586364061
transform 1 0 7360 0 -1 183328
box -38 -48 1142 592
use scs8hd_decap_3  PHY_665
timestamp 1586364061
transform -1 0 8832 0 -1 183328
box -38 -48 314 592
use scs8hd_fill_1  FILLER_332_80
timestamp 1586364061
transform 1 0 8464 0 -1 183328
box -38 -48 130 592
use scs8hd_decap_3  PHY_666
timestamp 1586364061
transform 1 0 1104 0 1 183328
box -38 -48 314 592
use scs8hd_decap_12  FILLER_333_3
timestamp 1586364061
transform 1 0 1380 0 1 183328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_333_15
timestamp 1586364061
transform 1 0 2484 0 1 183328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_333_27
timestamp 1586364061
transform 1 0 3588 0 1 183328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_333_39
timestamp 1586364061
transform 1 0 4692 0 1 183328
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_333_51
timestamp 1586364061
transform 1 0 5796 0 1 183328
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1542
timestamp 1586364061
transform 1 0 6716 0 1 183328
box -38 -48 130 592
use scs8hd_fill_2  FILLER_333_59
timestamp 1586364061
transform 1 0 6532 0 1 183328
box -38 -48 222 592
use scs8hd_decap_12  FILLER_333_62
timestamp 1586364061
transform 1 0 6808 0 1 183328
box -38 -48 1142 592
use scs8hd_decap_3  PHY_667
timestamp 1586364061
transform -1 0 8832 0 1 183328
box -38 -48 314 592
use scs8hd_decap_6  FILLER_333_74
timestamp 1586364061
transform 1 0 7912 0 1 183328
box -38 -48 590 592
use scs8hd_fill_1  FILLER_333_80
timestamp 1586364061
transform 1 0 8464 0 1 183328
box -38 -48 130 592
use scs8hd_decap_3  PHY_668
timestamp 1586364061
transform 1 0 1104 0 -1 184416
box -38 -48 314 592
use scs8hd_decap_12  FILLER_334_3
timestamp 1586364061
transform 1 0 1380 0 -1 184416
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_334_15
timestamp 1586364061
transform 1 0 2484 0 -1 184416
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1543
timestamp 1586364061
transform 1 0 3956 0 -1 184416
box -38 -48 130 592
use scs8hd_decap_4  FILLER_334_27
timestamp 1586364061
transform 1 0 3588 0 -1 184416
box -38 -48 406 592
use scs8hd_decap_12  FILLER_334_32
timestamp 1586364061
transform 1 0 4048 0 -1 184416
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_334_44
timestamp 1586364061
transform 1 0 5152 0 -1 184416
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_334_56
timestamp 1586364061
transform 1 0 6256 0 -1 184416
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_334_68
timestamp 1586364061
transform 1 0 7360 0 -1 184416
box -38 -48 1142 592
use scs8hd_decap_3  PHY_669
timestamp 1586364061
transform -1 0 8832 0 -1 184416
box -38 -48 314 592
use scs8hd_fill_1  FILLER_334_80
timestamp 1586364061
transform 1 0 8464 0 -1 184416
box -38 -48 130 592
use scs8hd_decap_3  PHY_670
timestamp 1586364061
transform 1 0 1104 0 1 184416
box -38 -48 314 592
use scs8hd_decap_12  FILLER_335_3
timestamp 1586364061
transform 1 0 1380 0 1 184416
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_335_15
timestamp 1586364061
transform 1 0 2484 0 1 184416
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_335_27
timestamp 1586364061
transform 1 0 3588 0 1 184416
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_335_39
timestamp 1586364061
transform 1 0 4692 0 1 184416
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_335_51
timestamp 1586364061
transform 1 0 5796 0 1 184416
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1544
timestamp 1586364061
transform 1 0 6716 0 1 184416
box -38 -48 130 592
use scs8hd_fill_2  FILLER_335_59
timestamp 1586364061
transform 1 0 6532 0 1 184416
box -38 -48 222 592
use scs8hd_decap_12  FILLER_335_62
timestamp 1586364061
transform 1 0 6808 0 1 184416
box -38 -48 1142 592
use scs8hd_decap_3  PHY_671
timestamp 1586364061
transform -1 0 8832 0 1 184416
box -38 -48 314 592
use scs8hd_decap_6  FILLER_335_74
timestamp 1586364061
transform 1 0 7912 0 1 184416
box -38 -48 590 592
use scs8hd_fill_1  FILLER_335_80
timestamp 1586364061
transform 1 0 8464 0 1 184416
box -38 -48 130 592
use scs8hd_decap_3  PHY_672
timestamp 1586364061
transform 1 0 1104 0 -1 185504
box -38 -48 314 592
use scs8hd_decap_12  FILLER_336_3
timestamp 1586364061
transform 1 0 1380 0 -1 185504
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_336_15
timestamp 1586364061
transform 1 0 2484 0 -1 185504
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1545
timestamp 1586364061
transform 1 0 3956 0 -1 185504
box -38 -48 130 592
use scs8hd_decap_4  FILLER_336_27
timestamp 1586364061
transform 1 0 3588 0 -1 185504
box -38 -48 406 592
use scs8hd_decap_12  FILLER_336_32
timestamp 1586364061
transform 1 0 4048 0 -1 185504
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_336_44
timestamp 1586364061
transform 1 0 5152 0 -1 185504
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_336_56
timestamp 1586364061
transform 1 0 6256 0 -1 185504
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_336_68
timestamp 1586364061
transform 1 0 7360 0 -1 185504
box -38 -48 1142 592
use scs8hd_decap_3  PHY_673
timestamp 1586364061
transform -1 0 8832 0 -1 185504
box -38 -48 314 592
use scs8hd_fill_1  FILLER_336_80
timestamp 1586364061
transform 1 0 8464 0 -1 185504
box -38 -48 130 592
use scs8hd_decap_3  PHY_674
timestamp 1586364061
transform 1 0 1104 0 1 185504
box -38 -48 314 592
use scs8hd_decap_3  PHY_676
timestamp 1586364061
transform 1 0 1104 0 -1 186592
box -38 -48 314 592
use scs8hd_decap_12  FILLER_337_3
timestamp 1586364061
transform 1 0 1380 0 1 185504
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_337_15
timestamp 1586364061
transform 1 0 2484 0 1 185504
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_338_3
timestamp 1586364061
transform 1 0 1380 0 -1 186592
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_338_15
timestamp 1586364061
transform 1 0 2484 0 -1 186592
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1547
timestamp 1586364061
transform 1 0 3956 0 -1 186592
box -38 -48 130 592
use scs8hd_decap_12  FILLER_337_27
timestamp 1586364061
transform 1 0 3588 0 1 185504
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_338_27
timestamp 1586364061
transform 1 0 3588 0 -1 186592
box -38 -48 406 592
use scs8hd_decap_12  FILLER_338_32
timestamp 1586364061
transform 1 0 4048 0 -1 186592
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_337_39
timestamp 1586364061
transform 1 0 4692 0 1 185504
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_337_51
timestamp 1586364061
transform 1 0 5796 0 1 185504
box -38 -48 774 592
use scs8hd_decap_12  FILLER_338_44
timestamp 1586364061
transform 1 0 5152 0 -1 186592
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1546
timestamp 1586364061
transform 1 0 6716 0 1 185504
box -38 -48 130 592
use scs8hd_fill_2  FILLER_337_59
timestamp 1586364061
transform 1 0 6532 0 1 185504
box -38 -48 222 592
use scs8hd_decap_12  FILLER_337_62
timestamp 1586364061
transform 1 0 6808 0 1 185504
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_338_56
timestamp 1586364061
transform 1 0 6256 0 -1 186592
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_338_68
timestamp 1586364061
transform 1 0 7360 0 -1 186592
box -38 -48 1142 592
use scs8hd_decap_3  PHY_675
timestamp 1586364061
transform -1 0 8832 0 1 185504
box -38 -48 314 592
use scs8hd_decap_3  PHY_677
timestamp 1586364061
transform -1 0 8832 0 -1 186592
box -38 -48 314 592
use scs8hd_decap_6  FILLER_337_74
timestamp 1586364061
transform 1 0 7912 0 1 185504
box -38 -48 590 592
use scs8hd_fill_1  FILLER_337_80
timestamp 1586364061
transform 1 0 8464 0 1 185504
box -38 -48 130 592
use scs8hd_fill_1  FILLER_338_80
timestamp 1586364061
transform 1 0 8464 0 -1 186592
box -38 -48 130 592
use scs8hd_decap_3  PHY_678
timestamp 1586364061
transform 1 0 1104 0 1 186592
box -38 -48 314 592
use scs8hd_decap_12  FILLER_339_3
timestamp 1586364061
transform 1 0 1380 0 1 186592
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_339_15
timestamp 1586364061
transform 1 0 2484 0 1 186592
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_339_27
timestamp 1586364061
transform 1 0 3588 0 1 186592
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_339_39
timestamp 1586364061
transform 1 0 4692 0 1 186592
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_339_51
timestamp 1586364061
transform 1 0 5796 0 1 186592
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1548
timestamp 1586364061
transform 1 0 6716 0 1 186592
box -38 -48 130 592
use scs8hd_fill_2  FILLER_339_59
timestamp 1586364061
transform 1 0 6532 0 1 186592
box -38 -48 222 592
use scs8hd_decap_12  FILLER_339_62
timestamp 1586364061
transform 1 0 6808 0 1 186592
box -38 -48 1142 592
use scs8hd_decap_3  PHY_679
timestamp 1586364061
transform -1 0 8832 0 1 186592
box -38 -48 314 592
use scs8hd_decap_6  FILLER_339_74
timestamp 1586364061
transform 1 0 7912 0 1 186592
box -38 -48 590 592
use scs8hd_fill_1  FILLER_339_80
timestamp 1586364061
transform 1 0 8464 0 1 186592
box -38 -48 130 592
use scs8hd_decap_3  PHY_680
timestamp 1586364061
transform 1 0 1104 0 -1 187680
box -38 -48 314 592
use scs8hd_decap_12  FILLER_340_3
timestamp 1586364061
transform 1 0 1380 0 -1 187680
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_340_15
timestamp 1586364061
transform 1 0 2484 0 -1 187680
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1549
timestamp 1586364061
transform 1 0 3956 0 -1 187680
box -38 -48 130 592
use scs8hd_decap_4  FILLER_340_27
timestamp 1586364061
transform 1 0 3588 0 -1 187680
box -38 -48 406 592
use scs8hd_decap_12  FILLER_340_32
timestamp 1586364061
transform 1 0 4048 0 -1 187680
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_340_44
timestamp 1586364061
transform 1 0 5152 0 -1 187680
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_340_56
timestamp 1586364061
transform 1 0 6256 0 -1 187680
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_340_68
timestamp 1586364061
transform 1 0 7360 0 -1 187680
box -38 -48 1142 592
use scs8hd_decap_3  PHY_681
timestamp 1586364061
transform -1 0 8832 0 -1 187680
box -38 -48 314 592
use scs8hd_fill_1  FILLER_340_80
timestamp 1586364061
transform 1 0 8464 0 -1 187680
box -38 -48 130 592
use scs8hd_decap_3  PHY_682
timestamp 1586364061
transform 1 0 1104 0 1 187680
box -38 -48 314 592
use scs8hd_decap_12  FILLER_341_3
timestamp 1586364061
transform 1 0 1380 0 1 187680
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_341_15
timestamp 1586364061
transform 1 0 2484 0 1 187680
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_341_27
timestamp 1586364061
transform 1 0 3588 0 1 187680
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_341_39
timestamp 1586364061
transform 1 0 4692 0 1 187680
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_341_51
timestamp 1586364061
transform 1 0 5796 0 1 187680
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1550
timestamp 1586364061
transform 1 0 6716 0 1 187680
box -38 -48 130 592
use scs8hd_fill_2  FILLER_341_59
timestamp 1586364061
transform 1 0 6532 0 1 187680
box -38 -48 222 592
use scs8hd_decap_12  FILLER_341_62
timestamp 1586364061
transform 1 0 6808 0 1 187680
box -38 -48 1142 592
use scs8hd_decap_3  PHY_683
timestamp 1586364061
transform -1 0 8832 0 1 187680
box -38 -48 314 592
use scs8hd_decap_6  FILLER_341_74
timestamp 1586364061
transform 1 0 7912 0 1 187680
box -38 -48 590 592
use scs8hd_fill_1  FILLER_341_80
timestamp 1586364061
transform 1 0 8464 0 1 187680
box -38 -48 130 592
use scs8hd_decap_3  PHY_684
timestamp 1586364061
transform 1 0 1104 0 -1 188768
box -38 -48 314 592
use scs8hd_decap_12  FILLER_342_3
timestamp 1586364061
transform 1 0 1380 0 -1 188768
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_342_15
timestamp 1586364061
transform 1 0 2484 0 -1 188768
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1551
timestamp 1586364061
transform 1 0 3956 0 -1 188768
box -38 -48 130 592
use scs8hd_decap_4  FILLER_342_27
timestamp 1586364061
transform 1 0 3588 0 -1 188768
box -38 -48 406 592
use scs8hd_decap_12  FILLER_342_32
timestamp 1586364061
transform 1 0 4048 0 -1 188768
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_342_44
timestamp 1586364061
transform 1 0 5152 0 -1 188768
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_342_56
timestamp 1586364061
transform 1 0 6256 0 -1 188768
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_342_68
timestamp 1586364061
transform 1 0 7360 0 -1 188768
box -38 -48 1142 592
use scs8hd_decap_3  PHY_685
timestamp 1586364061
transform -1 0 8832 0 -1 188768
box -38 -48 314 592
use scs8hd_fill_1  FILLER_342_80
timestamp 1586364061
transform 1 0 8464 0 -1 188768
box -38 -48 130 592
use scs8hd_decap_3  PHY_686
timestamp 1586364061
transform 1 0 1104 0 1 188768
box -38 -48 314 592
use scs8hd_decap_3  PHY_688
timestamp 1586364061
transform 1 0 1104 0 -1 189856
box -38 -48 314 592
use scs8hd_decap_12  FILLER_343_3
timestamp 1586364061
transform 1 0 1380 0 1 188768
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_343_15
timestamp 1586364061
transform 1 0 2484 0 1 188768
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_344_3
timestamp 1586364061
transform 1 0 1380 0 -1 189856
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_344_15
timestamp 1586364061
transform 1 0 2484 0 -1 189856
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1553
timestamp 1586364061
transform 1 0 3956 0 -1 189856
box -38 -48 130 592
use scs8hd_decap_12  FILLER_343_27
timestamp 1586364061
transform 1 0 3588 0 1 188768
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_344_27
timestamp 1586364061
transform 1 0 3588 0 -1 189856
box -38 -48 406 592
use scs8hd_decap_12  FILLER_344_32
timestamp 1586364061
transform 1 0 4048 0 -1 189856
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_343_39
timestamp 1586364061
transform 1 0 4692 0 1 188768
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_343_51
timestamp 1586364061
transform 1 0 5796 0 1 188768
box -38 -48 774 592
use scs8hd_decap_12  FILLER_344_44
timestamp 1586364061
transform 1 0 5152 0 -1 189856
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1552
timestamp 1586364061
transform 1 0 6716 0 1 188768
box -38 -48 130 592
use scs8hd_fill_2  FILLER_343_59
timestamp 1586364061
transform 1 0 6532 0 1 188768
box -38 -48 222 592
use scs8hd_decap_12  FILLER_343_62
timestamp 1586364061
transform 1 0 6808 0 1 188768
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_344_56
timestamp 1586364061
transform 1 0 6256 0 -1 189856
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_344_68
timestamp 1586364061
transform 1 0 7360 0 -1 189856
box -38 -48 1142 592
use scs8hd_decap_3  PHY_687
timestamp 1586364061
transform -1 0 8832 0 1 188768
box -38 -48 314 592
use scs8hd_decap_3  PHY_689
timestamp 1586364061
transform -1 0 8832 0 -1 189856
box -38 -48 314 592
use scs8hd_decap_6  FILLER_343_74
timestamp 1586364061
transform 1 0 7912 0 1 188768
box -38 -48 590 592
use scs8hd_fill_1  FILLER_343_80
timestamp 1586364061
transform 1 0 8464 0 1 188768
box -38 -48 130 592
use scs8hd_fill_1  FILLER_344_80
timestamp 1586364061
transform 1 0 8464 0 -1 189856
box -38 -48 130 592
use scs8hd_decap_3  PHY_690
timestamp 1586364061
transform 1 0 1104 0 1 189856
box -38 -48 314 592
use scs8hd_decap_12  FILLER_345_3
timestamp 1586364061
transform 1 0 1380 0 1 189856
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_345_15
timestamp 1586364061
transform 1 0 2484 0 1 189856
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_345_27
timestamp 1586364061
transform 1 0 3588 0 1 189856
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_345_39
timestamp 1586364061
transform 1 0 4692 0 1 189856
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_345_51
timestamp 1586364061
transform 1 0 5796 0 1 189856
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1554
timestamp 1586364061
transform 1 0 6716 0 1 189856
box -38 -48 130 592
use scs8hd_fill_2  FILLER_345_59
timestamp 1586364061
transform 1 0 6532 0 1 189856
box -38 -48 222 592
use scs8hd_decap_12  FILLER_345_62
timestamp 1586364061
transform 1 0 6808 0 1 189856
box -38 -48 1142 592
use scs8hd_decap_3  PHY_691
timestamp 1586364061
transform -1 0 8832 0 1 189856
box -38 -48 314 592
use scs8hd_decap_6  FILLER_345_74
timestamp 1586364061
transform 1 0 7912 0 1 189856
box -38 -48 590 592
use scs8hd_fill_1  FILLER_345_80
timestamp 1586364061
transform 1 0 8464 0 1 189856
box -38 -48 130 592
use scs8hd_decap_3  PHY_692
timestamp 1586364061
transform 1 0 1104 0 -1 190944
box -38 -48 314 592
use scs8hd_decap_12  FILLER_346_3
timestamp 1586364061
transform 1 0 1380 0 -1 190944
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_346_15
timestamp 1586364061
transform 1 0 2484 0 -1 190944
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1555
timestamp 1586364061
transform 1 0 3956 0 -1 190944
box -38 -48 130 592
use scs8hd_decap_4  FILLER_346_27
timestamp 1586364061
transform 1 0 3588 0 -1 190944
box -38 -48 406 592
use scs8hd_decap_12  FILLER_346_32
timestamp 1586364061
transform 1 0 4048 0 -1 190944
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_346_44
timestamp 1586364061
transform 1 0 5152 0 -1 190944
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_346_56
timestamp 1586364061
transform 1 0 6256 0 -1 190944
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_346_68
timestamp 1586364061
transform 1 0 7360 0 -1 190944
box -38 -48 1142 592
use scs8hd_decap_3  PHY_693
timestamp 1586364061
transform -1 0 8832 0 -1 190944
box -38 -48 314 592
use scs8hd_fill_1  FILLER_346_80
timestamp 1586364061
transform 1 0 8464 0 -1 190944
box -38 -48 130 592
use scs8hd_decap_3  PHY_694
timestamp 1586364061
transform 1 0 1104 0 1 190944
box -38 -48 314 592
use scs8hd_decap_12  FILLER_347_3
timestamp 1586364061
transform 1 0 1380 0 1 190944
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_347_15
timestamp 1586364061
transform 1 0 2484 0 1 190944
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_347_27
timestamp 1586364061
transform 1 0 3588 0 1 190944
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_347_39
timestamp 1586364061
transform 1 0 4692 0 1 190944
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_347_51
timestamp 1586364061
transform 1 0 5796 0 1 190944
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1556
timestamp 1586364061
transform 1 0 6716 0 1 190944
box -38 -48 130 592
use scs8hd_fill_2  FILLER_347_59
timestamp 1586364061
transform 1 0 6532 0 1 190944
box -38 -48 222 592
use scs8hd_decap_12  FILLER_347_62
timestamp 1586364061
transform 1 0 6808 0 1 190944
box -38 -48 1142 592
use scs8hd_decap_3  PHY_695
timestamp 1586364061
transform -1 0 8832 0 1 190944
box -38 -48 314 592
use scs8hd_decap_6  FILLER_347_74
timestamp 1586364061
transform 1 0 7912 0 1 190944
box -38 -48 590 592
use scs8hd_fill_1  FILLER_347_80
timestamp 1586364061
transform 1 0 8464 0 1 190944
box -38 -48 130 592
use scs8hd_decap_3  PHY_696
timestamp 1586364061
transform 1 0 1104 0 -1 192032
box -38 -48 314 592
use scs8hd_decap_12  FILLER_348_3
timestamp 1586364061
transform 1 0 1380 0 -1 192032
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_348_15
timestamp 1586364061
transform 1 0 2484 0 -1 192032
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1557
timestamp 1586364061
transform 1 0 3956 0 -1 192032
box -38 -48 130 592
use scs8hd_decap_4  FILLER_348_27
timestamp 1586364061
transform 1 0 3588 0 -1 192032
box -38 -48 406 592
use scs8hd_decap_12  FILLER_348_32
timestamp 1586364061
transform 1 0 4048 0 -1 192032
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_348_44
timestamp 1586364061
transform 1 0 5152 0 -1 192032
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_348_56
timestamp 1586364061
transform 1 0 6256 0 -1 192032
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_348_68
timestamp 1586364061
transform 1 0 7360 0 -1 192032
box -38 -48 1142 592
use scs8hd_decap_3  PHY_697
timestamp 1586364061
transform -1 0 8832 0 -1 192032
box -38 -48 314 592
use scs8hd_fill_1  FILLER_348_80
timestamp 1586364061
transform 1 0 8464 0 -1 192032
box -38 -48 130 592
use scs8hd_decap_3  PHY_698
timestamp 1586364061
transform 1 0 1104 0 1 192032
box -38 -48 314 592
use scs8hd_decap_12  FILLER_349_3
timestamp 1586364061
transform 1 0 1380 0 1 192032
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_349_15
timestamp 1586364061
transform 1 0 2484 0 1 192032
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_349_27
timestamp 1586364061
transform 1 0 3588 0 1 192032
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_349_39
timestamp 1586364061
transform 1 0 4692 0 1 192032
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_349_51
timestamp 1586364061
transform 1 0 5796 0 1 192032
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1558
timestamp 1586364061
transform 1 0 6716 0 1 192032
box -38 -48 130 592
use scs8hd_fill_2  FILLER_349_59
timestamp 1586364061
transform 1 0 6532 0 1 192032
box -38 -48 222 592
use scs8hd_decap_12  FILLER_349_62
timestamp 1586364061
transform 1 0 6808 0 1 192032
box -38 -48 1142 592
use scs8hd_decap_3  PHY_699
timestamp 1586364061
transform -1 0 8832 0 1 192032
box -38 -48 314 592
use scs8hd_decap_6  FILLER_349_74
timestamp 1586364061
transform 1 0 7912 0 1 192032
box -38 -48 590 592
use scs8hd_fill_1  FILLER_349_80
timestamp 1586364061
transform 1 0 8464 0 1 192032
box -38 -48 130 592
use scs8hd_decap_3  PHY_700
timestamp 1586364061
transform 1 0 1104 0 -1 193120
box -38 -48 314 592
use scs8hd_decap_3  PHY_702
timestamp 1586364061
transform 1 0 1104 0 1 193120
box -38 -48 314 592
use scs8hd_decap_12  FILLER_350_3
timestamp 1586364061
transform 1 0 1380 0 -1 193120
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_350_15
timestamp 1586364061
transform 1 0 2484 0 -1 193120
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_351_3
timestamp 1586364061
transform 1 0 1380 0 1 193120
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_351_15
timestamp 1586364061
transform 1 0 2484 0 1 193120
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1559
timestamp 1586364061
transform 1 0 3956 0 -1 193120
box -38 -48 130 592
use scs8hd_decap_4  FILLER_350_27
timestamp 1586364061
transform 1 0 3588 0 -1 193120
box -38 -48 406 592
use scs8hd_decap_12  FILLER_350_32
timestamp 1586364061
transform 1 0 4048 0 -1 193120
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_351_27
timestamp 1586364061
transform 1 0 3588 0 1 193120
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_350_44
timestamp 1586364061
transform 1 0 5152 0 -1 193120
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_351_39
timestamp 1586364061
transform 1 0 4692 0 1 193120
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_351_51
timestamp 1586364061
transform 1 0 5796 0 1 193120
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1560
timestamp 1586364061
transform 1 0 6716 0 1 193120
box -38 -48 130 592
use scs8hd_decap_12  FILLER_350_56
timestamp 1586364061
transform 1 0 6256 0 -1 193120
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_350_68
timestamp 1586364061
transform 1 0 7360 0 -1 193120
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_351_59
timestamp 1586364061
transform 1 0 6532 0 1 193120
box -38 -48 222 592
use scs8hd_decap_12  FILLER_351_62
timestamp 1586364061
transform 1 0 6808 0 1 193120
box -38 -48 1142 592
use scs8hd_decap_3  PHY_701
timestamp 1586364061
transform -1 0 8832 0 -1 193120
box -38 -48 314 592
use scs8hd_decap_3  PHY_703
timestamp 1586364061
transform -1 0 8832 0 1 193120
box -38 -48 314 592
use scs8hd_fill_1  FILLER_350_80
timestamp 1586364061
transform 1 0 8464 0 -1 193120
box -38 -48 130 592
use scs8hd_decap_6  FILLER_351_74
timestamp 1586364061
transform 1 0 7912 0 1 193120
box -38 -48 590 592
use scs8hd_fill_1  FILLER_351_80
timestamp 1586364061
transform 1 0 8464 0 1 193120
box -38 -48 130 592
use scs8hd_decap_3  PHY_704
timestamp 1586364061
transform 1 0 1104 0 -1 194208
box -38 -48 314 592
use scs8hd_decap_12  FILLER_352_3
timestamp 1586364061
transform 1 0 1380 0 -1 194208
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_352_15
timestamp 1586364061
transform 1 0 2484 0 -1 194208
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1561
timestamp 1586364061
transform 1 0 3956 0 -1 194208
box -38 -48 130 592
use scs8hd_decap_4  FILLER_352_27
timestamp 1586364061
transform 1 0 3588 0 -1 194208
box -38 -48 406 592
use scs8hd_decap_12  FILLER_352_32
timestamp 1586364061
transform 1 0 4048 0 -1 194208
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_352_44
timestamp 1586364061
transform 1 0 5152 0 -1 194208
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_352_56
timestamp 1586364061
transform 1 0 6256 0 -1 194208
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_352_68
timestamp 1586364061
transform 1 0 7360 0 -1 194208
box -38 -48 1142 592
use scs8hd_decap_3  PHY_705
timestamp 1586364061
transform -1 0 8832 0 -1 194208
box -38 -48 314 592
use scs8hd_fill_1  FILLER_352_80
timestamp 1586364061
transform 1 0 8464 0 -1 194208
box -38 -48 130 592
use scs8hd_decap_3  PHY_706
timestamp 1586364061
transform 1 0 1104 0 1 194208
box -38 -48 314 592
use scs8hd_decap_12  FILLER_353_3
timestamp 1586364061
transform 1 0 1380 0 1 194208
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_353_15
timestamp 1586364061
transform 1 0 2484 0 1 194208
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_353_27
timestamp 1586364061
transform 1 0 3588 0 1 194208
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_353_39
timestamp 1586364061
transform 1 0 4692 0 1 194208
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_353_51
timestamp 1586364061
transform 1 0 5796 0 1 194208
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1562
timestamp 1586364061
transform 1 0 6716 0 1 194208
box -38 -48 130 592
use scs8hd_fill_2  FILLER_353_59
timestamp 1586364061
transform 1 0 6532 0 1 194208
box -38 -48 222 592
use scs8hd_decap_12  FILLER_353_62
timestamp 1586364061
transform 1 0 6808 0 1 194208
box -38 -48 1142 592
use scs8hd_decap_3  PHY_707
timestamp 1586364061
transform -1 0 8832 0 1 194208
box -38 -48 314 592
use scs8hd_decap_6  FILLER_353_74
timestamp 1586364061
transform 1 0 7912 0 1 194208
box -38 -48 590 592
use scs8hd_fill_1  FILLER_353_80
timestamp 1586364061
transform 1 0 8464 0 1 194208
box -38 -48 130 592
use scs8hd_decap_3  PHY_708
timestamp 1586364061
transform 1 0 1104 0 -1 195296
box -38 -48 314 592
use scs8hd_decap_12  FILLER_354_3
timestamp 1586364061
transform 1 0 1380 0 -1 195296
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_354_15
timestamp 1586364061
transform 1 0 2484 0 -1 195296
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1563
timestamp 1586364061
transform 1 0 3956 0 -1 195296
box -38 -48 130 592
use scs8hd_decap_4  FILLER_354_27
timestamp 1586364061
transform 1 0 3588 0 -1 195296
box -38 -48 406 592
use scs8hd_decap_12  FILLER_354_32
timestamp 1586364061
transform 1 0 4048 0 -1 195296
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_354_44
timestamp 1586364061
transform 1 0 5152 0 -1 195296
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_354_56
timestamp 1586364061
transform 1 0 6256 0 -1 195296
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_354_68
timestamp 1586364061
transform 1 0 7360 0 -1 195296
box -38 -48 1142 592
use scs8hd_decap_3  PHY_709
timestamp 1586364061
transform -1 0 8832 0 -1 195296
box -38 -48 314 592
use scs8hd_fill_1  FILLER_354_80
timestamp 1586364061
transform 1 0 8464 0 -1 195296
box -38 -48 130 592
use scs8hd_decap_3  PHY_710
timestamp 1586364061
transform 1 0 1104 0 1 195296
box -38 -48 314 592
use scs8hd_decap_12  FILLER_355_3
timestamp 1586364061
transform 1 0 1380 0 1 195296
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_355_15
timestamp 1586364061
transform 1 0 2484 0 1 195296
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_355_27
timestamp 1586364061
transform 1 0 3588 0 1 195296
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_355_39
timestamp 1586364061
transform 1 0 4692 0 1 195296
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_355_51
timestamp 1586364061
transform 1 0 5796 0 1 195296
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1564
timestamp 1586364061
transform 1 0 6716 0 1 195296
box -38 -48 130 592
use scs8hd_fill_2  FILLER_355_59
timestamp 1586364061
transform 1 0 6532 0 1 195296
box -38 -48 222 592
use scs8hd_decap_12  FILLER_355_62
timestamp 1586364061
transform 1 0 6808 0 1 195296
box -38 -48 1142 592
use scs8hd_decap_3  PHY_711
timestamp 1586364061
transform -1 0 8832 0 1 195296
box -38 -48 314 592
use scs8hd_decap_6  FILLER_355_74
timestamp 1586364061
transform 1 0 7912 0 1 195296
box -38 -48 590 592
use scs8hd_fill_1  FILLER_355_80
timestamp 1586364061
transform 1 0 8464 0 1 195296
box -38 -48 130 592
use scs8hd_decap_3  PHY_712
timestamp 1586364061
transform 1 0 1104 0 -1 196384
box -38 -48 314 592
use scs8hd_decap_3  PHY_714
timestamp 1586364061
transform 1 0 1104 0 1 196384
box -38 -48 314 592
use scs8hd_decap_12  FILLER_356_3
timestamp 1586364061
transform 1 0 1380 0 -1 196384
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_356_15
timestamp 1586364061
transform 1 0 2484 0 -1 196384
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_357_3
timestamp 1586364061
transform 1 0 1380 0 1 196384
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_357_15
timestamp 1586364061
transform 1 0 2484 0 1 196384
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1565
timestamp 1586364061
transform 1 0 3956 0 -1 196384
box -38 -48 130 592
use scs8hd_decap_4  FILLER_356_27
timestamp 1586364061
transform 1 0 3588 0 -1 196384
box -38 -48 406 592
use scs8hd_decap_12  FILLER_356_32
timestamp 1586364061
transform 1 0 4048 0 -1 196384
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_357_27
timestamp 1586364061
transform 1 0 3588 0 1 196384
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_356_44
timestamp 1586364061
transform 1 0 5152 0 -1 196384
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_357_39
timestamp 1586364061
transform 1 0 4692 0 1 196384
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_357_51
timestamp 1586364061
transform 1 0 5796 0 1 196384
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1566
timestamp 1586364061
transform 1 0 6716 0 1 196384
box -38 -48 130 592
use scs8hd_decap_12  FILLER_356_56
timestamp 1586364061
transform 1 0 6256 0 -1 196384
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_356_68
timestamp 1586364061
transform 1 0 7360 0 -1 196384
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_357_59
timestamp 1586364061
transform 1 0 6532 0 1 196384
box -38 -48 222 592
use scs8hd_decap_12  FILLER_357_62
timestamp 1586364061
transform 1 0 6808 0 1 196384
box -38 -48 1142 592
use scs8hd_decap_3  PHY_713
timestamp 1586364061
transform -1 0 8832 0 -1 196384
box -38 -48 314 592
use scs8hd_decap_3  PHY_715
timestamp 1586364061
transform -1 0 8832 0 1 196384
box -38 -48 314 592
use scs8hd_fill_1  FILLER_356_80
timestamp 1586364061
transform 1 0 8464 0 -1 196384
box -38 -48 130 592
use scs8hd_decap_6  FILLER_357_74
timestamp 1586364061
transform 1 0 7912 0 1 196384
box -38 -48 590 592
use scs8hd_fill_1  FILLER_357_80
timestamp 1586364061
transform 1 0 8464 0 1 196384
box -38 -48 130 592
use scs8hd_decap_3  PHY_716
timestamp 1586364061
transform 1 0 1104 0 -1 197472
box -38 -48 314 592
use scs8hd_decap_12  FILLER_358_3
timestamp 1586364061
transform 1 0 1380 0 -1 197472
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_358_15
timestamp 1586364061
transform 1 0 2484 0 -1 197472
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1567
timestamp 1586364061
transform 1 0 3956 0 -1 197472
box -38 -48 130 592
use scs8hd_decap_4  FILLER_358_27
timestamp 1586364061
transform 1 0 3588 0 -1 197472
box -38 -48 406 592
use scs8hd_decap_12  FILLER_358_32
timestamp 1586364061
transform 1 0 4048 0 -1 197472
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_358_44
timestamp 1586364061
transform 1 0 5152 0 -1 197472
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_358_56
timestamp 1586364061
transform 1 0 6256 0 -1 197472
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_358_68
timestamp 1586364061
transform 1 0 7360 0 -1 197472
box -38 -48 1142 592
use scs8hd_decap_3  PHY_717
timestamp 1586364061
transform -1 0 8832 0 -1 197472
box -38 -48 314 592
use scs8hd_fill_1  FILLER_358_80
timestamp 1586364061
transform 1 0 8464 0 -1 197472
box -38 -48 130 592
use scs8hd_decap_3  PHY_718
timestamp 1586364061
transform 1 0 1104 0 1 197472
box -38 -48 314 592
use scs8hd_decap_12  FILLER_359_3
timestamp 1586364061
transform 1 0 1380 0 1 197472
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_359_15
timestamp 1586364061
transform 1 0 2484 0 1 197472
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_359_27
timestamp 1586364061
transform 1 0 3588 0 1 197472
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_359_39
timestamp 1586364061
transform 1 0 4692 0 1 197472
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_359_51
timestamp 1586364061
transform 1 0 5796 0 1 197472
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1568
timestamp 1586364061
transform 1 0 6716 0 1 197472
box -38 -48 130 592
use scs8hd_fill_2  FILLER_359_59
timestamp 1586364061
transform 1 0 6532 0 1 197472
box -38 -48 222 592
use scs8hd_decap_12  FILLER_359_62
timestamp 1586364061
transform 1 0 6808 0 1 197472
box -38 -48 1142 592
use scs8hd_decap_3  PHY_719
timestamp 1586364061
transform -1 0 8832 0 1 197472
box -38 -48 314 592
use scs8hd_decap_6  FILLER_359_74
timestamp 1586364061
transform 1 0 7912 0 1 197472
box -38 -48 590 592
use scs8hd_fill_1  FILLER_359_80
timestamp 1586364061
transform 1 0 8464 0 1 197472
box -38 -48 130 592
use scs8hd_decap_3  PHY_720
timestamp 1586364061
transform 1 0 1104 0 -1 198560
box -38 -48 314 592
use scs8hd_decap_12  FILLER_360_3
timestamp 1586364061
transform 1 0 1380 0 -1 198560
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_360_15
timestamp 1586364061
transform 1 0 2484 0 -1 198560
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1569
timestamp 1586364061
transform 1 0 3956 0 -1 198560
box -38 -48 130 592
use scs8hd_decap_4  FILLER_360_27
timestamp 1586364061
transform 1 0 3588 0 -1 198560
box -38 -48 406 592
use scs8hd_decap_12  FILLER_360_32
timestamp 1586364061
transform 1 0 4048 0 -1 198560
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_360_44
timestamp 1586364061
transform 1 0 5152 0 -1 198560
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_360_56
timestamp 1586364061
transform 1 0 6256 0 -1 198560
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_360_68
timestamp 1586364061
transform 1 0 7360 0 -1 198560
box -38 -48 1142 592
use scs8hd_decap_3  PHY_721
timestamp 1586364061
transform -1 0 8832 0 -1 198560
box -38 -48 314 592
use scs8hd_fill_1  FILLER_360_80
timestamp 1586364061
transform 1 0 8464 0 -1 198560
box -38 -48 130 592
use scs8hd_decap_3  PHY_722
timestamp 1586364061
transform 1 0 1104 0 1 198560
box -38 -48 314 592
use scs8hd_decap_12  FILLER_361_3
timestamp 1586364061
transform 1 0 1380 0 1 198560
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_361_15
timestamp 1586364061
transform 1 0 2484 0 1 198560
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_361_27
timestamp 1586364061
transform 1 0 3588 0 1 198560
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_361_39
timestamp 1586364061
transform 1 0 4692 0 1 198560
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_361_51
timestamp 1586364061
transform 1 0 5796 0 1 198560
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1570
timestamp 1586364061
transform 1 0 6716 0 1 198560
box -38 -48 130 592
use scs8hd_fill_2  FILLER_361_59
timestamp 1586364061
transform 1 0 6532 0 1 198560
box -38 -48 222 592
use scs8hd_decap_12  FILLER_361_62
timestamp 1586364061
transform 1 0 6808 0 1 198560
box -38 -48 1142 592
use scs8hd_decap_3  PHY_723
timestamp 1586364061
transform -1 0 8832 0 1 198560
box -38 -48 314 592
use scs8hd_decap_6  FILLER_361_74
timestamp 1586364061
transform 1 0 7912 0 1 198560
box -38 -48 590 592
use scs8hd_fill_1  FILLER_361_80
timestamp 1586364061
transform 1 0 8464 0 1 198560
box -38 -48 130 592
use scs8hd_decap_3  PHY_724
timestamp 1586364061
transform 1 0 1104 0 -1 199648
box -38 -48 314 592
use scs8hd_decap_12  FILLER_362_3
timestamp 1586364061
transform 1 0 1380 0 -1 199648
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_362_15
timestamp 1586364061
transform 1 0 2484 0 -1 199648
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1571
timestamp 1586364061
transform 1 0 3956 0 -1 199648
box -38 -48 130 592
use scs8hd_decap_4  FILLER_362_27
timestamp 1586364061
transform 1 0 3588 0 -1 199648
box -38 -48 406 592
use scs8hd_decap_12  FILLER_362_32
timestamp 1586364061
transform 1 0 4048 0 -1 199648
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_362_44
timestamp 1586364061
transform 1 0 5152 0 -1 199648
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_362_56
timestamp 1586364061
transform 1 0 6256 0 -1 199648
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_362_68
timestamp 1586364061
transform 1 0 7360 0 -1 199648
box -38 -48 1142 592
use scs8hd_decap_3  PHY_725
timestamp 1586364061
transform -1 0 8832 0 -1 199648
box -38 -48 314 592
use scs8hd_fill_1  FILLER_362_80
timestamp 1586364061
transform 1 0 8464 0 -1 199648
box -38 -48 130 592
use scs8hd_decap_3  PHY_726
timestamp 1586364061
transform 1 0 1104 0 1 199648
box -38 -48 314 592
use scs8hd_decap_3  PHY_728
timestamp 1586364061
transform 1 0 1104 0 -1 200736
box -38 -48 314 592
use scs8hd_decap_12  FILLER_363_3
timestamp 1586364061
transform 1 0 1380 0 1 199648
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_363_15
timestamp 1586364061
transform 1 0 2484 0 1 199648
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_364_3
timestamp 1586364061
transform 1 0 1380 0 -1 200736
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_364_15
timestamp 1586364061
transform 1 0 2484 0 -1 200736
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1573
timestamp 1586364061
transform 1 0 3956 0 -1 200736
box -38 -48 130 592
use scs8hd_decap_12  FILLER_363_27
timestamp 1586364061
transform 1 0 3588 0 1 199648
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_364_27
timestamp 1586364061
transform 1 0 3588 0 -1 200736
box -38 -48 406 592
use scs8hd_decap_12  FILLER_364_32
timestamp 1586364061
transform 1 0 4048 0 -1 200736
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_363_39
timestamp 1586364061
transform 1 0 4692 0 1 199648
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_363_51
timestamp 1586364061
transform 1 0 5796 0 1 199648
box -38 -48 774 592
use scs8hd_decap_12  FILLER_364_44
timestamp 1586364061
transform 1 0 5152 0 -1 200736
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1572
timestamp 1586364061
transform 1 0 6716 0 1 199648
box -38 -48 130 592
use scs8hd_fill_2  FILLER_363_59
timestamp 1586364061
transform 1 0 6532 0 1 199648
box -38 -48 222 592
use scs8hd_decap_12  FILLER_363_62
timestamp 1586364061
transform 1 0 6808 0 1 199648
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_364_56
timestamp 1586364061
transform 1 0 6256 0 -1 200736
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_364_68
timestamp 1586364061
transform 1 0 7360 0 -1 200736
box -38 -48 1142 592
use scs8hd_decap_3  PHY_727
timestamp 1586364061
transform -1 0 8832 0 1 199648
box -38 -48 314 592
use scs8hd_decap_3  PHY_729
timestamp 1586364061
transform -1 0 8832 0 -1 200736
box -38 -48 314 592
use scs8hd_decap_6  FILLER_363_74
timestamp 1586364061
transform 1 0 7912 0 1 199648
box -38 -48 590 592
use scs8hd_fill_1  FILLER_363_80
timestamp 1586364061
transform 1 0 8464 0 1 199648
box -38 -48 130 592
use scs8hd_fill_1  FILLER_364_80
timestamp 1586364061
transform 1 0 8464 0 -1 200736
box -38 -48 130 592
use scs8hd_decap_3  PHY_730
timestamp 1586364061
transform 1 0 1104 0 1 200736
box -38 -48 314 592
use scs8hd_decap_12  FILLER_365_3
timestamp 1586364061
transform 1 0 1380 0 1 200736
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_365_15
timestamp 1586364061
transform 1 0 2484 0 1 200736
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_365_27
timestamp 1586364061
transform 1 0 3588 0 1 200736
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_365_39
timestamp 1586364061
transform 1 0 4692 0 1 200736
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_365_51
timestamp 1586364061
transform 1 0 5796 0 1 200736
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1574
timestamp 1586364061
transform 1 0 6716 0 1 200736
box -38 -48 130 592
use scs8hd_fill_2  FILLER_365_59
timestamp 1586364061
transform 1 0 6532 0 1 200736
box -38 -48 222 592
use scs8hd_decap_12  FILLER_365_62
timestamp 1586364061
transform 1 0 6808 0 1 200736
box -38 -48 1142 592
use scs8hd_decap_3  PHY_731
timestamp 1586364061
transform -1 0 8832 0 1 200736
box -38 -48 314 592
use scs8hd_decap_6  FILLER_365_74
timestamp 1586364061
transform 1 0 7912 0 1 200736
box -38 -48 590 592
use scs8hd_fill_1  FILLER_365_80
timestamp 1586364061
transform 1 0 8464 0 1 200736
box -38 -48 130 592
use scs8hd_decap_3  PHY_732
timestamp 1586364061
transform 1 0 1104 0 -1 201824
box -38 -48 314 592
use scs8hd_decap_12  FILLER_366_3
timestamp 1586364061
transform 1 0 1380 0 -1 201824
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_366_15
timestamp 1586364061
transform 1 0 2484 0 -1 201824
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1575
timestamp 1586364061
transform 1 0 3956 0 -1 201824
box -38 -48 130 592
use scs8hd_decap_4  FILLER_366_27
timestamp 1586364061
transform 1 0 3588 0 -1 201824
box -38 -48 406 592
use scs8hd_decap_12  FILLER_366_32
timestamp 1586364061
transform 1 0 4048 0 -1 201824
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_366_44
timestamp 1586364061
transform 1 0 5152 0 -1 201824
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_366_56
timestamp 1586364061
transform 1 0 6256 0 -1 201824
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_366_68
timestamp 1586364061
transform 1 0 7360 0 -1 201824
box -38 -48 1142 592
use scs8hd_decap_3  PHY_733
timestamp 1586364061
transform -1 0 8832 0 -1 201824
box -38 -48 314 592
use scs8hd_fill_1  FILLER_366_80
timestamp 1586364061
transform 1 0 8464 0 -1 201824
box -38 -48 130 592
use scs8hd_decap_3  PHY_734
timestamp 1586364061
transform 1 0 1104 0 1 201824
box -38 -48 314 592
use scs8hd_decap_12  FILLER_367_3
timestamp 1586364061
transform 1 0 1380 0 1 201824
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_367_15
timestamp 1586364061
transform 1 0 2484 0 1 201824
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_367_27
timestamp 1586364061
transform 1 0 3588 0 1 201824
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_367_39
timestamp 1586364061
transform 1 0 4692 0 1 201824
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_367_51
timestamp 1586364061
transform 1 0 5796 0 1 201824
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1576
timestamp 1586364061
transform 1 0 6716 0 1 201824
box -38 -48 130 592
use scs8hd_fill_2  FILLER_367_59
timestamp 1586364061
transform 1 0 6532 0 1 201824
box -38 -48 222 592
use scs8hd_decap_12  FILLER_367_62
timestamp 1586364061
transform 1 0 6808 0 1 201824
box -38 -48 1142 592
use scs8hd_decap_3  PHY_735
timestamp 1586364061
transform -1 0 8832 0 1 201824
box -38 -48 314 592
use scs8hd_decap_6  FILLER_367_74
timestamp 1586364061
transform 1 0 7912 0 1 201824
box -38 -48 590 592
use scs8hd_fill_1  FILLER_367_80
timestamp 1586364061
transform 1 0 8464 0 1 201824
box -38 -48 130 592
use scs8hd_decap_3  PHY_736
timestamp 1586364061
transform 1 0 1104 0 -1 202912
box -38 -48 314 592
use scs8hd_decap_12  FILLER_368_3
timestamp 1586364061
transform 1 0 1380 0 -1 202912
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_368_15
timestamp 1586364061
transform 1 0 2484 0 -1 202912
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1577
timestamp 1586364061
transform 1 0 3956 0 -1 202912
box -38 -48 130 592
use scs8hd_decap_4  FILLER_368_27
timestamp 1586364061
transform 1 0 3588 0 -1 202912
box -38 -48 406 592
use scs8hd_decap_12  FILLER_368_32
timestamp 1586364061
transform 1 0 4048 0 -1 202912
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_368_44
timestamp 1586364061
transform 1 0 5152 0 -1 202912
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_368_56
timestamp 1586364061
transform 1 0 6256 0 -1 202912
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_368_68
timestamp 1586364061
transform 1 0 7360 0 -1 202912
box -38 -48 1142 592
use scs8hd_decap_3  PHY_737
timestamp 1586364061
transform -1 0 8832 0 -1 202912
box -38 -48 314 592
use scs8hd_fill_1  FILLER_368_80
timestamp 1586364061
transform 1 0 8464 0 -1 202912
box -38 -48 130 592
use scs8hd_decap_3  PHY_738
timestamp 1586364061
transform 1 0 1104 0 1 202912
box -38 -48 314 592
use scs8hd_decap_12  FILLER_369_3
timestamp 1586364061
transform 1 0 1380 0 1 202912
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_369_15
timestamp 1586364061
transform 1 0 2484 0 1 202912
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_369_27
timestamp 1586364061
transform 1 0 3588 0 1 202912
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_369_39
timestamp 1586364061
transform 1 0 4692 0 1 202912
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_369_51
timestamp 1586364061
transform 1 0 5796 0 1 202912
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1578
timestamp 1586364061
transform 1 0 6716 0 1 202912
box -38 -48 130 592
use scs8hd_fill_2  FILLER_369_59
timestamp 1586364061
transform 1 0 6532 0 1 202912
box -38 -48 222 592
use scs8hd_decap_12  FILLER_369_62
timestamp 1586364061
transform 1 0 6808 0 1 202912
box -38 -48 1142 592
use scs8hd_decap_3  PHY_739
timestamp 1586364061
transform -1 0 8832 0 1 202912
box -38 -48 314 592
use scs8hd_decap_6  FILLER_369_74
timestamp 1586364061
transform 1 0 7912 0 1 202912
box -38 -48 590 592
use scs8hd_fill_1  FILLER_369_80
timestamp 1586364061
transform 1 0 8464 0 1 202912
box -38 -48 130 592
use scs8hd_decap_3  PHY_740
timestamp 1586364061
transform 1 0 1104 0 -1 204000
box -38 -48 314 592
use scs8hd_decap_3  PHY_742
timestamp 1586364061
transform 1 0 1104 0 1 204000
box -38 -48 314 592
use scs8hd_decap_12  FILLER_370_3
timestamp 1586364061
transform 1 0 1380 0 -1 204000
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_370_15
timestamp 1586364061
transform 1 0 2484 0 -1 204000
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_371_3
timestamp 1586364061
transform 1 0 1380 0 1 204000
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_371_15
timestamp 1586364061
transform 1 0 2484 0 1 204000
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1579
timestamp 1586364061
transform 1 0 3956 0 -1 204000
box -38 -48 130 592
use scs8hd_decap_4  FILLER_370_27
timestamp 1586364061
transform 1 0 3588 0 -1 204000
box -38 -48 406 592
use scs8hd_decap_12  FILLER_370_32
timestamp 1586364061
transform 1 0 4048 0 -1 204000
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_371_27
timestamp 1586364061
transform 1 0 3588 0 1 204000
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_370_44
timestamp 1586364061
transform 1 0 5152 0 -1 204000
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_371_39
timestamp 1586364061
transform 1 0 4692 0 1 204000
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_371_51
timestamp 1586364061
transform 1 0 5796 0 1 204000
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1580
timestamp 1586364061
transform 1 0 6716 0 1 204000
box -38 -48 130 592
use scs8hd_decap_12  FILLER_370_56
timestamp 1586364061
transform 1 0 6256 0 -1 204000
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_370_68
timestamp 1586364061
transform 1 0 7360 0 -1 204000
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_371_59
timestamp 1586364061
transform 1 0 6532 0 1 204000
box -38 -48 222 592
use scs8hd_decap_12  FILLER_371_62
timestamp 1586364061
transform 1 0 6808 0 1 204000
box -38 -48 1142 592
use scs8hd_decap_3  PHY_741
timestamp 1586364061
transform -1 0 8832 0 -1 204000
box -38 -48 314 592
use scs8hd_decap_3  PHY_743
timestamp 1586364061
transform -1 0 8832 0 1 204000
box -38 -48 314 592
use scs8hd_fill_1  FILLER_370_80
timestamp 1586364061
transform 1 0 8464 0 -1 204000
box -38 -48 130 592
use scs8hd_decap_6  FILLER_371_74
timestamp 1586364061
transform 1 0 7912 0 1 204000
box -38 -48 590 592
use scs8hd_fill_1  FILLER_371_80
timestamp 1586364061
transform 1 0 8464 0 1 204000
box -38 -48 130 592
use scs8hd_decap_3  PHY_744
timestamp 1586364061
transform 1 0 1104 0 -1 205088
box -38 -48 314 592
use scs8hd_decap_12  FILLER_372_3
timestamp 1586364061
transform 1 0 1380 0 -1 205088
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_372_15
timestamp 1586364061
transform 1 0 2484 0 -1 205088
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1581
timestamp 1586364061
transform 1 0 3956 0 -1 205088
box -38 -48 130 592
use scs8hd_decap_4  FILLER_372_27
timestamp 1586364061
transform 1 0 3588 0 -1 205088
box -38 -48 406 592
use scs8hd_decap_12  FILLER_372_32
timestamp 1586364061
transform 1 0 4048 0 -1 205088
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_372_44
timestamp 1586364061
transform 1 0 5152 0 -1 205088
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_372_56
timestamp 1586364061
transform 1 0 6256 0 -1 205088
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_372_68
timestamp 1586364061
transform 1 0 7360 0 -1 205088
box -38 -48 1142 592
use scs8hd_decap_3  PHY_745
timestamp 1586364061
transform -1 0 8832 0 -1 205088
box -38 -48 314 592
use scs8hd_fill_1  FILLER_372_80
timestamp 1586364061
transform 1 0 8464 0 -1 205088
box -38 -48 130 592
use scs8hd_decap_3  PHY_746
timestamp 1586364061
transform 1 0 1104 0 1 205088
box -38 -48 314 592
use scs8hd_decap_12  FILLER_373_3
timestamp 1586364061
transform 1 0 1380 0 1 205088
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_373_15
timestamp 1586364061
transform 1 0 2484 0 1 205088
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_373_27
timestamp 1586364061
transform 1 0 3588 0 1 205088
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_373_39
timestamp 1586364061
transform 1 0 4692 0 1 205088
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_373_51
timestamp 1586364061
transform 1 0 5796 0 1 205088
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1582
timestamp 1586364061
transform 1 0 6716 0 1 205088
box -38 -48 130 592
use scs8hd_fill_2  FILLER_373_59
timestamp 1586364061
transform 1 0 6532 0 1 205088
box -38 -48 222 592
use scs8hd_decap_12  FILLER_373_62
timestamp 1586364061
transform 1 0 6808 0 1 205088
box -38 -48 1142 592
use scs8hd_decap_3  PHY_747
timestamp 1586364061
transform -1 0 8832 0 1 205088
box -38 -48 314 592
use scs8hd_decap_6  FILLER_373_74
timestamp 1586364061
transform 1 0 7912 0 1 205088
box -38 -48 590 592
use scs8hd_fill_1  FILLER_373_80
timestamp 1586364061
transform 1 0 8464 0 1 205088
box -38 -48 130 592
use scs8hd_decap_3  PHY_748
timestamp 1586364061
transform 1 0 1104 0 -1 206176
box -38 -48 314 592
use scs8hd_decap_12  FILLER_374_3
timestamp 1586364061
transform 1 0 1380 0 -1 206176
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_374_15
timestamp 1586364061
transform 1 0 2484 0 -1 206176
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1583
timestamp 1586364061
transform 1 0 3956 0 -1 206176
box -38 -48 130 592
use scs8hd_decap_4  FILLER_374_27
timestamp 1586364061
transform 1 0 3588 0 -1 206176
box -38 -48 406 592
use scs8hd_decap_12  FILLER_374_32
timestamp 1586364061
transform 1 0 4048 0 -1 206176
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_374_44
timestamp 1586364061
transform 1 0 5152 0 -1 206176
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_374_56
timestamp 1586364061
transform 1 0 6256 0 -1 206176
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_374_68
timestamp 1586364061
transform 1 0 7360 0 -1 206176
box -38 -48 1142 592
use scs8hd_decap_3  PHY_749
timestamp 1586364061
transform -1 0 8832 0 -1 206176
box -38 -48 314 592
use scs8hd_fill_1  FILLER_374_80
timestamp 1586364061
transform 1 0 8464 0 -1 206176
box -38 -48 130 592
use scs8hd_decap_3  PHY_750
timestamp 1586364061
transform 1 0 1104 0 1 206176
box -38 -48 314 592
use scs8hd_decap_12  FILLER_375_3
timestamp 1586364061
transform 1 0 1380 0 1 206176
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_375_15
timestamp 1586364061
transform 1 0 2484 0 1 206176
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_375_27
timestamp 1586364061
transform 1 0 3588 0 1 206176
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_375_39
timestamp 1586364061
transform 1 0 4692 0 1 206176
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_375_51
timestamp 1586364061
transform 1 0 5796 0 1 206176
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1584
timestamp 1586364061
transform 1 0 6716 0 1 206176
box -38 -48 130 592
use scs8hd_fill_2  FILLER_375_59
timestamp 1586364061
transform 1 0 6532 0 1 206176
box -38 -48 222 592
use scs8hd_decap_12  FILLER_375_62
timestamp 1586364061
transform 1 0 6808 0 1 206176
box -38 -48 1142 592
use scs8hd_decap_3  PHY_751
timestamp 1586364061
transform -1 0 8832 0 1 206176
box -38 -48 314 592
use scs8hd_decap_6  FILLER_375_74
timestamp 1586364061
transform 1 0 7912 0 1 206176
box -38 -48 590 592
use scs8hd_fill_1  FILLER_375_80
timestamp 1586364061
transform 1 0 8464 0 1 206176
box -38 -48 130 592
use scs8hd_decap_3  PHY_752
timestamp 1586364061
transform 1 0 1104 0 -1 207264
box -38 -48 314 592
use scs8hd_decap_3  PHY_754
timestamp 1586364061
transform 1 0 1104 0 1 207264
box -38 -48 314 592
use scs8hd_decap_12  FILLER_376_3
timestamp 1586364061
transform 1 0 1380 0 -1 207264
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_376_15
timestamp 1586364061
transform 1 0 2484 0 -1 207264
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_377_3
timestamp 1586364061
transform 1 0 1380 0 1 207264
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_377_15
timestamp 1586364061
transform 1 0 2484 0 1 207264
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1585
timestamp 1586364061
transform 1 0 3956 0 -1 207264
box -38 -48 130 592
use scs8hd_decap_4  FILLER_376_27
timestamp 1586364061
transform 1 0 3588 0 -1 207264
box -38 -48 406 592
use scs8hd_decap_12  FILLER_376_32
timestamp 1586364061
transform 1 0 4048 0 -1 207264
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_377_27
timestamp 1586364061
transform 1 0 3588 0 1 207264
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_376_44
timestamp 1586364061
transform 1 0 5152 0 -1 207264
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_377_39
timestamp 1586364061
transform 1 0 4692 0 1 207264
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_377_51
timestamp 1586364061
transform 1 0 5796 0 1 207264
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1586
timestamp 1586364061
transform 1 0 6716 0 1 207264
box -38 -48 130 592
use scs8hd_decap_12  FILLER_376_56
timestamp 1586364061
transform 1 0 6256 0 -1 207264
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_376_68
timestamp 1586364061
transform 1 0 7360 0 -1 207264
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_377_59
timestamp 1586364061
transform 1 0 6532 0 1 207264
box -38 -48 222 592
use scs8hd_decap_12  FILLER_377_62
timestamp 1586364061
transform 1 0 6808 0 1 207264
box -38 -48 1142 592
use scs8hd_decap_3  PHY_753
timestamp 1586364061
transform -1 0 8832 0 -1 207264
box -38 -48 314 592
use scs8hd_decap_3  PHY_755
timestamp 1586364061
transform -1 0 8832 0 1 207264
box -38 -48 314 592
use scs8hd_fill_1  FILLER_376_80
timestamp 1586364061
transform 1 0 8464 0 -1 207264
box -38 -48 130 592
use scs8hd_decap_6  FILLER_377_74
timestamp 1586364061
transform 1 0 7912 0 1 207264
box -38 -48 590 592
use scs8hd_fill_1  FILLER_377_80
timestamp 1586364061
transform 1 0 8464 0 1 207264
box -38 -48 130 592
use scs8hd_decap_3  PHY_756
timestamp 1586364061
transform 1 0 1104 0 -1 208352
box -38 -48 314 592
use scs8hd_decap_12  FILLER_378_3
timestamp 1586364061
transform 1 0 1380 0 -1 208352
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_378_15
timestamp 1586364061
transform 1 0 2484 0 -1 208352
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_1587
timestamp 1586364061
transform 1 0 3956 0 -1 208352
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2760 0 -1 208352
box -38 -48 222 592
use scs8hd_decap_8  FILLER_378_20
timestamp 1586364061
transform 1 0 2944 0 -1 208352
box -38 -48 774 592
use scs8hd_decap_3  FILLER_378_28
timestamp 1586364061
transform 1 0 3680 0 -1 208352
box -38 -48 314 592
use scs8hd_decap_12  FILLER_378_32
timestamp 1586364061
transform 1 0 4048 0 -1 208352
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_378_44
timestamp 1586364061
transform 1 0 5152 0 -1 208352
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_378_56
timestamp 1586364061
transform 1 0 6256 0 -1 208352
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_378_68
timestamp 1586364061
transform 1 0 7360 0 -1 208352
box -38 -48 1142 592
use scs8hd_decap_3  PHY_757
timestamp 1586364061
transform -1 0 8832 0 -1 208352
box -38 -48 314 592
use scs8hd_fill_1  FILLER_378_80
timestamp 1586364061
transform 1 0 8464 0 -1 208352
box -38 -48 130 592
use scs8hd_decap_3  PHY_758
timestamp 1586364061
transform 1 0 1104 0 1 208352
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2576 0 1 208352
box -38 -48 222 592
use scs8hd_decap_12  FILLER_379_3
timestamp 1586364061
transform 1 0 1380 0 1 208352
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_379_15
timestamp 1586364061
transform 1 0 2484 0 1 208352
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2760 0 1 208352
box -38 -48 1050 592
use scs8hd_decap_12  FILLER_379_29
timestamp 1586364061
transform 1 0 3772 0 1 208352
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_379_41
timestamp 1586364061
transform 1 0 4876 0 1 208352
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_379_53
timestamp 1586364061
transform 1 0 5980 0 1 208352
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1588
timestamp 1586364061
transform 1 0 6716 0 1 208352
box -38 -48 130 592
use scs8hd_decap_12  FILLER_379_62
timestamp 1586364061
transform 1 0 6808 0 1 208352
box -38 -48 1142 592
use scs8hd_decap_3  PHY_759
timestamp 1586364061
transform -1 0 8832 0 1 208352
box -38 -48 314 592
use scs8hd_decap_6  FILLER_379_74
timestamp 1586364061
transform 1 0 7912 0 1 208352
box -38 -48 590 592
use scs8hd_fill_1  FILLER_379_80
timestamp 1586364061
transform 1 0 8464 0 1 208352
box -38 -48 130 592
use scs8hd_decap_3  PHY_760
timestamp 1586364061
transform 1 0 1104 0 -1 209440
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 2668 0 -1 209440
box -38 -48 222 592
use scs8hd_decap_12  FILLER_380_3
timestamp 1586364061
transform 1 0 1380 0 -1 209440
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_380_15
timestamp 1586364061
transform 1 0 2484 0 -1 209440
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_1589
timestamp 1586364061
transform 1 0 3956 0 -1 209440
box -38 -48 130 592
use scs8hd_decap_12  FILLER_380_19
timestamp 1586364061
transform 1 0 2852 0 -1 209440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_380_32
timestamp 1586364061
transform 1 0 4048 0 -1 209440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_380_44
timestamp 1586364061
transform 1 0 5152 0 -1 209440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_380_56
timestamp 1586364061
transform 1 0 6256 0 -1 209440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_380_68
timestamp 1586364061
transform 1 0 7360 0 -1 209440
box -38 -48 1142 592
use scs8hd_decap_3  PHY_761
timestamp 1586364061
transform -1 0 8832 0 -1 209440
box -38 -48 314 592
use scs8hd_fill_1  FILLER_380_80
timestamp 1586364061
transform 1 0 8464 0 -1 209440
box -38 -48 130 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2668 0 1 209440
box -38 -48 774 592
use scs8hd_decap_3  PHY_762
timestamp 1586364061
transform 1 0 1104 0 1 209440
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 2484 0 1 209440
box -38 -48 222 592
use scs8hd_decap_12  FILLER_381_3
timestamp 1586364061
transform 1 0 1380 0 1 209440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_381_25
timestamp 1586364061
transform 1 0 3404 0 1 209440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_381_37
timestamp 1586364061
transform 1 0 4508 0 1 209440
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_381_49
timestamp 1586364061
transform 1 0 5612 0 1 209440
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1590
timestamp 1586364061
transform 1 0 6716 0 1 209440
box -38 -48 130 592
use scs8hd_decap_12  FILLER_381_62
timestamp 1586364061
transform 1 0 6808 0 1 209440
box -38 -48 1142 592
use scs8hd_decap_3  PHY_763
timestamp 1586364061
transform -1 0 8832 0 1 209440
box -38 -48 314 592
use scs8hd_decap_6  FILLER_381_74
timestamp 1586364061
transform 1 0 7912 0 1 209440
box -38 -48 590 592
use scs8hd_fill_1  FILLER_381_80
timestamp 1586364061
transform 1 0 8464 0 1 209440
box -38 -48 130 592
use scs8hd_decap_3  PHY_764
timestamp 1586364061
transform 1 0 1104 0 -1 210528
box -38 -48 314 592
use scs8hd_decap_12  FILLER_382_3
timestamp 1586364061
transform 1 0 1380 0 -1 210528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_382_15
timestamp 1586364061
transform 1 0 2484 0 -1 210528
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1591
timestamp 1586364061
transform 1 0 3956 0 -1 210528
box -38 -48 130 592
use scs8hd_decap_4  FILLER_382_27
timestamp 1586364061
transform 1 0 3588 0 -1 210528
box -38 -48 406 592
use scs8hd_decap_12  FILLER_382_32
timestamp 1586364061
transform 1 0 4048 0 -1 210528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_382_44
timestamp 1586364061
transform 1 0 5152 0 -1 210528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_382_56
timestamp 1586364061
transform 1 0 6256 0 -1 210528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_382_68
timestamp 1586364061
transform 1 0 7360 0 -1 210528
box -38 -48 1142 592
use scs8hd_decap_3  PHY_765
timestamp 1586364061
transform -1 0 8832 0 -1 210528
box -38 -48 314 592
use scs8hd_fill_1  FILLER_382_80
timestamp 1586364061
transform 1 0 8464 0 -1 210528
box -38 -48 130 592
use scs8hd_decap_3  PHY_766
timestamp 1586364061
transform 1 0 1104 0 1 210528
box -38 -48 314 592
use scs8hd_decap_3  PHY_768
timestamp 1586364061
transform 1 0 1104 0 -1 211616
box -38 -48 314 592
use scs8hd_decap_12  FILLER_383_3
timestamp 1586364061
transform 1 0 1380 0 1 210528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_383_15
timestamp 1586364061
transform 1 0 2484 0 1 210528
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_384_3
timestamp 1586364061
transform 1 0 1380 0 -1 211616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_384_15
timestamp 1586364061
transform 1 0 2484 0 -1 211616
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1593
timestamp 1586364061
transform 1 0 3956 0 -1 211616
box -38 -48 130 592
use scs8hd_decap_12  FILLER_383_27
timestamp 1586364061
transform 1 0 3588 0 1 210528
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_384_27
timestamp 1586364061
transform 1 0 3588 0 -1 211616
box -38 -48 406 592
use scs8hd_decap_4  FILLER_384_32
timestamp 1586364061
transform 1 0 4048 0 -1 211616
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 4416 0 -1 211616
box -38 -48 222 592
use scs8hd_decap_12  FILLER_383_39
timestamp 1586364061
transform 1 0 4692 0 1 210528
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_383_51
timestamp 1586364061
transform 1 0 5796 0 1 210528
box -38 -48 774 592
use scs8hd_decap_12  FILLER_384_38
timestamp 1586364061
transform 1 0 4600 0 -1 211616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_384_50
timestamp 1586364061
transform 1 0 5704 0 -1 211616
box -38 -48 1142 592
use scs8hd_buf_2  _20_
timestamp 1586364061
transform 1 0 6808 0 1 210528
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_1592
timestamp 1586364061
transform 1 0 6716 0 1 210528
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__20__A
timestamp 1586364061
transform 1 0 7360 0 1 210528
box -38 -48 222 592
use scs8hd_fill_2  FILLER_383_59
timestamp 1586364061
transform 1 0 6532 0 1 210528
box -38 -48 222 592
use scs8hd_fill_2  FILLER_383_66
timestamp 1586364061
transform 1 0 7176 0 1 210528
box -38 -48 222 592
use scs8hd_decap_8  FILLER_383_70
timestamp 1586364061
transform 1 0 7544 0 1 210528
box -38 -48 774 592
use scs8hd_decap_12  FILLER_384_62
timestamp 1586364061
transform 1 0 6808 0 -1 211616
box -38 -48 1142 592
use scs8hd_decap_3  PHY_767
timestamp 1586364061
transform -1 0 8832 0 1 210528
box -38 -48 314 592
use scs8hd_decap_3  PHY_769
timestamp 1586364061
transform -1 0 8832 0 -1 211616
box -38 -48 314 592
use scs8hd_decap_3  FILLER_383_78
timestamp 1586364061
transform 1 0 8280 0 1 210528
box -38 -48 314 592
use scs8hd_decap_6  FILLER_384_74
timestamp 1586364061
transform 1 0 7912 0 -1 211616
box -38 -48 590 592
use scs8hd_fill_1  FILLER_384_80
timestamp 1586364061
transform 1 0 8464 0 -1 211616
box -38 -48 130 592
use scs8hd_decap_3  PHY_770
timestamp 1586364061
transform 1 0 1104 0 1 211616
box -38 -48 314 592
use scs8hd_decap_12  FILLER_385_3
timestamp 1586364061
transform 1 0 1380 0 1 211616
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_385_15
timestamp 1586364061
transform 1 0 2484 0 1 211616
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 4232 0 1 211616
box -38 -48 222 592
use scs8hd_decap_6  FILLER_385_27
timestamp 1586364061
transform 1 0 3588 0 1 211616
box -38 -48 590 592
use scs8hd_fill_1  FILLER_385_33
timestamp 1586364061
transform 1 0 4140 0 1 211616
box -38 -48 130 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 4416 0 1 211616
box -38 -48 774 592
use scs8hd_decap_12  FILLER_385_44
timestamp 1586364061
transform 1 0 5152 0 1 211616
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1594
timestamp 1586364061
transform 1 0 6716 0 1 211616
box -38 -48 130 592
use scs8hd_decap_4  FILLER_385_56
timestamp 1586364061
transform 1 0 6256 0 1 211616
box -38 -48 406 592
use scs8hd_fill_1  FILLER_385_60
timestamp 1586364061
transform 1 0 6624 0 1 211616
box -38 -48 130 592
use scs8hd_decap_12  FILLER_385_62
timestamp 1586364061
transform 1 0 6808 0 1 211616
box -38 -48 1142 592
use scs8hd_decap_3  PHY_771
timestamp 1586364061
transform -1 0 8832 0 1 211616
box -38 -48 314 592
use scs8hd_decap_6  FILLER_385_74
timestamp 1586364061
transform 1 0 7912 0 1 211616
box -38 -48 590 592
use scs8hd_fill_1  FILLER_385_80
timestamp 1586364061
transform 1 0 8464 0 1 211616
box -38 -48 130 592
use scs8hd_decap_3  PHY_772
timestamp 1586364061
transform 1 0 1104 0 -1 212704
box -38 -48 314 592
use scs8hd_decap_12  FILLER_386_3
timestamp 1586364061
transform 1 0 1380 0 -1 212704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_386_15
timestamp 1586364061
transform 1 0 2484 0 -1 212704
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1595
timestamp 1586364061
transform 1 0 3956 0 -1 212704
box -38 -48 130 592
use scs8hd_decap_4  FILLER_386_27
timestamp 1586364061
transform 1 0 3588 0 -1 212704
box -38 -48 406 592
use scs8hd_decap_12  FILLER_386_32
timestamp 1586364061
transform 1 0 4048 0 -1 212704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_386_44
timestamp 1586364061
transform 1 0 5152 0 -1 212704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_386_56
timestamp 1586364061
transform 1 0 6256 0 -1 212704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_386_68
timestamp 1586364061
transform 1 0 7360 0 -1 212704
box -38 -48 1142 592
use scs8hd_decap_3  PHY_773
timestamp 1586364061
transform -1 0 8832 0 -1 212704
box -38 -48 314 592
use scs8hd_fill_1  FILLER_386_80
timestamp 1586364061
transform 1 0 8464 0 -1 212704
box -38 -48 130 592
use scs8hd_decap_3  PHY_774
timestamp 1586364061
transform 1 0 1104 0 1 212704
box -38 -48 314 592
use scs8hd_decap_12  FILLER_387_3
timestamp 1586364061
transform 1 0 1380 0 1 212704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_387_15
timestamp 1586364061
transform 1 0 2484 0 1 212704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_387_27
timestamp 1586364061
transform 1 0 3588 0 1 212704
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_387_39
timestamp 1586364061
transform 1 0 4692 0 1 212704
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_387_51
timestamp 1586364061
transform 1 0 5796 0 1 212704
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1596
timestamp 1586364061
transform 1 0 6716 0 1 212704
box -38 -48 130 592
use scs8hd_fill_2  FILLER_387_59
timestamp 1586364061
transform 1 0 6532 0 1 212704
box -38 -48 222 592
use scs8hd_decap_12  FILLER_387_62
timestamp 1586364061
transform 1 0 6808 0 1 212704
box -38 -48 1142 592
use scs8hd_decap_3  PHY_775
timestamp 1586364061
transform -1 0 8832 0 1 212704
box -38 -48 314 592
use scs8hd_decap_6  FILLER_387_74
timestamp 1586364061
transform 1 0 7912 0 1 212704
box -38 -48 590 592
use scs8hd_fill_1  FILLER_387_80
timestamp 1586364061
transform 1 0 8464 0 1 212704
box -38 -48 130 592
use scs8hd_decap_3  PHY_776
timestamp 1586364061
transform 1 0 1104 0 -1 213792
box -38 -48 314 592
use scs8hd_decap_12  FILLER_388_3
timestamp 1586364061
transform 1 0 1380 0 -1 213792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_388_15
timestamp 1586364061
transform 1 0 2484 0 -1 213792
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1597
timestamp 1586364061
transform 1 0 3956 0 -1 213792
box -38 -48 130 592
use scs8hd_decap_4  FILLER_388_27
timestamp 1586364061
transform 1 0 3588 0 -1 213792
box -38 -48 406 592
use scs8hd_decap_12  FILLER_388_32
timestamp 1586364061
transform 1 0 4048 0 -1 213792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_388_44
timestamp 1586364061
transform 1 0 5152 0 -1 213792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_388_56
timestamp 1586364061
transform 1 0 6256 0 -1 213792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_388_68
timestamp 1586364061
transform 1 0 7360 0 -1 213792
box -38 -48 1142 592
use scs8hd_decap_3  PHY_777
timestamp 1586364061
transform -1 0 8832 0 -1 213792
box -38 -48 314 592
use scs8hd_fill_1  FILLER_388_80
timestamp 1586364061
transform 1 0 8464 0 -1 213792
box -38 -48 130 592
use scs8hd_decap_3  PHY_778
timestamp 1586364061
transform 1 0 1104 0 1 213792
box -38 -48 314 592
use scs8hd_decap_3  PHY_780
timestamp 1586364061
transform 1 0 1104 0 -1 214880
box -38 -48 314 592
use scs8hd_decap_12  FILLER_389_3
timestamp 1586364061
transform 1 0 1380 0 1 213792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_389_15
timestamp 1586364061
transform 1 0 2484 0 1 213792
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_390_3
timestamp 1586364061
transform 1 0 1380 0 -1 214880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_390_15
timestamp 1586364061
transform 1 0 2484 0 -1 214880
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1599
timestamp 1586364061
transform 1 0 3956 0 -1 214880
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3588 0 -1 214880
box -38 -48 222 592
use scs8hd_decap_12  FILLER_389_27
timestamp 1586364061
transform 1 0 3588 0 1 213792
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_390_29
timestamp 1586364061
transform 1 0 3772 0 -1 214880
box -38 -48 222 592
use scs8hd_decap_12  FILLER_390_32
timestamp 1586364061
transform 1 0 4048 0 -1 214880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_389_39
timestamp 1586364061
transform 1 0 4692 0 1 213792
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_389_51
timestamp 1586364061
transform 1 0 5796 0 1 213792
box -38 -48 774 592
use scs8hd_decap_12  FILLER_390_44
timestamp 1586364061
transform 1 0 5152 0 -1 214880
box -38 -48 1142 592
use scs8hd_buf_2  _17_
timestamp 1586364061
transform 1 0 7452 0 1 213792
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_1598
timestamp 1586364061
transform 1 0 6716 0 1 213792
box -38 -48 130 592
use scs8hd_fill_2  FILLER_389_59
timestamp 1586364061
transform 1 0 6532 0 1 213792
box -38 -48 222 592
use scs8hd_decap_6  FILLER_389_62
timestamp 1586364061
transform 1 0 6808 0 1 213792
box -38 -48 590 592
use scs8hd_fill_1  FILLER_389_68
timestamp 1586364061
transform 1 0 7360 0 1 213792
box -38 -48 130 592
use scs8hd_decap_12  FILLER_390_56
timestamp 1586364061
transform 1 0 6256 0 -1 214880
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_390_68
timestamp 1586364061
transform 1 0 7360 0 -1 214880
box -38 -48 1142 592
use scs8hd_decap_3  PHY_779
timestamp 1586364061
transform -1 0 8832 0 1 213792
box -38 -48 314 592
use scs8hd_decap_3  PHY_781
timestamp 1586364061
transform -1 0 8832 0 -1 214880
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__17__A
timestamp 1586364061
transform 1 0 8004 0 1 213792
box -38 -48 222 592
use scs8hd_fill_2  FILLER_389_73
timestamp 1586364061
transform 1 0 7820 0 1 213792
box -38 -48 222 592
use scs8hd_decap_4  FILLER_389_77
timestamp 1586364061
transform 1 0 8188 0 1 213792
box -38 -48 406 592
use scs8hd_fill_1  FILLER_390_80
timestamp 1586364061
transform 1 0 8464 0 -1 214880
box -38 -48 130 592
use scs8hd_decap_3  PHY_782
timestamp 1586364061
transform 1 0 1104 0 1 214880
box -38 -48 314 592
use scs8hd_decap_12  FILLER_391_3
timestamp 1586364061
transform 1 0 1380 0 1 214880
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_391_15
timestamp 1586364061
transform 1 0 2484 0 1 214880
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 3588 0 1 214880
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3404 0 1 214880
box -38 -48 222 592
use scs8hd_fill_2  FILLER_391_23
timestamp 1586364061
transform 1 0 3220 0 1 214880
box -38 -48 222 592
use scs8hd_decap_12  FILLER_391_38
timestamp 1586364061
transform 1 0 4600 0 1 214880
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_391_50
timestamp 1586364061
transform 1 0 5704 0 1 214880
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1600
timestamp 1586364061
transform 1 0 6716 0 1 214880
box -38 -48 130 592
use scs8hd_decap_3  FILLER_391_58
timestamp 1586364061
transform 1 0 6440 0 1 214880
box -38 -48 314 592
use scs8hd_decap_12  FILLER_391_62
timestamp 1586364061
transform 1 0 6808 0 1 214880
box -38 -48 1142 592
use scs8hd_decap_3  PHY_783
timestamp 1586364061
transform -1 0 8832 0 1 214880
box -38 -48 314 592
use scs8hd_decap_6  FILLER_391_74
timestamp 1586364061
transform 1 0 7912 0 1 214880
box -38 -48 590 592
use scs8hd_fill_1  FILLER_391_80
timestamp 1586364061
transform 1 0 8464 0 1 214880
box -38 -48 130 592
use scs8hd_decap_3  PHY_784
timestamp 1586364061
transform 1 0 1104 0 -1 215968
box -38 -48 314 592
use scs8hd_decap_12  FILLER_392_3
timestamp 1586364061
transform 1 0 1380 0 -1 215968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_392_15
timestamp 1586364061
transform 1 0 2484 0 -1 215968
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1601
timestamp 1586364061
transform 1 0 3956 0 -1 215968
box -38 -48 130 592
use scs8hd_decap_4  FILLER_392_27
timestamp 1586364061
transform 1 0 3588 0 -1 215968
box -38 -48 406 592
use scs8hd_decap_12  FILLER_392_32
timestamp 1586364061
transform 1 0 4048 0 -1 215968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_392_44
timestamp 1586364061
transform 1 0 5152 0 -1 215968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_392_56
timestamp 1586364061
transform 1 0 6256 0 -1 215968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_392_68
timestamp 1586364061
transform 1 0 7360 0 -1 215968
box -38 -48 1142 592
use scs8hd_decap_3  PHY_785
timestamp 1586364061
transform -1 0 8832 0 -1 215968
box -38 -48 314 592
use scs8hd_fill_1  FILLER_392_80
timestamp 1586364061
transform 1 0 8464 0 -1 215968
box -38 -48 130 592
use scs8hd_decap_3  PHY_786
timestamp 1586364061
transform 1 0 1104 0 1 215968
box -38 -48 314 592
use scs8hd_decap_12  FILLER_393_3
timestamp 1586364061
transform 1 0 1380 0 1 215968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_393_15
timestamp 1586364061
transform 1 0 2484 0 1 215968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_393_27
timestamp 1586364061
transform 1 0 3588 0 1 215968
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_393_39
timestamp 1586364061
transform 1 0 4692 0 1 215968
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_393_51
timestamp 1586364061
transform 1 0 5796 0 1 215968
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1602
timestamp 1586364061
transform 1 0 6716 0 1 215968
box -38 -48 130 592
use scs8hd_fill_2  FILLER_393_59
timestamp 1586364061
transform 1 0 6532 0 1 215968
box -38 -48 222 592
use scs8hd_decap_12  FILLER_393_62
timestamp 1586364061
transform 1 0 6808 0 1 215968
box -38 -48 1142 592
use scs8hd_decap_3  PHY_787
timestamp 1586364061
transform -1 0 8832 0 1 215968
box -38 -48 314 592
use scs8hd_decap_6  FILLER_393_74
timestamp 1586364061
transform 1 0 7912 0 1 215968
box -38 -48 590 592
use scs8hd_fill_1  FILLER_393_80
timestamp 1586364061
transform 1 0 8464 0 1 215968
box -38 -48 130 592
use scs8hd_decap_3  PHY_788
timestamp 1586364061
transform 1 0 1104 0 -1 217056
box -38 -48 314 592
use scs8hd_decap_12  FILLER_394_3
timestamp 1586364061
transform 1 0 1380 0 -1 217056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_394_15
timestamp 1586364061
transform 1 0 2484 0 -1 217056
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1603
timestamp 1586364061
transform 1 0 3956 0 -1 217056
box -38 -48 130 592
use scs8hd_decap_4  FILLER_394_27
timestamp 1586364061
transform 1 0 3588 0 -1 217056
box -38 -48 406 592
use scs8hd_decap_12  FILLER_394_32
timestamp 1586364061
transform 1 0 4048 0 -1 217056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_394_44
timestamp 1586364061
transform 1 0 5152 0 -1 217056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_394_56
timestamp 1586364061
transform 1 0 6256 0 -1 217056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_394_68
timestamp 1586364061
transform 1 0 7360 0 -1 217056
box -38 -48 1142 592
use scs8hd_decap_3  PHY_789
timestamp 1586364061
transform -1 0 8832 0 -1 217056
box -38 -48 314 592
use scs8hd_fill_1  FILLER_394_80
timestamp 1586364061
transform 1 0 8464 0 -1 217056
box -38 -48 130 592
use scs8hd_decap_3  PHY_790
timestamp 1586364061
transform 1 0 1104 0 1 217056
box -38 -48 314 592
use scs8hd_decap_12  FILLER_395_3
timestamp 1586364061
transform 1 0 1380 0 1 217056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_395_15
timestamp 1586364061
transform 1 0 2484 0 1 217056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_395_27
timestamp 1586364061
transform 1 0 3588 0 1 217056
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_395_39
timestamp 1586364061
transform 1 0 4692 0 1 217056
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_395_51
timestamp 1586364061
transform 1 0 5796 0 1 217056
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1604
timestamp 1586364061
transform 1 0 6716 0 1 217056
box -38 -48 130 592
use scs8hd_fill_2  FILLER_395_59
timestamp 1586364061
transform 1 0 6532 0 1 217056
box -38 -48 222 592
use scs8hd_decap_12  FILLER_395_62
timestamp 1586364061
transform 1 0 6808 0 1 217056
box -38 -48 1142 592
use scs8hd_decap_3  PHY_791
timestamp 1586364061
transform -1 0 8832 0 1 217056
box -38 -48 314 592
use scs8hd_decap_6  FILLER_395_74
timestamp 1586364061
transform 1 0 7912 0 1 217056
box -38 -48 590 592
use scs8hd_fill_1  FILLER_395_80
timestamp 1586364061
transform 1 0 8464 0 1 217056
box -38 -48 130 592
use scs8hd_decap_3  PHY_792
timestamp 1586364061
transform 1 0 1104 0 -1 218144
box -38 -48 314 592
use scs8hd_decap_3  PHY_794
timestamp 1586364061
transform 1 0 1104 0 1 218144
box -38 -48 314 592
use scs8hd_decap_12  FILLER_396_3
timestamp 1586364061
transform 1 0 1380 0 -1 218144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_396_15
timestamp 1586364061
transform 1 0 2484 0 -1 218144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_397_3
timestamp 1586364061
transform 1 0 1380 0 1 218144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_397_15
timestamp 1586364061
transform 1 0 2484 0 1 218144
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1605
timestamp 1586364061
transform 1 0 3956 0 -1 218144
box -38 -48 130 592
use scs8hd_decap_4  FILLER_396_27
timestamp 1586364061
transform 1 0 3588 0 -1 218144
box -38 -48 406 592
use scs8hd_decap_12  FILLER_396_32
timestamp 1586364061
transform 1 0 4048 0 -1 218144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_397_27
timestamp 1586364061
transform 1 0 3588 0 1 218144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_396_44
timestamp 1586364061
transform 1 0 5152 0 -1 218144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_397_39
timestamp 1586364061
transform 1 0 4692 0 1 218144
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_397_51
timestamp 1586364061
transform 1 0 5796 0 1 218144
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1606
timestamp 1586364061
transform 1 0 6716 0 1 218144
box -38 -48 130 592
use scs8hd_decap_12  FILLER_396_56
timestamp 1586364061
transform 1 0 6256 0 -1 218144
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_396_68
timestamp 1586364061
transform 1 0 7360 0 -1 218144
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_397_59
timestamp 1586364061
transform 1 0 6532 0 1 218144
box -38 -48 222 592
use scs8hd_decap_12  FILLER_397_62
timestamp 1586364061
transform 1 0 6808 0 1 218144
box -38 -48 1142 592
use scs8hd_decap_3  PHY_793
timestamp 1586364061
transform -1 0 8832 0 -1 218144
box -38 -48 314 592
use scs8hd_decap_3  PHY_795
timestamp 1586364061
transform -1 0 8832 0 1 218144
box -38 -48 314 592
use scs8hd_fill_1  FILLER_396_80
timestamp 1586364061
transform 1 0 8464 0 -1 218144
box -38 -48 130 592
use scs8hd_decap_6  FILLER_397_74
timestamp 1586364061
transform 1 0 7912 0 1 218144
box -38 -48 590 592
use scs8hd_fill_1  FILLER_397_80
timestamp 1586364061
transform 1 0 8464 0 1 218144
box -38 -48 130 592
use scs8hd_decap_3  PHY_796
timestamp 1586364061
transform 1 0 1104 0 -1 219232
box -38 -48 314 592
use scs8hd_decap_12  FILLER_398_3
timestamp 1586364061
transform 1 0 1380 0 -1 219232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_398_15
timestamp 1586364061
transform 1 0 2484 0 -1 219232
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1607
timestamp 1586364061
transform 1 0 3956 0 -1 219232
box -38 -48 130 592
use scs8hd_decap_4  FILLER_398_27
timestamp 1586364061
transform 1 0 3588 0 -1 219232
box -38 -48 406 592
use scs8hd_decap_12  FILLER_398_32
timestamp 1586364061
transform 1 0 4048 0 -1 219232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_398_44
timestamp 1586364061
transform 1 0 5152 0 -1 219232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_398_56
timestamp 1586364061
transform 1 0 6256 0 -1 219232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_398_68
timestamp 1586364061
transform 1 0 7360 0 -1 219232
box -38 -48 1142 592
use scs8hd_decap_3  PHY_797
timestamp 1586364061
transform -1 0 8832 0 -1 219232
box -38 -48 314 592
use scs8hd_fill_1  FILLER_398_80
timestamp 1586364061
transform 1 0 8464 0 -1 219232
box -38 -48 130 592
use scs8hd_decap_3  PHY_798
timestamp 1586364061
transform 1 0 1104 0 1 219232
box -38 -48 314 592
use scs8hd_decap_12  FILLER_399_3
timestamp 1586364061
transform 1 0 1380 0 1 219232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_399_15
timestamp 1586364061
transform 1 0 2484 0 1 219232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_399_27
timestamp 1586364061
transform 1 0 3588 0 1 219232
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_399_39
timestamp 1586364061
transform 1 0 4692 0 1 219232
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_399_51
timestamp 1586364061
transform 1 0 5796 0 1 219232
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1608
timestamp 1586364061
transform 1 0 6716 0 1 219232
box -38 -48 130 592
use scs8hd_fill_2  FILLER_399_59
timestamp 1586364061
transform 1 0 6532 0 1 219232
box -38 -48 222 592
use scs8hd_decap_12  FILLER_399_62
timestamp 1586364061
transform 1 0 6808 0 1 219232
box -38 -48 1142 592
use scs8hd_decap_3  PHY_799
timestamp 1586364061
transform -1 0 8832 0 1 219232
box -38 -48 314 592
use scs8hd_decap_6  FILLER_399_74
timestamp 1586364061
transform 1 0 7912 0 1 219232
box -38 -48 590 592
use scs8hd_fill_1  FILLER_399_80
timestamp 1586364061
transform 1 0 8464 0 1 219232
box -38 -48 130 592
use scs8hd_decap_3  PHY_800
timestamp 1586364061
transform 1 0 1104 0 -1 220320
box -38 -48 314 592
use scs8hd_decap_12  FILLER_400_3
timestamp 1586364061
transform 1 0 1380 0 -1 220320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_400_15
timestamp 1586364061
transform 1 0 2484 0 -1 220320
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1609
timestamp 1586364061
transform 1 0 3956 0 -1 220320
box -38 -48 130 592
use scs8hd_decap_4  FILLER_400_27
timestamp 1586364061
transform 1 0 3588 0 -1 220320
box -38 -48 406 592
use scs8hd_decap_12  FILLER_400_32
timestamp 1586364061
transform 1 0 4048 0 -1 220320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_400_44
timestamp 1586364061
transform 1 0 5152 0 -1 220320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_400_56
timestamp 1586364061
transform 1 0 6256 0 -1 220320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_400_68
timestamp 1586364061
transform 1 0 7360 0 -1 220320
box -38 -48 1142 592
use scs8hd_decap_3  PHY_801
timestamp 1586364061
transform -1 0 8832 0 -1 220320
box -38 -48 314 592
use scs8hd_fill_1  FILLER_400_80
timestamp 1586364061
transform 1 0 8464 0 -1 220320
box -38 -48 130 592
use scs8hd_decap_3  PHY_802
timestamp 1586364061
transform 1 0 1104 0 1 220320
box -38 -48 314 592
use scs8hd_decap_12  FILLER_401_3
timestamp 1586364061
transform 1 0 1380 0 1 220320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_401_15
timestamp 1586364061
transform 1 0 2484 0 1 220320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_401_27
timestamp 1586364061
transform 1 0 3588 0 1 220320
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_401_39
timestamp 1586364061
transform 1 0 4692 0 1 220320
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_401_51
timestamp 1586364061
transform 1 0 5796 0 1 220320
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1610
timestamp 1586364061
transform 1 0 6716 0 1 220320
box -38 -48 130 592
use scs8hd_fill_2  FILLER_401_59
timestamp 1586364061
transform 1 0 6532 0 1 220320
box -38 -48 222 592
use scs8hd_decap_12  FILLER_401_62
timestamp 1586364061
transform 1 0 6808 0 1 220320
box -38 -48 1142 592
use scs8hd_decap_3  PHY_803
timestamp 1586364061
transform -1 0 8832 0 1 220320
box -38 -48 314 592
use scs8hd_decap_6  FILLER_401_74
timestamp 1586364061
transform 1 0 7912 0 1 220320
box -38 -48 590 592
use scs8hd_fill_1  FILLER_401_80
timestamp 1586364061
transform 1 0 8464 0 1 220320
box -38 -48 130 592
use scs8hd_decap_3  PHY_804
timestamp 1586364061
transform 1 0 1104 0 -1 221408
box -38 -48 314 592
use scs8hd_decap_12  FILLER_402_3
timestamp 1586364061
transform 1 0 1380 0 -1 221408
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_402_15
timestamp 1586364061
transform 1 0 2484 0 -1 221408
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_1611
timestamp 1586364061
transform 1 0 3956 0 -1 221408
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__07__D
timestamp 1586364061
transform 1 0 2944 0 -1 221408
box -38 -48 222 592
use scs8hd_fill_1  FILLER_402_19
timestamp 1586364061
transform 1 0 2852 0 -1 221408
box -38 -48 130 592
use scs8hd_decap_8  FILLER_402_22
timestamp 1586364061
transform 1 0 3128 0 -1 221408
box -38 -48 774 592
use scs8hd_fill_1  FILLER_402_30
timestamp 1586364061
transform 1 0 3864 0 -1 221408
box -38 -48 130 592
use scs8hd_decap_12  FILLER_402_32
timestamp 1586364061
transform 1 0 4048 0 -1 221408
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_402_44
timestamp 1586364061
transform 1 0 5152 0 -1 221408
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_402_56
timestamp 1586364061
transform 1 0 6256 0 -1 221408
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_402_68
timestamp 1586364061
transform 1 0 7360 0 -1 221408
box -38 -48 1142 592
use scs8hd_decap_3  PHY_805
timestamp 1586364061
transform -1 0 8832 0 -1 221408
box -38 -48 314 592
use scs8hd_fill_1  FILLER_402_80
timestamp 1586364061
transform 1 0 8464 0 -1 221408
box -38 -48 130 592
use scs8hd_decap_3  PHY_806
timestamp 1586364061
transform 1 0 1104 0 1 221408
box -38 -48 314 592
use scs8hd_decap_3  PHY_808
timestamp 1586364061
transform 1 0 1104 0 -1 222496
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__07__C
timestamp 1586364061
transform 1 0 2392 0 1 221408
box -38 -48 222 592
use scs8hd_decap_8  FILLER_403_3
timestamp 1586364061
transform 1 0 1380 0 1 221408
box -38 -48 774 592
use scs8hd_decap_3  FILLER_403_11
timestamp 1586364061
transform 1 0 2116 0 1 221408
box -38 -48 314 592
use scs8hd_fill_2  FILLER_403_16
timestamp 1586364061
transform 1 0 2576 0 1 221408
box -38 -48 222 592
use scs8hd_decap_12  FILLER_404_3
timestamp 1586364061
transform 1 0 1380 0 -1 222496
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_404_15
timestamp 1586364061
transform 1 0 2484 0 -1 222496
box -38 -48 406 592
use scs8hd_decap_8  FILLER_404_22
timestamp 1586364061
transform 1 0 3128 0 -1 222496
box -38 -48 774 592
use scs8hd_fill_1  FILLER_404_19
timestamp 1586364061
transform 1 0 2852 0 -1 222496
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__07__A
timestamp 1586364061
transform 1 0 2944 0 -1 222496
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__07__B
timestamp 1586364061
transform 1 0 2760 0 1 221408
box -38 -48 222 592
use scs8hd_fill_1  FILLER_404_30
timestamp 1586364061
transform 1 0 3864 0 -1 222496
box -38 -48 130 592
use scs8hd_decap_6  FILLER_403_29
timestamp 1586364061
transform 1 0 3772 0 1 221408
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__11__A
timestamp 1586364061
transform 1 0 4324 0 1 221408
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_1613
timestamp 1586364061
transform 1 0 3956 0 -1 222496
box -38 -48 130 592
use scs8hd_decap_12  FILLER_404_32
timestamp 1586364061
transform 1 0 4048 0 -1 222496
box -38 -48 1142 592
use scs8hd_and4_4  _07_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2944 0 1 221408
box -38 -48 866 592
use scs8hd_inv_8  _11_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4508 0 1 221408
box -38 -48 866 592
use scs8hd_decap_12  FILLER_403_46
timestamp 1586364061
transform 1 0 5336 0 1 221408
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_404_44
timestamp 1586364061
transform 1 0 5152 0 -1 222496
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1612
timestamp 1586364061
transform 1 0 6716 0 1 221408
box -38 -48 130 592
use scs8hd_decap_3  FILLER_403_58
timestamp 1586364061
transform 1 0 6440 0 1 221408
box -38 -48 314 592
use scs8hd_decap_12  FILLER_403_62
timestamp 1586364061
transform 1 0 6808 0 1 221408
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_404_56
timestamp 1586364061
transform 1 0 6256 0 -1 222496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_404_68
timestamp 1586364061
transform 1 0 7360 0 -1 222496
box -38 -48 1142 592
use scs8hd_decap_3  PHY_807
timestamp 1586364061
transform -1 0 8832 0 1 221408
box -38 -48 314 592
use scs8hd_decap_3  PHY_809
timestamp 1586364061
transform -1 0 8832 0 -1 222496
box -38 -48 314 592
use scs8hd_decap_6  FILLER_403_74
timestamp 1586364061
transform 1 0 7912 0 1 221408
box -38 -48 590 592
use scs8hd_fill_1  FILLER_403_80
timestamp 1586364061
transform 1 0 8464 0 1 221408
box -38 -48 130 592
use scs8hd_fill_1  FILLER_404_80
timestamp 1586364061
transform 1 0 8464 0 -1 222496
box -38 -48 130 592
use scs8hd_decap_3  PHY_810
timestamp 1586364061
transform 1 0 1104 0 1 222496
box -38 -48 314 592
use scs8hd_decap_12  FILLER_405_3
timestamp 1586364061
transform 1 0 1380 0 1 222496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_405_15
timestamp 1586364061
transform 1 0 2484 0 1 222496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_405_27
timestamp 1586364061
transform 1 0 3588 0 1 222496
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_405_39
timestamp 1586364061
transform 1 0 4692 0 1 222496
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_405_51
timestamp 1586364061
transform 1 0 5796 0 1 222496
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1614
timestamp 1586364061
transform 1 0 6716 0 1 222496
box -38 -48 130 592
use scs8hd_fill_2  FILLER_405_59
timestamp 1586364061
transform 1 0 6532 0 1 222496
box -38 -48 222 592
use scs8hd_decap_12  FILLER_405_62
timestamp 1586364061
transform 1 0 6808 0 1 222496
box -38 -48 1142 592
use scs8hd_decap_3  PHY_811
timestamp 1586364061
transform -1 0 8832 0 1 222496
box -38 -48 314 592
use scs8hd_decap_6  FILLER_405_74
timestamp 1586364061
transform 1 0 7912 0 1 222496
box -38 -48 590 592
use scs8hd_fill_1  FILLER_405_80
timestamp 1586364061
transform 1 0 8464 0 1 222496
box -38 -48 130 592
use scs8hd_decap_3  PHY_812
timestamp 1586364061
transform 1 0 1104 0 -1 223584
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__14__C
timestamp 1586364061
transform 1 0 2576 0 -1 223584
box -38 -48 222 592
use scs8hd_decap_12  FILLER_406_3
timestamp 1586364061
transform 1 0 1380 0 -1 223584
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_406_15
timestamp 1586364061
transform 1 0 2484 0 -1 223584
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_1615
timestamp 1586364061
transform 1 0 3956 0 -1 223584
box -38 -48 130 592
use scs8hd_decap_12  FILLER_406_18
timestamp 1586364061
transform 1 0 2760 0 -1 223584
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_406_30
timestamp 1586364061
transform 1 0 3864 0 -1 223584
box -38 -48 130 592
use scs8hd_decap_12  FILLER_406_32
timestamp 1586364061
transform 1 0 4048 0 -1 223584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_406_44
timestamp 1586364061
transform 1 0 5152 0 -1 223584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_406_56
timestamp 1586364061
transform 1 0 6256 0 -1 223584
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_406_68
timestamp 1586364061
transform 1 0 7360 0 -1 223584
box -38 -48 1142 592
use scs8hd_decap_3  PHY_813
timestamp 1586364061
transform -1 0 8832 0 -1 223584
box -38 -48 314 592
use scs8hd_fill_1  FILLER_406_80
timestamp 1586364061
transform 1 0 8464 0 -1 223584
box -38 -48 130 592
use scs8hd_nor4_4  _14_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2576 0 1 223584
box -38 -48 1602 592
use scs8hd_decap_3  PHY_814
timestamp 1586364061
transform 1 0 1104 0 1 223584
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__14__D
timestamp 1586364061
transform 1 0 2392 0 1 223584
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__14__B
timestamp 1586364061
transform 1 0 2024 0 1 223584
box -38 -48 222 592
use scs8hd_decap_6  FILLER_407_3
timestamp 1586364061
transform 1 0 1380 0 1 223584
box -38 -48 590 592
use scs8hd_fill_1  FILLER_407_9
timestamp 1586364061
transform 1 0 1932 0 1 223584
box -38 -48 130 592
use scs8hd_fill_2  FILLER_407_12
timestamp 1586364061
transform 1 0 2208 0 1 223584
box -38 -48 222 592
use scs8hd_decap_12  FILLER_407_33
timestamp 1586364061
transform 1 0 4140 0 1 223584
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 5796 0 1 223584
box -38 -48 222 592
use scs8hd_decap_6  FILLER_407_45
timestamp 1586364061
transform 1 0 5244 0 1 223584
box -38 -48 590 592
use scs8hd_fill_2  FILLER_407_53
timestamp 1586364061
transform 1 0 5980 0 1 223584
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_1616
timestamp 1586364061
transform 1 0 6716 0 1 223584
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 6164 0 1 223584
box -38 -48 222 592
use scs8hd_decap_4  FILLER_407_57
timestamp 1586364061
transform 1 0 6348 0 1 223584
box -38 -48 406 592
use scs8hd_decap_12  FILLER_407_62
timestamp 1586364061
transform 1 0 6808 0 1 223584
box -38 -48 1142 592
use scs8hd_decap_3  PHY_815
timestamp 1586364061
transform -1 0 8832 0 1 223584
box -38 -48 314 592
use scs8hd_decap_6  FILLER_407_74
timestamp 1586364061
transform 1 0 7912 0 1 223584
box -38 -48 590 592
use scs8hd_fill_1  FILLER_407_80
timestamp 1586364061
transform 1 0 8464 0 1 223584
box -38 -48 130 592
use scs8hd_decap_3  PHY_816
timestamp 1586364061
transform 1 0 1104 0 -1 224672
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__14__A
timestamp 1586364061
transform 1 0 2576 0 -1 224672
box -38 -48 222 592
use scs8hd_decap_12  FILLER_408_3
timestamp 1586364061
transform 1 0 1380 0 -1 224672
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_408_15
timestamp 1586364061
transform 1 0 2484 0 -1 224672
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_1617
timestamp 1586364061
transform 1 0 3956 0 -1 224672
box -38 -48 130 592
use scs8hd_decap_12  FILLER_408_18
timestamp 1586364061
transform 1 0 2760 0 -1 224672
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_408_30
timestamp 1586364061
transform 1 0 3864 0 -1 224672
box -38 -48 130 592
use scs8hd_decap_12  FILLER_408_32
timestamp 1586364061
transform 1 0 4048 0 -1 224672
box -38 -48 1142 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 5796 0 -1 224672
box -38 -48 774 592
use scs8hd_decap_6  FILLER_408_44
timestamp 1586364061
transform 1 0 5152 0 -1 224672
box -38 -48 590 592
use scs8hd_fill_1  FILLER_408_50
timestamp 1586364061
transform 1 0 5704 0 -1 224672
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 6808 0 -1 224672
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 7176 0 -1 224672
box -38 -48 222 592
use scs8hd_decap_3  FILLER_408_59
timestamp 1586364061
transform 1 0 6532 0 -1 224672
box -38 -48 314 592
use scs8hd_fill_2  FILLER_408_64
timestamp 1586364061
transform 1 0 6992 0 -1 224672
box -38 -48 222 592
use scs8hd_decap_12  FILLER_408_68
timestamp 1586364061
transform 1 0 7360 0 -1 224672
box -38 -48 1142 592
use scs8hd_decap_3  PHY_817
timestamp 1586364061
transform -1 0 8832 0 -1 224672
box -38 -48 314 592
use scs8hd_fill_1  FILLER_408_80
timestamp 1586364061
transform 1 0 8464 0 -1 224672
box -38 -48 130 592
use scs8hd_decap_3  PHY_818
timestamp 1586364061
transform 1 0 1104 0 1 224672
box -38 -48 314 592
use scs8hd_decap_3  PHY_820
timestamp 1586364061
transform 1 0 1104 0 -1 225760
box -38 -48 314 592
use scs8hd_decap_12  FILLER_409_3
timestamp 1586364061
transform 1 0 1380 0 1 224672
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_409_15
timestamp 1586364061
transform 1 0 2484 0 1 224672
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_410_3
timestamp 1586364061
transform 1 0 1380 0 -1 225760
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_410_15
timestamp 1586364061
transform 1 0 2484 0 -1 225760
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1619
timestamp 1586364061
transform 1 0 3956 0 -1 225760
box -38 -48 130 592
use scs8hd_decap_8  FILLER_409_27
timestamp 1586364061
transform 1 0 3588 0 1 224672
box -38 -48 774 592
use scs8hd_fill_1  FILLER_409_35
timestamp 1586364061
transform 1 0 4324 0 1 224672
box -38 -48 130 592
use scs8hd_decap_4  FILLER_410_27
timestamp 1586364061
transform 1 0 3588 0 -1 225760
box -38 -48 406 592
use scs8hd_decap_4  FILLER_410_32
timestamp 1586364061
transform 1 0 4048 0 -1 225760
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4416 0 -1 225760
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4416 0 1 224672
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4784 0 1 224672
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 5888 0 1 224672
box -38 -48 222 592
use scs8hd_fill_2  FILLER_409_38
timestamp 1586364061
transform 1 0 4600 0 1 224672
box -38 -48 222 592
use scs8hd_decap_8  FILLER_409_42
timestamp 1586364061
transform 1 0 4968 0 1 224672
box -38 -48 774 592
use scs8hd_fill_2  FILLER_409_50
timestamp 1586364061
transform 1 0 5704 0 1 224672
box -38 -48 222 592
use scs8hd_decap_8  FILLER_410_47
timestamp 1586364061
transform 1 0 5428 0 -1 225760
box -38 -48 774 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 6808 0 1 224672
box -38 -48 774 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 6256 0 -1 225760
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1618
timestamp 1586364061
transform 1 0 6716 0 1 224672
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 6256 0 1 224672
box -38 -48 222 592
use scs8hd_fill_2  FILLER_409_54
timestamp 1586364061
transform 1 0 6072 0 1 224672
box -38 -48 222 592
use scs8hd_decap_3  FILLER_409_58
timestamp 1586364061
transform 1 0 6440 0 1 224672
box -38 -48 314 592
use scs8hd_decap_8  FILLER_409_70
timestamp 1586364061
transform 1 0 7544 0 1 224672
box -38 -48 774 592
use scs8hd_fill_1  FILLER_410_55
timestamp 1586364061
transform 1 0 6164 0 -1 225760
box -38 -48 130 592
use scs8hd_decap_12  FILLER_410_64
timestamp 1586364061
transform 1 0 6992 0 -1 225760
box -38 -48 1142 592
use scs8hd_decap_3  PHY_819
timestamp 1586364061
transform -1 0 8832 0 1 224672
box -38 -48 314 592
use scs8hd_decap_3  PHY_821
timestamp 1586364061
transform -1 0 8832 0 -1 225760
box -38 -48 314 592
use scs8hd_decap_3  FILLER_409_78
timestamp 1586364061
transform 1 0 8280 0 1 224672
box -38 -48 314 592
use scs8hd_decap_4  FILLER_410_76
timestamp 1586364061
transform 1 0 8096 0 -1 225760
box -38 -48 406 592
use scs8hd_fill_1  FILLER_410_80
timestamp 1586364061
transform 1 0 8464 0 -1 225760
box -38 -48 130 592
use scs8hd_decap_3  PHY_822
timestamp 1586364061
transform 1 0 1104 0 1 225760
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__08__A
timestamp 1586364061
transform 1 0 2392 0 1 225760
box -38 -48 222 592
use scs8hd_decap_8  FILLER_411_3
timestamp 1586364061
transform 1 0 1380 0 1 225760
box -38 -48 774 592
use scs8hd_decap_3  FILLER_411_11
timestamp 1586364061
transform 1 0 2116 0 1 225760
box -38 -48 314 592
use scs8hd_decap_8  FILLER_411_16
timestamp 1586364061
transform 1 0 2576 0 1 225760
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4232 0 1 225760
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3864 0 1 225760
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3496 0 1 225760
box -38 -48 222 592
use scs8hd_fill_2  FILLER_411_24
timestamp 1586364061
transform 1 0 3312 0 1 225760
box -38 -48 222 592
use scs8hd_fill_2  FILLER_411_28
timestamp 1586364061
transform 1 0 3680 0 1 225760
box -38 -48 222 592
use scs8hd_fill_2  FILLER_411_32
timestamp 1586364061
transform 1 0 4048 0 1 225760
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4416 0 1 225760
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5612 0 1 225760
box -38 -48 222 592
use scs8hd_fill_2  FILLER_411_47
timestamp 1586364061
transform 1 0 5428 0 1 225760
box -38 -48 222 592
use scs8hd_decap_8  FILLER_411_51
timestamp 1586364061
transform 1 0 5796 0 1 225760
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1620
timestamp 1586364061
transform 1 0 6716 0 1 225760
box -38 -48 130 592
use scs8hd_fill_2  FILLER_411_59
timestamp 1586364061
transform 1 0 6532 0 1 225760
box -38 -48 222 592
use scs8hd_decap_12  FILLER_411_62
timestamp 1586364061
transform 1 0 6808 0 1 225760
box -38 -48 1142 592
use scs8hd_decap_3  PHY_823
timestamp 1586364061
transform -1 0 8832 0 1 225760
box -38 -48 314 592
use scs8hd_decap_6  FILLER_411_74
timestamp 1586364061
transform 1 0 7912 0 1 225760
box -38 -48 590 592
use scs8hd_fill_1  FILLER_411_80
timestamp 1586364061
transform 1 0 8464 0 1 225760
box -38 -48 130 592
use scs8hd_inv_8  _08_
timestamp 1586364061
transform 1 0 2392 0 -1 226848
box -38 -48 866 592
use scs8hd_decap_3  PHY_824
timestamp 1586364061
transform 1 0 1104 0 -1 226848
box -38 -48 314 592
use scs8hd_decap_8  FILLER_412_3
timestamp 1586364061
transform 1 0 1380 0 -1 226848
box -38 -48 774 592
use scs8hd_decap_3  FILLER_412_11
timestamp 1586364061
transform 1 0 2116 0 -1 226848
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_1621
timestamp 1586364061
transform 1 0 3956 0 -1 226848
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__15__C
timestamp 1586364061
transform 1 0 3404 0 -1 226848
box -38 -48 222 592
use scs8hd_fill_2  FILLER_412_23
timestamp 1586364061
transform 1 0 3220 0 -1 226848
box -38 -48 222 592
use scs8hd_decap_4  FILLER_412_27
timestamp 1586364061
transform 1 0 3588 0 -1 226848
box -38 -48 406 592
use scs8hd_decap_4  FILLER_412_32
timestamp 1586364061
transform 1 0 4048 0 -1 226848
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4416 0 -1 226848
box -38 -48 1050 592
use scs8hd_decap_12  FILLER_412_47
timestamp 1586364061
transform 1 0 5428 0 -1 226848
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_412_59
timestamp 1586364061
transform 1 0 6532 0 -1 226848
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_412_71
timestamp 1586364061
transform 1 0 7636 0 -1 226848
box -38 -48 774 592
use scs8hd_decap_3  PHY_825
timestamp 1586364061
transform -1 0 8832 0 -1 226848
box -38 -48 314 592
use scs8hd_fill_2  FILLER_412_79
timestamp 1586364061
transform 1 0 8372 0 -1 226848
box -38 -48 222 592
use scs8hd_decap_3  PHY_826
timestamp 1586364061
transform 1 0 1104 0 1 226848
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__15__A
timestamp 1586364061
transform 1 0 2668 0 1 226848
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__15__D
timestamp 1586364061
transform 1 0 2300 0 1 226848
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__04__A
timestamp 1586364061
transform 1 0 1932 0 1 226848
box -38 -48 222 592
use scs8hd_decap_6  FILLER_413_3
timestamp 1586364061
transform 1 0 1380 0 1 226848
box -38 -48 590 592
use scs8hd_fill_2  FILLER_413_11
timestamp 1586364061
transform 1 0 2116 0 1 226848
box -38 -48 222 592
use scs8hd_fill_2  FILLER_413_15
timestamp 1586364061
transform 1 0 2484 0 1 226848
box -38 -48 222 592
use scs8hd_nor4_4  _15_
timestamp 1586364061
transform 1 0 2852 0 1 226848
box -38 -48 1602 592
use scs8hd_decap_12  FILLER_413_36
timestamp 1586364061
transform 1 0 4416 0 1 226848
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_413_48
timestamp 1586364061
transform 1 0 5520 0 1 226848
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1622
timestamp 1586364061
transform 1 0 6716 0 1 226848
box -38 -48 130 592
use scs8hd_fill_1  FILLER_413_60
timestamp 1586364061
transform 1 0 6624 0 1 226848
box -38 -48 130 592
use scs8hd_decap_12  FILLER_413_62
timestamp 1586364061
transform 1 0 6808 0 1 226848
box -38 -48 1142 592
use scs8hd_decap_3  PHY_827
timestamp 1586364061
transform -1 0 8832 0 1 226848
box -38 -48 314 592
use scs8hd_decap_6  FILLER_413_74
timestamp 1586364061
transform 1 0 7912 0 1 226848
box -38 -48 590 592
use scs8hd_fill_1  FILLER_413_80
timestamp 1586364061
transform 1 0 8464 0 1 226848
box -38 -48 130 592
use scs8hd_decap_3  PHY_828
timestamp 1586364061
transform 1 0 1104 0 -1 227936
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__10__B
timestamp 1586364061
transform 1 0 2392 0 -1 227936
box -38 -48 222 592
use scs8hd_decap_8  FILLER_414_3
timestamp 1586364061
transform 1 0 1380 0 -1 227936
box -38 -48 774 592
use scs8hd_decap_3  FILLER_414_11
timestamp 1586364061
transform 1 0 2116 0 -1 227936
box -38 -48 314 592
use scs8hd_decap_3  FILLER_414_16
timestamp 1586364061
transform 1 0 2576 0 -1 227936
box -38 -48 314 592
use scs8hd_buf_1  _04_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2852 0 -1 227936
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_1623
timestamp 1586364061
transform 1 0 3956 0 -1 227936
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__05__D
timestamp 1586364061
transform 1 0 3312 0 -1 227936
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__15__B
timestamp 1586364061
transform 1 0 3680 0 -1 227936
box -38 -48 222 592
use scs8hd_fill_2  FILLER_414_22
timestamp 1586364061
transform 1 0 3128 0 -1 227936
box -38 -48 222 592
use scs8hd_fill_2  FILLER_414_26
timestamp 1586364061
transform 1 0 3496 0 -1 227936
box -38 -48 222 592
use scs8hd_fill_1  FILLER_414_30
timestamp 1586364061
transform 1 0 3864 0 -1 227936
box -38 -48 130 592
use scs8hd_decap_12  FILLER_414_32
timestamp 1586364061
transform 1 0 4048 0 -1 227936
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_414_44
timestamp 1586364061
transform 1 0 5152 0 -1 227936
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_414_56
timestamp 1586364061
transform 1 0 6256 0 -1 227936
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_414_68
timestamp 1586364061
transform 1 0 7360 0 -1 227936
box -38 -48 1142 592
use scs8hd_decap_3  PHY_829
timestamp 1586364061
transform -1 0 8832 0 -1 227936
box -38 -48 314 592
use scs8hd_fill_1  FILLER_414_80
timestamp 1586364061
transform 1 0 8464 0 -1 227936
box -38 -48 130 592
use scs8hd_decap_3  PHY_830
timestamp 1586364061
transform 1 0 1104 0 1 227936
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__05__B
timestamp 1586364061
transform 1 0 2392 0 1 227936
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__10__C
timestamp 1586364061
transform 1 0 2024 0 1 227936
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__10__A
timestamp 1586364061
transform 1 0 1656 0 1 227936
box -38 -48 222 592
use scs8hd_decap_3  FILLER_415_3
timestamp 1586364061
transform 1 0 1380 0 1 227936
box -38 -48 314 592
use scs8hd_fill_2  FILLER_415_8
timestamp 1586364061
transform 1 0 1840 0 1 227936
box -38 -48 222 592
use scs8hd_fill_2  FILLER_415_12
timestamp 1586364061
transform 1 0 2208 0 1 227936
box -38 -48 222 592
use scs8hd_fill_2  FILLER_415_16
timestamp 1586364061
transform 1 0 2576 0 1 227936
box -38 -48 222 592
use scs8hd_and4_4  _05_
timestamp 1586364061
transform 1 0 2944 0 1 227936
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__06__A
timestamp 1586364061
transform 1 0 4048 0 1 227936
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__05__C
timestamp 1586364061
transform 1 0 2760 0 1 227936
box -38 -48 222 592
use scs8hd_decap_3  FILLER_415_29
timestamp 1586364061
transform 1 0 3772 0 1 227936
box -38 -48 314 592
use scs8hd_decap_12  FILLER_415_34
timestamp 1586364061
transform 1 0 4232 0 1 227936
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_415_46
timestamp 1586364061
transform 1 0 5336 0 1 227936
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1624
timestamp 1586364061
transform 1 0 6716 0 1 227936
box -38 -48 130 592
use scs8hd_decap_3  FILLER_415_58
timestamp 1586364061
transform 1 0 6440 0 1 227936
box -38 -48 314 592
use scs8hd_decap_12  FILLER_415_62
timestamp 1586364061
transform 1 0 6808 0 1 227936
box -38 -48 1142 592
use scs8hd_decap_3  PHY_831
timestamp 1586364061
transform -1 0 8832 0 1 227936
box -38 -48 314 592
use scs8hd_decap_6  FILLER_415_74
timestamp 1586364061
transform 1 0 7912 0 1 227936
box -38 -48 590 592
use scs8hd_fill_1  FILLER_415_80
timestamp 1586364061
transform 1 0 8464 0 1 227936
box -38 -48 130 592
use scs8hd_decap_6  FILLER_417_3
timestamp 1586364061
transform 1 0 1380 0 1 229024
box -38 -48 590 592
use scs8hd_decap_8  FILLER_416_3
timestamp 1586364061
transform 1 0 1380 0 -1 229024
box -38 -48 774 592
use scs8hd_decap_3  PHY_834
timestamp 1586364061
transform 1 0 1104 0 1 229024
box -38 -48 314 592
use scs8hd_decap_3  PHY_832
timestamp 1586364061
transform 1 0 1104 0 -1 229024
box -38 -48 314 592
use scs8hd_fill_2  FILLER_417_15
timestamp 1586364061
transform 1 0 2484 0 1 229024
box -38 -48 222 592
use scs8hd_fill_2  FILLER_417_11
timestamp 1586364061
transform 1 0 2116 0 1 229024
box -38 -48 222 592
use scs8hd_fill_1  FILLER_416_11
timestamp 1586364061
transform 1 0 2116 0 -1 229024
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__12__B
timestamp 1586364061
transform 1 0 1932 0 1 229024
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__10__D
timestamp 1586364061
transform 1 0 2208 0 -1 229024
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__12__A
timestamp 1586364061
transform 1 0 2300 0 1 229024
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__12__C
timestamp 1586364061
transform 1 0 2668 0 1 229024
box -38 -48 222 592
use scs8hd_and4_4  _10_
timestamp 1586364061
transform 1 0 2392 0 -1 229024
box -38 -48 866 592
use scs8hd_inv_8  _06_
timestamp 1586364061
transform 1 0 4048 0 -1 229024
box -38 -48 866 592
use scs8hd_nor4_4  _12_
timestamp 1586364061
transform 1 0 2852 0 1 229024
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_1625
timestamp 1586364061
transform 1 0 3956 0 -1 229024
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__05__A
timestamp 1586364061
transform 1 0 3404 0 -1 229024
box -38 -48 222 592
use scs8hd_fill_2  FILLER_416_23
timestamp 1586364061
transform 1 0 3220 0 -1 229024
box -38 -48 222 592
use scs8hd_decap_4  FILLER_416_27
timestamp 1586364061
transform 1 0 3588 0 -1 229024
box -38 -48 406 592
use scs8hd_fill_2  FILLER_417_44
timestamp 1586364061
transform 1 0 5152 0 1 229024
box -38 -48 222 592
use scs8hd_fill_2  FILLER_417_40
timestamp 1586364061
transform 1 0 4784 0 1 229024
box -38 -48 222 592
use scs8hd_fill_2  FILLER_417_36
timestamp 1586364061
transform 1 0 4416 0 1 229024
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__09__C
timestamp 1586364061
transform 1 0 4968 0 1 229024
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__09__A
timestamp 1586364061
transform 1 0 4600 0 1 229024
box -38 -48 222 592
use scs8hd_decap_8  FILLER_417_52
timestamp 1586364061
transform 1 0 5888 0 1 229024
box -38 -48 774 592
use scs8hd_fill_2  FILLER_417_48
timestamp 1586364061
transform 1 0 5520 0 1 229024
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__09__D
timestamp 1586364061
transform 1 0 5704 0 1 229024
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__09__B
timestamp 1586364061
transform 1 0 5336 0 1 229024
box -38 -48 222 592
use scs8hd_decap_12  FILLER_416_53
timestamp 1586364061
transform 1 0 5980 0 -1 229024
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_416_41
timestamp 1586364061
transform 1 0 4876 0 -1 229024
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1626
timestamp 1586364061
transform 1 0 6716 0 1 229024
box -38 -48 130 592
use scs8hd_decap_12  FILLER_416_65
timestamp 1586364061
transform 1 0 7084 0 -1 229024
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_417_60
timestamp 1586364061
transform 1 0 6624 0 1 229024
box -38 -48 130 592
use scs8hd_decap_12  FILLER_417_62
timestamp 1586364061
transform 1 0 6808 0 1 229024
box -38 -48 1142 592
use scs8hd_decap_3  PHY_833
timestamp 1586364061
transform -1 0 8832 0 -1 229024
box -38 -48 314 592
use scs8hd_decap_3  PHY_835
timestamp 1586364061
transform -1 0 8832 0 1 229024
box -38 -48 314 592
use scs8hd_decap_4  FILLER_416_77
timestamp 1586364061
transform 1 0 8188 0 -1 229024
box -38 -48 406 592
use scs8hd_decap_6  FILLER_417_74
timestamp 1586364061
transform 1 0 7912 0 1 229024
box -38 -48 590 592
use scs8hd_fill_1  FILLER_417_80
timestamp 1586364061
transform 1 0 8464 0 1 229024
box -38 -48 130 592
use scs8hd_decap_3  PHY_836
timestamp 1586364061
transform 1 0 1104 0 -1 230112
box -38 -48 314 592
use scs8hd_decap_12  FILLER_418_3
timestamp 1586364061
transform 1 0 1380 0 -1 230112
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_418_15
timestamp 1586364061
transform 1 0 2484 0 -1 230112
box -38 -48 406 592
use scs8hd_and4_4  _09_
timestamp 1586364061
transform 1 0 4048 0 -1 230112
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_1627
timestamp 1586364061
transform 1 0 3956 0 -1 230112
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__13__C
timestamp 1586364061
transform 1 0 2852 0 -1 230112
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__12__D
timestamp 1586364061
transform 1 0 3220 0 -1 230112
box -38 -48 222 592
use scs8hd_fill_2  FILLER_418_21
timestamp 1586364061
transform 1 0 3036 0 -1 230112
box -38 -48 222 592
use scs8hd_decap_6  FILLER_418_25
timestamp 1586364061
transform 1 0 3404 0 -1 230112
box -38 -48 590 592
use scs8hd_decap_12  FILLER_418_41
timestamp 1586364061
transform 1 0 4876 0 -1 230112
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_418_53
timestamp 1586364061
transform 1 0 5980 0 -1 230112
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_418_65
timestamp 1586364061
transform 1 0 7084 0 -1 230112
box -38 -48 1142 592
use scs8hd_decap_3  PHY_837
timestamp 1586364061
transform -1 0 8832 0 -1 230112
box -38 -48 314 592
use scs8hd_decap_4  FILLER_418_77
timestamp 1586364061
transform 1 0 8188 0 -1 230112
box -38 -48 406 592
use scs8hd_decap_3  PHY_838
timestamp 1586364061
transform 1 0 1104 0 1 230112
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__13__A
timestamp 1586364061
transform 1 0 2668 0 1 230112
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__13__B
timestamp 1586364061
transform 1 0 2300 0 1 230112
box -38 -48 222 592
use scs8hd_decap_8  FILLER_419_3
timestamp 1586364061
transform 1 0 1380 0 1 230112
box -38 -48 774 592
use scs8hd_fill_2  FILLER_419_11
timestamp 1586364061
transform 1 0 2116 0 1 230112
box -38 -48 222 592
use scs8hd_fill_2  FILLER_419_15
timestamp 1586364061
transform 1 0 2484 0 1 230112
box -38 -48 222 592
use scs8hd_nor4_4  _13_
timestamp 1586364061
transform 1 0 2852 0 1 230112
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4600 0 1 230112
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4968 0 1 230112
box -38 -48 222 592
use scs8hd_fill_2  FILLER_419_36
timestamp 1586364061
transform 1 0 4416 0 1 230112
box -38 -48 222 592
use scs8hd_fill_2  FILLER_419_40
timestamp 1586364061
transform 1 0 4784 0 1 230112
box -38 -48 222 592
use scs8hd_decap_12  FILLER_419_44
timestamp 1586364061
transform 1 0 5152 0 1 230112
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1628
timestamp 1586364061
transform 1 0 6716 0 1 230112
box -38 -48 130 592
use scs8hd_decap_4  FILLER_419_56
timestamp 1586364061
transform 1 0 6256 0 1 230112
box -38 -48 406 592
use scs8hd_fill_1  FILLER_419_60
timestamp 1586364061
transform 1 0 6624 0 1 230112
box -38 -48 130 592
use scs8hd_decap_12  FILLER_419_62
timestamp 1586364061
transform 1 0 6808 0 1 230112
box -38 -48 1142 592
use scs8hd_decap_3  PHY_839
timestamp 1586364061
transform -1 0 8832 0 1 230112
box -38 -48 314 592
use scs8hd_decap_6  FILLER_419_74
timestamp 1586364061
transform 1 0 7912 0 1 230112
box -38 -48 590 592
use scs8hd_fill_1  FILLER_419_80
timestamp 1586364061
transform 1 0 8464 0 1 230112
box -38 -48 130 592
use scs8hd_decap_3  PHY_840
timestamp 1586364061
transform 1 0 1104 0 -1 231200
box -38 -48 314 592
use scs8hd_decap_12  FILLER_420_3
timestamp 1586364061
transform 1 0 1380 0 -1 231200
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_420_15
timestamp 1586364061
transform 1 0 2484 0 -1 231200
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_1629
timestamp 1586364061
transform 1 0 3956 0 -1 231200
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__13__D
timestamp 1586364061
transform 1 0 2852 0 -1 231200
box -38 -48 222 592
use scs8hd_decap_8  FILLER_420_21
timestamp 1586364061
transform 1 0 3036 0 -1 231200
box -38 -48 774 592
use scs8hd_fill_2  FILLER_420_29
timestamp 1586364061
transform 1 0 3772 0 -1 231200
box -38 -48 222 592
use scs8hd_decap_4  FILLER_420_32
timestamp 1586364061
transform 1 0 4048 0 -1 231200
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4416 0 -1 231200
box -38 -48 1050 592
use scs8hd_decap_12  FILLER_420_47
timestamp 1586364061
transform 1 0 5428 0 -1 231200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_420_59
timestamp 1586364061
transform 1 0 6532 0 -1 231200
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_420_71
timestamp 1586364061
transform 1 0 7636 0 -1 231200
box -38 -48 774 592
use scs8hd_decap_3  PHY_841
timestamp 1586364061
transform -1 0 8832 0 -1 231200
box -38 -48 314 592
use scs8hd_fill_2  FILLER_420_79
timestamp 1586364061
transform 1 0 8372 0 -1 231200
box -38 -48 222 592
use scs8hd_decap_3  PHY_842
timestamp 1586364061
transform 1 0 1104 0 1 231200
box -38 -48 314 592
use scs8hd_decap_12  FILLER_421_3
timestamp 1586364061
transform 1 0 1380 0 1 231200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_421_15
timestamp 1586364061
transform 1 0 2484 0 1 231200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_421_27
timestamp 1586364061
transform 1 0 3588 0 1 231200
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_421_39
timestamp 1586364061
transform 1 0 4692 0 1 231200
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_421_51
timestamp 1586364061
transform 1 0 5796 0 1 231200
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1630
timestamp 1586364061
transform 1 0 6716 0 1 231200
box -38 -48 130 592
use scs8hd_fill_2  FILLER_421_59
timestamp 1586364061
transform 1 0 6532 0 1 231200
box -38 -48 222 592
use scs8hd_decap_12  FILLER_421_62
timestamp 1586364061
transform 1 0 6808 0 1 231200
box -38 -48 1142 592
use scs8hd_decap_3  PHY_843
timestamp 1586364061
transform -1 0 8832 0 1 231200
box -38 -48 314 592
use scs8hd_decap_6  FILLER_421_74
timestamp 1586364061
transform 1 0 7912 0 1 231200
box -38 -48 590 592
use scs8hd_fill_1  FILLER_421_80
timestamp 1586364061
transform 1 0 8464 0 1 231200
box -38 -48 130 592
use scs8hd_decap_3  PHY_844
timestamp 1586364061
transform 1 0 1104 0 -1 232288
box -38 -48 314 592
use scs8hd_decap_3  PHY_846
timestamp 1586364061
transform 1 0 1104 0 1 232288
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2668 0 1 232288
box -38 -48 222 592
use scs8hd_decap_12  FILLER_422_3
timestamp 1586364061
transform 1 0 1380 0 -1 232288
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_422_15
timestamp 1586364061
transform 1 0 2484 0 -1 232288
box -38 -48 406 592
use scs8hd_decap_12  FILLER_423_3
timestamp 1586364061
transform 1 0 1380 0 1 232288
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_423_15
timestamp 1586364061
transform 1 0 2484 0 1 232288
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 2852 0 1 232288
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_1631
timestamp 1586364061
transform 1 0 3956 0 -1 232288
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2852 0 -1 232288
box -38 -48 222 592
use scs8hd_decap_8  FILLER_422_21
timestamp 1586364061
transform 1 0 3036 0 -1 232288
box -38 -48 774 592
use scs8hd_fill_2  FILLER_422_29
timestamp 1586364061
transform 1 0 3772 0 -1 232288
box -38 -48 222 592
use scs8hd_decap_12  FILLER_422_32
timestamp 1586364061
transform 1 0 4048 0 -1 232288
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_423_30
timestamp 1586364061
transform 1 0 3864 0 1 232288
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_422_44
timestamp 1586364061
transform 1 0 5152 0 -1 232288
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_423_42
timestamp 1586364061
transform 1 0 4968 0 1 232288
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1632
timestamp 1586364061
transform 1 0 6716 0 1 232288
box -38 -48 130 592
use scs8hd_decap_12  FILLER_422_56
timestamp 1586364061
transform 1 0 6256 0 -1 232288
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_422_68
timestamp 1586364061
transform 1 0 7360 0 -1 232288
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_423_54
timestamp 1586364061
transform 1 0 6072 0 1 232288
box -38 -48 590 592
use scs8hd_fill_1  FILLER_423_60
timestamp 1586364061
transform 1 0 6624 0 1 232288
box -38 -48 130 592
use scs8hd_decap_12  FILLER_423_62
timestamp 1586364061
transform 1 0 6808 0 1 232288
box -38 -48 1142 592
use scs8hd_decap_3  PHY_845
timestamp 1586364061
transform -1 0 8832 0 -1 232288
box -38 -48 314 592
use scs8hd_decap_3  PHY_847
timestamp 1586364061
transform -1 0 8832 0 1 232288
box -38 -48 314 592
use scs8hd_fill_1  FILLER_422_80
timestamp 1586364061
transform 1 0 8464 0 -1 232288
box -38 -48 130 592
use scs8hd_decap_6  FILLER_423_74
timestamp 1586364061
transform 1 0 7912 0 1 232288
box -38 -48 590 592
use scs8hd_fill_1  FILLER_423_80
timestamp 1586364061
transform 1 0 8464 0 1 232288
box -38 -48 130 592
use scs8hd_decap_3  PHY_848
timestamp 1586364061
transform 1 0 1104 0 -1 233376
box -38 -48 314 592
use scs8hd_decap_12  FILLER_424_3
timestamp 1586364061
transform 1 0 1380 0 -1 233376
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_424_15
timestamp 1586364061
transform 1 0 2484 0 -1 233376
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1633
timestamp 1586364061
transform 1 0 3956 0 -1 233376
box -38 -48 130 592
use scs8hd_decap_4  FILLER_424_27
timestamp 1586364061
transform 1 0 3588 0 -1 233376
box -38 -48 406 592
use scs8hd_decap_4  FILLER_424_32
timestamp 1586364061
transform 1 0 4048 0 -1 233376
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 4416 0 -1 233376
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 4784 0 -1 233376
box -38 -48 222 592
use scs8hd_fill_2  FILLER_424_38
timestamp 1586364061
transform 1 0 4600 0 -1 233376
box -38 -48 222 592
use scs8hd_decap_12  FILLER_424_42
timestamp 1586364061
transform 1 0 4968 0 -1 233376
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_424_54
timestamp 1586364061
transform 1 0 6072 0 -1 233376
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_424_66
timestamp 1586364061
transform 1 0 7176 0 -1 233376
box -38 -48 1142 592
use scs8hd_decap_3  PHY_849
timestamp 1586364061
transform -1 0 8832 0 -1 233376
box -38 -48 314 592
use scs8hd_decap_3  FILLER_424_78
timestamp 1586364061
transform 1 0 8280 0 -1 233376
box -38 -48 314 592
use scs8hd_decap_3  PHY_850
timestamp 1586364061
transform 1 0 1104 0 1 233376
box -38 -48 314 592
use scs8hd_decap_12  FILLER_425_3
timestamp 1586364061
transform 1 0 1380 0 1 233376
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_425_15
timestamp 1586364061
transform 1 0 2484 0 1 233376
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4048 0 1 233376
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3680 0 1 233376
box -38 -48 222 592
use scs8hd_fill_1  FILLER_425_27
timestamp 1586364061
transform 1 0 3588 0 1 233376
box -38 -48 130 592
use scs8hd_fill_2  FILLER_425_30
timestamp 1586364061
transform 1 0 3864 0 1 233376
box -38 -48 222 592
use scs8hd_fill_2  FILLER_425_34
timestamp 1586364061
transform 1 0 4232 0 1 233376
box -38 -48 222 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 4416 0 1 233376
box -38 -48 774 592
use scs8hd_decap_12  FILLER_425_44
timestamp 1586364061
transform 1 0 5152 0 1 233376
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1634
timestamp 1586364061
transform 1 0 6716 0 1 233376
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 6992 0 1 233376
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 7360 0 1 233376
box -38 -48 222 592
use scs8hd_decap_4  FILLER_425_56
timestamp 1586364061
transform 1 0 6256 0 1 233376
box -38 -48 406 592
use scs8hd_fill_1  FILLER_425_60
timestamp 1586364061
transform 1 0 6624 0 1 233376
box -38 -48 130 592
use scs8hd_fill_2  FILLER_425_62
timestamp 1586364061
transform 1 0 6808 0 1 233376
box -38 -48 222 592
use scs8hd_fill_2  FILLER_425_66
timestamp 1586364061
transform 1 0 7176 0 1 233376
box -38 -48 222 592
use scs8hd_decap_8  FILLER_425_70
timestamp 1586364061
transform 1 0 7544 0 1 233376
box -38 -48 774 592
use scs8hd_decap_3  PHY_851
timestamp 1586364061
transform -1 0 8832 0 1 233376
box -38 -48 314 592
use scs8hd_decap_3  FILLER_425_78
timestamp 1586364061
transform 1 0 8280 0 1 233376
box -38 -48 314 592
use scs8hd_decap_3  PHY_852
timestamp 1586364061
transform 1 0 1104 0 -1 234464
box -38 -48 314 592
use scs8hd_decap_12  FILLER_426_3
timestamp 1586364061
transform 1 0 1380 0 -1 234464
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_426_15
timestamp 1586364061
transform 1 0 2484 0 -1 234464
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 234464
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_1635
timestamp 1586364061
transform 1 0 3956 0 -1 234464
box -38 -48 130 592
use scs8hd_decap_4  FILLER_426_27
timestamp 1586364061
transform 1 0 3588 0 -1 234464
box -38 -48 406 592
use scs8hd_decap_12  FILLER_426_43
timestamp 1586364061
transform 1 0 5060 0 -1 234464
box -38 -48 1142 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 6716 0 -1 234464
box -38 -48 774 592
use scs8hd_decap_6  FILLER_426_55
timestamp 1586364061
transform 1 0 6164 0 -1 234464
box -38 -48 590 592
use scs8hd_decap_12  FILLER_426_69
timestamp 1586364061
transform 1 0 7452 0 -1 234464
box -38 -48 1142 592
use scs8hd_decap_3  PHY_853
timestamp 1586364061
transform -1 0 8832 0 -1 234464
box -38 -48 314 592
use scs8hd_decap_3  PHY_854
timestamp 1586364061
transform 1 0 1104 0 1 234464
box -38 -48 314 592
use scs8hd_decap_12  FILLER_427_3
timestamp 1586364061
transform 1 0 1380 0 1 234464
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_427_15
timestamp 1586364061
transform 1 0 2484 0 1 234464
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_427_27
timestamp 1586364061
transform 1 0 3588 0 1 234464
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_427_39
timestamp 1586364061
transform 1 0 4692 0 1 234464
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_427_51
timestamp 1586364061
transform 1 0 5796 0 1 234464
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1636
timestamp 1586364061
transform 1 0 6716 0 1 234464
box -38 -48 130 592
use scs8hd_fill_2  FILLER_427_59
timestamp 1586364061
transform 1 0 6532 0 1 234464
box -38 -48 222 592
use scs8hd_decap_12  FILLER_427_62
timestamp 1586364061
transform 1 0 6808 0 1 234464
box -38 -48 1142 592
use scs8hd_decap_3  PHY_855
timestamp 1586364061
transform -1 0 8832 0 1 234464
box -38 -48 314 592
use scs8hd_decap_6  FILLER_427_74
timestamp 1586364061
transform 1 0 7912 0 1 234464
box -38 -48 590 592
use scs8hd_fill_1  FILLER_427_80
timestamp 1586364061
transform 1 0 8464 0 1 234464
box -38 -48 130 592
use scs8hd_decap_3  PHY_856
timestamp 1586364061
transform 1 0 1104 0 -1 235552
box -38 -48 314 592
use scs8hd_decap_12  FILLER_428_3
timestamp 1586364061
transform 1 0 1380 0 -1 235552
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_428_15
timestamp 1586364061
transform 1 0 2484 0 -1 235552
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1637
timestamp 1586364061
transform 1 0 3956 0 -1 235552
box -38 -48 130 592
use scs8hd_decap_4  FILLER_428_27
timestamp 1586364061
transform 1 0 3588 0 -1 235552
box -38 -48 406 592
use scs8hd_decap_12  FILLER_428_32
timestamp 1586364061
transform 1 0 4048 0 -1 235552
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_428_44
timestamp 1586364061
transform 1 0 5152 0 -1 235552
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_428_56
timestamp 1586364061
transform 1 0 6256 0 -1 235552
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_428_68
timestamp 1586364061
transform 1 0 7360 0 -1 235552
box -38 -48 1142 592
use scs8hd_decap_3  PHY_857
timestamp 1586364061
transform -1 0 8832 0 -1 235552
box -38 -48 314 592
use scs8hd_fill_1  FILLER_428_80
timestamp 1586364061
transform 1 0 8464 0 -1 235552
box -38 -48 130 592
use scs8hd_decap_3  PHY_858
timestamp 1586364061
transform 1 0 1104 0 1 235552
box -38 -48 314 592
use scs8hd_decap_3  PHY_860
timestamp 1586364061
transform 1 0 1104 0 -1 236640
box -38 -48 314 592
use scs8hd_decap_12  FILLER_429_3
timestamp 1586364061
transform 1 0 1380 0 1 235552
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_429_15
timestamp 1586364061
transform 1 0 2484 0 1 235552
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_430_3
timestamp 1586364061
transform 1 0 1380 0 -1 236640
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_430_15
timestamp 1586364061
transform 1 0 2484 0 -1 236640
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1639
timestamp 1586364061
transform 1 0 3956 0 -1 236640
box -38 -48 130 592
use scs8hd_decap_12  FILLER_429_27
timestamp 1586364061
transform 1 0 3588 0 1 235552
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_430_27
timestamp 1586364061
transform 1 0 3588 0 -1 236640
box -38 -48 406 592
use scs8hd_decap_12  FILLER_430_32
timestamp 1586364061
transform 1 0 4048 0 -1 236640
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_429_39
timestamp 1586364061
transform 1 0 4692 0 1 235552
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_429_51
timestamp 1586364061
transform 1 0 5796 0 1 235552
box -38 -48 774 592
use scs8hd_decap_12  FILLER_430_44
timestamp 1586364061
transform 1 0 5152 0 -1 236640
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1638
timestamp 1586364061
transform 1 0 6716 0 1 235552
box -38 -48 130 592
use scs8hd_fill_2  FILLER_429_59
timestamp 1586364061
transform 1 0 6532 0 1 235552
box -38 -48 222 592
use scs8hd_decap_12  FILLER_429_62
timestamp 1586364061
transform 1 0 6808 0 1 235552
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_430_56
timestamp 1586364061
transform 1 0 6256 0 -1 236640
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_430_68
timestamp 1586364061
transform 1 0 7360 0 -1 236640
box -38 -48 1142 592
use scs8hd_decap_3  PHY_859
timestamp 1586364061
transform -1 0 8832 0 1 235552
box -38 -48 314 592
use scs8hd_decap_3  PHY_861
timestamp 1586364061
transform -1 0 8832 0 -1 236640
box -38 -48 314 592
use scs8hd_decap_6  FILLER_429_74
timestamp 1586364061
transform 1 0 7912 0 1 235552
box -38 -48 590 592
use scs8hd_fill_1  FILLER_429_80
timestamp 1586364061
transform 1 0 8464 0 1 235552
box -38 -48 130 592
use scs8hd_fill_1  FILLER_430_80
timestamp 1586364061
transform 1 0 8464 0 -1 236640
box -38 -48 130 592
use scs8hd_decap_3  PHY_862
timestamp 1586364061
transform 1 0 1104 0 1 236640
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 2484 0 1 236640
box -38 -48 222 592
use scs8hd_decap_12  FILLER_431_3
timestamp 1586364061
transform 1 0 1380 0 1 236640
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_431_17
timestamp 1586364061
transform 1 0 2668 0 1 236640
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 2852 0 1 236640
box -38 -48 222 592
use scs8hd_decap_12  FILLER_431_21
timestamp 1586364061
transform 1 0 3036 0 1 236640
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_431_33
timestamp 1586364061
transform 1 0 4140 0 1 236640
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_431_45
timestamp 1586364061
transform 1 0 5244 0 1 236640
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1640
timestamp 1586364061
transform 1 0 6716 0 1 236640
box -38 -48 130 592
use scs8hd_decap_4  FILLER_431_57
timestamp 1586364061
transform 1 0 6348 0 1 236640
box -38 -48 406 592
use scs8hd_decap_12  FILLER_431_62
timestamp 1586364061
transform 1 0 6808 0 1 236640
box -38 -48 1142 592
use scs8hd_decap_3  PHY_863
timestamp 1586364061
transform -1 0 8832 0 1 236640
box -38 -48 314 592
use scs8hd_decap_6  FILLER_431_74
timestamp 1586364061
transform 1 0 7912 0 1 236640
box -38 -48 590 592
use scs8hd_fill_1  FILLER_431_80
timestamp 1586364061
transform 1 0 8464 0 1 236640
box -38 -48 130 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 2484 0 -1 237728
box -38 -48 774 592
use scs8hd_decap_3  PHY_864
timestamp 1586364061
transform 1 0 1104 0 -1 237728
box -38 -48 314 592
use scs8hd_decap_12  FILLER_432_3
timestamp 1586364061
transform 1 0 1380 0 -1 237728
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1641
timestamp 1586364061
transform 1 0 3956 0 -1 237728
box -38 -48 130 592
use scs8hd_decap_8  FILLER_432_23
timestamp 1586364061
transform 1 0 3220 0 -1 237728
box -38 -48 774 592
use scs8hd_decap_12  FILLER_432_32
timestamp 1586364061
transform 1 0 4048 0 -1 237728
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_432_44
timestamp 1586364061
transform 1 0 5152 0 -1 237728
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_432_56
timestamp 1586364061
transform 1 0 6256 0 -1 237728
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_432_68
timestamp 1586364061
transform 1 0 7360 0 -1 237728
box -38 -48 1142 592
use scs8hd_decap_3  PHY_865
timestamp 1586364061
transform -1 0 8832 0 -1 237728
box -38 -48 314 592
use scs8hd_fill_1  FILLER_432_80
timestamp 1586364061
transform 1 0 8464 0 -1 237728
box -38 -48 130 592
use scs8hd_decap_3  PHY_866
timestamp 1586364061
transform 1 0 1104 0 1 237728
box -38 -48 314 592
use scs8hd_decap_12  FILLER_433_3
timestamp 1586364061
transform 1 0 1380 0 1 237728
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_433_15
timestamp 1586364061
transform 1 0 2484 0 1 237728
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_433_27
timestamp 1586364061
transform 1 0 3588 0 1 237728
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_433_39
timestamp 1586364061
transform 1 0 4692 0 1 237728
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_433_51
timestamp 1586364061
transform 1 0 5796 0 1 237728
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1642
timestamp 1586364061
transform 1 0 6716 0 1 237728
box -38 -48 130 592
use scs8hd_fill_2  FILLER_433_59
timestamp 1586364061
transform 1 0 6532 0 1 237728
box -38 -48 222 592
use scs8hd_decap_12  FILLER_433_62
timestamp 1586364061
transform 1 0 6808 0 1 237728
box -38 -48 1142 592
use scs8hd_decap_3  PHY_867
timestamp 1586364061
transform -1 0 8832 0 1 237728
box -38 -48 314 592
use scs8hd_decap_6  FILLER_433_74
timestamp 1586364061
transform 1 0 7912 0 1 237728
box -38 -48 590 592
use scs8hd_fill_1  FILLER_433_80
timestamp 1586364061
transform 1 0 8464 0 1 237728
box -38 -48 130 592
use scs8hd_decap_3  PHY_868
timestamp 1586364061
transform 1 0 1104 0 -1 238816
box -38 -48 314 592
use scs8hd_decap_12  FILLER_434_3
timestamp 1586364061
transform 1 0 1380 0 -1 238816
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_434_15
timestamp 1586364061
transform 1 0 2484 0 -1 238816
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1643
timestamp 1586364061
transform 1 0 3956 0 -1 238816
box -38 -48 130 592
use scs8hd_decap_4  FILLER_434_27
timestamp 1586364061
transform 1 0 3588 0 -1 238816
box -38 -48 406 592
use scs8hd_decap_12  FILLER_434_32
timestamp 1586364061
transform 1 0 4048 0 -1 238816
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_434_44
timestamp 1586364061
transform 1 0 5152 0 -1 238816
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_434_56
timestamp 1586364061
transform 1 0 6256 0 -1 238816
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_434_68
timestamp 1586364061
transform 1 0 7360 0 -1 238816
box -38 -48 1142 592
use scs8hd_decap_3  PHY_869
timestamp 1586364061
transform -1 0 8832 0 -1 238816
box -38 -48 314 592
use scs8hd_fill_1  FILLER_434_80
timestamp 1586364061
transform 1 0 8464 0 -1 238816
box -38 -48 130 592
use scs8hd_decap_3  PHY_870
timestamp 1586364061
transform 1 0 1104 0 1 238816
box -38 -48 314 592
use scs8hd_decap_12  FILLER_435_3
timestamp 1586364061
transform 1 0 1380 0 1 238816
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_435_15
timestamp 1586364061
transform 1 0 2484 0 1 238816
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_435_27
timestamp 1586364061
transform 1 0 3588 0 1 238816
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_435_39
timestamp 1586364061
transform 1 0 4692 0 1 238816
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_435_51
timestamp 1586364061
transform 1 0 5796 0 1 238816
box -38 -48 774 592
use scs8hd_buf_2  _21_
timestamp 1586364061
transform 1 0 6808 0 1 238816
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_1644
timestamp 1586364061
transform 1 0 6716 0 1 238816
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__21__A
timestamp 1586364061
transform 1 0 7360 0 1 238816
box -38 -48 222 592
use scs8hd_fill_2  FILLER_435_59
timestamp 1586364061
transform 1 0 6532 0 1 238816
box -38 -48 222 592
use scs8hd_fill_2  FILLER_435_66
timestamp 1586364061
transform 1 0 7176 0 1 238816
box -38 -48 222 592
use scs8hd_decap_8  FILLER_435_70
timestamp 1586364061
transform 1 0 7544 0 1 238816
box -38 -48 774 592
use scs8hd_decap_3  PHY_871
timestamp 1586364061
transform -1 0 8832 0 1 238816
box -38 -48 314 592
use scs8hd_decap_3  FILLER_435_78
timestamp 1586364061
transform 1 0 8280 0 1 238816
box -38 -48 314 592
use scs8hd_decap_3  PHY_872
timestamp 1586364061
transform 1 0 1104 0 -1 239904
box -38 -48 314 592
use scs8hd_decap_3  PHY_874
timestamp 1586364061
transform 1 0 1104 0 1 239904
box -38 -48 314 592
use scs8hd_decap_12  FILLER_436_3
timestamp 1586364061
transform 1 0 1380 0 -1 239904
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_436_15
timestamp 1586364061
transform 1 0 2484 0 -1 239904
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_437_3
timestamp 1586364061
transform 1 0 1380 0 1 239904
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_437_15
timestamp 1586364061
transform 1 0 2484 0 1 239904
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1645
timestamp 1586364061
transform 1 0 3956 0 -1 239904
box -38 -48 130 592
use scs8hd_decap_4  FILLER_436_27
timestamp 1586364061
transform 1 0 3588 0 -1 239904
box -38 -48 406 592
use scs8hd_decap_12  FILLER_436_32
timestamp 1586364061
transform 1 0 4048 0 -1 239904
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_437_27
timestamp 1586364061
transform 1 0 3588 0 1 239904
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_436_44
timestamp 1586364061
transform 1 0 5152 0 -1 239904
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_437_39
timestamp 1586364061
transform 1 0 4692 0 1 239904
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_437_51
timestamp 1586364061
transform 1 0 5796 0 1 239904
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1646
timestamp 1586364061
transform 1 0 6716 0 1 239904
box -38 -48 130 592
use scs8hd_decap_12  FILLER_436_56
timestamp 1586364061
transform 1 0 6256 0 -1 239904
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_436_68
timestamp 1586364061
transform 1 0 7360 0 -1 239904
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_437_59
timestamp 1586364061
transform 1 0 6532 0 1 239904
box -38 -48 222 592
use scs8hd_decap_12  FILLER_437_62
timestamp 1586364061
transform 1 0 6808 0 1 239904
box -38 -48 1142 592
use scs8hd_decap_3  PHY_873
timestamp 1586364061
transform -1 0 8832 0 -1 239904
box -38 -48 314 592
use scs8hd_decap_3  PHY_875
timestamp 1586364061
transform -1 0 8832 0 1 239904
box -38 -48 314 592
use scs8hd_fill_1  FILLER_436_80
timestamp 1586364061
transform 1 0 8464 0 -1 239904
box -38 -48 130 592
use scs8hd_decap_6  FILLER_437_74
timestamp 1586364061
transform 1 0 7912 0 1 239904
box -38 -48 590 592
use scs8hd_fill_1  FILLER_437_80
timestamp 1586364061
transform 1 0 8464 0 1 239904
box -38 -48 130 592
use scs8hd_decap_3  PHY_876
timestamp 1586364061
transform 1 0 1104 0 -1 240992
box -38 -48 314 592
use scs8hd_decap_12  FILLER_438_3
timestamp 1586364061
transform 1 0 1380 0 -1 240992
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_438_15
timestamp 1586364061
transform 1 0 2484 0 -1 240992
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1647
timestamp 1586364061
transform 1 0 3956 0 -1 240992
box -38 -48 130 592
use scs8hd_decap_4  FILLER_438_27
timestamp 1586364061
transform 1 0 3588 0 -1 240992
box -38 -48 406 592
use scs8hd_decap_12  FILLER_438_32
timestamp 1586364061
transform 1 0 4048 0 -1 240992
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_438_44
timestamp 1586364061
transform 1 0 5152 0 -1 240992
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_438_56
timestamp 1586364061
transform 1 0 6256 0 -1 240992
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_438_68
timestamp 1586364061
transform 1 0 7360 0 -1 240992
box -38 -48 1142 592
use scs8hd_decap_3  PHY_877
timestamp 1586364061
transform -1 0 8832 0 -1 240992
box -38 -48 314 592
use scs8hd_fill_1  FILLER_438_80
timestamp 1586364061
transform 1 0 8464 0 -1 240992
box -38 -48 130 592
use scs8hd_decap_3  PHY_878
timestamp 1586364061
transform 1 0 1104 0 1 240992
box -38 -48 314 592
use scs8hd_decap_12  FILLER_439_3
timestamp 1586364061
transform 1 0 1380 0 1 240992
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_439_15
timestamp 1586364061
transform 1 0 2484 0 1 240992
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_439_27
timestamp 1586364061
transform 1 0 3588 0 1 240992
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_439_39
timestamp 1586364061
transform 1 0 4692 0 1 240992
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_439_51
timestamp 1586364061
transform 1 0 5796 0 1 240992
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1648
timestamp 1586364061
transform 1 0 6716 0 1 240992
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__22__A
timestamp 1586364061
transform 1 0 7452 0 1 240992
box -38 -48 222 592
use scs8hd_fill_2  FILLER_439_59
timestamp 1586364061
transform 1 0 6532 0 1 240992
box -38 -48 222 592
use scs8hd_decap_6  FILLER_439_62
timestamp 1586364061
transform 1 0 6808 0 1 240992
box -38 -48 590 592
use scs8hd_fill_1  FILLER_439_68
timestamp 1586364061
transform 1 0 7360 0 1 240992
box -38 -48 130 592
use scs8hd_decap_8  FILLER_439_71
timestamp 1586364061
transform 1 0 7636 0 1 240992
box -38 -48 774 592
use scs8hd_decap_3  PHY_879
timestamp 1586364061
transform -1 0 8832 0 1 240992
box -38 -48 314 592
use scs8hd_fill_2  FILLER_439_79
timestamp 1586364061
transform 1 0 8372 0 1 240992
box -38 -48 222 592
use scs8hd_decap_3  PHY_880
timestamp 1586364061
transform 1 0 1104 0 -1 242080
box -38 -48 314 592
use scs8hd_decap_12  FILLER_440_3
timestamp 1586364061
transform 1 0 1380 0 -1 242080
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_440_15
timestamp 1586364061
transform 1 0 2484 0 -1 242080
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1649
timestamp 1586364061
transform 1 0 3956 0 -1 242080
box -38 -48 130 592
use scs8hd_decap_4  FILLER_440_27
timestamp 1586364061
transform 1 0 3588 0 -1 242080
box -38 -48 406 592
use scs8hd_decap_12  FILLER_440_32
timestamp 1586364061
transform 1 0 4048 0 -1 242080
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_440_44
timestamp 1586364061
transform 1 0 5152 0 -1 242080
box -38 -48 1142 592
use scs8hd_buf_2  _22_
timestamp 1586364061
transform 1 0 7452 0 -1 242080
box -38 -48 406 592
use scs8hd_decap_12  FILLER_440_56
timestamp 1586364061
transform 1 0 6256 0 -1 242080
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_440_68
timestamp 1586364061
transform 1 0 7360 0 -1 242080
box -38 -48 130 592
use scs8hd_decap_3  PHY_881
timestamp 1586364061
transform -1 0 8832 0 -1 242080
box -38 -48 314 592
use scs8hd_decap_8  FILLER_440_73
timestamp 1586364061
transform 1 0 7820 0 -1 242080
box -38 -48 774 592
use scs8hd_decap_3  PHY_882
timestamp 1586364061
transform 1 0 1104 0 1 242080
box -38 -48 314 592
use scs8hd_decap_12  FILLER_441_3
timestamp 1586364061
transform 1 0 1380 0 1 242080
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_441_15
timestamp 1586364061
transform 1 0 2484 0 1 242080
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_441_27
timestamp 1586364061
transform 1 0 3588 0 1 242080
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_441_39
timestamp 1586364061
transform 1 0 4692 0 1 242080
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_441_51
timestamp 1586364061
transform 1 0 5796 0 1 242080
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1650
timestamp 1586364061
transform 1 0 6716 0 1 242080
box -38 -48 130 592
use scs8hd_fill_2  FILLER_441_59
timestamp 1586364061
transform 1 0 6532 0 1 242080
box -38 -48 222 592
use scs8hd_decap_12  FILLER_441_62
timestamp 1586364061
transform 1 0 6808 0 1 242080
box -38 -48 1142 592
use scs8hd_decap_3  PHY_883
timestamp 1586364061
transform -1 0 8832 0 1 242080
box -38 -48 314 592
use scs8hd_decap_6  FILLER_441_74
timestamp 1586364061
transform 1 0 7912 0 1 242080
box -38 -48 590 592
use scs8hd_fill_1  FILLER_441_80
timestamp 1586364061
transform 1 0 8464 0 1 242080
box -38 -48 130 592
use scs8hd_decap_3  PHY_884
timestamp 1586364061
transform 1 0 1104 0 -1 243168
box -38 -48 314 592
use scs8hd_decap_3  PHY_886
timestamp 1586364061
transform 1 0 1104 0 1 243168
box -38 -48 314 592
use scs8hd_decap_12  FILLER_442_3
timestamp 1586364061
transform 1 0 1380 0 -1 243168
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_442_15
timestamp 1586364061
transform 1 0 2484 0 -1 243168
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_443_3
timestamp 1586364061
transform 1 0 1380 0 1 243168
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_443_15
timestamp 1586364061
transform 1 0 2484 0 1 243168
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1651
timestamp 1586364061
transform 1 0 3956 0 -1 243168
box -38 -48 130 592
use scs8hd_decap_4  FILLER_442_27
timestamp 1586364061
transform 1 0 3588 0 -1 243168
box -38 -48 406 592
use scs8hd_decap_12  FILLER_442_32
timestamp 1586364061
transform 1 0 4048 0 -1 243168
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_443_27
timestamp 1586364061
transform 1 0 3588 0 1 243168
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_442_44
timestamp 1586364061
transform 1 0 5152 0 -1 243168
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_443_39
timestamp 1586364061
transform 1 0 4692 0 1 243168
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_443_51
timestamp 1586364061
transform 1 0 5796 0 1 243168
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1652
timestamp 1586364061
transform 1 0 6716 0 1 243168
box -38 -48 130 592
use scs8hd_decap_12  FILLER_442_56
timestamp 1586364061
transform 1 0 6256 0 -1 243168
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_442_68
timestamp 1586364061
transform 1 0 7360 0 -1 243168
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_443_59
timestamp 1586364061
transform 1 0 6532 0 1 243168
box -38 -48 222 592
use scs8hd_decap_12  FILLER_443_62
timestamp 1586364061
transform 1 0 6808 0 1 243168
box -38 -48 1142 592
use scs8hd_decap_3  PHY_885
timestamp 1586364061
transform -1 0 8832 0 -1 243168
box -38 -48 314 592
use scs8hd_decap_3  PHY_887
timestamp 1586364061
transform -1 0 8832 0 1 243168
box -38 -48 314 592
use scs8hd_fill_1  FILLER_442_80
timestamp 1586364061
transform 1 0 8464 0 -1 243168
box -38 -48 130 592
use scs8hd_decap_6  FILLER_443_74
timestamp 1586364061
transform 1 0 7912 0 1 243168
box -38 -48 590 592
use scs8hd_fill_1  FILLER_443_80
timestamp 1586364061
transform 1 0 8464 0 1 243168
box -38 -48 130 592
use scs8hd_decap_3  PHY_888
timestamp 1586364061
transform 1 0 1104 0 -1 244256
box -38 -48 314 592
use scs8hd_decap_12  FILLER_444_3
timestamp 1586364061
transform 1 0 1380 0 -1 244256
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_444_15
timestamp 1586364061
transform 1 0 2484 0 -1 244256
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1653
timestamp 1586364061
transform 1 0 3956 0 -1 244256
box -38 -48 130 592
use scs8hd_decap_4  FILLER_444_27
timestamp 1586364061
transform 1 0 3588 0 -1 244256
box -38 -48 406 592
use scs8hd_decap_12  FILLER_444_32
timestamp 1586364061
transform 1 0 4048 0 -1 244256
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_444_44
timestamp 1586364061
transform 1 0 5152 0 -1 244256
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_444_56
timestamp 1586364061
transform 1 0 6256 0 -1 244256
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_444_68
timestamp 1586364061
transform 1 0 7360 0 -1 244256
box -38 -48 1142 592
use scs8hd_decap_3  PHY_889
timestamp 1586364061
transform -1 0 8832 0 -1 244256
box -38 -48 314 592
use scs8hd_fill_1  FILLER_444_80
timestamp 1586364061
transform 1 0 8464 0 -1 244256
box -38 -48 130 592
use scs8hd_buf_2  _18_
timestamp 1586364061
transform 1 0 2024 0 1 244256
box -38 -48 406 592
use scs8hd_decap_3  PHY_890
timestamp 1586364061
transform 1 0 1104 0 1 244256
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__18__A
timestamp 1586364061
transform 1 0 2576 0 1 244256
box -38 -48 222 592
use scs8hd_decap_6  FILLER_445_3
timestamp 1586364061
transform 1 0 1380 0 1 244256
box -38 -48 590 592
use scs8hd_fill_1  FILLER_445_9
timestamp 1586364061
transform 1 0 1932 0 1 244256
box -38 -48 130 592
use scs8hd_fill_2  FILLER_445_14
timestamp 1586364061
transform 1 0 2392 0 1 244256
box -38 -48 222 592
use scs8hd_decap_12  FILLER_445_18
timestamp 1586364061
transform 1 0 2760 0 1 244256
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_445_30
timestamp 1586364061
transform 1 0 3864 0 1 244256
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_445_42
timestamp 1586364061
transform 1 0 4968 0 1 244256
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1654
timestamp 1586364061
transform 1 0 6716 0 1 244256
box -38 -48 130 592
use scs8hd_decap_6  FILLER_445_54
timestamp 1586364061
transform 1 0 6072 0 1 244256
box -38 -48 590 592
use scs8hd_fill_1  FILLER_445_60
timestamp 1586364061
transform 1 0 6624 0 1 244256
box -38 -48 130 592
use scs8hd_decap_12  FILLER_445_62
timestamp 1586364061
transform 1 0 6808 0 1 244256
box -38 -48 1142 592
use scs8hd_decap_3  PHY_891
timestamp 1586364061
transform -1 0 8832 0 1 244256
box -38 -48 314 592
use scs8hd_decap_6  FILLER_445_74
timestamp 1586364061
transform 1 0 7912 0 1 244256
box -38 -48 590 592
use scs8hd_fill_1  FILLER_445_80
timestamp 1586364061
transform 1 0 8464 0 1 244256
box -38 -48 130 592
use scs8hd_decap_3  PHY_892
timestamp 1586364061
transform 1 0 1104 0 -1 245344
box -38 -48 314 592
use scs8hd_decap_12  FILLER_446_3
timestamp 1586364061
transform 1 0 1380 0 -1 245344
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_446_15
timestamp 1586364061
transform 1 0 2484 0 -1 245344
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1655
timestamp 1586364061
transform 1 0 3956 0 -1 245344
box -38 -48 130 592
use scs8hd_decap_4  FILLER_446_27
timestamp 1586364061
transform 1 0 3588 0 -1 245344
box -38 -48 406 592
use scs8hd_decap_12  FILLER_446_32
timestamp 1586364061
transform 1 0 4048 0 -1 245344
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_446_44
timestamp 1586364061
transform 1 0 5152 0 -1 245344
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_446_56
timestamp 1586364061
transform 1 0 6256 0 -1 245344
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_446_68
timestamp 1586364061
transform 1 0 7360 0 -1 245344
box -38 -48 1142 592
use scs8hd_decap_3  PHY_893
timestamp 1586364061
transform -1 0 8832 0 -1 245344
box -38 -48 314 592
use scs8hd_fill_1  FILLER_446_80
timestamp 1586364061
transform 1 0 8464 0 -1 245344
box -38 -48 130 592
use scs8hd_decap_3  PHY_894
timestamp 1586364061
transform 1 0 1104 0 1 245344
box -38 -48 314 592
use scs8hd_decap_12  FILLER_447_3
timestamp 1586364061
transform 1 0 1380 0 1 245344
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_447_15
timestamp 1586364061
transform 1 0 2484 0 1 245344
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_447_27
timestamp 1586364061
transform 1 0 3588 0 1 245344
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_447_39
timestamp 1586364061
transform 1 0 4692 0 1 245344
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_447_51
timestamp 1586364061
transform 1 0 5796 0 1 245344
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1656
timestamp 1586364061
transform 1 0 6716 0 1 245344
box -38 -48 130 592
use scs8hd_fill_2  FILLER_447_59
timestamp 1586364061
transform 1 0 6532 0 1 245344
box -38 -48 222 592
use scs8hd_decap_12  FILLER_447_62
timestamp 1586364061
transform 1 0 6808 0 1 245344
box -38 -48 1142 592
use scs8hd_decap_3  PHY_895
timestamp 1586364061
transform -1 0 8832 0 1 245344
box -38 -48 314 592
use scs8hd_decap_6  FILLER_447_74
timestamp 1586364061
transform 1 0 7912 0 1 245344
box -38 -48 590 592
use scs8hd_fill_1  FILLER_447_80
timestamp 1586364061
transform 1 0 8464 0 1 245344
box -38 -48 130 592
use scs8hd_decap_3  PHY_896
timestamp 1586364061
transform 1 0 1104 0 -1 246432
box -38 -48 314 592
use scs8hd_decap_12  FILLER_448_3
timestamp 1586364061
transform 1 0 1380 0 -1 246432
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_448_15
timestamp 1586364061
transform 1 0 2484 0 -1 246432
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1657
timestamp 1586364061
transform 1 0 3956 0 -1 246432
box -38 -48 130 592
use scs8hd_decap_4  FILLER_448_27
timestamp 1586364061
transform 1 0 3588 0 -1 246432
box -38 -48 406 592
use scs8hd_decap_12  FILLER_448_32
timestamp 1586364061
transform 1 0 4048 0 -1 246432
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_448_44
timestamp 1586364061
transform 1 0 5152 0 -1 246432
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_448_56
timestamp 1586364061
transform 1 0 6256 0 -1 246432
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_448_68
timestamp 1586364061
transform 1 0 7360 0 -1 246432
box -38 -48 1142 592
use scs8hd_decap_3  PHY_897
timestamp 1586364061
transform -1 0 8832 0 -1 246432
box -38 -48 314 592
use scs8hd_fill_1  FILLER_448_80
timestamp 1586364061
transform 1 0 8464 0 -1 246432
box -38 -48 130 592
use scs8hd_decap_3  PHY_898
timestamp 1586364061
transform 1 0 1104 0 1 246432
box -38 -48 314 592
use scs8hd_decap_3  PHY_900
timestamp 1586364061
transform 1 0 1104 0 -1 247520
box -38 -48 314 592
use scs8hd_decap_12  FILLER_449_3
timestamp 1586364061
transform 1 0 1380 0 1 246432
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_449_15
timestamp 1586364061
transform 1 0 2484 0 1 246432
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_450_3
timestamp 1586364061
transform 1 0 1380 0 -1 247520
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_450_15
timestamp 1586364061
transform 1 0 2484 0 -1 247520
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1659
timestamp 1586364061
transform 1 0 3956 0 -1 247520
box -38 -48 130 592
use scs8hd_decap_12  FILLER_449_27
timestamp 1586364061
transform 1 0 3588 0 1 246432
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_450_27
timestamp 1586364061
transform 1 0 3588 0 -1 247520
box -38 -48 406 592
use scs8hd_decap_12  FILLER_450_32
timestamp 1586364061
transform 1 0 4048 0 -1 247520
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_449_39
timestamp 1586364061
transform 1 0 4692 0 1 246432
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_449_51
timestamp 1586364061
transform 1 0 5796 0 1 246432
box -38 -48 774 592
use scs8hd_decap_12  FILLER_450_44
timestamp 1586364061
transform 1 0 5152 0 -1 247520
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1658
timestamp 1586364061
transform 1 0 6716 0 1 246432
box -38 -48 130 592
use scs8hd_fill_2  FILLER_449_59
timestamp 1586364061
transform 1 0 6532 0 1 246432
box -38 -48 222 592
use scs8hd_decap_12  FILLER_449_62
timestamp 1586364061
transform 1 0 6808 0 1 246432
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_450_56
timestamp 1586364061
transform 1 0 6256 0 -1 247520
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_450_68
timestamp 1586364061
transform 1 0 7360 0 -1 247520
box -38 -48 1142 592
use scs8hd_decap_3  PHY_899
timestamp 1586364061
transform -1 0 8832 0 1 246432
box -38 -48 314 592
use scs8hd_decap_3  PHY_901
timestamp 1586364061
transform -1 0 8832 0 -1 247520
box -38 -48 314 592
use scs8hd_decap_6  FILLER_449_74
timestamp 1586364061
transform 1 0 7912 0 1 246432
box -38 -48 590 592
use scs8hd_fill_1  FILLER_449_80
timestamp 1586364061
transform 1 0 8464 0 1 246432
box -38 -48 130 592
use scs8hd_fill_1  FILLER_450_80
timestamp 1586364061
transform 1 0 8464 0 -1 247520
box -38 -48 130 592
use scs8hd_decap_3  PHY_902
timestamp 1586364061
transform 1 0 1104 0 1 247520
box -38 -48 314 592
use scs8hd_decap_12  FILLER_451_3
timestamp 1586364061
transform 1 0 1380 0 1 247520
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_451_15
timestamp 1586364061
transform 1 0 2484 0 1 247520
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_451_27
timestamp 1586364061
transform 1 0 3588 0 1 247520
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_451_39
timestamp 1586364061
transform 1 0 4692 0 1 247520
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_451_51
timestamp 1586364061
transform 1 0 5796 0 1 247520
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1660
timestamp 1586364061
transform 1 0 6716 0 1 247520
box -38 -48 130 592
use scs8hd_fill_2  FILLER_451_59
timestamp 1586364061
transform 1 0 6532 0 1 247520
box -38 -48 222 592
use scs8hd_decap_12  FILLER_451_62
timestamp 1586364061
transform 1 0 6808 0 1 247520
box -38 -48 1142 592
use scs8hd_decap_3  PHY_903
timestamp 1586364061
transform -1 0 8832 0 1 247520
box -38 -48 314 592
use scs8hd_decap_6  FILLER_451_74
timestamp 1586364061
transform 1 0 7912 0 1 247520
box -38 -48 590 592
use scs8hd_fill_1  FILLER_451_80
timestamp 1586364061
transform 1 0 8464 0 1 247520
box -38 -48 130 592
use scs8hd_decap_3  PHY_904
timestamp 1586364061
transform 1 0 1104 0 -1 248608
box -38 -48 314 592
use scs8hd_decap_12  FILLER_452_3
timestamp 1586364061
transform 1 0 1380 0 -1 248608
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_452_15
timestamp 1586364061
transform 1 0 2484 0 -1 248608
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1661
timestamp 1586364061
transform 1 0 3956 0 -1 248608
box -38 -48 130 592
use scs8hd_decap_4  FILLER_452_27
timestamp 1586364061
transform 1 0 3588 0 -1 248608
box -38 -48 406 592
use scs8hd_decap_12  FILLER_452_32
timestamp 1586364061
transform 1 0 4048 0 -1 248608
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_452_44
timestamp 1586364061
transform 1 0 5152 0 -1 248608
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_452_56
timestamp 1586364061
transform 1 0 6256 0 -1 248608
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_452_68
timestamp 1586364061
transform 1 0 7360 0 -1 248608
box -38 -48 1142 592
use scs8hd_decap_3  PHY_905
timestamp 1586364061
transform -1 0 8832 0 -1 248608
box -38 -48 314 592
use scs8hd_fill_1  FILLER_452_80
timestamp 1586364061
transform 1 0 8464 0 -1 248608
box -38 -48 130 592
use scs8hd_decap_3  PHY_906
timestamp 1586364061
transform 1 0 1104 0 1 248608
box -38 -48 314 592
use scs8hd_decap_12  FILLER_453_3
timestamp 1586364061
transform 1 0 1380 0 1 248608
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_453_15
timestamp 1586364061
transform 1 0 2484 0 1 248608
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_453_27
timestamp 1586364061
transform 1 0 3588 0 1 248608
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_453_39
timestamp 1586364061
transform 1 0 4692 0 1 248608
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_453_51
timestamp 1586364061
transform 1 0 5796 0 1 248608
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1662
timestamp 1586364061
transform 1 0 6716 0 1 248608
box -38 -48 130 592
use scs8hd_fill_2  FILLER_453_59
timestamp 1586364061
transform 1 0 6532 0 1 248608
box -38 -48 222 592
use scs8hd_decap_12  FILLER_453_62
timestamp 1586364061
transform 1 0 6808 0 1 248608
box -38 -48 1142 592
use scs8hd_decap_3  PHY_907
timestamp 1586364061
transform -1 0 8832 0 1 248608
box -38 -48 314 592
use scs8hd_decap_6  FILLER_453_74
timestamp 1586364061
transform 1 0 7912 0 1 248608
box -38 -48 590 592
use scs8hd_fill_1  FILLER_453_80
timestamp 1586364061
transform 1 0 8464 0 1 248608
box -38 -48 130 592
use scs8hd_decap_3  PHY_908
timestamp 1586364061
transform 1 0 1104 0 -1 249696
box -38 -48 314 592
use scs8hd_decap_12  FILLER_454_3
timestamp 1586364061
transform 1 0 1380 0 -1 249696
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_454_15
timestamp 1586364061
transform 1 0 2484 0 -1 249696
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1663
timestamp 1586364061
transform 1 0 3956 0 -1 249696
box -38 -48 130 592
use scs8hd_decap_4  FILLER_454_27
timestamp 1586364061
transform 1 0 3588 0 -1 249696
box -38 -48 406 592
use scs8hd_decap_12  FILLER_454_32
timestamp 1586364061
transform 1 0 4048 0 -1 249696
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_454_44
timestamp 1586364061
transform 1 0 5152 0 -1 249696
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_454_56
timestamp 1586364061
transform 1 0 6256 0 -1 249696
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_454_68
timestamp 1586364061
transform 1 0 7360 0 -1 249696
box -38 -48 1142 592
use scs8hd_decap_3  PHY_909
timestamp 1586364061
transform -1 0 8832 0 -1 249696
box -38 -48 314 592
use scs8hd_fill_1  FILLER_454_80
timestamp 1586364061
transform 1 0 8464 0 -1 249696
box -38 -48 130 592
use scs8hd_decap_3  PHY_910
timestamp 1586364061
transform 1 0 1104 0 1 249696
box -38 -48 314 592
use scs8hd_decap_3  PHY_912
timestamp 1586364061
transform 1 0 1104 0 -1 250784
box -38 -48 314 592
use scs8hd_decap_12  FILLER_455_3
timestamp 1586364061
transform 1 0 1380 0 1 249696
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_455_15
timestamp 1586364061
transform 1 0 2484 0 1 249696
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_456_3
timestamp 1586364061
transform 1 0 1380 0 -1 250784
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_456_15
timestamp 1586364061
transform 1 0 2484 0 -1 250784
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1665
timestamp 1586364061
transform 1 0 3956 0 -1 250784
box -38 -48 130 592
use scs8hd_decap_12  FILLER_455_27
timestamp 1586364061
transform 1 0 3588 0 1 249696
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_456_27
timestamp 1586364061
transform 1 0 3588 0 -1 250784
box -38 -48 406 592
use scs8hd_decap_12  FILLER_456_32
timestamp 1586364061
transform 1 0 4048 0 -1 250784
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_455_39
timestamp 1586364061
transform 1 0 4692 0 1 249696
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_455_51
timestamp 1586364061
transform 1 0 5796 0 1 249696
box -38 -48 774 592
use scs8hd_decap_12  FILLER_456_44
timestamp 1586364061
transform 1 0 5152 0 -1 250784
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1664
timestamp 1586364061
transform 1 0 6716 0 1 249696
box -38 -48 130 592
use scs8hd_fill_2  FILLER_455_59
timestamp 1586364061
transform 1 0 6532 0 1 249696
box -38 -48 222 592
use scs8hd_decap_12  FILLER_455_62
timestamp 1586364061
transform 1 0 6808 0 1 249696
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_456_56
timestamp 1586364061
transform 1 0 6256 0 -1 250784
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_456_68
timestamp 1586364061
transform 1 0 7360 0 -1 250784
box -38 -48 1142 592
use scs8hd_decap_3  PHY_911
timestamp 1586364061
transform -1 0 8832 0 1 249696
box -38 -48 314 592
use scs8hd_decap_3  PHY_913
timestamp 1586364061
transform -1 0 8832 0 -1 250784
box -38 -48 314 592
use scs8hd_decap_6  FILLER_455_74
timestamp 1586364061
transform 1 0 7912 0 1 249696
box -38 -48 590 592
use scs8hd_fill_1  FILLER_455_80
timestamp 1586364061
transform 1 0 8464 0 1 249696
box -38 -48 130 592
use scs8hd_fill_1  FILLER_456_80
timestamp 1586364061
transform 1 0 8464 0 -1 250784
box -38 -48 130 592
use scs8hd_decap_3  PHY_914
timestamp 1586364061
transform 1 0 1104 0 1 250784
box -38 -48 314 592
use scs8hd_decap_12  FILLER_457_3
timestamp 1586364061
transform 1 0 1380 0 1 250784
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_457_15
timestamp 1586364061
transform 1 0 2484 0 1 250784
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_457_27
timestamp 1586364061
transform 1 0 3588 0 1 250784
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_457_39
timestamp 1586364061
transform 1 0 4692 0 1 250784
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_457_51
timestamp 1586364061
transform 1 0 5796 0 1 250784
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1666
timestamp 1586364061
transform 1 0 6716 0 1 250784
box -38 -48 130 592
use scs8hd_fill_2  FILLER_457_59
timestamp 1586364061
transform 1 0 6532 0 1 250784
box -38 -48 222 592
use scs8hd_decap_12  FILLER_457_62
timestamp 1586364061
transform 1 0 6808 0 1 250784
box -38 -48 1142 592
use scs8hd_decap_3  PHY_915
timestamp 1586364061
transform -1 0 8832 0 1 250784
box -38 -48 314 592
use scs8hd_decap_6  FILLER_457_74
timestamp 1586364061
transform 1 0 7912 0 1 250784
box -38 -48 590 592
use scs8hd_fill_1  FILLER_457_80
timestamp 1586364061
transform 1 0 8464 0 1 250784
box -38 -48 130 592
use scs8hd_decap_3  PHY_916
timestamp 1586364061
transform 1 0 1104 0 -1 251872
box -38 -48 314 592
use scs8hd_decap_12  FILLER_458_3
timestamp 1586364061
transform 1 0 1380 0 -1 251872
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_458_15
timestamp 1586364061
transform 1 0 2484 0 -1 251872
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1667
timestamp 1586364061
transform 1 0 3956 0 -1 251872
box -38 -48 130 592
use scs8hd_decap_4  FILLER_458_27
timestamp 1586364061
transform 1 0 3588 0 -1 251872
box -38 -48 406 592
use scs8hd_decap_12  FILLER_458_32
timestamp 1586364061
transform 1 0 4048 0 -1 251872
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_458_44
timestamp 1586364061
transform 1 0 5152 0 -1 251872
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_458_56
timestamp 1586364061
transform 1 0 6256 0 -1 251872
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_458_68
timestamp 1586364061
transform 1 0 7360 0 -1 251872
box -38 -48 1142 592
use scs8hd_decap_3  PHY_917
timestamp 1586364061
transform -1 0 8832 0 -1 251872
box -38 -48 314 592
use scs8hd_fill_1  FILLER_458_80
timestamp 1586364061
transform 1 0 8464 0 -1 251872
box -38 -48 130 592
use scs8hd_decap_3  PHY_918
timestamp 1586364061
transform 1 0 1104 0 1 251872
box -38 -48 314 592
use scs8hd_decap_12  FILLER_459_3
timestamp 1586364061
transform 1 0 1380 0 1 251872
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_459_15
timestamp 1586364061
transform 1 0 2484 0 1 251872
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_459_27
timestamp 1586364061
transform 1 0 3588 0 1 251872
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_459_39
timestamp 1586364061
transform 1 0 4692 0 1 251872
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_459_51
timestamp 1586364061
transform 1 0 5796 0 1 251872
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1668
timestamp 1586364061
transform 1 0 6716 0 1 251872
box -38 -48 130 592
use scs8hd_fill_2  FILLER_459_59
timestamp 1586364061
transform 1 0 6532 0 1 251872
box -38 -48 222 592
use scs8hd_decap_12  FILLER_459_62
timestamp 1586364061
transform 1 0 6808 0 1 251872
box -38 -48 1142 592
use scs8hd_decap_3  PHY_919
timestamp 1586364061
transform -1 0 8832 0 1 251872
box -38 -48 314 592
use scs8hd_decap_6  FILLER_459_74
timestamp 1586364061
transform 1 0 7912 0 1 251872
box -38 -48 590 592
use scs8hd_fill_1  FILLER_459_80
timestamp 1586364061
transform 1 0 8464 0 1 251872
box -38 -48 130 592
use scs8hd_decap_3  PHY_920
timestamp 1586364061
transform 1 0 1104 0 -1 252960
box -38 -48 314 592
use scs8hd_decap_12  FILLER_460_3
timestamp 1586364061
transform 1 0 1380 0 -1 252960
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_460_15
timestamp 1586364061
transform 1 0 2484 0 -1 252960
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1669
timestamp 1586364061
transform 1 0 3956 0 -1 252960
box -38 -48 130 592
use scs8hd_decap_4  FILLER_460_27
timestamp 1586364061
transform 1 0 3588 0 -1 252960
box -38 -48 406 592
use scs8hd_decap_12  FILLER_460_32
timestamp 1586364061
transform 1 0 4048 0 -1 252960
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_460_44
timestamp 1586364061
transform 1 0 5152 0 -1 252960
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_460_56
timestamp 1586364061
transform 1 0 6256 0 -1 252960
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_460_68
timestamp 1586364061
transform 1 0 7360 0 -1 252960
box -38 -48 1142 592
use scs8hd_decap_3  PHY_921
timestamp 1586364061
transform -1 0 8832 0 -1 252960
box -38 -48 314 592
use scs8hd_fill_1  FILLER_460_80
timestamp 1586364061
transform 1 0 8464 0 -1 252960
box -38 -48 130 592
use scs8hd_decap_3  PHY_922
timestamp 1586364061
transform 1 0 1104 0 1 252960
box -38 -48 314 592
use scs8hd_decap_12  FILLER_461_3
timestamp 1586364061
transform 1 0 1380 0 1 252960
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_461_15
timestamp 1586364061
transform 1 0 2484 0 1 252960
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_461_27
timestamp 1586364061
transform 1 0 3588 0 1 252960
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_461_39
timestamp 1586364061
transform 1 0 4692 0 1 252960
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_461_51
timestamp 1586364061
transform 1 0 5796 0 1 252960
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1670
timestamp 1586364061
transform 1 0 6716 0 1 252960
box -38 -48 130 592
use scs8hd_fill_2  FILLER_461_59
timestamp 1586364061
transform 1 0 6532 0 1 252960
box -38 -48 222 592
use scs8hd_decap_12  FILLER_461_62
timestamp 1586364061
transform 1 0 6808 0 1 252960
box -38 -48 1142 592
use scs8hd_decap_3  PHY_923
timestamp 1586364061
transform -1 0 8832 0 1 252960
box -38 -48 314 592
use scs8hd_decap_6  FILLER_461_74
timestamp 1586364061
transform 1 0 7912 0 1 252960
box -38 -48 590 592
use scs8hd_fill_1  FILLER_461_80
timestamp 1586364061
transform 1 0 8464 0 1 252960
box -38 -48 130 592
use scs8hd_decap_3  PHY_924
timestamp 1586364061
transform 1 0 1104 0 -1 254048
box -38 -48 314 592
use scs8hd_decap_3  PHY_926
timestamp 1586364061
transform 1 0 1104 0 1 254048
box -38 -48 314 592
use scs8hd_decap_12  FILLER_462_3
timestamp 1586364061
transform 1 0 1380 0 -1 254048
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_462_15
timestamp 1586364061
transform 1 0 2484 0 -1 254048
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_463_3
timestamp 1586364061
transform 1 0 1380 0 1 254048
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_463_15
timestamp 1586364061
transform 1 0 2484 0 1 254048
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1671
timestamp 1586364061
transform 1 0 3956 0 -1 254048
box -38 -48 130 592
use scs8hd_decap_4  FILLER_462_27
timestamp 1586364061
transform 1 0 3588 0 -1 254048
box -38 -48 406 592
use scs8hd_decap_12  FILLER_462_32
timestamp 1586364061
transform 1 0 4048 0 -1 254048
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_463_27
timestamp 1586364061
transform 1 0 3588 0 1 254048
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_462_44
timestamp 1586364061
transform 1 0 5152 0 -1 254048
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_463_39
timestamp 1586364061
transform 1 0 4692 0 1 254048
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_463_51
timestamp 1586364061
transform 1 0 5796 0 1 254048
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1672
timestamp 1586364061
transform 1 0 6716 0 1 254048
box -38 -48 130 592
use scs8hd_decap_12  FILLER_462_56
timestamp 1586364061
transform 1 0 6256 0 -1 254048
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_462_68
timestamp 1586364061
transform 1 0 7360 0 -1 254048
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_463_59
timestamp 1586364061
transform 1 0 6532 0 1 254048
box -38 -48 222 592
use scs8hd_decap_12  FILLER_463_62
timestamp 1586364061
transform 1 0 6808 0 1 254048
box -38 -48 1142 592
use scs8hd_decap_3  PHY_925
timestamp 1586364061
transform -1 0 8832 0 -1 254048
box -38 -48 314 592
use scs8hd_decap_3  PHY_927
timestamp 1586364061
transform -1 0 8832 0 1 254048
box -38 -48 314 592
use scs8hd_fill_1  FILLER_462_80
timestamp 1586364061
transform 1 0 8464 0 -1 254048
box -38 -48 130 592
use scs8hd_decap_6  FILLER_463_74
timestamp 1586364061
transform 1 0 7912 0 1 254048
box -38 -48 590 592
use scs8hd_fill_1  FILLER_463_80
timestamp 1586364061
transform 1 0 8464 0 1 254048
box -38 -48 130 592
use scs8hd_decap_3  PHY_928
timestamp 1586364061
transform 1 0 1104 0 -1 255136
box -38 -48 314 592
use scs8hd_decap_12  FILLER_464_3
timestamp 1586364061
transform 1 0 1380 0 -1 255136
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_464_15
timestamp 1586364061
transform 1 0 2484 0 -1 255136
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1673
timestamp 1586364061
transform 1 0 3956 0 -1 255136
box -38 -48 130 592
use scs8hd_decap_4  FILLER_464_27
timestamp 1586364061
transform 1 0 3588 0 -1 255136
box -38 -48 406 592
use scs8hd_decap_12  FILLER_464_32
timestamp 1586364061
transform 1 0 4048 0 -1 255136
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_464_44
timestamp 1586364061
transform 1 0 5152 0 -1 255136
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_464_56
timestamp 1586364061
transform 1 0 6256 0 -1 255136
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_464_68
timestamp 1586364061
transform 1 0 7360 0 -1 255136
box -38 -48 1142 592
use scs8hd_decap_3  PHY_929
timestamp 1586364061
transform -1 0 8832 0 -1 255136
box -38 -48 314 592
use scs8hd_fill_1  FILLER_464_80
timestamp 1586364061
transform 1 0 8464 0 -1 255136
box -38 -48 130 592
use scs8hd_decap_3  PHY_930
timestamp 1586364061
transform 1 0 1104 0 1 255136
box -38 -48 314 592
use scs8hd_decap_12  FILLER_465_3
timestamp 1586364061
transform 1 0 1380 0 1 255136
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_465_15
timestamp 1586364061
transform 1 0 2484 0 1 255136
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_465_27
timestamp 1586364061
transform 1 0 3588 0 1 255136
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_465_39
timestamp 1586364061
transform 1 0 4692 0 1 255136
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_465_51
timestamp 1586364061
transform 1 0 5796 0 1 255136
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1674
timestamp 1586364061
transform 1 0 6716 0 1 255136
box -38 -48 130 592
use scs8hd_fill_2  FILLER_465_59
timestamp 1586364061
transform 1 0 6532 0 1 255136
box -38 -48 222 592
use scs8hd_decap_12  FILLER_465_62
timestamp 1586364061
transform 1 0 6808 0 1 255136
box -38 -48 1142 592
use scs8hd_decap_3  PHY_931
timestamp 1586364061
transform -1 0 8832 0 1 255136
box -38 -48 314 592
use scs8hd_decap_6  FILLER_465_74
timestamp 1586364061
transform 1 0 7912 0 1 255136
box -38 -48 590 592
use scs8hd_fill_1  FILLER_465_80
timestamp 1586364061
transform 1 0 8464 0 1 255136
box -38 -48 130 592
use scs8hd_decap_3  PHY_932
timestamp 1586364061
transform 1 0 1104 0 -1 256224
box -38 -48 314 592
use scs8hd_decap_12  FILLER_466_3
timestamp 1586364061
transform 1 0 1380 0 -1 256224
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_466_15
timestamp 1586364061
transform 1 0 2484 0 -1 256224
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1675
timestamp 1586364061
transform 1 0 3956 0 -1 256224
box -38 -48 130 592
use scs8hd_decap_4  FILLER_466_27
timestamp 1586364061
transform 1 0 3588 0 -1 256224
box -38 -48 406 592
use scs8hd_decap_12  FILLER_466_32
timestamp 1586364061
transform 1 0 4048 0 -1 256224
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_466_44
timestamp 1586364061
transform 1 0 5152 0 -1 256224
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_466_56
timestamp 1586364061
transform 1 0 6256 0 -1 256224
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_466_68
timestamp 1586364061
transform 1 0 7360 0 -1 256224
box -38 -48 1142 592
use scs8hd_decap_3  PHY_933
timestamp 1586364061
transform -1 0 8832 0 -1 256224
box -38 -48 314 592
use scs8hd_fill_1  FILLER_466_80
timestamp 1586364061
transform 1 0 8464 0 -1 256224
box -38 -48 130 592
use scs8hd_decap_3  PHY_934
timestamp 1586364061
transform 1 0 1104 0 1 256224
box -38 -48 314 592
use scs8hd_decap_12  FILLER_467_3
timestamp 1586364061
transform 1 0 1380 0 1 256224
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_467_15
timestamp 1586364061
transform 1 0 2484 0 1 256224
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_467_27
timestamp 1586364061
transform 1 0 3588 0 1 256224
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_467_39
timestamp 1586364061
transform 1 0 4692 0 1 256224
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_467_51
timestamp 1586364061
transform 1 0 5796 0 1 256224
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1676
timestamp 1586364061
transform 1 0 6716 0 1 256224
box -38 -48 130 592
use scs8hd_fill_2  FILLER_467_59
timestamp 1586364061
transform 1 0 6532 0 1 256224
box -38 -48 222 592
use scs8hd_decap_12  FILLER_467_62
timestamp 1586364061
transform 1 0 6808 0 1 256224
box -38 -48 1142 592
use scs8hd_decap_3  PHY_935
timestamp 1586364061
transform -1 0 8832 0 1 256224
box -38 -48 314 592
use scs8hd_decap_6  FILLER_467_74
timestamp 1586364061
transform 1 0 7912 0 1 256224
box -38 -48 590 592
use scs8hd_fill_1  FILLER_467_80
timestamp 1586364061
transform 1 0 8464 0 1 256224
box -38 -48 130 592
use scs8hd_decap_3  PHY_936
timestamp 1586364061
transform 1 0 1104 0 -1 257312
box -38 -48 314 592
use scs8hd_decap_12  FILLER_468_3
timestamp 1586364061
transform 1 0 1380 0 -1 257312
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_468_15
timestamp 1586364061
transform 1 0 2484 0 -1 257312
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1677
timestamp 1586364061
transform 1 0 3956 0 -1 257312
box -38 -48 130 592
use scs8hd_decap_4  FILLER_468_27
timestamp 1586364061
transform 1 0 3588 0 -1 257312
box -38 -48 406 592
use scs8hd_decap_12  FILLER_468_32
timestamp 1586364061
transform 1 0 4048 0 -1 257312
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_468_44
timestamp 1586364061
transform 1 0 5152 0 -1 257312
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_468_56
timestamp 1586364061
transform 1 0 6256 0 -1 257312
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_468_68
timestamp 1586364061
transform 1 0 7360 0 -1 257312
box -38 -48 1142 592
use scs8hd_decap_3  PHY_937
timestamp 1586364061
transform -1 0 8832 0 -1 257312
box -38 -48 314 592
use scs8hd_fill_1  FILLER_468_80
timestamp 1586364061
transform 1 0 8464 0 -1 257312
box -38 -48 130 592
use scs8hd_decap_3  PHY_938
timestamp 1586364061
transform 1 0 1104 0 1 257312
box -38 -48 314 592
use scs8hd_decap_3  PHY_940
timestamp 1586364061
transform 1 0 1104 0 -1 258400
box -38 -48 314 592
use scs8hd_decap_12  FILLER_469_3
timestamp 1586364061
transform 1 0 1380 0 1 257312
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_469_15
timestamp 1586364061
transform 1 0 2484 0 1 257312
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_470_3
timestamp 1586364061
transform 1 0 1380 0 -1 258400
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_470_15
timestamp 1586364061
transform 1 0 2484 0 -1 258400
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1679
timestamp 1586364061
transform 1 0 3956 0 -1 258400
box -38 -48 130 592
use scs8hd_decap_12  FILLER_469_27
timestamp 1586364061
transform 1 0 3588 0 1 257312
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_470_27
timestamp 1586364061
transform 1 0 3588 0 -1 258400
box -38 -48 406 592
use scs8hd_decap_12  FILLER_470_32
timestamp 1586364061
transform 1 0 4048 0 -1 258400
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_469_39
timestamp 1586364061
transform 1 0 4692 0 1 257312
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_469_51
timestamp 1586364061
transform 1 0 5796 0 1 257312
box -38 -48 774 592
use scs8hd_decap_12  FILLER_470_44
timestamp 1586364061
transform 1 0 5152 0 -1 258400
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1678
timestamp 1586364061
transform 1 0 6716 0 1 257312
box -38 -48 130 592
use scs8hd_fill_2  FILLER_469_59
timestamp 1586364061
transform 1 0 6532 0 1 257312
box -38 -48 222 592
use scs8hd_decap_12  FILLER_469_62
timestamp 1586364061
transform 1 0 6808 0 1 257312
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_470_56
timestamp 1586364061
transform 1 0 6256 0 -1 258400
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_470_68
timestamp 1586364061
transform 1 0 7360 0 -1 258400
box -38 -48 1142 592
use scs8hd_decap_3  PHY_939
timestamp 1586364061
transform -1 0 8832 0 1 257312
box -38 -48 314 592
use scs8hd_decap_3  PHY_941
timestamp 1586364061
transform -1 0 8832 0 -1 258400
box -38 -48 314 592
use scs8hd_decap_6  FILLER_469_74
timestamp 1586364061
transform 1 0 7912 0 1 257312
box -38 -48 590 592
use scs8hd_fill_1  FILLER_469_80
timestamp 1586364061
transform 1 0 8464 0 1 257312
box -38 -48 130 592
use scs8hd_fill_1  FILLER_470_80
timestamp 1586364061
transform 1 0 8464 0 -1 258400
box -38 -48 130 592
use scs8hd_decap_3  PHY_942
timestamp 1586364061
transform 1 0 1104 0 1 258400
box -38 -48 314 592
use scs8hd_decap_12  FILLER_471_3
timestamp 1586364061
transform 1 0 1380 0 1 258400
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_471_15
timestamp 1586364061
transform 1 0 2484 0 1 258400
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_471_27
timestamp 1586364061
transform 1 0 3588 0 1 258400
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_471_39
timestamp 1586364061
transform 1 0 4692 0 1 258400
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_471_51
timestamp 1586364061
transform 1 0 5796 0 1 258400
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1680
timestamp 1586364061
transform 1 0 6716 0 1 258400
box -38 -48 130 592
use scs8hd_fill_2  FILLER_471_59
timestamp 1586364061
transform 1 0 6532 0 1 258400
box -38 -48 222 592
use scs8hd_decap_12  FILLER_471_62
timestamp 1586364061
transform 1 0 6808 0 1 258400
box -38 -48 1142 592
use scs8hd_decap_3  PHY_943
timestamp 1586364061
transform -1 0 8832 0 1 258400
box -38 -48 314 592
use scs8hd_decap_6  FILLER_471_74
timestamp 1586364061
transform 1 0 7912 0 1 258400
box -38 -48 590 592
use scs8hd_fill_1  FILLER_471_80
timestamp 1586364061
transform 1 0 8464 0 1 258400
box -38 -48 130 592
use scs8hd_decap_3  PHY_944
timestamp 1586364061
transform 1 0 1104 0 -1 259488
box -38 -48 314 592
use scs8hd_decap_12  FILLER_472_3
timestamp 1586364061
transform 1 0 1380 0 -1 259488
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_472_15
timestamp 1586364061
transform 1 0 2484 0 -1 259488
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1681
timestamp 1586364061
transform 1 0 3956 0 -1 259488
box -38 -48 130 592
use scs8hd_decap_4  FILLER_472_27
timestamp 1586364061
transform 1 0 3588 0 -1 259488
box -38 -48 406 592
use scs8hd_decap_12  FILLER_472_32
timestamp 1586364061
transform 1 0 4048 0 -1 259488
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_472_44
timestamp 1586364061
transform 1 0 5152 0 -1 259488
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_472_56
timestamp 1586364061
transform 1 0 6256 0 -1 259488
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_472_68
timestamp 1586364061
transform 1 0 7360 0 -1 259488
box -38 -48 1142 592
use scs8hd_decap_3  PHY_945
timestamp 1586364061
transform -1 0 8832 0 -1 259488
box -38 -48 314 592
use scs8hd_fill_1  FILLER_472_80
timestamp 1586364061
transform 1 0 8464 0 -1 259488
box -38 -48 130 592
use scs8hd_decap_3  PHY_946
timestamp 1586364061
transform 1 0 1104 0 1 259488
box -38 -48 314 592
use scs8hd_decap_12  FILLER_473_3
timestamp 1586364061
transform 1 0 1380 0 1 259488
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_473_15
timestamp 1586364061
transform 1 0 2484 0 1 259488
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_473_27
timestamp 1586364061
transform 1 0 3588 0 1 259488
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_473_39
timestamp 1586364061
transform 1 0 4692 0 1 259488
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_473_51
timestamp 1586364061
transform 1 0 5796 0 1 259488
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1682
timestamp 1586364061
transform 1 0 6716 0 1 259488
box -38 -48 130 592
use scs8hd_fill_2  FILLER_473_59
timestamp 1586364061
transform 1 0 6532 0 1 259488
box -38 -48 222 592
use scs8hd_decap_12  FILLER_473_62
timestamp 1586364061
transform 1 0 6808 0 1 259488
box -38 -48 1142 592
use scs8hd_decap_3  PHY_947
timestamp 1586364061
transform -1 0 8832 0 1 259488
box -38 -48 314 592
use scs8hd_decap_6  FILLER_473_74
timestamp 1586364061
transform 1 0 7912 0 1 259488
box -38 -48 590 592
use scs8hd_fill_1  FILLER_473_80
timestamp 1586364061
transform 1 0 8464 0 1 259488
box -38 -48 130 592
use scs8hd_decap_3  PHY_948
timestamp 1586364061
transform 1 0 1104 0 -1 260576
box -38 -48 314 592
use scs8hd_decap_12  FILLER_474_3
timestamp 1586364061
transform 1 0 1380 0 -1 260576
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_474_15
timestamp 1586364061
transform 1 0 2484 0 -1 260576
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1683
timestamp 1586364061
transform 1 0 3956 0 -1 260576
box -38 -48 130 592
use scs8hd_decap_4  FILLER_474_27
timestamp 1586364061
transform 1 0 3588 0 -1 260576
box -38 -48 406 592
use scs8hd_decap_12  FILLER_474_32
timestamp 1586364061
transform 1 0 4048 0 -1 260576
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_474_44
timestamp 1586364061
transform 1 0 5152 0 -1 260576
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_474_56
timestamp 1586364061
transform 1 0 6256 0 -1 260576
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_474_68
timestamp 1586364061
transform 1 0 7360 0 -1 260576
box -38 -48 1142 592
use scs8hd_decap_3  PHY_949
timestamp 1586364061
transform -1 0 8832 0 -1 260576
box -38 -48 314 592
use scs8hd_fill_1  FILLER_474_80
timestamp 1586364061
transform 1 0 8464 0 -1 260576
box -38 -48 130 592
use scs8hd_decap_3  PHY_950
timestamp 1586364061
transform 1 0 1104 0 1 260576
box -38 -48 314 592
use scs8hd_decap_3  PHY_952
timestamp 1586364061
transform 1 0 1104 0 -1 261664
box -38 -48 314 592
use scs8hd_decap_12  FILLER_475_3
timestamp 1586364061
transform 1 0 1380 0 1 260576
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_475_15
timestamp 1586364061
transform 1 0 2484 0 1 260576
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_476_3
timestamp 1586364061
transform 1 0 1380 0 -1 261664
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_476_15
timestamp 1586364061
transform 1 0 2484 0 -1 261664
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1685
timestamp 1586364061
transform 1 0 3956 0 -1 261664
box -38 -48 130 592
use scs8hd_decap_12  FILLER_475_27
timestamp 1586364061
transform 1 0 3588 0 1 260576
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_476_27
timestamp 1586364061
transform 1 0 3588 0 -1 261664
box -38 -48 406 592
use scs8hd_decap_12  FILLER_476_32
timestamp 1586364061
transform 1 0 4048 0 -1 261664
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_475_39
timestamp 1586364061
transform 1 0 4692 0 1 260576
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_475_51
timestamp 1586364061
transform 1 0 5796 0 1 260576
box -38 -48 774 592
use scs8hd_decap_12  FILLER_476_44
timestamp 1586364061
transform 1 0 5152 0 -1 261664
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1684
timestamp 1586364061
transform 1 0 6716 0 1 260576
box -38 -48 130 592
use scs8hd_fill_2  FILLER_475_59
timestamp 1586364061
transform 1 0 6532 0 1 260576
box -38 -48 222 592
use scs8hd_decap_12  FILLER_475_62
timestamp 1586364061
transform 1 0 6808 0 1 260576
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_476_56
timestamp 1586364061
transform 1 0 6256 0 -1 261664
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_476_68
timestamp 1586364061
transform 1 0 7360 0 -1 261664
box -38 -48 1142 592
use scs8hd_decap_3  PHY_951
timestamp 1586364061
transform -1 0 8832 0 1 260576
box -38 -48 314 592
use scs8hd_decap_3  PHY_953
timestamp 1586364061
transform -1 0 8832 0 -1 261664
box -38 -48 314 592
use scs8hd_decap_6  FILLER_475_74
timestamp 1586364061
transform 1 0 7912 0 1 260576
box -38 -48 590 592
use scs8hd_fill_1  FILLER_475_80
timestamp 1586364061
transform 1 0 8464 0 1 260576
box -38 -48 130 592
use scs8hd_fill_1  FILLER_476_80
timestamp 1586364061
transform 1 0 8464 0 -1 261664
box -38 -48 130 592
use scs8hd_decap_3  PHY_954
timestamp 1586364061
transform 1 0 1104 0 1 261664
box -38 -48 314 592
use scs8hd_decap_12  FILLER_477_3
timestamp 1586364061
transform 1 0 1380 0 1 261664
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_477_15
timestamp 1586364061
transform 1 0 2484 0 1 261664
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_477_27
timestamp 1586364061
transform 1 0 3588 0 1 261664
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_477_39
timestamp 1586364061
transform 1 0 4692 0 1 261664
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_477_51
timestamp 1586364061
transform 1 0 5796 0 1 261664
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1686
timestamp 1586364061
transform 1 0 6716 0 1 261664
box -38 -48 130 592
use scs8hd_fill_2  FILLER_477_59
timestamp 1586364061
transform 1 0 6532 0 1 261664
box -38 -48 222 592
use scs8hd_decap_12  FILLER_477_62
timestamp 1586364061
transform 1 0 6808 0 1 261664
box -38 -48 1142 592
use scs8hd_decap_3  PHY_955
timestamp 1586364061
transform -1 0 8832 0 1 261664
box -38 -48 314 592
use scs8hd_decap_6  FILLER_477_74
timestamp 1586364061
transform 1 0 7912 0 1 261664
box -38 -48 590 592
use scs8hd_fill_1  FILLER_477_80
timestamp 1586364061
transform 1 0 8464 0 1 261664
box -38 -48 130 592
use scs8hd_decap_3  PHY_956
timestamp 1586364061
transform 1 0 1104 0 -1 262752
box -38 -48 314 592
use scs8hd_decap_12  FILLER_478_3
timestamp 1586364061
transform 1 0 1380 0 -1 262752
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_478_15
timestamp 1586364061
transform 1 0 2484 0 -1 262752
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1687
timestamp 1586364061
transform 1 0 3956 0 -1 262752
box -38 -48 130 592
use scs8hd_decap_4  FILLER_478_27
timestamp 1586364061
transform 1 0 3588 0 -1 262752
box -38 -48 406 592
use scs8hd_decap_12  FILLER_478_32
timestamp 1586364061
transform 1 0 4048 0 -1 262752
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_478_44
timestamp 1586364061
transform 1 0 5152 0 -1 262752
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_478_56
timestamp 1586364061
transform 1 0 6256 0 -1 262752
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_478_68
timestamp 1586364061
transform 1 0 7360 0 -1 262752
box -38 -48 1142 592
use scs8hd_decap_3  PHY_957
timestamp 1586364061
transform -1 0 8832 0 -1 262752
box -38 -48 314 592
use scs8hd_fill_1  FILLER_478_80
timestamp 1586364061
transform 1 0 8464 0 -1 262752
box -38 -48 130 592
use scs8hd_decap_3  PHY_958
timestamp 1586364061
transform 1 0 1104 0 1 262752
box -38 -48 314 592
use scs8hd_decap_12  FILLER_479_3
timestamp 1586364061
transform 1 0 1380 0 1 262752
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_479_15
timestamp 1586364061
transform 1 0 2484 0 1 262752
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_479_27
timestamp 1586364061
transform 1 0 3588 0 1 262752
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_479_39
timestamp 1586364061
transform 1 0 4692 0 1 262752
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_479_51
timestamp 1586364061
transform 1 0 5796 0 1 262752
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1688
timestamp 1586364061
transform 1 0 6716 0 1 262752
box -38 -48 130 592
use scs8hd_fill_2  FILLER_479_59
timestamp 1586364061
transform 1 0 6532 0 1 262752
box -38 -48 222 592
use scs8hd_decap_12  FILLER_479_62
timestamp 1586364061
transform 1 0 6808 0 1 262752
box -38 -48 1142 592
use scs8hd_decap_3  PHY_959
timestamp 1586364061
transform -1 0 8832 0 1 262752
box -38 -48 314 592
use scs8hd_decap_6  FILLER_479_74
timestamp 1586364061
transform 1 0 7912 0 1 262752
box -38 -48 590 592
use scs8hd_fill_1  FILLER_479_80
timestamp 1586364061
transform 1 0 8464 0 1 262752
box -38 -48 130 592
use scs8hd_decap_3  PHY_960
timestamp 1586364061
transform 1 0 1104 0 -1 263840
box -38 -48 314 592
use scs8hd_decap_12  FILLER_480_3
timestamp 1586364061
transform 1 0 1380 0 -1 263840
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_480_15
timestamp 1586364061
transform 1 0 2484 0 -1 263840
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1689
timestamp 1586364061
transform 1 0 3956 0 -1 263840
box -38 -48 130 592
use scs8hd_decap_4  FILLER_480_27
timestamp 1586364061
transform 1 0 3588 0 -1 263840
box -38 -48 406 592
use scs8hd_decap_12  FILLER_480_32
timestamp 1586364061
transform 1 0 4048 0 -1 263840
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_480_44
timestamp 1586364061
transform 1 0 5152 0 -1 263840
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_480_56
timestamp 1586364061
transform 1 0 6256 0 -1 263840
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_480_68
timestamp 1586364061
transform 1 0 7360 0 -1 263840
box -38 -48 1142 592
use scs8hd_decap_3  PHY_961
timestamp 1586364061
transform -1 0 8832 0 -1 263840
box -38 -48 314 592
use scs8hd_fill_1  FILLER_480_80
timestamp 1586364061
transform 1 0 8464 0 -1 263840
box -38 -48 130 592
use scs8hd_decap_3  PHY_962
timestamp 1586364061
transform 1 0 1104 0 1 263840
box -38 -48 314 592
use scs8hd_decap_12  FILLER_481_3
timestamp 1586364061
transform 1 0 1380 0 1 263840
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_481_15
timestamp 1586364061
transform 1 0 2484 0 1 263840
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_481_27
timestamp 1586364061
transform 1 0 3588 0 1 263840
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_481_39
timestamp 1586364061
transform 1 0 4692 0 1 263840
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_481_51
timestamp 1586364061
transform 1 0 5796 0 1 263840
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1690
timestamp 1586364061
transform 1 0 6716 0 1 263840
box -38 -48 130 592
use scs8hd_fill_2  FILLER_481_59
timestamp 1586364061
transform 1 0 6532 0 1 263840
box -38 -48 222 592
use scs8hd_decap_12  FILLER_481_62
timestamp 1586364061
transform 1 0 6808 0 1 263840
box -38 -48 1142 592
use scs8hd_decap_3  PHY_963
timestamp 1586364061
transform -1 0 8832 0 1 263840
box -38 -48 314 592
use scs8hd_decap_6  FILLER_481_74
timestamp 1586364061
transform 1 0 7912 0 1 263840
box -38 -48 590 592
use scs8hd_fill_1  FILLER_481_80
timestamp 1586364061
transform 1 0 8464 0 1 263840
box -38 -48 130 592
use scs8hd_decap_3  PHY_964
timestamp 1586364061
transform 1 0 1104 0 -1 264928
box -38 -48 314 592
use scs8hd_decap_3  PHY_966
timestamp 1586364061
transform 1 0 1104 0 1 264928
box -38 -48 314 592
use scs8hd_decap_12  FILLER_482_3
timestamp 1586364061
transform 1 0 1380 0 -1 264928
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_482_15
timestamp 1586364061
transform 1 0 2484 0 -1 264928
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_483_3
timestamp 1586364061
transform 1 0 1380 0 1 264928
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_483_15
timestamp 1586364061
transform 1 0 2484 0 1 264928
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1691
timestamp 1586364061
transform 1 0 3956 0 -1 264928
box -38 -48 130 592
use scs8hd_decap_4  FILLER_482_27
timestamp 1586364061
transform 1 0 3588 0 -1 264928
box -38 -48 406 592
use scs8hd_decap_12  FILLER_482_32
timestamp 1586364061
transform 1 0 4048 0 -1 264928
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_483_27
timestamp 1586364061
transform 1 0 3588 0 1 264928
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_482_44
timestamp 1586364061
transform 1 0 5152 0 -1 264928
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_483_39
timestamp 1586364061
transform 1 0 4692 0 1 264928
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_483_51
timestamp 1586364061
transform 1 0 5796 0 1 264928
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1692
timestamp 1586364061
transform 1 0 6716 0 1 264928
box -38 -48 130 592
use scs8hd_decap_12  FILLER_482_56
timestamp 1586364061
transform 1 0 6256 0 -1 264928
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_482_68
timestamp 1586364061
transform 1 0 7360 0 -1 264928
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_483_59
timestamp 1586364061
transform 1 0 6532 0 1 264928
box -38 -48 222 592
use scs8hd_decap_12  FILLER_483_62
timestamp 1586364061
transform 1 0 6808 0 1 264928
box -38 -48 1142 592
use scs8hd_decap_3  PHY_965
timestamp 1586364061
transform -1 0 8832 0 -1 264928
box -38 -48 314 592
use scs8hd_decap_3  PHY_967
timestamp 1586364061
transform -1 0 8832 0 1 264928
box -38 -48 314 592
use scs8hd_fill_1  FILLER_482_80
timestamp 1586364061
transform 1 0 8464 0 -1 264928
box -38 -48 130 592
use scs8hd_decap_6  FILLER_483_74
timestamp 1586364061
transform 1 0 7912 0 1 264928
box -38 -48 590 592
use scs8hd_fill_1  FILLER_483_80
timestamp 1586364061
transform 1 0 8464 0 1 264928
box -38 -48 130 592
use scs8hd_decap_3  PHY_968
timestamp 1586364061
transform 1 0 1104 0 -1 266016
box -38 -48 314 592
use scs8hd_decap_12  FILLER_484_3
timestamp 1586364061
transform 1 0 1380 0 -1 266016
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_484_15
timestamp 1586364061
transform 1 0 2484 0 -1 266016
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1693
timestamp 1586364061
transform 1 0 3956 0 -1 266016
box -38 -48 130 592
use scs8hd_decap_4  FILLER_484_27
timestamp 1586364061
transform 1 0 3588 0 -1 266016
box -38 -48 406 592
use scs8hd_decap_12  FILLER_484_32
timestamp 1586364061
transform 1 0 4048 0 -1 266016
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_484_44
timestamp 1586364061
transform 1 0 5152 0 -1 266016
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_484_56
timestamp 1586364061
transform 1 0 6256 0 -1 266016
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_484_68
timestamp 1586364061
transform 1 0 7360 0 -1 266016
box -38 -48 1142 592
use scs8hd_decap_3  PHY_969
timestamp 1586364061
transform -1 0 8832 0 -1 266016
box -38 -48 314 592
use scs8hd_fill_1  FILLER_484_80
timestamp 1586364061
transform 1 0 8464 0 -1 266016
box -38 -48 130 592
use scs8hd_decap_3  PHY_970
timestamp 1586364061
transform 1 0 1104 0 1 266016
box -38 -48 314 592
use scs8hd_decap_12  FILLER_485_3
timestamp 1586364061
transform 1 0 1380 0 1 266016
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_485_15
timestamp 1586364061
transform 1 0 2484 0 1 266016
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_485_27
timestamp 1586364061
transform 1 0 3588 0 1 266016
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_485_39
timestamp 1586364061
transform 1 0 4692 0 1 266016
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_485_51
timestamp 1586364061
transform 1 0 5796 0 1 266016
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1694
timestamp 1586364061
transform 1 0 6716 0 1 266016
box -38 -48 130 592
use scs8hd_fill_2  FILLER_485_59
timestamp 1586364061
transform 1 0 6532 0 1 266016
box -38 -48 222 592
use scs8hd_decap_12  FILLER_485_62
timestamp 1586364061
transform 1 0 6808 0 1 266016
box -38 -48 1142 592
use scs8hd_decap_3  PHY_971
timestamp 1586364061
transform -1 0 8832 0 1 266016
box -38 -48 314 592
use scs8hd_decap_6  FILLER_485_74
timestamp 1586364061
transform 1 0 7912 0 1 266016
box -38 -48 590 592
use scs8hd_fill_1  FILLER_485_80
timestamp 1586364061
transform 1 0 8464 0 1 266016
box -38 -48 130 592
use scs8hd_decap_3  PHY_972
timestamp 1586364061
transform 1 0 1104 0 -1 267104
box -38 -48 314 592
use scs8hd_decap_12  FILLER_486_3
timestamp 1586364061
transform 1 0 1380 0 -1 267104
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_486_15
timestamp 1586364061
transform 1 0 2484 0 -1 267104
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1695
timestamp 1586364061
transform 1 0 3956 0 -1 267104
box -38 -48 130 592
use scs8hd_decap_4  FILLER_486_27
timestamp 1586364061
transform 1 0 3588 0 -1 267104
box -38 -48 406 592
use scs8hd_decap_12  FILLER_486_32
timestamp 1586364061
transform 1 0 4048 0 -1 267104
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_486_44
timestamp 1586364061
transform 1 0 5152 0 -1 267104
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_486_56
timestamp 1586364061
transform 1 0 6256 0 -1 267104
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_486_68
timestamp 1586364061
transform 1 0 7360 0 -1 267104
box -38 -48 1142 592
use scs8hd_decap_3  PHY_973
timestamp 1586364061
transform -1 0 8832 0 -1 267104
box -38 -48 314 592
use scs8hd_fill_1  FILLER_486_80
timestamp 1586364061
transform 1 0 8464 0 -1 267104
box -38 -48 130 592
use scs8hd_decap_3  PHY_974
timestamp 1586364061
transform 1 0 1104 0 1 267104
box -38 -48 314 592
use scs8hd_decap_12  FILLER_487_3
timestamp 1586364061
transform 1 0 1380 0 1 267104
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_487_15
timestamp 1586364061
transform 1 0 2484 0 1 267104
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_487_27
timestamp 1586364061
transform 1 0 3588 0 1 267104
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_487_39
timestamp 1586364061
transform 1 0 4692 0 1 267104
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_487_51
timestamp 1586364061
transform 1 0 5796 0 1 267104
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1696
timestamp 1586364061
transform 1 0 6716 0 1 267104
box -38 -48 130 592
use scs8hd_fill_2  FILLER_487_59
timestamp 1586364061
transform 1 0 6532 0 1 267104
box -38 -48 222 592
use scs8hd_decap_12  FILLER_487_62
timestamp 1586364061
transform 1 0 6808 0 1 267104
box -38 -48 1142 592
use scs8hd_decap_3  PHY_975
timestamp 1586364061
transform -1 0 8832 0 1 267104
box -38 -48 314 592
use scs8hd_decap_6  FILLER_487_74
timestamp 1586364061
transform 1 0 7912 0 1 267104
box -38 -48 590 592
use scs8hd_fill_1  FILLER_487_80
timestamp 1586364061
transform 1 0 8464 0 1 267104
box -38 -48 130 592
use scs8hd_decap_3  PHY_976
timestamp 1586364061
transform 1 0 1104 0 -1 268192
box -38 -48 314 592
use scs8hd_decap_12  FILLER_488_3
timestamp 1586364061
transform 1 0 1380 0 -1 268192
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_488_15
timestamp 1586364061
transform 1 0 2484 0 -1 268192
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1697
timestamp 1586364061
transform 1 0 3956 0 -1 268192
box -38 -48 130 592
use scs8hd_decap_4  FILLER_488_27
timestamp 1586364061
transform 1 0 3588 0 -1 268192
box -38 -48 406 592
use scs8hd_decap_12  FILLER_488_32
timestamp 1586364061
transform 1 0 4048 0 -1 268192
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_488_44
timestamp 1586364061
transform 1 0 5152 0 -1 268192
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_488_56
timestamp 1586364061
transform 1 0 6256 0 -1 268192
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_488_68
timestamp 1586364061
transform 1 0 7360 0 -1 268192
box -38 -48 1142 592
use scs8hd_decap_3  PHY_977
timestamp 1586364061
transform -1 0 8832 0 -1 268192
box -38 -48 314 592
use scs8hd_fill_1  FILLER_488_80
timestamp 1586364061
transform 1 0 8464 0 -1 268192
box -38 -48 130 592
use scs8hd_decap_3  PHY_978
timestamp 1586364061
transform 1 0 1104 0 1 268192
box -38 -48 314 592
use scs8hd_decap_3  PHY_980
timestamp 1586364061
transform 1 0 1104 0 -1 269280
box -38 -48 314 592
use scs8hd_decap_12  FILLER_489_3
timestamp 1586364061
transform 1 0 1380 0 1 268192
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_489_15
timestamp 1586364061
transform 1 0 2484 0 1 268192
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_490_3
timestamp 1586364061
transform 1 0 1380 0 -1 269280
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_490_15
timestamp 1586364061
transform 1 0 2484 0 -1 269280
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1699
timestamp 1586364061
transform 1 0 3956 0 -1 269280
box -38 -48 130 592
use scs8hd_decap_12  FILLER_489_27
timestamp 1586364061
transform 1 0 3588 0 1 268192
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_490_27
timestamp 1586364061
transform 1 0 3588 0 -1 269280
box -38 -48 406 592
use scs8hd_decap_12  FILLER_490_32
timestamp 1586364061
transform 1 0 4048 0 -1 269280
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_489_39
timestamp 1586364061
transform 1 0 4692 0 1 268192
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_489_51
timestamp 1586364061
transform 1 0 5796 0 1 268192
box -38 -48 774 592
use scs8hd_decap_12  FILLER_490_44
timestamp 1586364061
transform 1 0 5152 0 -1 269280
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1698
timestamp 1586364061
transform 1 0 6716 0 1 268192
box -38 -48 130 592
use scs8hd_fill_2  FILLER_489_59
timestamp 1586364061
transform 1 0 6532 0 1 268192
box -38 -48 222 592
use scs8hd_decap_12  FILLER_489_62
timestamp 1586364061
transform 1 0 6808 0 1 268192
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_490_56
timestamp 1586364061
transform 1 0 6256 0 -1 269280
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_490_68
timestamp 1586364061
transform 1 0 7360 0 -1 269280
box -38 -48 1142 592
use scs8hd_decap_3  PHY_979
timestamp 1586364061
transform -1 0 8832 0 1 268192
box -38 -48 314 592
use scs8hd_decap_3  PHY_981
timestamp 1586364061
transform -1 0 8832 0 -1 269280
box -38 -48 314 592
use scs8hd_decap_6  FILLER_489_74
timestamp 1586364061
transform 1 0 7912 0 1 268192
box -38 -48 590 592
use scs8hd_fill_1  FILLER_489_80
timestamp 1586364061
transform 1 0 8464 0 1 268192
box -38 -48 130 592
use scs8hd_fill_1  FILLER_490_80
timestamp 1586364061
transform 1 0 8464 0 -1 269280
box -38 -48 130 592
use scs8hd_decap_3  PHY_982
timestamp 1586364061
transform 1 0 1104 0 1 269280
box -38 -48 314 592
use scs8hd_decap_12  FILLER_491_3
timestamp 1586364061
transform 1 0 1380 0 1 269280
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_491_15
timestamp 1586364061
transform 1 0 2484 0 1 269280
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_491_27
timestamp 1586364061
transform 1 0 3588 0 1 269280
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_491_39
timestamp 1586364061
transform 1 0 4692 0 1 269280
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_491_51
timestamp 1586364061
transform 1 0 5796 0 1 269280
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1700
timestamp 1586364061
transform 1 0 6716 0 1 269280
box -38 -48 130 592
use scs8hd_fill_2  FILLER_491_59
timestamp 1586364061
transform 1 0 6532 0 1 269280
box -38 -48 222 592
use scs8hd_decap_12  FILLER_491_62
timestamp 1586364061
transform 1 0 6808 0 1 269280
box -38 -48 1142 592
use scs8hd_decap_3  PHY_983
timestamp 1586364061
transform -1 0 8832 0 1 269280
box -38 -48 314 592
use scs8hd_decap_6  FILLER_491_74
timestamp 1586364061
transform 1 0 7912 0 1 269280
box -38 -48 590 592
use scs8hd_fill_1  FILLER_491_80
timestamp 1586364061
transform 1 0 8464 0 1 269280
box -38 -48 130 592
use scs8hd_decap_3  PHY_984
timestamp 1586364061
transform 1 0 1104 0 -1 270368
box -38 -48 314 592
use scs8hd_decap_12  FILLER_492_3
timestamp 1586364061
transform 1 0 1380 0 -1 270368
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_492_15
timestamp 1586364061
transform 1 0 2484 0 -1 270368
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1701
timestamp 1586364061
transform 1 0 3956 0 -1 270368
box -38 -48 130 592
use scs8hd_decap_4  FILLER_492_27
timestamp 1586364061
transform 1 0 3588 0 -1 270368
box -38 -48 406 592
use scs8hd_decap_12  FILLER_492_32
timestamp 1586364061
transform 1 0 4048 0 -1 270368
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_492_44
timestamp 1586364061
transform 1 0 5152 0 -1 270368
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_492_56
timestamp 1586364061
transform 1 0 6256 0 -1 270368
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_492_68
timestamp 1586364061
transform 1 0 7360 0 -1 270368
box -38 -48 1142 592
use scs8hd_decap_3  PHY_985
timestamp 1586364061
transform -1 0 8832 0 -1 270368
box -38 -48 314 592
use scs8hd_fill_1  FILLER_492_80
timestamp 1586364061
transform 1 0 8464 0 -1 270368
box -38 -48 130 592
use scs8hd_decap_3  PHY_986
timestamp 1586364061
transform 1 0 1104 0 1 270368
box -38 -48 314 592
use scs8hd_decap_12  FILLER_493_3
timestamp 1586364061
transform 1 0 1380 0 1 270368
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_493_15
timestamp 1586364061
transform 1 0 2484 0 1 270368
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_493_27
timestamp 1586364061
transform 1 0 3588 0 1 270368
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_493_39
timestamp 1586364061
transform 1 0 4692 0 1 270368
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_493_51
timestamp 1586364061
transform 1 0 5796 0 1 270368
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1702
timestamp 1586364061
transform 1 0 6716 0 1 270368
box -38 -48 130 592
use scs8hd_fill_2  FILLER_493_59
timestamp 1586364061
transform 1 0 6532 0 1 270368
box -38 -48 222 592
use scs8hd_decap_12  FILLER_493_62
timestamp 1586364061
transform 1 0 6808 0 1 270368
box -38 -48 1142 592
use scs8hd_decap_3  PHY_987
timestamp 1586364061
transform -1 0 8832 0 1 270368
box -38 -48 314 592
use scs8hd_decap_6  FILLER_493_74
timestamp 1586364061
transform 1 0 7912 0 1 270368
box -38 -48 590 592
use scs8hd_fill_1  FILLER_493_80
timestamp 1586364061
transform 1 0 8464 0 1 270368
box -38 -48 130 592
use scs8hd_decap_3  PHY_988
timestamp 1586364061
transform 1 0 1104 0 -1 271456
box -38 -48 314 592
use scs8hd_decap_12  FILLER_494_3
timestamp 1586364061
transform 1 0 1380 0 -1 271456
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_494_15
timestamp 1586364061
transform 1 0 2484 0 -1 271456
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1703
timestamp 1586364061
transform 1 0 3956 0 -1 271456
box -38 -48 130 592
use scs8hd_decap_4  FILLER_494_27
timestamp 1586364061
transform 1 0 3588 0 -1 271456
box -38 -48 406 592
use scs8hd_decap_12  FILLER_494_32
timestamp 1586364061
transform 1 0 4048 0 -1 271456
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_494_44
timestamp 1586364061
transform 1 0 5152 0 -1 271456
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_494_56
timestamp 1586364061
transform 1 0 6256 0 -1 271456
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_494_68
timestamp 1586364061
transform 1 0 7360 0 -1 271456
box -38 -48 1142 592
use scs8hd_decap_3  PHY_989
timestamp 1586364061
transform -1 0 8832 0 -1 271456
box -38 -48 314 592
use scs8hd_fill_1  FILLER_494_80
timestamp 1586364061
transform 1 0 8464 0 -1 271456
box -38 -48 130 592
use scs8hd_decap_3  PHY_990
timestamp 1586364061
transform 1 0 1104 0 1 271456
box -38 -48 314 592
use scs8hd_decap_3  PHY_992
timestamp 1586364061
transform 1 0 1104 0 -1 272544
box -38 -48 314 592
use scs8hd_decap_12  FILLER_495_3
timestamp 1586364061
transform 1 0 1380 0 1 271456
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_495_15
timestamp 1586364061
transform 1 0 2484 0 1 271456
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_496_3
timestamp 1586364061
transform 1 0 1380 0 -1 272544
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_496_15
timestamp 1586364061
transform 1 0 2484 0 -1 272544
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1705
timestamp 1586364061
transform 1 0 3956 0 -1 272544
box -38 -48 130 592
use scs8hd_decap_12  FILLER_495_27
timestamp 1586364061
transform 1 0 3588 0 1 271456
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_496_27
timestamp 1586364061
transform 1 0 3588 0 -1 272544
box -38 -48 406 592
use scs8hd_decap_12  FILLER_496_32
timestamp 1586364061
transform 1 0 4048 0 -1 272544
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_495_39
timestamp 1586364061
transform 1 0 4692 0 1 271456
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_495_51
timestamp 1586364061
transform 1 0 5796 0 1 271456
box -38 -48 774 592
use scs8hd_decap_12  FILLER_496_44
timestamp 1586364061
transform 1 0 5152 0 -1 272544
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1704
timestamp 1586364061
transform 1 0 6716 0 1 271456
box -38 -48 130 592
use scs8hd_fill_2  FILLER_495_59
timestamp 1586364061
transform 1 0 6532 0 1 271456
box -38 -48 222 592
use scs8hd_decap_12  FILLER_495_62
timestamp 1586364061
transform 1 0 6808 0 1 271456
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_496_56
timestamp 1586364061
transform 1 0 6256 0 -1 272544
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_496_68
timestamp 1586364061
transform 1 0 7360 0 -1 272544
box -38 -48 1142 592
use scs8hd_decap_3  PHY_991
timestamp 1586364061
transform -1 0 8832 0 1 271456
box -38 -48 314 592
use scs8hd_decap_3  PHY_993
timestamp 1586364061
transform -1 0 8832 0 -1 272544
box -38 -48 314 592
use scs8hd_decap_6  FILLER_495_74
timestamp 1586364061
transform 1 0 7912 0 1 271456
box -38 -48 590 592
use scs8hd_fill_1  FILLER_495_80
timestamp 1586364061
transform 1 0 8464 0 1 271456
box -38 -48 130 592
use scs8hd_fill_1  FILLER_496_80
timestamp 1586364061
transform 1 0 8464 0 -1 272544
box -38 -48 130 592
use scs8hd_decap_3  PHY_994
timestamp 1586364061
transform 1 0 1104 0 1 272544
box -38 -48 314 592
use scs8hd_decap_12  FILLER_497_3
timestamp 1586364061
transform 1 0 1380 0 1 272544
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_497_15
timestamp 1586364061
transform 1 0 2484 0 1 272544
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_497_27
timestamp 1586364061
transform 1 0 3588 0 1 272544
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_497_39
timestamp 1586364061
transform 1 0 4692 0 1 272544
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_497_51
timestamp 1586364061
transform 1 0 5796 0 1 272544
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1706
timestamp 1586364061
transform 1 0 6716 0 1 272544
box -38 -48 130 592
use scs8hd_fill_2  FILLER_497_59
timestamp 1586364061
transform 1 0 6532 0 1 272544
box -38 -48 222 592
use scs8hd_decap_12  FILLER_497_62
timestamp 1586364061
transform 1 0 6808 0 1 272544
box -38 -48 1142 592
use scs8hd_decap_3  PHY_995
timestamp 1586364061
transform -1 0 8832 0 1 272544
box -38 -48 314 592
use scs8hd_decap_6  FILLER_497_74
timestamp 1586364061
transform 1 0 7912 0 1 272544
box -38 -48 590 592
use scs8hd_fill_1  FILLER_497_80
timestamp 1586364061
transform 1 0 8464 0 1 272544
box -38 -48 130 592
use scs8hd_decap_3  PHY_996
timestamp 1586364061
transform 1 0 1104 0 -1 273632
box -38 -48 314 592
use scs8hd_decap_12  FILLER_498_3
timestamp 1586364061
transform 1 0 1380 0 -1 273632
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_498_15
timestamp 1586364061
transform 1 0 2484 0 -1 273632
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1707
timestamp 1586364061
transform 1 0 3956 0 -1 273632
box -38 -48 130 592
use scs8hd_decap_4  FILLER_498_27
timestamp 1586364061
transform 1 0 3588 0 -1 273632
box -38 -48 406 592
use scs8hd_decap_12  FILLER_498_32
timestamp 1586364061
transform 1 0 4048 0 -1 273632
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_498_44
timestamp 1586364061
transform 1 0 5152 0 -1 273632
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_498_56
timestamp 1586364061
transform 1 0 6256 0 -1 273632
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_498_68
timestamp 1586364061
transform 1 0 7360 0 -1 273632
box -38 -48 1142 592
use scs8hd_decap_3  PHY_997
timestamp 1586364061
transform -1 0 8832 0 -1 273632
box -38 -48 314 592
use scs8hd_fill_1  FILLER_498_80
timestamp 1586364061
transform 1 0 8464 0 -1 273632
box -38 -48 130 592
use scs8hd_decap_3  PHY_998
timestamp 1586364061
transform 1 0 1104 0 1 273632
box -38 -48 314 592
use scs8hd_decap_12  FILLER_499_3
timestamp 1586364061
transform 1 0 1380 0 1 273632
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_499_15
timestamp 1586364061
transform 1 0 2484 0 1 273632
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_499_27
timestamp 1586364061
transform 1 0 3588 0 1 273632
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_499_39
timestamp 1586364061
transform 1 0 4692 0 1 273632
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_499_51
timestamp 1586364061
transform 1 0 5796 0 1 273632
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1708
timestamp 1586364061
transform 1 0 6716 0 1 273632
box -38 -48 130 592
use scs8hd_fill_2  FILLER_499_59
timestamp 1586364061
transform 1 0 6532 0 1 273632
box -38 -48 222 592
use scs8hd_decap_12  FILLER_499_62
timestamp 1586364061
transform 1 0 6808 0 1 273632
box -38 -48 1142 592
use scs8hd_decap_3  PHY_999
timestamp 1586364061
transform -1 0 8832 0 1 273632
box -38 -48 314 592
use scs8hd_decap_6  FILLER_499_74
timestamp 1586364061
transform 1 0 7912 0 1 273632
box -38 -48 590 592
use scs8hd_fill_1  FILLER_499_80
timestamp 1586364061
transform 1 0 8464 0 1 273632
box -38 -48 130 592
use scs8hd_decap_3  PHY_1000
timestamp 1586364061
transform 1 0 1104 0 -1 274720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_500_3
timestamp 1586364061
transform 1 0 1380 0 -1 274720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_500_15
timestamp 1586364061
transform 1 0 2484 0 -1 274720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1709
timestamp 1586364061
transform 1 0 3956 0 -1 274720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_500_27
timestamp 1586364061
transform 1 0 3588 0 -1 274720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_500_32
timestamp 1586364061
transform 1 0 4048 0 -1 274720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_500_44
timestamp 1586364061
transform 1 0 5152 0 -1 274720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_500_56
timestamp 1586364061
transform 1 0 6256 0 -1 274720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_500_68
timestamp 1586364061
transform 1 0 7360 0 -1 274720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1001
timestamp 1586364061
transform -1 0 8832 0 -1 274720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_500_80
timestamp 1586364061
transform 1 0 8464 0 -1 274720
box -38 -48 130 592
use scs8hd_decap_3  PHY_1002
timestamp 1586364061
transform 1 0 1104 0 1 274720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_501_3
timestamp 1586364061
transform 1 0 1380 0 1 274720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_501_15
timestamp 1586364061
transform 1 0 2484 0 1 274720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_501_27
timestamp 1586364061
transform 1 0 3588 0 1 274720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_501_39
timestamp 1586364061
transform 1 0 4692 0 1 274720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_501_51
timestamp 1586364061
transform 1 0 5796 0 1 274720
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1710
timestamp 1586364061
transform 1 0 6716 0 1 274720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_501_59
timestamp 1586364061
transform 1 0 6532 0 1 274720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_501_62
timestamp 1586364061
transform 1 0 6808 0 1 274720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1003
timestamp 1586364061
transform -1 0 8832 0 1 274720
box -38 -48 314 592
use scs8hd_decap_6  FILLER_501_74
timestamp 1586364061
transform 1 0 7912 0 1 274720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_501_80
timestamp 1586364061
transform 1 0 8464 0 1 274720
box -38 -48 130 592
use scs8hd_decap_3  PHY_1004
timestamp 1586364061
transform 1 0 1104 0 -1 275808
box -38 -48 314 592
use scs8hd_decap_3  PHY_1006
timestamp 1586364061
transform 1 0 1104 0 1 275808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_502_3
timestamp 1586364061
transform 1 0 1380 0 -1 275808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_502_15
timestamp 1586364061
transform 1 0 2484 0 -1 275808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_503_3
timestamp 1586364061
transform 1 0 1380 0 1 275808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_503_15
timestamp 1586364061
transform 1 0 2484 0 1 275808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1711
timestamp 1586364061
transform 1 0 3956 0 -1 275808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_502_27
timestamp 1586364061
transform 1 0 3588 0 -1 275808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_502_32
timestamp 1586364061
transform 1 0 4048 0 -1 275808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_503_27
timestamp 1586364061
transform 1 0 3588 0 1 275808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_502_44
timestamp 1586364061
transform 1 0 5152 0 -1 275808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_503_39
timestamp 1586364061
transform 1 0 4692 0 1 275808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_503_51
timestamp 1586364061
transform 1 0 5796 0 1 275808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1712
timestamp 1586364061
transform 1 0 6716 0 1 275808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_502_56
timestamp 1586364061
transform 1 0 6256 0 -1 275808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_502_68
timestamp 1586364061
transform 1 0 7360 0 -1 275808
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_503_59
timestamp 1586364061
transform 1 0 6532 0 1 275808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_503_62
timestamp 1586364061
transform 1 0 6808 0 1 275808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1005
timestamp 1586364061
transform -1 0 8832 0 -1 275808
box -38 -48 314 592
use scs8hd_decap_3  PHY_1007
timestamp 1586364061
transform -1 0 8832 0 1 275808
box -38 -48 314 592
use scs8hd_fill_1  FILLER_502_80
timestamp 1586364061
transform 1 0 8464 0 -1 275808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_503_74
timestamp 1586364061
transform 1 0 7912 0 1 275808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_503_80
timestamp 1586364061
transform 1 0 8464 0 1 275808
box -38 -48 130 592
use scs8hd_decap_3  PHY_1008
timestamp 1586364061
transform 1 0 1104 0 -1 276896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_504_3
timestamp 1586364061
transform 1 0 1380 0 -1 276896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_504_15
timestamp 1586364061
transform 1 0 2484 0 -1 276896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1713
timestamp 1586364061
transform 1 0 3956 0 -1 276896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_504_27
timestamp 1586364061
transform 1 0 3588 0 -1 276896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_504_32
timestamp 1586364061
transform 1 0 4048 0 -1 276896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_504_44
timestamp 1586364061
transform 1 0 5152 0 -1 276896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_504_56
timestamp 1586364061
transform 1 0 6256 0 -1 276896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_504_68
timestamp 1586364061
transform 1 0 7360 0 -1 276896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1009
timestamp 1586364061
transform -1 0 8832 0 -1 276896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_504_80
timestamp 1586364061
transform 1 0 8464 0 -1 276896
box -38 -48 130 592
use scs8hd_decap_3  PHY_1010
timestamp 1586364061
transform 1 0 1104 0 1 276896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_505_3
timestamp 1586364061
transform 1 0 1380 0 1 276896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_505_15
timestamp 1586364061
transform 1 0 2484 0 1 276896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_505_27
timestamp 1586364061
transform 1 0 3588 0 1 276896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_505_39
timestamp 1586364061
transform 1 0 4692 0 1 276896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_505_51
timestamp 1586364061
transform 1 0 5796 0 1 276896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1714
timestamp 1586364061
transform 1 0 6716 0 1 276896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_505_59
timestamp 1586364061
transform 1 0 6532 0 1 276896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_505_62
timestamp 1586364061
transform 1 0 6808 0 1 276896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1011
timestamp 1586364061
transform -1 0 8832 0 1 276896
box -38 -48 314 592
use scs8hd_decap_6  FILLER_505_74
timestamp 1586364061
transform 1 0 7912 0 1 276896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_505_80
timestamp 1586364061
transform 1 0 8464 0 1 276896
box -38 -48 130 592
use scs8hd_decap_3  PHY_1012
timestamp 1586364061
transform 1 0 1104 0 -1 277984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_506_3
timestamp 1586364061
transform 1 0 1380 0 -1 277984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_506_15
timestamp 1586364061
transform 1 0 2484 0 -1 277984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1715
timestamp 1586364061
transform 1 0 3956 0 -1 277984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_506_27
timestamp 1586364061
transform 1 0 3588 0 -1 277984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_506_32
timestamp 1586364061
transform 1 0 4048 0 -1 277984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_506_44
timestamp 1586364061
transform 1 0 5152 0 -1 277984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_506_56
timestamp 1586364061
transform 1 0 6256 0 -1 277984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_506_68
timestamp 1586364061
transform 1 0 7360 0 -1 277984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1013
timestamp 1586364061
transform -1 0 8832 0 -1 277984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_506_80
timestamp 1586364061
transform 1 0 8464 0 -1 277984
box -38 -48 130 592
use scs8hd_decap_3  PHY_1014
timestamp 1586364061
transform 1 0 1104 0 1 277984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_507_3
timestamp 1586364061
transform 1 0 1380 0 1 277984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_507_15
timestamp 1586364061
transform 1 0 2484 0 1 277984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_507_27
timestamp 1586364061
transform 1 0 3588 0 1 277984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_507_39
timestamp 1586364061
transform 1 0 4692 0 1 277984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_507_51
timestamp 1586364061
transform 1 0 5796 0 1 277984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1716
timestamp 1586364061
transform 1 0 6716 0 1 277984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_507_59
timestamp 1586364061
transform 1 0 6532 0 1 277984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_507_62
timestamp 1586364061
transform 1 0 6808 0 1 277984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1015
timestamp 1586364061
transform -1 0 8832 0 1 277984
box -38 -48 314 592
use scs8hd_decap_6  FILLER_507_74
timestamp 1586364061
transform 1 0 7912 0 1 277984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_507_80
timestamp 1586364061
transform 1 0 8464 0 1 277984
box -38 -48 130 592
use scs8hd_decap_3  PHY_1016
timestamp 1586364061
transform 1 0 1104 0 -1 279072
box -38 -48 314 592
use scs8hd_decap_3  PHY_1018
timestamp 1586364061
transform 1 0 1104 0 1 279072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_508_3
timestamp 1586364061
transform 1 0 1380 0 -1 279072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_508_15
timestamp 1586364061
transform 1 0 2484 0 -1 279072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_509_3
timestamp 1586364061
transform 1 0 1380 0 1 279072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_509_15
timestamp 1586364061
transform 1 0 2484 0 1 279072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1717
timestamp 1586364061
transform 1 0 3956 0 -1 279072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_508_27
timestamp 1586364061
transform 1 0 3588 0 -1 279072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_508_32
timestamp 1586364061
transform 1 0 4048 0 -1 279072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_509_27
timestamp 1586364061
transform 1 0 3588 0 1 279072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_508_44
timestamp 1586364061
transform 1 0 5152 0 -1 279072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_509_39
timestamp 1586364061
transform 1 0 4692 0 1 279072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_509_51
timestamp 1586364061
transform 1 0 5796 0 1 279072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1718
timestamp 1586364061
transform 1 0 6716 0 1 279072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_508_56
timestamp 1586364061
transform 1 0 6256 0 -1 279072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_508_68
timestamp 1586364061
transform 1 0 7360 0 -1 279072
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_509_59
timestamp 1586364061
transform 1 0 6532 0 1 279072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_509_62
timestamp 1586364061
transform 1 0 6808 0 1 279072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1017
timestamp 1586364061
transform -1 0 8832 0 -1 279072
box -38 -48 314 592
use scs8hd_decap_3  PHY_1019
timestamp 1586364061
transform -1 0 8832 0 1 279072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_508_80
timestamp 1586364061
transform 1 0 8464 0 -1 279072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_509_74
timestamp 1586364061
transform 1 0 7912 0 1 279072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_509_80
timestamp 1586364061
transform 1 0 8464 0 1 279072
box -38 -48 130 592
use scs8hd_decap_3  PHY_1020
timestamp 1586364061
transform 1 0 1104 0 -1 280160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_510_3
timestamp 1586364061
transform 1 0 1380 0 -1 280160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_510_15
timestamp 1586364061
transform 1 0 2484 0 -1 280160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1719
timestamp 1586364061
transform 1 0 3956 0 -1 280160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_510_27
timestamp 1586364061
transform 1 0 3588 0 -1 280160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_510_32
timestamp 1586364061
transform 1 0 4048 0 -1 280160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_510_44
timestamp 1586364061
transform 1 0 5152 0 -1 280160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_510_56
timestamp 1586364061
transform 1 0 6256 0 -1 280160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_510_68
timestamp 1586364061
transform 1 0 7360 0 -1 280160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1021
timestamp 1586364061
transform -1 0 8832 0 -1 280160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_510_80
timestamp 1586364061
transform 1 0 8464 0 -1 280160
box -38 -48 130 592
use scs8hd_decap_3  PHY_1022
timestamp 1586364061
transform 1 0 1104 0 1 280160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_511_3
timestamp 1586364061
transform 1 0 1380 0 1 280160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_511_15
timestamp 1586364061
transform 1 0 2484 0 1 280160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_511_27
timestamp 1586364061
transform 1 0 3588 0 1 280160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_511_39
timestamp 1586364061
transform 1 0 4692 0 1 280160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_511_51
timestamp 1586364061
transform 1 0 5796 0 1 280160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1720
timestamp 1586364061
transform 1 0 6716 0 1 280160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_511_59
timestamp 1586364061
transform 1 0 6532 0 1 280160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_511_62
timestamp 1586364061
transform 1 0 6808 0 1 280160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1023
timestamp 1586364061
transform -1 0 8832 0 1 280160
box -38 -48 314 592
use scs8hd_decap_6  FILLER_511_74
timestamp 1586364061
transform 1 0 7912 0 1 280160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_511_80
timestamp 1586364061
transform 1 0 8464 0 1 280160
box -38 -48 130 592
use scs8hd_decap_3  PHY_1024
timestamp 1586364061
transform 1 0 1104 0 -1 281248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_512_3
timestamp 1586364061
transform 1 0 1380 0 -1 281248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_512_15
timestamp 1586364061
transform 1 0 2484 0 -1 281248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1721
timestamp 1586364061
transform 1 0 3956 0 -1 281248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_512_27
timestamp 1586364061
transform 1 0 3588 0 -1 281248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_512_32
timestamp 1586364061
transform 1 0 4048 0 -1 281248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_512_44
timestamp 1586364061
transform 1 0 5152 0 -1 281248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_512_56
timestamp 1586364061
transform 1 0 6256 0 -1 281248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_512_68
timestamp 1586364061
transform 1 0 7360 0 -1 281248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1025
timestamp 1586364061
transform -1 0 8832 0 -1 281248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_512_80
timestamp 1586364061
transform 1 0 8464 0 -1 281248
box -38 -48 130 592
use scs8hd_decap_3  PHY_1026
timestamp 1586364061
transform 1 0 1104 0 1 281248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_513_3
timestamp 1586364061
transform 1 0 1380 0 1 281248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_513_15
timestamp 1586364061
transform 1 0 2484 0 1 281248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_513_27
timestamp 1586364061
transform 1 0 3588 0 1 281248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_513_39
timestamp 1586364061
transform 1 0 4692 0 1 281248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_513_51
timestamp 1586364061
transform 1 0 5796 0 1 281248
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1722
timestamp 1586364061
transform 1 0 6716 0 1 281248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_513_59
timestamp 1586364061
transform 1 0 6532 0 1 281248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_513_62
timestamp 1586364061
transform 1 0 6808 0 1 281248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1027
timestamp 1586364061
transform -1 0 8832 0 1 281248
box -38 -48 314 592
use scs8hd_decap_6  FILLER_513_74
timestamp 1586364061
transform 1 0 7912 0 1 281248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_513_80
timestamp 1586364061
transform 1 0 8464 0 1 281248
box -38 -48 130 592
use scs8hd_decap_3  PHY_1028
timestamp 1586364061
transform 1 0 1104 0 -1 282336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_514_3
timestamp 1586364061
transform 1 0 1380 0 -1 282336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_514_15
timestamp 1586364061
transform 1 0 2484 0 -1 282336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1723
timestamp 1586364061
transform 1 0 3956 0 -1 282336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_514_27
timestamp 1586364061
transform 1 0 3588 0 -1 282336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_514_32
timestamp 1586364061
transform 1 0 4048 0 -1 282336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_514_44
timestamp 1586364061
transform 1 0 5152 0 -1 282336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_514_56
timestamp 1586364061
transform 1 0 6256 0 -1 282336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_514_68
timestamp 1586364061
transform 1 0 7360 0 -1 282336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1029
timestamp 1586364061
transform -1 0 8832 0 -1 282336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_514_80
timestamp 1586364061
transform 1 0 8464 0 -1 282336
box -38 -48 130 592
use scs8hd_decap_3  PHY_1030
timestamp 1586364061
transform 1 0 1104 0 1 282336
box -38 -48 314 592
use scs8hd_decap_3  PHY_1032
timestamp 1586364061
transform 1 0 1104 0 -1 283424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_515_3
timestamp 1586364061
transform 1 0 1380 0 1 282336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_515_15
timestamp 1586364061
transform 1 0 2484 0 1 282336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_516_3
timestamp 1586364061
transform 1 0 1380 0 -1 283424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_516_15
timestamp 1586364061
transform 1 0 2484 0 -1 283424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1725
timestamp 1586364061
transform 1 0 3956 0 -1 283424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_515_27
timestamp 1586364061
transform 1 0 3588 0 1 282336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_516_27
timestamp 1586364061
transform 1 0 3588 0 -1 283424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_516_32
timestamp 1586364061
transform 1 0 4048 0 -1 283424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_515_39
timestamp 1586364061
transform 1 0 4692 0 1 282336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_515_51
timestamp 1586364061
transform 1 0 5796 0 1 282336
box -38 -48 774 592
use scs8hd_decap_12  FILLER_516_44
timestamp 1586364061
transform 1 0 5152 0 -1 283424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1724
timestamp 1586364061
transform 1 0 6716 0 1 282336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_515_59
timestamp 1586364061
transform 1 0 6532 0 1 282336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_515_62
timestamp 1586364061
transform 1 0 6808 0 1 282336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_516_56
timestamp 1586364061
transform 1 0 6256 0 -1 283424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_516_68
timestamp 1586364061
transform 1 0 7360 0 -1 283424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1031
timestamp 1586364061
transform -1 0 8832 0 1 282336
box -38 -48 314 592
use scs8hd_decap_3  PHY_1033
timestamp 1586364061
transform -1 0 8832 0 -1 283424
box -38 -48 314 592
use scs8hd_decap_6  FILLER_515_74
timestamp 1586364061
transform 1 0 7912 0 1 282336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_515_80
timestamp 1586364061
transform 1 0 8464 0 1 282336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_516_80
timestamp 1586364061
transform 1 0 8464 0 -1 283424
box -38 -48 130 592
use scs8hd_decap_3  PHY_1034
timestamp 1586364061
transform 1 0 1104 0 1 283424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_517_3
timestamp 1586364061
transform 1 0 1380 0 1 283424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_517_15
timestamp 1586364061
transform 1 0 2484 0 1 283424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_517_27
timestamp 1586364061
transform 1 0 3588 0 1 283424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_517_39
timestamp 1586364061
transform 1 0 4692 0 1 283424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_517_51
timestamp 1586364061
transform 1 0 5796 0 1 283424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1726
timestamp 1586364061
transform 1 0 6716 0 1 283424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_517_59
timestamp 1586364061
transform 1 0 6532 0 1 283424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_517_62
timestamp 1586364061
transform 1 0 6808 0 1 283424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1035
timestamp 1586364061
transform -1 0 8832 0 1 283424
box -38 -48 314 592
use scs8hd_decap_6  FILLER_517_74
timestamp 1586364061
transform 1 0 7912 0 1 283424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_517_80
timestamp 1586364061
transform 1 0 8464 0 1 283424
box -38 -48 130 592
use scs8hd_decap_3  PHY_1036
timestamp 1586364061
transform 1 0 1104 0 -1 284512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_518_3
timestamp 1586364061
transform 1 0 1380 0 -1 284512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_518_15
timestamp 1586364061
transform 1 0 2484 0 -1 284512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1727
timestamp 1586364061
transform 1 0 3956 0 -1 284512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_518_27
timestamp 1586364061
transform 1 0 3588 0 -1 284512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_518_32
timestamp 1586364061
transform 1 0 4048 0 -1 284512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_518_44
timestamp 1586364061
transform 1 0 5152 0 -1 284512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_518_56
timestamp 1586364061
transform 1 0 6256 0 -1 284512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_518_68
timestamp 1586364061
transform 1 0 7360 0 -1 284512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1037
timestamp 1586364061
transform -1 0 8832 0 -1 284512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_518_80
timestamp 1586364061
transform 1 0 8464 0 -1 284512
box -38 -48 130 592
use scs8hd_decap_3  PHY_1038
timestamp 1586364061
transform 1 0 1104 0 1 284512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_519_3
timestamp 1586364061
transform 1 0 1380 0 1 284512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_519_15
timestamp 1586364061
transform 1 0 2484 0 1 284512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_519_27
timestamp 1586364061
transform 1 0 3588 0 1 284512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_519_39
timestamp 1586364061
transform 1 0 4692 0 1 284512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_519_51
timestamp 1586364061
transform 1 0 5796 0 1 284512
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1728
timestamp 1586364061
transform 1 0 6716 0 1 284512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_519_59
timestamp 1586364061
transform 1 0 6532 0 1 284512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_519_62
timestamp 1586364061
transform 1 0 6808 0 1 284512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1039
timestamp 1586364061
transform -1 0 8832 0 1 284512
box -38 -48 314 592
use scs8hd_decap_6  FILLER_519_74
timestamp 1586364061
transform 1 0 7912 0 1 284512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_519_80
timestamp 1586364061
transform 1 0 8464 0 1 284512
box -38 -48 130 592
use scs8hd_decap_3  PHY_1040
timestamp 1586364061
transform 1 0 1104 0 -1 285600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_520_3
timestamp 1586364061
transform 1 0 1380 0 -1 285600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_520_15
timestamp 1586364061
transform 1 0 2484 0 -1 285600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1729
timestamp 1586364061
transform 1 0 3956 0 -1 285600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_520_27
timestamp 1586364061
transform 1 0 3588 0 -1 285600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_520_32
timestamp 1586364061
transform 1 0 4048 0 -1 285600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_520_44
timestamp 1586364061
transform 1 0 5152 0 -1 285600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_520_56
timestamp 1586364061
transform 1 0 6256 0 -1 285600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_520_68
timestamp 1586364061
transform 1 0 7360 0 -1 285600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1041
timestamp 1586364061
transform -1 0 8832 0 -1 285600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_520_80
timestamp 1586364061
transform 1 0 8464 0 -1 285600
box -38 -48 130 592
use scs8hd_decap_3  PHY_1042
timestamp 1586364061
transform 1 0 1104 0 1 285600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_521_3
timestamp 1586364061
transform 1 0 1380 0 1 285600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_521_15
timestamp 1586364061
transform 1 0 2484 0 1 285600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_521_27
timestamp 1586364061
transform 1 0 3588 0 1 285600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_521_39
timestamp 1586364061
transform 1 0 4692 0 1 285600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_521_51
timestamp 1586364061
transform 1 0 5796 0 1 285600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1730
timestamp 1586364061
transform 1 0 6716 0 1 285600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_521_59
timestamp 1586364061
transform 1 0 6532 0 1 285600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_521_62
timestamp 1586364061
transform 1 0 6808 0 1 285600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1043
timestamp 1586364061
transform -1 0 8832 0 1 285600
box -38 -48 314 592
use scs8hd_decap_6  FILLER_521_74
timestamp 1586364061
transform 1 0 7912 0 1 285600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_521_80
timestamp 1586364061
transform 1 0 8464 0 1 285600
box -38 -48 130 592
use scs8hd_decap_3  PHY_1044
timestamp 1586364061
transform 1 0 1104 0 -1 286688
box -38 -48 314 592
use scs8hd_decap_3  PHY_1046
timestamp 1586364061
transform 1 0 1104 0 1 286688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_522_3
timestamp 1586364061
transform 1 0 1380 0 -1 286688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_522_15
timestamp 1586364061
transform 1 0 2484 0 -1 286688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_523_3
timestamp 1586364061
transform 1 0 1380 0 1 286688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_523_15
timestamp 1586364061
transform 1 0 2484 0 1 286688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1731
timestamp 1586364061
transform 1 0 3956 0 -1 286688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_522_27
timestamp 1586364061
transform 1 0 3588 0 -1 286688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_522_32
timestamp 1586364061
transform 1 0 4048 0 -1 286688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_523_27
timestamp 1586364061
transform 1 0 3588 0 1 286688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_522_44
timestamp 1586364061
transform 1 0 5152 0 -1 286688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_523_39
timestamp 1586364061
transform 1 0 4692 0 1 286688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_523_51
timestamp 1586364061
transform 1 0 5796 0 1 286688
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1732
timestamp 1586364061
transform 1 0 6716 0 1 286688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_522_56
timestamp 1586364061
transform 1 0 6256 0 -1 286688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_522_68
timestamp 1586364061
transform 1 0 7360 0 -1 286688
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_523_59
timestamp 1586364061
transform 1 0 6532 0 1 286688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_523_62
timestamp 1586364061
transform 1 0 6808 0 1 286688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1045
timestamp 1586364061
transform -1 0 8832 0 -1 286688
box -38 -48 314 592
use scs8hd_decap_3  PHY_1047
timestamp 1586364061
transform -1 0 8832 0 1 286688
box -38 -48 314 592
use scs8hd_fill_1  FILLER_522_80
timestamp 1586364061
transform 1 0 8464 0 -1 286688
box -38 -48 130 592
use scs8hd_decap_6  FILLER_523_74
timestamp 1586364061
transform 1 0 7912 0 1 286688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_523_80
timestamp 1586364061
transform 1 0 8464 0 1 286688
box -38 -48 130 592
use scs8hd_decap_3  PHY_1048
timestamp 1586364061
transform 1 0 1104 0 -1 287776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_524_3
timestamp 1586364061
transform 1 0 1380 0 -1 287776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_524_15
timestamp 1586364061
transform 1 0 2484 0 -1 287776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1733
timestamp 1586364061
transform 1 0 3956 0 -1 287776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_524_27
timestamp 1586364061
transform 1 0 3588 0 -1 287776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_524_32
timestamp 1586364061
transform 1 0 4048 0 -1 287776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_524_44
timestamp 1586364061
transform 1 0 5152 0 -1 287776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_524_56
timestamp 1586364061
transform 1 0 6256 0 -1 287776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_524_68
timestamp 1586364061
transform 1 0 7360 0 -1 287776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1049
timestamp 1586364061
transform -1 0 8832 0 -1 287776
box -38 -48 314 592
use scs8hd_fill_1  FILLER_524_80
timestamp 1586364061
transform 1 0 8464 0 -1 287776
box -38 -48 130 592
use scs8hd_decap_3  PHY_1050
timestamp 1586364061
transform 1 0 1104 0 1 287776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_525_3
timestamp 1586364061
transform 1 0 1380 0 1 287776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_525_15
timestamp 1586364061
transform 1 0 2484 0 1 287776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_525_27
timestamp 1586364061
transform 1 0 3588 0 1 287776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_525_39
timestamp 1586364061
transform 1 0 4692 0 1 287776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_525_51
timestamp 1586364061
transform 1 0 5796 0 1 287776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1734
timestamp 1586364061
transform 1 0 6716 0 1 287776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_525_59
timestamp 1586364061
transform 1 0 6532 0 1 287776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_525_62
timestamp 1586364061
transform 1 0 6808 0 1 287776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1051
timestamp 1586364061
transform -1 0 8832 0 1 287776
box -38 -48 314 592
use scs8hd_decap_6  FILLER_525_74
timestamp 1586364061
transform 1 0 7912 0 1 287776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_525_80
timestamp 1586364061
transform 1 0 8464 0 1 287776
box -38 -48 130 592
use scs8hd_decap_3  PHY_1052
timestamp 1586364061
transform 1 0 1104 0 -1 288864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_526_3
timestamp 1586364061
transform 1 0 1380 0 -1 288864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_526_15
timestamp 1586364061
transform 1 0 2484 0 -1 288864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1735
timestamp 1586364061
transform 1 0 3956 0 -1 288864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_526_27
timestamp 1586364061
transform 1 0 3588 0 -1 288864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_526_32
timestamp 1586364061
transform 1 0 4048 0 -1 288864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_526_44
timestamp 1586364061
transform 1 0 5152 0 -1 288864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_526_56
timestamp 1586364061
transform 1 0 6256 0 -1 288864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_526_68
timestamp 1586364061
transform 1 0 7360 0 -1 288864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1053
timestamp 1586364061
transform -1 0 8832 0 -1 288864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_526_80
timestamp 1586364061
transform 1 0 8464 0 -1 288864
box -38 -48 130 592
use scs8hd_decap_3  PHY_1054
timestamp 1586364061
transform 1 0 1104 0 1 288864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_527_3
timestamp 1586364061
transform 1 0 1380 0 1 288864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_527_15
timestamp 1586364061
transform 1 0 2484 0 1 288864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_527_27
timestamp 1586364061
transform 1 0 3588 0 1 288864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_527_39
timestamp 1586364061
transform 1 0 4692 0 1 288864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_527_51
timestamp 1586364061
transform 1 0 5796 0 1 288864
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1736
timestamp 1586364061
transform 1 0 6716 0 1 288864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_527_59
timestamp 1586364061
transform 1 0 6532 0 1 288864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_527_62
timestamp 1586364061
transform 1 0 6808 0 1 288864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1055
timestamp 1586364061
transform -1 0 8832 0 1 288864
box -38 -48 314 592
use scs8hd_decap_6  FILLER_527_74
timestamp 1586364061
transform 1 0 7912 0 1 288864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_527_80
timestamp 1586364061
transform 1 0 8464 0 1 288864
box -38 -48 130 592
use scs8hd_decap_3  PHY_1056
timestamp 1586364061
transform 1 0 1104 0 -1 289952
box -38 -48 314 592
use scs8hd_decap_3  PHY_1058
timestamp 1586364061
transform 1 0 1104 0 1 289952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_528_3
timestamp 1586364061
transform 1 0 1380 0 -1 289952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_528_15
timestamp 1586364061
transform 1 0 2484 0 -1 289952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_529_3
timestamp 1586364061
transform 1 0 1380 0 1 289952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_529_15
timestamp 1586364061
transform 1 0 2484 0 1 289952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1737
timestamp 1586364061
transform 1 0 3956 0 -1 289952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_528_27
timestamp 1586364061
transform 1 0 3588 0 -1 289952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_528_32
timestamp 1586364061
transform 1 0 4048 0 -1 289952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_529_27
timestamp 1586364061
transform 1 0 3588 0 1 289952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_528_44
timestamp 1586364061
transform 1 0 5152 0 -1 289952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_529_39
timestamp 1586364061
transform 1 0 4692 0 1 289952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_529_51
timestamp 1586364061
transform 1 0 5796 0 1 289952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1738
timestamp 1586364061
transform 1 0 6716 0 1 289952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_528_56
timestamp 1586364061
transform 1 0 6256 0 -1 289952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_528_68
timestamp 1586364061
transform 1 0 7360 0 -1 289952
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_529_59
timestamp 1586364061
transform 1 0 6532 0 1 289952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_529_62
timestamp 1586364061
transform 1 0 6808 0 1 289952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1057
timestamp 1586364061
transform -1 0 8832 0 -1 289952
box -38 -48 314 592
use scs8hd_decap_3  PHY_1059
timestamp 1586364061
transform -1 0 8832 0 1 289952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_528_80
timestamp 1586364061
transform 1 0 8464 0 -1 289952
box -38 -48 130 592
use scs8hd_decap_6  FILLER_529_74
timestamp 1586364061
transform 1 0 7912 0 1 289952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_529_80
timestamp 1586364061
transform 1 0 8464 0 1 289952
box -38 -48 130 592
use scs8hd_decap_3  PHY_1060
timestamp 1586364061
transform 1 0 1104 0 -1 291040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_530_3
timestamp 1586364061
transform 1 0 1380 0 -1 291040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_530_15
timestamp 1586364061
transform 1 0 2484 0 -1 291040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1739
timestamp 1586364061
transform 1 0 3956 0 -1 291040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_530_27
timestamp 1586364061
transform 1 0 3588 0 -1 291040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_530_32
timestamp 1586364061
transform 1 0 4048 0 -1 291040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_530_44
timestamp 1586364061
transform 1 0 5152 0 -1 291040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_530_56
timestamp 1586364061
transform 1 0 6256 0 -1 291040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_530_68
timestamp 1586364061
transform 1 0 7360 0 -1 291040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1061
timestamp 1586364061
transform -1 0 8832 0 -1 291040
box -38 -48 314 592
use scs8hd_fill_1  FILLER_530_80
timestamp 1586364061
transform 1 0 8464 0 -1 291040
box -38 -48 130 592
use scs8hd_decap_3  PHY_1062
timestamp 1586364061
transform 1 0 1104 0 1 291040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_531_3
timestamp 1586364061
transform 1 0 1380 0 1 291040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_531_15
timestamp 1586364061
transform 1 0 2484 0 1 291040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_531_27
timestamp 1586364061
transform 1 0 3588 0 1 291040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_531_39
timestamp 1586364061
transform 1 0 4692 0 1 291040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_531_51
timestamp 1586364061
transform 1 0 5796 0 1 291040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1740
timestamp 1586364061
transform 1 0 6716 0 1 291040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_531_59
timestamp 1586364061
transform 1 0 6532 0 1 291040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_531_62
timestamp 1586364061
transform 1 0 6808 0 1 291040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1063
timestamp 1586364061
transform -1 0 8832 0 1 291040
box -38 -48 314 592
use scs8hd_decap_6  FILLER_531_74
timestamp 1586364061
transform 1 0 7912 0 1 291040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_531_80
timestamp 1586364061
transform 1 0 8464 0 1 291040
box -38 -48 130 592
use scs8hd_decap_3  PHY_1064
timestamp 1586364061
transform 1 0 1104 0 -1 292128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_532_3
timestamp 1586364061
transform 1 0 1380 0 -1 292128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_532_15
timestamp 1586364061
transform 1 0 2484 0 -1 292128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1741
timestamp 1586364061
transform 1 0 3956 0 -1 292128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_532_27
timestamp 1586364061
transform 1 0 3588 0 -1 292128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_532_32
timestamp 1586364061
transform 1 0 4048 0 -1 292128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_532_44
timestamp 1586364061
transform 1 0 5152 0 -1 292128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_532_56
timestamp 1586364061
transform 1 0 6256 0 -1 292128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_532_68
timestamp 1586364061
transform 1 0 7360 0 -1 292128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1065
timestamp 1586364061
transform -1 0 8832 0 -1 292128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_532_80
timestamp 1586364061
transform 1 0 8464 0 -1 292128
box -38 -48 130 592
use scs8hd_decap_3  PHY_1066
timestamp 1586364061
transform 1 0 1104 0 1 292128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_533_3
timestamp 1586364061
transform 1 0 1380 0 1 292128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_533_15
timestamp 1586364061
transform 1 0 2484 0 1 292128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_533_27
timestamp 1586364061
transform 1 0 3588 0 1 292128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_533_39
timestamp 1586364061
transform 1 0 4692 0 1 292128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_533_51
timestamp 1586364061
transform 1 0 5796 0 1 292128
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1742
timestamp 1586364061
transform 1 0 6716 0 1 292128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_533_59
timestamp 1586364061
transform 1 0 6532 0 1 292128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_533_62
timestamp 1586364061
transform 1 0 6808 0 1 292128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1067
timestamp 1586364061
transform -1 0 8832 0 1 292128
box -38 -48 314 592
use scs8hd_decap_6  FILLER_533_74
timestamp 1586364061
transform 1 0 7912 0 1 292128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_533_80
timestamp 1586364061
transform 1 0 8464 0 1 292128
box -38 -48 130 592
use scs8hd_decap_3  PHY_1068
timestamp 1586364061
transform 1 0 1104 0 -1 293216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_534_3
timestamp 1586364061
transform 1 0 1380 0 -1 293216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_534_15
timestamp 1586364061
transform 1 0 2484 0 -1 293216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1743
timestamp 1586364061
transform 1 0 3956 0 -1 293216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_534_27
timestamp 1586364061
transform 1 0 3588 0 -1 293216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_534_32
timestamp 1586364061
transform 1 0 4048 0 -1 293216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_534_44
timestamp 1586364061
transform 1 0 5152 0 -1 293216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_534_56
timestamp 1586364061
transform 1 0 6256 0 -1 293216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_534_68
timestamp 1586364061
transform 1 0 7360 0 -1 293216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1069
timestamp 1586364061
transform -1 0 8832 0 -1 293216
box -38 -48 314 592
use scs8hd_fill_1  FILLER_534_80
timestamp 1586364061
transform 1 0 8464 0 -1 293216
box -38 -48 130 592
use scs8hd_decap_3  PHY_1070
timestamp 1586364061
transform 1 0 1104 0 1 293216
box -38 -48 314 592
use scs8hd_decap_3  PHY_1072
timestamp 1586364061
transform 1 0 1104 0 -1 294304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_535_3
timestamp 1586364061
transform 1 0 1380 0 1 293216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_535_15
timestamp 1586364061
transform 1 0 2484 0 1 293216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_536_3
timestamp 1586364061
transform 1 0 1380 0 -1 294304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_536_15
timestamp 1586364061
transform 1 0 2484 0 -1 294304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1745
timestamp 1586364061
transform 1 0 3956 0 -1 294304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_535_27
timestamp 1586364061
transform 1 0 3588 0 1 293216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_536_27
timestamp 1586364061
transform 1 0 3588 0 -1 294304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_536_32
timestamp 1586364061
transform 1 0 4048 0 -1 294304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_535_39
timestamp 1586364061
transform 1 0 4692 0 1 293216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_535_51
timestamp 1586364061
transform 1 0 5796 0 1 293216
box -38 -48 774 592
use scs8hd_decap_12  FILLER_536_44
timestamp 1586364061
transform 1 0 5152 0 -1 294304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1744
timestamp 1586364061
transform 1 0 6716 0 1 293216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_535_59
timestamp 1586364061
transform 1 0 6532 0 1 293216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_535_62
timestamp 1586364061
transform 1 0 6808 0 1 293216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_536_56
timestamp 1586364061
transform 1 0 6256 0 -1 294304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_536_68
timestamp 1586364061
transform 1 0 7360 0 -1 294304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1071
timestamp 1586364061
transform -1 0 8832 0 1 293216
box -38 -48 314 592
use scs8hd_decap_3  PHY_1073
timestamp 1586364061
transform -1 0 8832 0 -1 294304
box -38 -48 314 592
use scs8hd_decap_6  FILLER_535_74
timestamp 1586364061
transform 1 0 7912 0 1 293216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_535_80
timestamp 1586364061
transform 1 0 8464 0 1 293216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_536_80
timestamp 1586364061
transform 1 0 8464 0 -1 294304
box -38 -48 130 592
use scs8hd_decap_3  PHY_1074
timestamp 1586364061
transform 1 0 1104 0 1 294304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_537_3
timestamp 1586364061
transform 1 0 1380 0 1 294304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_537_15
timestamp 1586364061
transform 1 0 2484 0 1 294304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_537_27
timestamp 1586364061
transform 1 0 3588 0 1 294304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_537_39
timestamp 1586364061
transform 1 0 4692 0 1 294304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_537_51
timestamp 1586364061
transform 1 0 5796 0 1 294304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1746
timestamp 1586364061
transform 1 0 6716 0 1 294304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_537_59
timestamp 1586364061
transform 1 0 6532 0 1 294304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_537_62
timestamp 1586364061
transform 1 0 6808 0 1 294304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1075
timestamp 1586364061
transform -1 0 8832 0 1 294304
box -38 -48 314 592
use scs8hd_decap_6  FILLER_537_74
timestamp 1586364061
transform 1 0 7912 0 1 294304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_537_80
timestamp 1586364061
transform 1 0 8464 0 1 294304
box -38 -48 130 592
use scs8hd_decap_3  PHY_1076
timestamp 1586364061
transform 1 0 1104 0 -1 295392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_538_3
timestamp 1586364061
transform 1 0 1380 0 -1 295392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_538_15
timestamp 1586364061
transform 1 0 2484 0 -1 295392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1747
timestamp 1586364061
transform 1 0 3956 0 -1 295392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_538_27
timestamp 1586364061
transform 1 0 3588 0 -1 295392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_538_32
timestamp 1586364061
transform 1 0 4048 0 -1 295392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_538_44
timestamp 1586364061
transform 1 0 5152 0 -1 295392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_538_56
timestamp 1586364061
transform 1 0 6256 0 -1 295392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_538_68
timestamp 1586364061
transform 1 0 7360 0 -1 295392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1077
timestamp 1586364061
transform -1 0 8832 0 -1 295392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_538_80
timestamp 1586364061
transform 1 0 8464 0 -1 295392
box -38 -48 130 592
use scs8hd_decap_3  PHY_1078
timestamp 1586364061
transform 1 0 1104 0 1 295392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_539_3
timestamp 1586364061
transform 1 0 1380 0 1 295392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_539_15
timestamp 1586364061
transform 1 0 2484 0 1 295392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_539_27
timestamp 1586364061
transform 1 0 3588 0 1 295392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_539_39
timestamp 1586364061
transform 1 0 4692 0 1 295392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_539_51
timestamp 1586364061
transform 1 0 5796 0 1 295392
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1748
timestamp 1586364061
transform 1 0 6716 0 1 295392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_539_59
timestamp 1586364061
transform 1 0 6532 0 1 295392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_539_62
timestamp 1586364061
transform 1 0 6808 0 1 295392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1079
timestamp 1586364061
transform -1 0 8832 0 1 295392
box -38 -48 314 592
use scs8hd_decap_6  FILLER_539_74
timestamp 1586364061
transform 1 0 7912 0 1 295392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_539_80
timestamp 1586364061
transform 1 0 8464 0 1 295392
box -38 -48 130 592
use scs8hd_decap_3  PHY_1080
timestamp 1586364061
transform 1 0 1104 0 -1 296480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_540_3
timestamp 1586364061
transform 1 0 1380 0 -1 296480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_540_15
timestamp 1586364061
transform 1 0 2484 0 -1 296480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1749
timestamp 1586364061
transform 1 0 3956 0 -1 296480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_540_27
timestamp 1586364061
transform 1 0 3588 0 -1 296480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_540_32
timestamp 1586364061
transform 1 0 4048 0 -1 296480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_540_44
timestamp 1586364061
transform 1 0 5152 0 -1 296480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_540_56
timestamp 1586364061
transform 1 0 6256 0 -1 296480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_540_68
timestamp 1586364061
transform 1 0 7360 0 -1 296480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1081
timestamp 1586364061
transform -1 0 8832 0 -1 296480
box -38 -48 314 592
use scs8hd_fill_1  FILLER_540_80
timestamp 1586364061
transform 1 0 8464 0 -1 296480
box -38 -48 130 592
use scs8hd_decap_3  PHY_1082
timestamp 1586364061
transform 1 0 1104 0 1 296480
box -38 -48 314 592
use scs8hd_decap_3  PHY_1084
timestamp 1586364061
transform 1 0 1104 0 -1 297568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_541_3
timestamp 1586364061
transform 1 0 1380 0 1 296480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_541_15
timestamp 1586364061
transform 1 0 2484 0 1 296480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_542_3
timestamp 1586364061
transform 1 0 1380 0 -1 297568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_542_15
timestamp 1586364061
transform 1 0 2484 0 -1 297568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1751
timestamp 1586364061
transform 1 0 3956 0 -1 297568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_541_27
timestamp 1586364061
transform 1 0 3588 0 1 296480
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_542_27
timestamp 1586364061
transform 1 0 3588 0 -1 297568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_542_32
timestamp 1586364061
transform 1 0 4048 0 -1 297568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_541_39
timestamp 1586364061
transform 1 0 4692 0 1 296480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_541_51
timestamp 1586364061
transform 1 0 5796 0 1 296480
box -38 -48 774 592
use scs8hd_decap_12  FILLER_542_44
timestamp 1586364061
transform 1 0 5152 0 -1 297568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1750
timestamp 1586364061
transform 1 0 6716 0 1 296480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_541_59
timestamp 1586364061
transform 1 0 6532 0 1 296480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_541_62
timestamp 1586364061
transform 1 0 6808 0 1 296480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_542_56
timestamp 1586364061
transform 1 0 6256 0 -1 297568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_542_68
timestamp 1586364061
transform 1 0 7360 0 -1 297568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1083
timestamp 1586364061
transform -1 0 8832 0 1 296480
box -38 -48 314 592
use scs8hd_decap_3  PHY_1085
timestamp 1586364061
transform -1 0 8832 0 -1 297568
box -38 -48 314 592
use scs8hd_decap_6  FILLER_541_74
timestamp 1586364061
transform 1 0 7912 0 1 296480
box -38 -48 590 592
use scs8hd_fill_1  FILLER_541_80
timestamp 1586364061
transform 1 0 8464 0 1 296480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_542_80
timestamp 1586364061
transform 1 0 8464 0 -1 297568
box -38 -48 130 592
use scs8hd_decap_3  PHY_1086
timestamp 1586364061
transform 1 0 1104 0 1 297568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_543_3
timestamp 1586364061
transform 1 0 1380 0 1 297568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_543_15
timestamp 1586364061
transform 1 0 2484 0 1 297568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_543_27
timestamp 1586364061
transform 1 0 3588 0 1 297568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_543_39
timestamp 1586364061
transform 1 0 4692 0 1 297568
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_543_51
timestamp 1586364061
transform 1 0 5796 0 1 297568
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1752
timestamp 1586364061
transform 1 0 6716 0 1 297568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_543_59
timestamp 1586364061
transform 1 0 6532 0 1 297568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_543_62
timestamp 1586364061
transform 1 0 6808 0 1 297568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1087
timestamp 1586364061
transform -1 0 8832 0 1 297568
box -38 -48 314 592
use scs8hd_decap_6  FILLER_543_74
timestamp 1586364061
transform 1 0 7912 0 1 297568
box -38 -48 590 592
use scs8hd_fill_1  FILLER_543_80
timestamp 1586364061
transform 1 0 8464 0 1 297568
box -38 -48 130 592
use scs8hd_decap_3  PHY_1088
timestamp 1586364061
transform 1 0 1104 0 -1 298656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_544_3
timestamp 1586364061
transform 1 0 1380 0 -1 298656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_544_15
timestamp 1586364061
transform 1 0 2484 0 -1 298656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1753
timestamp 1586364061
transform 1 0 3956 0 -1 298656
box -38 -48 130 592
use scs8hd_decap_4  FILLER_544_27
timestamp 1586364061
transform 1 0 3588 0 -1 298656
box -38 -48 406 592
use scs8hd_decap_12  FILLER_544_32
timestamp 1586364061
transform 1 0 4048 0 -1 298656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_544_44
timestamp 1586364061
transform 1 0 5152 0 -1 298656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_544_56
timestamp 1586364061
transform 1 0 6256 0 -1 298656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_544_68
timestamp 1586364061
transform 1 0 7360 0 -1 298656
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1089
timestamp 1586364061
transform -1 0 8832 0 -1 298656
box -38 -48 314 592
use scs8hd_fill_1  FILLER_544_80
timestamp 1586364061
transform 1 0 8464 0 -1 298656
box -38 -48 130 592
use scs8hd_decap_3  PHY_1090
timestamp 1586364061
transform 1 0 1104 0 1 298656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_545_3
timestamp 1586364061
transform 1 0 1380 0 1 298656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_545_15
timestamp 1586364061
transform 1 0 2484 0 1 298656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_545_27
timestamp 1586364061
transform 1 0 3588 0 1 298656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_545_39
timestamp 1586364061
transform 1 0 4692 0 1 298656
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_545_51
timestamp 1586364061
transform 1 0 5796 0 1 298656
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1754
timestamp 1586364061
transform 1 0 6716 0 1 298656
box -38 -48 130 592
use scs8hd_fill_2  FILLER_545_59
timestamp 1586364061
transform 1 0 6532 0 1 298656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_545_62
timestamp 1586364061
transform 1 0 6808 0 1 298656
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1091
timestamp 1586364061
transform -1 0 8832 0 1 298656
box -38 -48 314 592
use scs8hd_decap_6  FILLER_545_74
timestamp 1586364061
transform 1 0 7912 0 1 298656
box -38 -48 590 592
use scs8hd_fill_1  FILLER_545_80
timestamp 1586364061
transform 1 0 8464 0 1 298656
box -38 -48 130 592
use scs8hd_decap_3  PHY_1092
timestamp 1586364061
transform 1 0 1104 0 -1 299744
box -38 -48 314 592
use scs8hd_decap_12  FILLER_546_3
timestamp 1586364061
transform 1 0 1380 0 -1 299744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_546_15
timestamp 1586364061
transform 1 0 2484 0 -1 299744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1755
timestamp 1586364061
transform 1 0 3956 0 -1 299744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_546_27
timestamp 1586364061
transform 1 0 3588 0 -1 299744
box -38 -48 406 592
use scs8hd_decap_12  FILLER_546_32
timestamp 1586364061
transform 1 0 4048 0 -1 299744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_546_44
timestamp 1586364061
transform 1 0 5152 0 -1 299744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_546_56
timestamp 1586364061
transform 1 0 6256 0 -1 299744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_546_68
timestamp 1586364061
transform 1 0 7360 0 -1 299744
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1093
timestamp 1586364061
transform -1 0 8832 0 -1 299744
box -38 -48 314 592
use scs8hd_fill_1  FILLER_546_80
timestamp 1586364061
transform 1 0 8464 0 -1 299744
box -38 -48 130 592
use scs8hd_decap_3  PHY_1094
timestamp 1586364061
transform 1 0 1104 0 1 299744
box -38 -48 314 592
use scs8hd_decap_12  FILLER_547_3
timestamp 1586364061
transform 1 0 1380 0 1 299744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_547_15
timestamp 1586364061
transform 1 0 2484 0 1 299744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_547_27
timestamp 1586364061
transform 1 0 3588 0 1 299744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_547_39
timestamp 1586364061
transform 1 0 4692 0 1 299744
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_547_51
timestamp 1586364061
transform 1 0 5796 0 1 299744
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1756
timestamp 1586364061
transform 1 0 6716 0 1 299744
box -38 -48 130 592
use scs8hd_fill_2  FILLER_547_59
timestamp 1586364061
transform 1 0 6532 0 1 299744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_547_62
timestamp 1586364061
transform 1 0 6808 0 1 299744
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1095
timestamp 1586364061
transform -1 0 8832 0 1 299744
box -38 -48 314 592
use scs8hd_decap_6  FILLER_547_74
timestamp 1586364061
transform 1 0 7912 0 1 299744
box -38 -48 590 592
use scs8hd_fill_1  FILLER_547_80
timestamp 1586364061
transform 1 0 8464 0 1 299744
box -38 -48 130 592
use scs8hd_decap_3  PHY_1096
timestamp 1586364061
transform 1 0 1104 0 -1 300832
box -38 -48 314 592
use scs8hd_decap_3  PHY_1098
timestamp 1586364061
transform 1 0 1104 0 1 300832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_548_3
timestamp 1586364061
transform 1 0 1380 0 -1 300832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_548_15
timestamp 1586364061
transform 1 0 2484 0 -1 300832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_549_3
timestamp 1586364061
transform 1 0 1380 0 1 300832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_549_15
timestamp 1586364061
transform 1 0 2484 0 1 300832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1757
timestamp 1586364061
transform 1 0 3956 0 -1 300832
box -38 -48 130 592
use scs8hd_decap_4  FILLER_548_27
timestamp 1586364061
transform 1 0 3588 0 -1 300832
box -38 -48 406 592
use scs8hd_decap_12  FILLER_548_32
timestamp 1586364061
transform 1 0 4048 0 -1 300832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_549_27
timestamp 1586364061
transform 1 0 3588 0 1 300832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_548_44
timestamp 1586364061
transform 1 0 5152 0 -1 300832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_549_39
timestamp 1586364061
transform 1 0 4692 0 1 300832
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_549_51
timestamp 1586364061
transform 1 0 5796 0 1 300832
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1758
timestamp 1586364061
transform 1 0 6716 0 1 300832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_548_56
timestamp 1586364061
transform 1 0 6256 0 -1 300832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_548_68
timestamp 1586364061
transform 1 0 7360 0 -1 300832
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_549_59
timestamp 1586364061
transform 1 0 6532 0 1 300832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_549_62
timestamp 1586364061
transform 1 0 6808 0 1 300832
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1097
timestamp 1586364061
transform -1 0 8832 0 -1 300832
box -38 -48 314 592
use scs8hd_decap_3  PHY_1099
timestamp 1586364061
transform -1 0 8832 0 1 300832
box -38 -48 314 592
use scs8hd_fill_1  FILLER_548_80
timestamp 1586364061
transform 1 0 8464 0 -1 300832
box -38 -48 130 592
use scs8hd_decap_6  FILLER_549_74
timestamp 1586364061
transform 1 0 7912 0 1 300832
box -38 -48 590 592
use scs8hd_fill_1  FILLER_549_80
timestamp 1586364061
transform 1 0 8464 0 1 300832
box -38 -48 130 592
use scs8hd_decap_3  PHY_1100
timestamp 1586364061
transform 1 0 1104 0 -1 301920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_550_3
timestamp 1586364061
transform 1 0 1380 0 -1 301920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_550_15
timestamp 1586364061
transform 1 0 2484 0 -1 301920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1759
timestamp 1586364061
transform 1 0 3956 0 -1 301920
box -38 -48 130 592
use scs8hd_decap_4  FILLER_550_27
timestamp 1586364061
transform 1 0 3588 0 -1 301920
box -38 -48 406 592
use scs8hd_decap_12  FILLER_550_32
timestamp 1586364061
transform 1 0 4048 0 -1 301920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_550_44
timestamp 1586364061
transform 1 0 5152 0 -1 301920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_550_56
timestamp 1586364061
transform 1 0 6256 0 -1 301920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_550_68
timestamp 1586364061
transform 1 0 7360 0 -1 301920
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1101
timestamp 1586364061
transform -1 0 8832 0 -1 301920
box -38 -48 314 592
use scs8hd_fill_1  FILLER_550_80
timestamp 1586364061
transform 1 0 8464 0 -1 301920
box -38 -48 130 592
use scs8hd_decap_3  PHY_1102
timestamp 1586364061
transform 1 0 1104 0 1 301920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_551_3
timestamp 1586364061
transform 1 0 1380 0 1 301920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_551_15
timestamp 1586364061
transform 1 0 2484 0 1 301920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_551_27
timestamp 1586364061
transform 1 0 3588 0 1 301920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_551_39
timestamp 1586364061
transform 1 0 4692 0 1 301920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_551_51
timestamp 1586364061
transform 1 0 5796 0 1 301920
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1760
timestamp 1586364061
transform 1 0 6716 0 1 301920
box -38 -48 130 592
use scs8hd_fill_2  FILLER_551_59
timestamp 1586364061
transform 1 0 6532 0 1 301920
box -38 -48 222 592
use scs8hd_decap_12  FILLER_551_62
timestamp 1586364061
transform 1 0 6808 0 1 301920
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1103
timestamp 1586364061
transform -1 0 8832 0 1 301920
box -38 -48 314 592
use scs8hd_decap_6  FILLER_551_74
timestamp 1586364061
transform 1 0 7912 0 1 301920
box -38 -48 590 592
use scs8hd_fill_1  FILLER_551_80
timestamp 1586364061
transform 1 0 8464 0 1 301920
box -38 -48 130 592
use scs8hd_decap_3  PHY_1104
timestamp 1586364061
transform 1 0 1104 0 -1 303008
box -38 -48 314 592
use scs8hd_decap_12  FILLER_552_3
timestamp 1586364061
transform 1 0 1380 0 -1 303008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_552_15
timestamp 1586364061
transform 1 0 2484 0 -1 303008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1761
timestamp 1586364061
transform 1 0 3956 0 -1 303008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_552_27
timestamp 1586364061
transform 1 0 3588 0 -1 303008
box -38 -48 406 592
use scs8hd_decap_12  FILLER_552_32
timestamp 1586364061
transform 1 0 4048 0 -1 303008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_552_44
timestamp 1586364061
transform 1 0 5152 0 -1 303008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_552_56
timestamp 1586364061
transform 1 0 6256 0 -1 303008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_552_68
timestamp 1586364061
transform 1 0 7360 0 -1 303008
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1105
timestamp 1586364061
transform -1 0 8832 0 -1 303008
box -38 -48 314 592
use scs8hd_fill_1  FILLER_552_80
timestamp 1586364061
transform 1 0 8464 0 -1 303008
box -38 -48 130 592
use scs8hd_decap_3  PHY_1106
timestamp 1586364061
transform 1 0 1104 0 1 303008
box -38 -48 314 592
use scs8hd_decap_12  FILLER_553_3
timestamp 1586364061
transform 1 0 1380 0 1 303008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_553_15
timestamp 1586364061
transform 1 0 2484 0 1 303008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_553_27
timestamp 1586364061
transform 1 0 3588 0 1 303008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_553_39
timestamp 1586364061
transform 1 0 4692 0 1 303008
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_553_51
timestamp 1586364061
transform 1 0 5796 0 1 303008
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1762
timestamp 1586364061
transform 1 0 6716 0 1 303008
box -38 -48 130 592
use scs8hd_fill_2  FILLER_553_59
timestamp 1586364061
transform 1 0 6532 0 1 303008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_553_62
timestamp 1586364061
transform 1 0 6808 0 1 303008
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1107
timestamp 1586364061
transform -1 0 8832 0 1 303008
box -38 -48 314 592
use scs8hd_decap_6  FILLER_553_74
timestamp 1586364061
transform 1 0 7912 0 1 303008
box -38 -48 590 592
use scs8hd_fill_1  FILLER_553_80
timestamp 1586364061
transform 1 0 8464 0 1 303008
box -38 -48 130 592
use scs8hd_decap_3  PHY_1108
timestamp 1586364061
transform 1 0 1104 0 -1 304096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_554_3
timestamp 1586364061
transform 1 0 1380 0 -1 304096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_554_15
timestamp 1586364061
transform 1 0 2484 0 -1 304096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1763
timestamp 1586364061
transform 1 0 3956 0 -1 304096
box -38 -48 130 592
use scs8hd_decap_4  FILLER_554_27
timestamp 1586364061
transform 1 0 3588 0 -1 304096
box -38 -48 406 592
use scs8hd_decap_12  FILLER_554_32
timestamp 1586364061
transform 1 0 4048 0 -1 304096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_554_44
timestamp 1586364061
transform 1 0 5152 0 -1 304096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_554_56
timestamp 1586364061
transform 1 0 6256 0 -1 304096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_554_68
timestamp 1586364061
transform 1 0 7360 0 -1 304096
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1109
timestamp 1586364061
transform -1 0 8832 0 -1 304096
box -38 -48 314 592
use scs8hd_fill_1  FILLER_554_80
timestamp 1586364061
transform 1 0 8464 0 -1 304096
box -38 -48 130 592
use scs8hd_decap_3  PHY_1110
timestamp 1586364061
transform 1 0 1104 0 1 304096
box -38 -48 314 592
use scs8hd_decap_3  PHY_1112
timestamp 1586364061
transform 1 0 1104 0 -1 305184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_555_3
timestamp 1586364061
transform 1 0 1380 0 1 304096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_555_15
timestamp 1586364061
transform 1 0 2484 0 1 304096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_556_3
timestamp 1586364061
transform 1 0 1380 0 -1 305184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_556_15
timestamp 1586364061
transform 1 0 2484 0 -1 305184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1765
timestamp 1586364061
transform 1 0 3956 0 -1 305184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_555_27
timestamp 1586364061
transform 1 0 3588 0 1 304096
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_556_27
timestamp 1586364061
transform 1 0 3588 0 -1 305184
box -38 -48 406 592
use scs8hd_decap_12  FILLER_556_32
timestamp 1586364061
transform 1 0 4048 0 -1 305184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_555_39
timestamp 1586364061
transform 1 0 4692 0 1 304096
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_555_51
timestamp 1586364061
transform 1 0 5796 0 1 304096
box -38 -48 774 592
use scs8hd_decap_12  FILLER_556_44
timestamp 1586364061
transform 1 0 5152 0 -1 305184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1764
timestamp 1586364061
transform 1 0 6716 0 1 304096
box -38 -48 130 592
use scs8hd_fill_2  FILLER_555_59
timestamp 1586364061
transform 1 0 6532 0 1 304096
box -38 -48 222 592
use scs8hd_decap_12  FILLER_555_62
timestamp 1586364061
transform 1 0 6808 0 1 304096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_556_56
timestamp 1586364061
transform 1 0 6256 0 -1 305184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_556_68
timestamp 1586364061
transform 1 0 7360 0 -1 305184
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1111
timestamp 1586364061
transform -1 0 8832 0 1 304096
box -38 -48 314 592
use scs8hd_decap_3  PHY_1113
timestamp 1586364061
transform -1 0 8832 0 -1 305184
box -38 -48 314 592
use scs8hd_decap_6  FILLER_555_74
timestamp 1586364061
transform 1 0 7912 0 1 304096
box -38 -48 590 592
use scs8hd_fill_1  FILLER_555_80
timestamp 1586364061
transform 1 0 8464 0 1 304096
box -38 -48 130 592
use scs8hd_fill_1  FILLER_556_80
timestamp 1586364061
transform 1 0 8464 0 -1 305184
box -38 -48 130 592
use scs8hd_decap_3  PHY_1114
timestamp 1586364061
transform 1 0 1104 0 1 305184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_557_3
timestamp 1586364061
transform 1 0 1380 0 1 305184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_557_15
timestamp 1586364061
transform 1 0 2484 0 1 305184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_557_27
timestamp 1586364061
transform 1 0 3588 0 1 305184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_557_39
timestamp 1586364061
transform 1 0 4692 0 1 305184
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_557_51
timestamp 1586364061
transform 1 0 5796 0 1 305184
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1766
timestamp 1586364061
transform 1 0 6716 0 1 305184
box -38 -48 130 592
use scs8hd_fill_2  FILLER_557_59
timestamp 1586364061
transform 1 0 6532 0 1 305184
box -38 -48 222 592
use scs8hd_decap_12  FILLER_557_62
timestamp 1586364061
transform 1 0 6808 0 1 305184
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1115
timestamp 1586364061
transform -1 0 8832 0 1 305184
box -38 -48 314 592
use scs8hd_decap_6  FILLER_557_74
timestamp 1586364061
transform 1 0 7912 0 1 305184
box -38 -48 590 592
use scs8hd_fill_1  FILLER_557_80
timestamp 1586364061
transform 1 0 8464 0 1 305184
box -38 -48 130 592
use scs8hd_decap_3  PHY_1116
timestamp 1586364061
transform 1 0 1104 0 -1 306272
box -38 -48 314 592
use scs8hd_decap_12  FILLER_558_3
timestamp 1586364061
transform 1 0 1380 0 -1 306272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_558_15
timestamp 1586364061
transform 1 0 2484 0 -1 306272
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1767
timestamp 1586364061
transform 1 0 3956 0 -1 306272
box -38 -48 130 592
use scs8hd_decap_4  FILLER_558_27
timestamp 1586364061
transform 1 0 3588 0 -1 306272
box -38 -48 406 592
use scs8hd_decap_12  FILLER_558_32
timestamp 1586364061
transform 1 0 4048 0 -1 306272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_558_44
timestamp 1586364061
transform 1 0 5152 0 -1 306272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_558_56
timestamp 1586364061
transform 1 0 6256 0 -1 306272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_558_68
timestamp 1586364061
transform 1 0 7360 0 -1 306272
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1117
timestamp 1586364061
transform -1 0 8832 0 -1 306272
box -38 -48 314 592
use scs8hd_fill_1  FILLER_558_80
timestamp 1586364061
transform 1 0 8464 0 -1 306272
box -38 -48 130 592
use scs8hd_decap_3  PHY_1118
timestamp 1586364061
transform 1 0 1104 0 1 306272
box -38 -48 314 592
use scs8hd_decap_12  FILLER_559_3
timestamp 1586364061
transform 1 0 1380 0 1 306272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_559_15
timestamp 1586364061
transform 1 0 2484 0 1 306272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_559_27
timestamp 1586364061
transform 1 0 3588 0 1 306272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_559_39
timestamp 1586364061
transform 1 0 4692 0 1 306272
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_559_51
timestamp 1586364061
transform 1 0 5796 0 1 306272
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1768
timestamp 1586364061
transform 1 0 6716 0 1 306272
box -38 -48 130 592
use scs8hd_fill_2  FILLER_559_59
timestamp 1586364061
transform 1 0 6532 0 1 306272
box -38 -48 222 592
use scs8hd_decap_12  FILLER_559_62
timestamp 1586364061
transform 1 0 6808 0 1 306272
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1119
timestamp 1586364061
transform -1 0 8832 0 1 306272
box -38 -48 314 592
use scs8hd_decap_6  FILLER_559_74
timestamp 1586364061
transform 1 0 7912 0 1 306272
box -38 -48 590 592
use scs8hd_fill_1  FILLER_559_80
timestamp 1586364061
transform 1 0 8464 0 1 306272
box -38 -48 130 592
use scs8hd_decap_3  PHY_1120
timestamp 1586364061
transform 1 0 1104 0 -1 307360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_560_3
timestamp 1586364061
transform 1 0 1380 0 -1 307360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_560_15
timestamp 1586364061
transform 1 0 2484 0 -1 307360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1769
timestamp 1586364061
transform 1 0 3956 0 -1 307360
box -38 -48 130 592
use scs8hd_decap_4  FILLER_560_27
timestamp 1586364061
transform 1 0 3588 0 -1 307360
box -38 -48 406 592
use scs8hd_decap_12  FILLER_560_32
timestamp 1586364061
transform 1 0 4048 0 -1 307360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_560_44
timestamp 1586364061
transform 1 0 5152 0 -1 307360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_560_56
timestamp 1586364061
transform 1 0 6256 0 -1 307360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_560_68
timestamp 1586364061
transform 1 0 7360 0 -1 307360
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1121
timestamp 1586364061
transform -1 0 8832 0 -1 307360
box -38 -48 314 592
use scs8hd_fill_1  FILLER_560_80
timestamp 1586364061
transform 1 0 8464 0 -1 307360
box -38 -48 130 592
use scs8hd_decap_3  PHY_1122
timestamp 1586364061
transform 1 0 1104 0 1 307360
box -38 -48 314 592
use scs8hd_decap_3  PHY_1124
timestamp 1586364061
transform 1 0 1104 0 -1 308448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_561_3
timestamp 1586364061
transform 1 0 1380 0 1 307360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_561_15
timestamp 1586364061
transform 1 0 2484 0 1 307360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_562_3
timestamp 1586364061
transform 1 0 1380 0 -1 308448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_562_15
timestamp 1586364061
transform 1 0 2484 0 -1 308448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1771
timestamp 1586364061
transform 1 0 3956 0 -1 308448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_561_27
timestamp 1586364061
transform 1 0 3588 0 1 307360
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_562_27
timestamp 1586364061
transform 1 0 3588 0 -1 308448
box -38 -48 406 592
use scs8hd_decap_12  FILLER_562_32
timestamp 1586364061
transform 1 0 4048 0 -1 308448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_561_39
timestamp 1586364061
transform 1 0 4692 0 1 307360
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_561_51
timestamp 1586364061
transform 1 0 5796 0 1 307360
box -38 -48 774 592
use scs8hd_decap_12  FILLER_562_44
timestamp 1586364061
transform 1 0 5152 0 -1 308448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1770
timestamp 1586364061
transform 1 0 6716 0 1 307360
box -38 -48 130 592
use scs8hd_fill_2  FILLER_561_59
timestamp 1586364061
transform 1 0 6532 0 1 307360
box -38 -48 222 592
use scs8hd_decap_12  FILLER_561_62
timestamp 1586364061
transform 1 0 6808 0 1 307360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_562_56
timestamp 1586364061
transform 1 0 6256 0 -1 308448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_562_68
timestamp 1586364061
transform 1 0 7360 0 -1 308448
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1123
timestamp 1586364061
transform -1 0 8832 0 1 307360
box -38 -48 314 592
use scs8hd_decap_3  PHY_1125
timestamp 1586364061
transform -1 0 8832 0 -1 308448
box -38 -48 314 592
use scs8hd_decap_6  FILLER_561_74
timestamp 1586364061
transform 1 0 7912 0 1 307360
box -38 -48 590 592
use scs8hd_fill_1  FILLER_561_80
timestamp 1586364061
transform 1 0 8464 0 1 307360
box -38 -48 130 592
use scs8hd_fill_1  FILLER_562_80
timestamp 1586364061
transform 1 0 8464 0 -1 308448
box -38 -48 130 592
use scs8hd_decap_3  PHY_1126
timestamp 1586364061
transform 1 0 1104 0 1 308448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_563_3
timestamp 1586364061
transform 1 0 1380 0 1 308448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_563_15
timestamp 1586364061
transform 1 0 2484 0 1 308448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_563_27
timestamp 1586364061
transform 1 0 3588 0 1 308448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_563_39
timestamp 1586364061
transform 1 0 4692 0 1 308448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_563_51
timestamp 1586364061
transform 1 0 5796 0 1 308448
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1772
timestamp 1586364061
transform 1 0 6716 0 1 308448
box -38 -48 130 592
use scs8hd_fill_2  FILLER_563_59
timestamp 1586364061
transform 1 0 6532 0 1 308448
box -38 -48 222 592
use scs8hd_decap_12  FILLER_563_62
timestamp 1586364061
transform 1 0 6808 0 1 308448
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1127
timestamp 1586364061
transform -1 0 8832 0 1 308448
box -38 -48 314 592
use scs8hd_decap_6  FILLER_563_74
timestamp 1586364061
transform 1 0 7912 0 1 308448
box -38 -48 590 592
use scs8hd_fill_1  FILLER_563_80
timestamp 1586364061
transform 1 0 8464 0 1 308448
box -38 -48 130 592
use scs8hd_decap_3  PHY_1128
timestamp 1586364061
transform 1 0 1104 0 -1 309536
box -38 -48 314 592
use scs8hd_decap_12  FILLER_564_3
timestamp 1586364061
transform 1 0 1380 0 -1 309536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_564_15
timestamp 1586364061
transform 1 0 2484 0 -1 309536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1773
timestamp 1586364061
transform 1 0 3956 0 -1 309536
box -38 -48 130 592
use scs8hd_decap_4  FILLER_564_27
timestamp 1586364061
transform 1 0 3588 0 -1 309536
box -38 -48 406 592
use scs8hd_decap_12  FILLER_564_32
timestamp 1586364061
transform 1 0 4048 0 -1 309536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_564_44
timestamp 1586364061
transform 1 0 5152 0 -1 309536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_564_56
timestamp 1586364061
transform 1 0 6256 0 -1 309536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_564_68
timestamp 1586364061
transform 1 0 7360 0 -1 309536
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1129
timestamp 1586364061
transform -1 0 8832 0 -1 309536
box -38 -48 314 592
use scs8hd_fill_1  FILLER_564_80
timestamp 1586364061
transform 1 0 8464 0 -1 309536
box -38 -48 130 592
use scs8hd_decap_3  PHY_1130
timestamp 1586364061
transform 1 0 1104 0 1 309536
box -38 -48 314 592
use scs8hd_decap_12  FILLER_565_3
timestamp 1586364061
transform 1 0 1380 0 1 309536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_565_15
timestamp 1586364061
transform 1 0 2484 0 1 309536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_565_27
timestamp 1586364061
transform 1 0 3588 0 1 309536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_565_39
timestamp 1586364061
transform 1 0 4692 0 1 309536
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_565_51
timestamp 1586364061
transform 1 0 5796 0 1 309536
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1774
timestamp 1586364061
transform 1 0 6716 0 1 309536
box -38 -48 130 592
use scs8hd_fill_2  FILLER_565_59
timestamp 1586364061
transform 1 0 6532 0 1 309536
box -38 -48 222 592
use scs8hd_decap_12  FILLER_565_62
timestamp 1586364061
transform 1 0 6808 0 1 309536
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1131
timestamp 1586364061
transform -1 0 8832 0 1 309536
box -38 -48 314 592
use scs8hd_decap_6  FILLER_565_74
timestamp 1586364061
transform 1 0 7912 0 1 309536
box -38 -48 590 592
use scs8hd_fill_1  FILLER_565_80
timestamp 1586364061
transform 1 0 8464 0 1 309536
box -38 -48 130 592
use scs8hd_decap_3  PHY_1132
timestamp 1586364061
transform 1 0 1104 0 -1 310624
box -38 -48 314 592
use scs8hd_decap_12  FILLER_566_3
timestamp 1586364061
transform 1 0 1380 0 -1 310624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_566_15
timestamp 1586364061
transform 1 0 2484 0 -1 310624
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1775
timestamp 1586364061
transform 1 0 3956 0 -1 310624
box -38 -48 130 592
use scs8hd_decap_4  FILLER_566_27
timestamp 1586364061
transform 1 0 3588 0 -1 310624
box -38 -48 406 592
use scs8hd_decap_12  FILLER_566_32
timestamp 1586364061
transform 1 0 4048 0 -1 310624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_566_44
timestamp 1586364061
transform 1 0 5152 0 -1 310624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_566_56
timestamp 1586364061
transform 1 0 6256 0 -1 310624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_566_68
timestamp 1586364061
transform 1 0 7360 0 -1 310624
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1133
timestamp 1586364061
transform -1 0 8832 0 -1 310624
box -38 -48 314 592
use scs8hd_fill_1  FILLER_566_80
timestamp 1586364061
transform 1 0 8464 0 -1 310624
box -38 -48 130 592
use scs8hd_decap_3  PHY_1134
timestamp 1586364061
transform 1 0 1104 0 1 310624
box -38 -48 314 592
use scs8hd_decap_12  FILLER_567_3
timestamp 1586364061
transform 1 0 1380 0 1 310624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_567_15
timestamp 1586364061
transform 1 0 2484 0 1 310624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_567_27
timestamp 1586364061
transform 1 0 3588 0 1 310624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_567_39
timestamp 1586364061
transform 1 0 4692 0 1 310624
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_567_51
timestamp 1586364061
transform 1 0 5796 0 1 310624
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1776
timestamp 1586364061
transform 1 0 6716 0 1 310624
box -38 -48 130 592
use scs8hd_fill_2  FILLER_567_59
timestamp 1586364061
transform 1 0 6532 0 1 310624
box -38 -48 222 592
use scs8hd_decap_12  FILLER_567_62
timestamp 1586364061
transform 1 0 6808 0 1 310624
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1135
timestamp 1586364061
transform -1 0 8832 0 1 310624
box -38 -48 314 592
use scs8hd_decap_6  FILLER_567_74
timestamp 1586364061
transform 1 0 7912 0 1 310624
box -38 -48 590 592
use scs8hd_fill_1  FILLER_567_80
timestamp 1586364061
transform 1 0 8464 0 1 310624
box -38 -48 130 592
use scs8hd_decap_3  PHY_1136
timestamp 1586364061
transform 1 0 1104 0 -1 311712
box -38 -48 314 592
use scs8hd_decap_3  PHY_1138
timestamp 1586364061
transform 1 0 1104 0 1 311712
box -38 -48 314 592
use scs8hd_decap_12  FILLER_568_3
timestamp 1586364061
transform 1 0 1380 0 -1 311712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_568_15
timestamp 1586364061
transform 1 0 2484 0 -1 311712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_569_3
timestamp 1586364061
transform 1 0 1380 0 1 311712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_569_15
timestamp 1586364061
transform 1 0 2484 0 1 311712
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1777
timestamp 1586364061
transform 1 0 3956 0 -1 311712
box -38 -48 130 592
use scs8hd_decap_4  FILLER_568_27
timestamp 1586364061
transform 1 0 3588 0 -1 311712
box -38 -48 406 592
use scs8hd_decap_12  FILLER_568_32
timestamp 1586364061
transform 1 0 4048 0 -1 311712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_569_27
timestamp 1586364061
transform 1 0 3588 0 1 311712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_568_44
timestamp 1586364061
transform 1 0 5152 0 -1 311712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_569_39
timestamp 1586364061
transform 1 0 4692 0 1 311712
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_569_51
timestamp 1586364061
transform 1 0 5796 0 1 311712
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1778
timestamp 1586364061
transform 1 0 6716 0 1 311712
box -38 -48 130 592
use scs8hd_decap_12  FILLER_568_56
timestamp 1586364061
transform 1 0 6256 0 -1 311712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_568_68
timestamp 1586364061
transform 1 0 7360 0 -1 311712
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_569_59
timestamp 1586364061
transform 1 0 6532 0 1 311712
box -38 -48 222 592
use scs8hd_decap_12  FILLER_569_62
timestamp 1586364061
transform 1 0 6808 0 1 311712
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1137
timestamp 1586364061
transform -1 0 8832 0 -1 311712
box -38 -48 314 592
use scs8hd_decap_3  PHY_1139
timestamp 1586364061
transform -1 0 8832 0 1 311712
box -38 -48 314 592
use scs8hd_fill_1  FILLER_568_80
timestamp 1586364061
transform 1 0 8464 0 -1 311712
box -38 -48 130 592
use scs8hd_decap_6  FILLER_569_74
timestamp 1586364061
transform 1 0 7912 0 1 311712
box -38 -48 590 592
use scs8hd_fill_1  FILLER_569_80
timestamp 1586364061
transform 1 0 8464 0 1 311712
box -38 -48 130 592
use scs8hd_decap_3  PHY_1140
timestamp 1586364061
transform 1 0 1104 0 -1 312800
box -38 -48 314 592
use scs8hd_decap_12  FILLER_570_3
timestamp 1586364061
transform 1 0 1380 0 -1 312800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_570_15
timestamp 1586364061
transform 1 0 2484 0 -1 312800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1779
timestamp 1586364061
transform 1 0 3956 0 -1 312800
box -38 -48 130 592
use scs8hd_decap_4  FILLER_570_27
timestamp 1586364061
transform 1 0 3588 0 -1 312800
box -38 -48 406 592
use scs8hd_decap_12  FILLER_570_32
timestamp 1586364061
transform 1 0 4048 0 -1 312800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_570_44
timestamp 1586364061
transform 1 0 5152 0 -1 312800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_570_56
timestamp 1586364061
transform 1 0 6256 0 -1 312800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_570_68
timestamp 1586364061
transform 1 0 7360 0 -1 312800
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1141
timestamp 1586364061
transform -1 0 8832 0 -1 312800
box -38 -48 314 592
use scs8hd_fill_1  FILLER_570_80
timestamp 1586364061
transform 1 0 8464 0 -1 312800
box -38 -48 130 592
use scs8hd_decap_3  PHY_1142
timestamp 1586364061
transform 1 0 1104 0 1 312800
box -38 -48 314 592
use scs8hd_decap_12  FILLER_571_3
timestamp 1586364061
transform 1 0 1380 0 1 312800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_571_15
timestamp 1586364061
transform 1 0 2484 0 1 312800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_571_27
timestamp 1586364061
transform 1 0 3588 0 1 312800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_571_39
timestamp 1586364061
transform 1 0 4692 0 1 312800
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_571_51
timestamp 1586364061
transform 1 0 5796 0 1 312800
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1780
timestamp 1586364061
transform 1 0 6716 0 1 312800
box -38 -48 130 592
use scs8hd_fill_2  FILLER_571_59
timestamp 1586364061
transform 1 0 6532 0 1 312800
box -38 -48 222 592
use scs8hd_decap_12  FILLER_571_62
timestamp 1586364061
transform 1 0 6808 0 1 312800
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1143
timestamp 1586364061
transform -1 0 8832 0 1 312800
box -38 -48 314 592
use scs8hd_decap_6  FILLER_571_74
timestamp 1586364061
transform 1 0 7912 0 1 312800
box -38 -48 590 592
use scs8hd_fill_1  FILLER_571_80
timestamp 1586364061
transform 1 0 8464 0 1 312800
box -38 -48 130 592
use scs8hd_decap_3  PHY_1144
timestamp 1586364061
transform 1 0 1104 0 -1 313888
box -38 -48 314 592
use scs8hd_decap_12  FILLER_572_3
timestamp 1586364061
transform 1 0 1380 0 -1 313888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_572_15
timestamp 1586364061
transform 1 0 2484 0 -1 313888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1781
timestamp 1586364061
transform 1 0 3956 0 -1 313888
box -38 -48 130 592
use scs8hd_decap_4  FILLER_572_27
timestamp 1586364061
transform 1 0 3588 0 -1 313888
box -38 -48 406 592
use scs8hd_decap_12  FILLER_572_32
timestamp 1586364061
transform 1 0 4048 0 -1 313888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_572_44
timestamp 1586364061
transform 1 0 5152 0 -1 313888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_572_56
timestamp 1586364061
transform 1 0 6256 0 -1 313888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_572_68
timestamp 1586364061
transform 1 0 7360 0 -1 313888
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1145
timestamp 1586364061
transform -1 0 8832 0 -1 313888
box -38 -48 314 592
use scs8hd_fill_1  FILLER_572_80
timestamp 1586364061
transform 1 0 8464 0 -1 313888
box -38 -48 130 592
use scs8hd_decap_3  PHY_1146
timestamp 1586364061
transform 1 0 1104 0 1 313888
box -38 -48 314 592
use scs8hd_decap_12  FILLER_573_3
timestamp 1586364061
transform 1 0 1380 0 1 313888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_573_15
timestamp 1586364061
transform 1 0 2484 0 1 313888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_573_27
timestamp 1586364061
transform 1 0 3588 0 1 313888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_573_39
timestamp 1586364061
transform 1 0 4692 0 1 313888
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_573_51
timestamp 1586364061
transform 1 0 5796 0 1 313888
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1782
timestamp 1586364061
transform 1 0 6716 0 1 313888
box -38 -48 130 592
use scs8hd_fill_2  FILLER_573_59
timestamp 1586364061
transform 1 0 6532 0 1 313888
box -38 -48 222 592
use scs8hd_decap_12  FILLER_573_62
timestamp 1586364061
transform 1 0 6808 0 1 313888
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1147
timestamp 1586364061
transform -1 0 8832 0 1 313888
box -38 -48 314 592
use scs8hd_decap_6  FILLER_573_74
timestamp 1586364061
transform 1 0 7912 0 1 313888
box -38 -48 590 592
use scs8hd_fill_1  FILLER_573_80
timestamp 1586364061
transform 1 0 8464 0 1 313888
box -38 -48 130 592
use scs8hd_decap_3  PHY_1148
timestamp 1586364061
transform 1 0 1104 0 -1 314976
box -38 -48 314 592
use scs8hd_decap_3  PHY_1150
timestamp 1586364061
transform 1 0 1104 0 1 314976
box -38 -48 314 592
use scs8hd_decap_12  FILLER_574_3
timestamp 1586364061
transform 1 0 1380 0 -1 314976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_574_15
timestamp 1586364061
transform 1 0 2484 0 -1 314976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_575_3
timestamp 1586364061
transform 1 0 1380 0 1 314976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_575_15
timestamp 1586364061
transform 1 0 2484 0 1 314976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1783
timestamp 1586364061
transform 1 0 3956 0 -1 314976
box -38 -48 130 592
use scs8hd_decap_4  FILLER_574_27
timestamp 1586364061
transform 1 0 3588 0 -1 314976
box -38 -48 406 592
use scs8hd_decap_12  FILLER_574_32
timestamp 1586364061
transform 1 0 4048 0 -1 314976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_575_27
timestamp 1586364061
transform 1 0 3588 0 1 314976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_574_44
timestamp 1586364061
transform 1 0 5152 0 -1 314976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_575_39
timestamp 1586364061
transform 1 0 4692 0 1 314976
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_575_51
timestamp 1586364061
transform 1 0 5796 0 1 314976
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1784
timestamp 1586364061
transform 1 0 6716 0 1 314976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_574_56
timestamp 1586364061
transform 1 0 6256 0 -1 314976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_574_68
timestamp 1586364061
transform 1 0 7360 0 -1 314976
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_575_59
timestamp 1586364061
transform 1 0 6532 0 1 314976
box -38 -48 222 592
use scs8hd_decap_12  FILLER_575_62
timestamp 1586364061
transform 1 0 6808 0 1 314976
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1149
timestamp 1586364061
transform -1 0 8832 0 -1 314976
box -38 -48 314 592
use scs8hd_decap_3  PHY_1151
timestamp 1586364061
transform -1 0 8832 0 1 314976
box -38 -48 314 592
use scs8hd_fill_1  FILLER_574_80
timestamp 1586364061
transform 1 0 8464 0 -1 314976
box -38 -48 130 592
use scs8hd_decap_6  FILLER_575_74
timestamp 1586364061
transform 1 0 7912 0 1 314976
box -38 -48 590 592
use scs8hd_fill_1  FILLER_575_80
timestamp 1586364061
transform 1 0 8464 0 1 314976
box -38 -48 130 592
use scs8hd_decap_3  PHY_1152
timestamp 1586364061
transform 1 0 1104 0 -1 316064
box -38 -48 314 592
use scs8hd_decap_12  FILLER_576_3
timestamp 1586364061
transform 1 0 1380 0 -1 316064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_576_15
timestamp 1586364061
transform 1 0 2484 0 -1 316064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1785
timestamp 1586364061
transform 1 0 3956 0 -1 316064
box -38 -48 130 592
use scs8hd_decap_4  FILLER_576_27
timestamp 1586364061
transform 1 0 3588 0 -1 316064
box -38 -48 406 592
use scs8hd_decap_12  FILLER_576_32
timestamp 1586364061
transform 1 0 4048 0 -1 316064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_576_44
timestamp 1586364061
transform 1 0 5152 0 -1 316064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_576_56
timestamp 1586364061
transform 1 0 6256 0 -1 316064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_576_68
timestamp 1586364061
transform 1 0 7360 0 -1 316064
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1153
timestamp 1586364061
transform -1 0 8832 0 -1 316064
box -38 -48 314 592
use scs8hd_fill_1  FILLER_576_80
timestamp 1586364061
transform 1 0 8464 0 -1 316064
box -38 -48 130 592
use scs8hd_decap_3  PHY_1154
timestamp 1586364061
transform 1 0 1104 0 1 316064
box -38 -48 314 592
use scs8hd_decap_12  FILLER_577_3
timestamp 1586364061
transform 1 0 1380 0 1 316064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_577_15
timestamp 1586364061
transform 1 0 2484 0 1 316064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_577_27
timestamp 1586364061
transform 1 0 3588 0 1 316064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_577_39
timestamp 1586364061
transform 1 0 4692 0 1 316064
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_577_51
timestamp 1586364061
transform 1 0 5796 0 1 316064
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1786
timestamp 1586364061
transform 1 0 6716 0 1 316064
box -38 -48 130 592
use scs8hd_fill_2  FILLER_577_59
timestamp 1586364061
transform 1 0 6532 0 1 316064
box -38 -48 222 592
use scs8hd_decap_12  FILLER_577_62
timestamp 1586364061
transform 1 0 6808 0 1 316064
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1155
timestamp 1586364061
transform -1 0 8832 0 1 316064
box -38 -48 314 592
use scs8hd_decap_6  FILLER_577_74
timestamp 1586364061
transform 1 0 7912 0 1 316064
box -38 -48 590 592
use scs8hd_fill_1  FILLER_577_80
timestamp 1586364061
transform 1 0 8464 0 1 316064
box -38 -48 130 592
use scs8hd_decap_3  PHY_1156
timestamp 1586364061
transform 1 0 1104 0 -1 317152
box -38 -48 314 592
use scs8hd_decap_12  FILLER_578_3
timestamp 1586364061
transform 1 0 1380 0 -1 317152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_578_15
timestamp 1586364061
transform 1 0 2484 0 -1 317152
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1787
timestamp 1586364061
transform 1 0 3956 0 -1 317152
box -38 -48 130 592
use scs8hd_decap_4  FILLER_578_27
timestamp 1586364061
transform 1 0 3588 0 -1 317152
box -38 -48 406 592
use scs8hd_decap_12  FILLER_578_32
timestamp 1586364061
transform 1 0 4048 0 -1 317152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_578_44
timestamp 1586364061
transform 1 0 5152 0 -1 317152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_578_56
timestamp 1586364061
transform 1 0 6256 0 -1 317152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_578_68
timestamp 1586364061
transform 1 0 7360 0 -1 317152
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1157
timestamp 1586364061
transform -1 0 8832 0 -1 317152
box -38 -48 314 592
use scs8hd_fill_1  FILLER_578_80
timestamp 1586364061
transform 1 0 8464 0 -1 317152
box -38 -48 130 592
use scs8hd_decap_3  PHY_1158
timestamp 1586364061
transform 1 0 1104 0 1 317152
box -38 -48 314 592
use scs8hd_decap_12  FILLER_579_3
timestamp 1586364061
transform 1 0 1380 0 1 317152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_579_15
timestamp 1586364061
transform 1 0 2484 0 1 317152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_579_27
timestamp 1586364061
transform 1 0 3588 0 1 317152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_579_39
timestamp 1586364061
transform 1 0 4692 0 1 317152
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_579_51
timestamp 1586364061
transform 1 0 5796 0 1 317152
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1788
timestamp 1586364061
transform 1 0 6716 0 1 317152
box -38 -48 130 592
use scs8hd_fill_2  FILLER_579_59
timestamp 1586364061
transform 1 0 6532 0 1 317152
box -38 -48 222 592
use scs8hd_decap_12  FILLER_579_62
timestamp 1586364061
transform 1 0 6808 0 1 317152
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1159
timestamp 1586364061
transform -1 0 8832 0 1 317152
box -38 -48 314 592
use scs8hd_decap_6  FILLER_579_74
timestamp 1586364061
transform 1 0 7912 0 1 317152
box -38 -48 590 592
use scs8hd_fill_1  FILLER_579_80
timestamp 1586364061
transform 1 0 8464 0 1 317152
box -38 -48 130 592
use scs8hd_decap_3  PHY_1160
timestamp 1586364061
transform 1 0 1104 0 -1 318240
box -38 -48 314 592
use scs8hd_decap_12  FILLER_580_3
timestamp 1586364061
transform 1 0 1380 0 -1 318240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_580_15
timestamp 1586364061
transform 1 0 2484 0 -1 318240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1789
timestamp 1586364061
transform 1 0 3956 0 -1 318240
box -38 -48 130 592
use scs8hd_decap_4  FILLER_580_27
timestamp 1586364061
transform 1 0 3588 0 -1 318240
box -38 -48 406 592
use scs8hd_decap_12  FILLER_580_32
timestamp 1586364061
transform 1 0 4048 0 -1 318240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_580_44
timestamp 1586364061
transform 1 0 5152 0 -1 318240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_580_56
timestamp 1586364061
transform 1 0 6256 0 -1 318240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_580_68
timestamp 1586364061
transform 1 0 7360 0 -1 318240
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1161
timestamp 1586364061
transform -1 0 8832 0 -1 318240
box -38 -48 314 592
use scs8hd_fill_1  FILLER_580_80
timestamp 1586364061
transform 1 0 8464 0 -1 318240
box -38 -48 130 592
use scs8hd_decap_3  PHY_1162
timestamp 1586364061
transform 1 0 1104 0 1 318240
box -38 -48 314 592
use scs8hd_decap_3  PHY_1164
timestamp 1586364061
transform 1 0 1104 0 -1 319328
box -38 -48 314 592
use scs8hd_decap_12  FILLER_581_3
timestamp 1586364061
transform 1 0 1380 0 1 318240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_581_15
timestamp 1586364061
transform 1 0 2484 0 1 318240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_582_3
timestamp 1586364061
transform 1 0 1380 0 -1 319328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_582_15
timestamp 1586364061
transform 1 0 2484 0 -1 319328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1791
timestamp 1586364061
transform 1 0 3956 0 -1 319328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_581_27
timestamp 1586364061
transform 1 0 3588 0 1 318240
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_582_27
timestamp 1586364061
transform 1 0 3588 0 -1 319328
box -38 -48 406 592
use scs8hd_decap_12  FILLER_582_32
timestamp 1586364061
transform 1 0 4048 0 -1 319328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_581_39
timestamp 1586364061
transform 1 0 4692 0 1 318240
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_581_51
timestamp 1586364061
transform 1 0 5796 0 1 318240
box -38 -48 774 592
use scs8hd_decap_12  FILLER_582_44
timestamp 1586364061
transform 1 0 5152 0 -1 319328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1790
timestamp 1586364061
transform 1 0 6716 0 1 318240
box -38 -48 130 592
use scs8hd_fill_2  FILLER_581_59
timestamp 1586364061
transform 1 0 6532 0 1 318240
box -38 -48 222 592
use scs8hd_decap_12  FILLER_581_62
timestamp 1586364061
transform 1 0 6808 0 1 318240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_582_56
timestamp 1586364061
transform 1 0 6256 0 -1 319328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_582_68
timestamp 1586364061
transform 1 0 7360 0 -1 319328
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1163
timestamp 1586364061
transform -1 0 8832 0 1 318240
box -38 -48 314 592
use scs8hd_decap_3  PHY_1165
timestamp 1586364061
transform -1 0 8832 0 -1 319328
box -38 -48 314 592
use scs8hd_decap_6  FILLER_581_74
timestamp 1586364061
transform 1 0 7912 0 1 318240
box -38 -48 590 592
use scs8hd_fill_1  FILLER_581_80
timestamp 1586364061
transform 1 0 8464 0 1 318240
box -38 -48 130 592
use scs8hd_fill_1  FILLER_582_80
timestamp 1586364061
transform 1 0 8464 0 -1 319328
box -38 -48 130 592
use scs8hd_decap_3  PHY_1166
timestamp 1586364061
transform 1 0 1104 0 1 319328
box -38 -48 314 592
use scs8hd_decap_12  FILLER_583_3
timestamp 1586364061
transform 1 0 1380 0 1 319328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_583_15
timestamp 1586364061
transform 1 0 2484 0 1 319328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_583_27
timestamp 1586364061
transform 1 0 3588 0 1 319328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_583_39
timestamp 1586364061
transform 1 0 4692 0 1 319328
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_583_51
timestamp 1586364061
transform 1 0 5796 0 1 319328
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1792
timestamp 1586364061
transform 1 0 6716 0 1 319328
box -38 -48 130 592
use scs8hd_fill_2  FILLER_583_59
timestamp 1586364061
transform 1 0 6532 0 1 319328
box -38 -48 222 592
use scs8hd_decap_12  FILLER_583_62
timestamp 1586364061
transform 1 0 6808 0 1 319328
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1167
timestamp 1586364061
transform -1 0 8832 0 1 319328
box -38 -48 314 592
use scs8hd_decap_6  FILLER_583_74
timestamp 1586364061
transform 1 0 7912 0 1 319328
box -38 -48 590 592
use scs8hd_fill_1  FILLER_583_80
timestamp 1586364061
transform 1 0 8464 0 1 319328
box -38 -48 130 592
use scs8hd_decap_3  PHY_1168
timestamp 1586364061
transform 1 0 1104 0 -1 320416
box -38 -48 314 592
use scs8hd_decap_12  FILLER_584_3
timestamp 1586364061
transform 1 0 1380 0 -1 320416
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_584_15
timestamp 1586364061
transform 1 0 2484 0 -1 320416
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1793
timestamp 1586364061
transform 1 0 3956 0 -1 320416
box -38 -48 130 592
use scs8hd_decap_4  FILLER_584_27
timestamp 1586364061
transform 1 0 3588 0 -1 320416
box -38 -48 406 592
use scs8hd_decap_12  FILLER_584_32
timestamp 1586364061
transform 1 0 4048 0 -1 320416
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_584_44
timestamp 1586364061
transform 1 0 5152 0 -1 320416
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_584_56
timestamp 1586364061
transform 1 0 6256 0 -1 320416
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_584_68
timestamp 1586364061
transform 1 0 7360 0 -1 320416
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1169
timestamp 1586364061
transform -1 0 8832 0 -1 320416
box -38 -48 314 592
use scs8hd_fill_1  FILLER_584_80
timestamp 1586364061
transform 1 0 8464 0 -1 320416
box -38 -48 130 592
use scs8hd_decap_3  PHY_1170
timestamp 1586364061
transform 1 0 1104 0 1 320416
box -38 -48 314 592
use scs8hd_decap_12  FILLER_585_3
timestamp 1586364061
transform 1 0 1380 0 1 320416
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_585_15
timestamp 1586364061
transform 1 0 2484 0 1 320416
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_585_27
timestamp 1586364061
transform 1 0 3588 0 1 320416
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_585_39
timestamp 1586364061
transform 1 0 4692 0 1 320416
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_585_51
timestamp 1586364061
transform 1 0 5796 0 1 320416
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1794
timestamp 1586364061
transform 1 0 6716 0 1 320416
box -38 -48 130 592
use scs8hd_fill_2  FILLER_585_59
timestamp 1586364061
transform 1 0 6532 0 1 320416
box -38 -48 222 592
use scs8hd_decap_12  FILLER_585_62
timestamp 1586364061
transform 1 0 6808 0 1 320416
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1171
timestamp 1586364061
transform -1 0 8832 0 1 320416
box -38 -48 314 592
use scs8hd_decap_6  FILLER_585_74
timestamp 1586364061
transform 1 0 7912 0 1 320416
box -38 -48 590 592
use scs8hd_fill_1  FILLER_585_80
timestamp 1586364061
transform 1 0 8464 0 1 320416
box -38 -48 130 592
use scs8hd_decap_3  PHY_1172
timestamp 1586364061
transform 1 0 1104 0 -1 321504
box -38 -48 314 592
use scs8hd_decap_12  FILLER_586_3
timestamp 1586364061
transform 1 0 1380 0 -1 321504
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_586_15
timestamp 1586364061
transform 1 0 2484 0 -1 321504
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1795
timestamp 1586364061
transform 1 0 3956 0 -1 321504
box -38 -48 130 592
use scs8hd_decap_4  FILLER_586_27
timestamp 1586364061
transform 1 0 3588 0 -1 321504
box -38 -48 406 592
use scs8hd_decap_12  FILLER_586_32
timestamp 1586364061
transform 1 0 4048 0 -1 321504
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_586_44
timestamp 1586364061
transform 1 0 5152 0 -1 321504
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_586_56
timestamp 1586364061
transform 1 0 6256 0 -1 321504
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_586_68
timestamp 1586364061
transform 1 0 7360 0 -1 321504
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1173
timestamp 1586364061
transform -1 0 8832 0 -1 321504
box -38 -48 314 592
use scs8hd_fill_1  FILLER_586_80
timestamp 1586364061
transform 1 0 8464 0 -1 321504
box -38 -48 130 592
use scs8hd_decap_3  PHY_1174
timestamp 1586364061
transform 1 0 1104 0 1 321504
box -38 -48 314 592
use scs8hd_decap_12  FILLER_587_3
timestamp 1586364061
transform 1 0 1380 0 1 321504
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_587_15
timestamp 1586364061
transform 1 0 2484 0 1 321504
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_587_27
timestamp 1586364061
transform 1 0 3588 0 1 321504
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_587_39
timestamp 1586364061
transform 1 0 4692 0 1 321504
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_587_51
timestamp 1586364061
transform 1 0 5796 0 1 321504
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1796
timestamp 1586364061
transform 1 0 6716 0 1 321504
box -38 -48 130 592
use scs8hd_fill_2  FILLER_587_59
timestamp 1586364061
transform 1 0 6532 0 1 321504
box -38 -48 222 592
use scs8hd_decap_12  FILLER_587_62
timestamp 1586364061
transform 1 0 6808 0 1 321504
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1175
timestamp 1586364061
transform -1 0 8832 0 1 321504
box -38 -48 314 592
use scs8hd_decap_6  FILLER_587_74
timestamp 1586364061
transform 1 0 7912 0 1 321504
box -38 -48 590 592
use scs8hd_fill_1  FILLER_587_80
timestamp 1586364061
transform 1 0 8464 0 1 321504
box -38 -48 130 592
use scs8hd_decap_3  PHY_1176
timestamp 1586364061
transform 1 0 1104 0 -1 322592
box -38 -48 314 592
use scs8hd_decap_3  PHY_1178
timestamp 1586364061
transform 1 0 1104 0 1 322592
box -38 -48 314 592
use scs8hd_decap_12  FILLER_588_3
timestamp 1586364061
transform 1 0 1380 0 -1 322592
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_588_15
timestamp 1586364061
transform 1 0 2484 0 -1 322592
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_589_3
timestamp 1586364061
transform 1 0 1380 0 1 322592
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_589_15
timestamp 1586364061
transform 1 0 2484 0 1 322592
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1797
timestamp 1586364061
transform 1 0 3956 0 -1 322592
box -38 -48 130 592
use scs8hd_decap_4  FILLER_588_27
timestamp 1586364061
transform 1 0 3588 0 -1 322592
box -38 -48 406 592
use scs8hd_decap_12  FILLER_588_32
timestamp 1586364061
transform 1 0 4048 0 -1 322592
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_589_27
timestamp 1586364061
transform 1 0 3588 0 1 322592
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_588_44
timestamp 1586364061
transform 1 0 5152 0 -1 322592
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_589_39
timestamp 1586364061
transform 1 0 4692 0 1 322592
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_589_51
timestamp 1586364061
transform 1 0 5796 0 1 322592
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1798
timestamp 1586364061
transform 1 0 6716 0 1 322592
box -38 -48 130 592
use scs8hd_decap_12  FILLER_588_56
timestamp 1586364061
transform 1 0 6256 0 -1 322592
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_588_68
timestamp 1586364061
transform 1 0 7360 0 -1 322592
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_589_59
timestamp 1586364061
transform 1 0 6532 0 1 322592
box -38 -48 222 592
use scs8hd_decap_12  FILLER_589_62
timestamp 1586364061
transform 1 0 6808 0 1 322592
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1177
timestamp 1586364061
transform -1 0 8832 0 -1 322592
box -38 -48 314 592
use scs8hd_decap_3  PHY_1179
timestamp 1586364061
transform -1 0 8832 0 1 322592
box -38 -48 314 592
use scs8hd_fill_1  FILLER_588_80
timestamp 1586364061
transform 1 0 8464 0 -1 322592
box -38 -48 130 592
use scs8hd_decap_6  FILLER_589_74
timestamp 1586364061
transform 1 0 7912 0 1 322592
box -38 -48 590 592
use scs8hd_fill_1  FILLER_589_80
timestamp 1586364061
transform 1 0 8464 0 1 322592
box -38 -48 130 592
use scs8hd_decap_3  PHY_1180
timestamp 1586364061
transform 1 0 1104 0 -1 323680
box -38 -48 314 592
use scs8hd_decap_12  FILLER_590_3
timestamp 1586364061
transform 1 0 1380 0 -1 323680
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_590_15
timestamp 1586364061
transform 1 0 2484 0 -1 323680
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1799
timestamp 1586364061
transform 1 0 3956 0 -1 323680
box -38 -48 130 592
use scs8hd_decap_4  FILLER_590_27
timestamp 1586364061
transform 1 0 3588 0 -1 323680
box -38 -48 406 592
use scs8hd_decap_12  FILLER_590_32
timestamp 1586364061
transform 1 0 4048 0 -1 323680
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_590_44
timestamp 1586364061
transform 1 0 5152 0 -1 323680
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_590_56
timestamp 1586364061
transform 1 0 6256 0 -1 323680
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_590_68
timestamp 1586364061
transform 1 0 7360 0 -1 323680
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1181
timestamp 1586364061
transform -1 0 8832 0 -1 323680
box -38 -48 314 592
use scs8hd_fill_1  FILLER_590_80
timestamp 1586364061
transform 1 0 8464 0 -1 323680
box -38 -48 130 592
use scs8hd_decap_3  PHY_1182
timestamp 1586364061
transform 1 0 1104 0 1 323680
box -38 -48 314 592
use scs8hd_decap_12  FILLER_591_3
timestamp 1586364061
transform 1 0 1380 0 1 323680
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_591_15
timestamp 1586364061
transform 1 0 2484 0 1 323680
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_591_27
timestamp 1586364061
transform 1 0 3588 0 1 323680
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_591_39
timestamp 1586364061
transform 1 0 4692 0 1 323680
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_591_51
timestamp 1586364061
transform 1 0 5796 0 1 323680
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1800
timestamp 1586364061
transform 1 0 6716 0 1 323680
box -38 -48 130 592
use scs8hd_fill_2  FILLER_591_59
timestamp 1586364061
transform 1 0 6532 0 1 323680
box -38 -48 222 592
use scs8hd_decap_12  FILLER_591_62
timestamp 1586364061
transform 1 0 6808 0 1 323680
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1183
timestamp 1586364061
transform -1 0 8832 0 1 323680
box -38 -48 314 592
use scs8hd_decap_6  FILLER_591_74
timestamp 1586364061
transform 1 0 7912 0 1 323680
box -38 -48 590 592
use scs8hd_fill_1  FILLER_591_80
timestamp 1586364061
transform 1 0 8464 0 1 323680
box -38 -48 130 592
use scs8hd_decap_3  PHY_1184
timestamp 1586364061
transform 1 0 1104 0 -1 324768
box -38 -48 314 592
use scs8hd_decap_12  FILLER_592_3
timestamp 1586364061
transform 1 0 1380 0 -1 324768
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_592_15
timestamp 1586364061
transform 1 0 2484 0 -1 324768
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1801
timestamp 1586364061
transform 1 0 3956 0 -1 324768
box -38 -48 130 592
use scs8hd_decap_4  FILLER_592_27
timestamp 1586364061
transform 1 0 3588 0 -1 324768
box -38 -48 406 592
use scs8hd_decap_12  FILLER_592_32
timestamp 1586364061
transform 1 0 4048 0 -1 324768
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_592_44
timestamp 1586364061
transform 1 0 5152 0 -1 324768
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_592_56
timestamp 1586364061
transform 1 0 6256 0 -1 324768
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_592_68
timestamp 1586364061
transform 1 0 7360 0 -1 324768
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1185
timestamp 1586364061
transform -1 0 8832 0 -1 324768
box -38 -48 314 592
use scs8hd_fill_1  FILLER_592_80
timestamp 1586364061
transform 1 0 8464 0 -1 324768
box -38 -48 130 592
use scs8hd_decap_3  PHY_1186
timestamp 1586364061
transform 1 0 1104 0 1 324768
box -38 -48 314 592
use scs8hd_decap_12  FILLER_593_3
timestamp 1586364061
transform 1 0 1380 0 1 324768
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_593_15
timestamp 1586364061
transform 1 0 2484 0 1 324768
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_593_27
timestamp 1586364061
transform 1 0 3588 0 1 324768
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_593_39
timestamp 1586364061
transform 1 0 4692 0 1 324768
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_593_51
timestamp 1586364061
transform 1 0 5796 0 1 324768
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1802
timestamp 1586364061
transform 1 0 6716 0 1 324768
box -38 -48 130 592
use scs8hd_fill_2  FILLER_593_59
timestamp 1586364061
transform 1 0 6532 0 1 324768
box -38 -48 222 592
use scs8hd_decap_12  FILLER_593_62
timestamp 1586364061
transform 1 0 6808 0 1 324768
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1187
timestamp 1586364061
transform -1 0 8832 0 1 324768
box -38 -48 314 592
use scs8hd_decap_6  FILLER_593_74
timestamp 1586364061
transform 1 0 7912 0 1 324768
box -38 -48 590 592
use scs8hd_fill_1  FILLER_593_80
timestamp 1586364061
transform 1 0 8464 0 1 324768
box -38 -48 130 592
use scs8hd_decap_3  PHY_1188
timestamp 1586364061
transform 1 0 1104 0 -1 325856
box -38 -48 314 592
use scs8hd_decap_3  PHY_1190
timestamp 1586364061
transform 1 0 1104 0 1 325856
box -38 -48 314 592
use scs8hd_decap_12  FILLER_594_3
timestamp 1586364061
transform 1 0 1380 0 -1 325856
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_594_15
timestamp 1586364061
transform 1 0 2484 0 -1 325856
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_595_3
timestamp 1586364061
transform 1 0 1380 0 1 325856
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_595_15
timestamp 1586364061
transform 1 0 2484 0 1 325856
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1803
timestamp 1586364061
transform 1 0 3956 0 -1 325856
box -38 -48 130 592
use scs8hd_decap_4  FILLER_594_27
timestamp 1586364061
transform 1 0 3588 0 -1 325856
box -38 -48 406 592
use scs8hd_decap_12  FILLER_594_32
timestamp 1586364061
transform 1 0 4048 0 -1 325856
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_595_27
timestamp 1586364061
transform 1 0 3588 0 1 325856
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_594_44
timestamp 1586364061
transform 1 0 5152 0 -1 325856
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_595_39
timestamp 1586364061
transform 1 0 4692 0 1 325856
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_595_51
timestamp 1586364061
transform 1 0 5796 0 1 325856
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1804
timestamp 1586364061
transform 1 0 6716 0 1 325856
box -38 -48 130 592
use scs8hd_decap_12  FILLER_594_56
timestamp 1586364061
transform 1 0 6256 0 -1 325856
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_594_68
timestamp 1586364061
transform 1 0 7360 0 -1 325856
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_595_59
timestamp 1586364061
transform 1 0 6532 0 1 325856
box -38 -48 222 592
use scs8hd_decap_12  FILLER_595_62
timestamp 1586364061
transform 1 0 6808 0 1 325856
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1189
timestamp 1586364061
transform -1 0 8832 0 -1 325856
box -38 -48 314 592
use scs8hd_decap_3  PHY_1191
timestamp 1586364061
transform -1 0 8832 0 1 325856
box -38 -48 314 592
use scs8hd_fill_1  FILLER_594_80
timestamp 1586364061
transform 1 0 8464 0 -1 325856
box -38 -48 130 592
use scs8hd_decap_6  FILLER_595_74
timestamp 1586364061
transform 1 0 7912 0 1 325856
box -38 -48 590 592
use scs8hd_fill_1  FILLER_595_80
timestamp 1586364061
transform 1 0 8464 0 1 325856
box -38 -48 130 592
use scs8hd_decap_3  PHY_1192
timestamp 1586364061
transform 1 0 1104 0 -1 326944
box -38 -48 314 592
use scs8hd_decap_12  FILLER_596_3
timestamp 1586364061
transform 1 0 1380 0 -1 326944
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_596_15
timestamp 1586364061
transform 1 0 2484 0 -1 326944
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1805
timestamp 1586364061
transform 1 0 3956 0 -1 326944
box -38 -48 130 592
use scs8hd_decap_4  FILLER_596_27
timestamp 1586364061
transform 1 0 3588 0 -1 326944
box -38 -48 406 592
use scs8hd_decap_12  FILLER_596_32
timestamp 1586364061
transform 1 0 4048 0 -1 326944
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_596_44
timestamp 1586364061
transform 1 0 5152 0 -1 326944
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_596_56
timestamp 1586364061
transform 1 0 6256 0 -1 326944
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_596_68
timestamp 1586364061
transform 1 0 7360 0 -1 326944
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1193
timestamp 1586364061
transform -1 0 8832 0 -1 326944
box -38 -48 314 592
use scs8hd_fill_1  FILLER_596_80
timestamp 1586364061
transform 1 0 8464 0 -1 326944
box -38 -48 130 592
use scs8hd_decap_3  PHY_1194
timestamp 1586364061
transform 1 0 1104 0 1 326944
box -38 -48 314 592
use scs8hd_decap_12  FILLER_597_3
timestamp 1586364061
transform 1 0 1380 0 1 326944
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_597_15
timestamp 1586364061
transform 1 0 2484 0 1 326944
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_597_27
timestamp 1586364061
transform 1 0 3588 0 1 326944
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_597_39
timestamp 1586364061
transform 1 0 4692 0 1 326944
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_597_51
timestamp 1586364061
transform 1 0 5796 0 1 326944
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1806
timestamp 1586364061
transform 1 0 6716 0 1 326944
box -38 -48 130 592
use scs8hd_fill_2  FILLER_597_59
timestamp 1586364061
transform 1 0 6532 0 1 326944
box -38 -48 222 592
use scs8hd_decap_12  FILLER_597_62
timestamp 1586364061
transform 1 0 6808 0 1 326944
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1195
timestamp 1586364061
transform -1 0 8832 0 1 326944
box -38 -48 314 592
use scs8hd_decap_6  FILLER_597_74
timestamp 1586364061
transform 1 0 7912 0 1 326944
box -38 -48 590 592
use scs8hd_fill_1  FILLER_597_80
timestamp 1586364061
transform 1 0 8464 0 1 326944
box -38 -48 130 592
use scs8hd_decap_3  PHY_1196
timestamp 1586364061
transform 1 0 1104 0 -1 328032
box -38 -48 314 592
use scs8hd_decap_12  FILLER_598_3
timestamp 1586364061
transform 1 0 1380 0 -1 328032
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_598_15
timestamp 1586364061
transform 1 0 2484 0 -1 328032
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1807
timestamp 1586364061
transform 1 0 3956 0 -1 328032
box -38 -48 130 592
use scs8hd_decap_4  FILLER_598_27
timestamp 1586364061
transform 1 0 3588 0 -1 328032
box -38 -48 406 592
use scs8hd_decap_12  FILLER_598_32
timestamp 1586364061
transform 1 0 4048 0 -1 328032
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_598_44
timestamp 1586364061
transform 1 0 5152 0 -1 328032
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_598_56
timestamp 1586364061
transform 1 0 6256 0 -1 328032
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_598_68
timestamp 1586364061
transform 1 0 7360 0 -1 328032
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1197
timestamp 1586364061
transform -1 0 8832 0 -1 328032
box -38 -48 314 592
use scs8hd_fill_1  FILLER_598_80
timestamp 1586364061
transform 1 0 8464 0 -1 328032
box -38 -48 130 592
use scs8hd_decap_3  PHY_1198
timestamp 1586364061
transform 1 0 1104 0 1 328032
box -38 -48 314 592
use scs8hd_decap_12  FILLER_599_3
timestamp 1586364061
transform 1 0 1380 0 1 328032
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_599_15
timestamp 1586364061
transform 1 0 2484 0 1 328032
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_599_27
timestamp 1586364061
transform 1 0 3588 0 1 328032
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_599_39
timestamp 1586364061
transform 1 0 4692 0 1 328032
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_599_51
timestamp 1586364061
transform 1 0 5796 0 1 328032
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_1808
timestamp 1586364061
transform 1 0 6716 0 1 328032
box -38 -48 130 592
use scs8hd_fill_2  FILLER_599_59
timestamp 1586364061
transform 1 0 6532 0 1 328032
box -38 -48 222 592
use scs8hd_decap_12  FILLER_599_62
timestamp 1586364061
transform 1 0 6808 0 1 328032
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1199
timestamp 1586364061
transform -1 0 8832 0 1 328032
box -38 -48 314 592
use scs8hd_decap_6  FILLER_599_74
timestamp 1586364061
transform 1 0 7912 0 1 328032
box -38 -48 590 592
use scs8hd_fill_1  FILLER_599_80
timestamp 1586364061
transform 1 0 8464 0 1 328032
box -38 -48 130 592
use scs8hd_decap_3  PHY_1200
timestamp 1586364061
transform 1 0 1104 0 -1 329120
box -38 -48 314 592
use scs8hd_decap_12  FILLER_600_3
timestamp 1586364061
transform 1 0 1380 0 -1 329120
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_600_15
timestamp 1586364061
transform 1 0 2484 0 -1 329120
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1809
timestamp 1586364061
transform 1 0 3956 0 -1 329120
box -38 -48 130 592
use scs8hd_decap_4  FILLER_600_27
timestamp 1586364061
transform 1 0 3588 0 -1 329120
box -38 -48 406 592
use scs8hd_decap_12  FILLER_600_32
timestamp 1586364061
transform 1 0 4048 0 -1 329120
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_600_44
timestamp 1586364061
transform 1 0 5152 0 -1 329120
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_600_56
timestamp 1586364061
transform 1 0 6256 0 -1 329120
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_600_68
timestamp 1586364061
transform 1 0 7360 0 -1 329120
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1201
timestamp 1586364061
transform -1 0 8832 0 -1 329120
box -38 -48 314 592
use scs8hd_fill_1  FILLER_600_80
timestamp 1586364061
transform 1 0 8464 0 -1 329120
box -38 -48 130 592
use scs8hd_decap_3  PHY_1202
timestamp 1586364061
transform 1 0 1104 0 1 329120
box -38 -48 314 592
use scs8hd_decap_3  PHY_1204
timestamp 1586364061
transform 1 0 1104 0 -1 330208
box -38 -48 314 592
use scs8hd_decap_12  FILLER_601_3
timestamp 1586364061
transform 1 0 1380 0 1 329120
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_601_15
timestamp 1586364061
transform 1 0 2484 0 1 329120
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_602_3
timestamp 1586364061
transform 1 0 1380 0 -1 330208
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_602_15
timestamp 1586364061
transform 1 0 2484 0 -1 330208
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1811
timestamp 1586364061
transform 1 0 3956 0 -1 330208
box -38 -48 130 592
use scs8hd_decap_12  FILLER_601_27
timestamp 1586364061
transform 1 0 3588 0 1 329120
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_602_27
timestamp 1586364061
transform 1 0 3588 0 -1 330208
box -38 -48 406 592
use scs8hd_decap_12  FILLER_602_32
timestamp 1586364061
transform 1 0 4048 0 -1 330208
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_601_39
timestamp 1586364061
transform 1 0 4692 0 1 329120
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_601_51
timestamp 1586364061
transform 1 0 5796 0 1 329120
box -38 -48 774 592
use scs8hd_decap_12  FILLER_602_44
timestamp 1586364061
transform 1 0 5152 0 -1 330208
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1810
timestamp 1586364061
transform 1 0 6716 0 1 329120
box -38 -48 130 592
use scs8hd_fill_2  FILLER_601_59
timestamp 1586364061
transform 1 0 6532 0 1 329120
box -38 -48 222 592
use scs8hd_decap_12  FILLER_601_62
timestamp 1586364061
transform 1 0 6808 0 1 329120
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_602_56
timestamp 1586364061
transform 1 0 6256 0 -1 330208
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_602_68
timestamp 1586364061
transform 1 0 7360 0 -1 330208
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1203
timestamp 1586364061
transform -1 0 8832 0 1 329120
box -38 -48 314 592
use scs8hd_decap_3  PHY_1205
timestamp 1586364061
transform -1 0 8832 0 -1 330208
box -38 -48 314 592
use scs8hd_decap_6  FILLER_601_74
timestamp 1586364061
transform 1 0 7912 0 1 329120
box -38 -48 590 592
use scs8hd_fill_1  FILLER_601_80
timestamp 1586364061
transform 1 0 8464 0 1 329120
box -38 -48 130 592
use scs8hd_fill_1  FILLER_602_80
timestamp 1586364061
transform 1 0 8464 0 -1 330208
box -38 -48 130 592
use scs8hd_decap_3  PHY_1206
timestamp 1586364061
transform 1 0 1104 0 1 330208
box -38 -48 314 592
use scs8hd_decap_12  FILLER_603_3
timestamp 1586364061
transform 1 0 1380 0 1 330208
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_603_15
timestamp 1586364061
transform 1 0 2484 0 1 330208
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1812
timestamp 1586364061
transform 1 0 3956 0 1 330208
box -38 -48 130 592
use scs8hd_decap_4  FILLER_603_27
timestamp 1586364061
transform 1 0 3588 0 1 330208
box -38 -48 406 592
use scs8hd_decap_12  FILLER_603_32
timestamp 1586364061
transform 1 0 4048 0 1 330208
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_603_44
timestamp 1586364061
transform 1 0 5152 0 1 330208
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_1813
timestamp 1586364061
transform 1 0 6808 0 1 330208
box -38 -48 130 592
use scs8hd_decap_6  FILLER_603_56
timestamp 1586364061
transform 1 0 6256 0 1 330208
box -38 -48 590 592
use scs8hd_decap_12  FILLER_603_63
timestamp 1586364061
transform 1 0 6900 0 1 330208
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1207
timestamp 1586364061
transform -1 0 8832 0 1 330208
box -38 -48 314 592
use scs8hd_decap_6  FILLER_603_75
timestamp 1586364061
transform 1 0 8004 0 1 330208
box -38 -48 590 592
<< labels >>
rlabel metal2 s 4894 0 4950 480 6 address[0]
port 0 nsew default input
rlabel metal3 s 9520 16600 10000 16720 6 address[1]
port 1 nsew default input
rlabel metal2 s 570 332520 626 333000 6 address[2]
port 2 nsew default input
rlabel metal2 s 1766 332520 1822 333000 6 address[3]
port 3 nsew default input
rlabel metal2 s 2870 0 2926 480 6 data_in
port 4 nsew default input
rlabel metal2 s 938 0 994 480 6 enable
port 5 nsew default input
rlabel metal3 s 9520 49784 10000 49904 6 gfpga_pad_GPIO_PAD[0]
port 6 nsew default bidirectional
rlabel metal2 s 3054 332520 3110 333000 6 gfpga_pad_GPIO_PAD[1]
port 7 nsew default bidirectional
rlabel metal3 s 0 23672 480 23792 6 gfpga_pad_GPIO_PAD[2]
port 8 nsew default bidirectional
rlabel metal3 s 9520 83104 10000 83224 6 gfpga_pad_GPIO_PAD[3]
port 9 nsew default bidirectional
rlabel metal2 s 6918 0 6974 480 6 gfpga_pad_GPIO_PAD[4]
port 10 nsew default bidirectional
rlabel metal3 s 0 71136 480 71256 6 gfpga_pad_GPIO_PAD[5]
port 11 nsew default bidirectional
rlabel metal3 s 9520 116424 10000 116544 6 gfpga_pad_GPIO_PAD[6]
port 12 nsew default bidirectional
rlabel metal3 s 9520 149744 10000 149864 6 gfpga_pad_GPIO_PAD[7]
port 13 nsew default bidirectional
rlabel metal2 s 4250 332520 4306 333000 6 left_width_0_height_0__pin_0_
port 14 nsew default input
rlabel metal3 s 9520 283024 10000 283144 6 left_width_0_height_0__pin_10_
port 15 nsew default input
rlabel metal2 s 8942 0 8998 480 6 left_width_0_height_0__pin_11_
port 16 nsew default tristate
rlabel metal3 s 0 213936 480 214056 6 left_width_0_height_0__pin_12_
port 17 nsew default input
rlabel metal3 s 9520 316344 10000 316464 6 left_width_0_height_0__pin_13_
port 18 nsew default tristate
rlabel metal3 s 0 261536 480 261656 6 left_width_0_height_0__pin_14_
port 19 nsew default input
rlabel metal3 s 0 309136 480 309256 6 left_width_0_height_0__pin_15_
port 20 nsew default tristate
rlabel metal3 s 9520 183064 10000 183184 6 left_width_0_height_0__pin_1_
port 21 nsew default tristate
rlabel metal3 s 0 118736 480 118856 6 left_width_0_height_0__pin_2_
port 22 nsew default input
rlabel metal3 s 9520 216384 10000 216504 6 left_width_0_height_0__pin_3_
port 23 nsew default tristate
rlabel metal2 s 5538 332520 5594 333000 6 left_width_0_height_0__pin_4_
port 24 nsew default input
rlabel metal3 s 9520 249704 10000 249824 6 left_width_0_height_0__pin_5_
port 25 nsew default tristate
rlabel metal2 s 6826 332520 6882 333000 6 left_width_0_height_0__pin_6_
port 26 nsew default input
rlabel metal2 s 8022 332520 8078 333000 6 left_width_0_height_0__pin_7_
port 27 nsew default tristate
rlabel metal2 s 9310 332520 9366 333000 6 left_width_0_height_0__pin_8_
port 28 nsew default input
rlabel metal3 s 0 166336 480 166456 6 left_width_0_height_0__pin_9_
port 29 nsew default tristate
rlabel metal4 s 2611 2128 2931 330800 6 vpwr
port 30 nsew default input
rlabel metal4 s 4277 2128 4597 330800 6 vgnd
port 31 nsew default input
<< end >>
