magic
tech sky130A
magscale 1 2
timestamp 1605110728
<< locali >>
rect 15485 11611 15519 11849
rect 7941 10455 7975 10693
<< viali >>
rect 4905 20553 4939 20587
rect 7021 20553 7055 20587
rect 8125 20553 8159 20587
rect 10149 20553 10183 20587
rect 18245 20553 18279 20587
rect 16681 20485 16715 20519
rect 25789 20485 25823 20519
rect 20545 20417 20579 20451
rect 4721 20349 4755 20383
rect 6837 20349 6871 20383
rect 7941 20349 7975 20383
rect 14105 20349 14139 20383
rect 14749 20349 14783 20383
rect 15393 20349 15427 20383
rect 16497 20349 16531 20383
rect 18061 20349 18095 20383
rect 19993 20349 20027 20383
rect 21097 20349 21131 20383
rect 21649 20349 21683 20383
rect 24225 20349 24259 20383
rect 24777 20349 24811 20383
rect 25605 20349 25639 20383
rect 26157 20349 26191 20383
rect 26709 20349 26743 20383
rect 7481 20281 7515 20315
rect 5365 20213 5399 20247
rect 8585 20213 8619 20247
rect 14289 20213 14323 20247
rect 15577 20213 15611 20247
rect 16037 20213 16071 20247
rect 17049 20213 17083 20247
rect 18705 20213 18739 20247
rect 20177 20213 20211 20247
rect 21281 20213 21315 20247
rect 24409 20213 24443 20247
rect 26893 20213 26927 20247
rect 27261 20213 27295 20247
rect 16589 20009 16623 20043
rect 26709 20009 26743 20043
rect 15301 19873 15335 19907
rect 16405 19873 16439 19907
rect 26525 19873 26559 19907
rect 15485 19737 15519 19771
rect 15393 19397 15427 19431
rect 16497 19329 16531 19363
rect 26525 19125 26559 19159
rect 8585 13345 8619 13379
rect 10057 13345 10091 13379
rect 11612 13345 11646 13379
rect 2513 13277 2547 13311
rect 10149 13277 10183 13311
rect 10241 13277 10275 13311
rect 11345 13277 11379 13311
rect 9689 13209 9723 13243
rect 11069 13209 11103 13243
rect 3065 13141 3099 13175
rect 9137 13141 9171 13175
rect 10701 13141 10735 13175
rect 12725 13141 12759 13175
rect 10425 12937 10459 12971
rect 13829 12937 13863 12971
rect 15117 12937 15151 12971
rect 10057 12869 10091 12903
rect 11621 12869 11655 12903
rect 3157 12801 3191 12835
rect 4077 12801 4111 12835
rect 9597 12801 9631 12835
rect 11161 12801 11195 12835
rect 12173 12801 12207 12835
rect 1409 12733 1443 12767
rect 2973 12733 3007 12767
rect 4261 12733 4295 12767
rect 4517 12733 4551 12767
rect 8953 12733 8987 12767
rect 9413 12733 9447 12767
rect 10977 12733 11011 12767
rect 12449 12733 12483 12767
rect 12716 12733 12750 12767
rect 15301 12733 15335 12767
rect 15557 12733 15591 12767
rect 2421 12665 2455 12699
rect 2881 12665 2915 12699
rect 11069 12665 11103 12699
rect 1593 12597 1627 12631
rect 1961 12597 1995 12631
rect 2513 12597 2547 12631
rect 5641 12597 5675 12631
rect 9045 12597 9079 12631
rect 9505 12597 9539 12631
rect 10609 12597 10643 12631
rect 14749 12597 14783 12631
rect 16681 12597 16715 12631
rect 1593 12393 1627 12427
rect 7941 12393 7975 12427
rect 8401 12393 8435 12427
rect 10977 12393 11011 12427
rect 11345 12393 11379 12427
rect 12449 12393 12483 12427
rect 5702 12325 5736 12359
rect 17570 12325 17604 12359
rect 2789 12257 2823 12291
rect 2881 12257 2915 12291
rect 10333 12257 10367 12291
rect 10425 12257 10459 12291
rect 17325 12257 17359 12291
rect 3065 12189 3099 12223
rect 4353 12189 4387 12223
rect 5457 12189 5491 12223
rect 8493 12189 8527 12223
rect 8585 12189 8619 12223
rect 10517 12189 10551 12223
rect 15301 12189 15335 12223
rect 15761 12189 15795 12223
rect 2237 12121 2271 12155
rect 2421 12053 2455 12087
rect 3433 12053 3467 12087
rect 3801 12053 3835 12087
rect 6837 12053 6871 12087
rect 8033 12053 8067 12087
rect 9137 12053 9171 12087
rect 9505 12053 9539 12087
rect 9965 12053 9999 12087
rect 14289 12053 14323 12087
rect 18705 12053 18739 12087
rect 2053 11849 2087 11883
rect 8125 11849 8159 11883
rect 15485 11849 15519 11883
rect 15577 11849 15611 11883
rect 17693 11849 17727 11883
rect 1685 11781 1719 11815
rect 7389 11781 7423 11815
rect 8493 11781 8527 11815
rect 2605 11713 2639 11747
rect 2697 11713 2731 11747
rect 3249 11713 3283 11747
rect 3617 11713 3651 11747
rect 4261 11713 4295 11747
rect 9045 11713 9079 11747
rect 9597 11713 9631 11747
rect 10609 11713 10643 11747
rect 14749 11713 14783 11747
rect 15301 11713 15335 11747
rect 4169 11645 4203 11679
rect 5549 11645 5583 11679
rect 8861 11645 8895 11679
rect 14565 11645 14599 11679
rect 15761 11781 15795 11815
rect 17417 11781 17451 11815
rect 16405 11713 16439 11747
rect 16129 11645 16163 11679
rect 26433 11645 26467 11679
rect 26985 11645 27019 11679
rect 4077 11577 4111 11611
rect 4721 11577 4755 11611
rect 7757 11577 7791 11611
rect 8953 11577 8987 11611
rect 10425 11577 10459 11611
rect 11437 11577 11471 11611
rect 14105 11577 14139 11611
rect 15485 11577 15519 11611
rect 16221 11577 16255 11611
rect 2145 11509 2179 11543
rect 2513 11509 2547 11543
rect 3709 11509 3743 11543
rect 5917 11509 5951 11543
rect 9873 11509 9907 11543
rect 10057 11509 10091 11543
rect 10517 11509 10551 11543
rect 11069 11509 11103 11543
rect 14197 11509 14231 11543
rect 14657 11509 14691 11543
rect 26617 11509 26651 11543
rect 2237 11305 2271 11339
rect 3617 11305 3651 11339
rect 8677 11305 8711 11339
rect 9045 11305 9079 11339
rect 9505 11305 9539 11339
rect 10425 11305 10459 11339
rect 14289 11305 14323 11339
rect 15301 11305 15335 11339
rect 15669 11305 15703 11339
rect 18429 11305 18463 11339
rect 26709 11305 26743 11339
rect 6898 11237 6932 11271
rect 10149 11237 10183 11271
rect 1777 11169 1811 11203
rect 2605 11169 2639 11203
rect 10793 11169 10827 11203
rect 26525 11169 26559 11203
rect 2697 11101 2731 11135
rect 2789 11101 2823 11135
rect 6653 11101 6687 11135
rect 10885 11101 10919 11135
rect 10977 11101 11011 11135
rect 15761 11101 15795 11135
rect 15945 11101 15979 11135
rect 18521 11101 18555 11135
rect 18613 11101 18647 11135
rect 11437 11033 11471 11067
rect 16865 11033 16899 11067
rect 18061 11033 18095 11067
rect 2145 10965 2179 10999
rect 3341 10965 3375 10999
rect 8033 10965 8067 10999
rect 16405 10965 16439 10999
rect 1593 10761 1627 10795
rect 2513 10761 2547 10795
rect 7021 10761 7055 10795
rect 8125 10761 8159 10795
rect 9597 10761 9631 10795
rect 10701 10761 10735 10795
rect 12173 10761 12207 10795
rect 15301 10761 15335 10795
rect 15853 10761 15887 10795
rect 17877 10761 17911 10795
rect 19165 10761 19199 10795
rect 27353 10761 27387 10795
rect 2053 10693 2087 10727
rect 7941 10693 7975 10727
rect 16313 10693 16347 10727
rect 3157 10625 3191 10659
rect 4721 10625 4755 10659
rect 1409 10557 1443 10591
rect 3985 10557 4019 10591
rect 2973 10489 3007 10523
rect 3617 10489 3651 10523
rect 11253 10625 11287 10659
rect 13829 10625 13863 10659
rect 16865 10625 16899 10659
rect 17049 10625 17083 10659
rect 18613 10625 18647 10659
rect 19441 10625 19475 10659
rect 19809 10625 19843 10659
rect 8217 10557 8251 10591
rect 8473 10557 8507 10591
rect 13921 10557 13955 10591
rect 14188 10557 14222 10591
rect 17509 10557 17543 10591
rect 26433 10557 26467 10591
rect 26985 10557 27019 10591
rect 10241 10489 10275 10523
rect 11069 10489 11103 10523
rect 16773 10489 16807 10523
rect 2421 10421 2455 10455
rect 2881 10421 2915 10455
rect 4077 10421 4111 10455
rect 4445 10421 4479 10455
rect 4537 10421 4571 10455
rect 7389 10421 7423 10455
rect 7941 10421 7975 10455
rect 10517 10421 10551 10455
rect 11161 10421 11195 10455
rect 11805 10421 11839 10455
rect 16405 10421 16439 10455
rect 18061 10421 18095 10455
rect 18429 10421 18463 10455
rect 18521 10421 18555 10455
rect 26617 10421 26651 10455
rect 1961 10217 1995 10251
rect 2421 10217 2455 10251
rect 2881 10217 2915 10251
rect 3525 10217 3559 10251
rect 10333 10217 10367 10251
rect 10517 10217 10551 10251
rect 13921 10217 13955 10251
rect 14381 10217 14415 10251
rect 16589 10217 16623 10251
rect 17233 10217 17267 10251
rect 2329 10149 2363 10183
rect 2789 10081 2823 10115
rect 5181 10081 5215 10115
rect 5448 10081 5482 10115
rect 10885 10081 10919 10115
rect 14749 10081 14783 10115
rect 16497 10081 16531 10115
rect 18245 10081 18279 10115
rect 18337 10081 18371 10115
rect 2973 10013 3007 10047
rect 4261 10013 4295 10047
rect 10977 10013 11011 10047
rect 11069 10013 11103 10047
rect 16681 10013 16715 10047
rect 18521 10013 18555 10047
rect 14565 9945 14599 9979
rect 18889 9945 18923 9979
rect 6561 9877 6595 9911
rect 8217 9877 8251 9911
rect 15485 9877 15519 9911
rect 16129 9877 16163 9911
rect 17877 9877 17911 9911
rect 2881 9673 2915 9707
rect 10517 9673 10551 9707
rect 11253 9673 11287 9707
rect 16497 9673 16531 9707
rect 1593 9605 1627 9639
rect 2513 9605 2547 9639
rect 2973 9605 3007 9639
rect 4537 9605 4571 9639
rect 15853 9605 15887 9639
rect 18061 9605 18095 9639
rect 2053 9537 2087 9571
rect 3433 9537 3467 9571
rect 3617 9537 3651 9571
rect 5089 9537 5123 9571
rect 5549 9537 5583 9571
rect 14841 9537 14875 9571
rect 14933 9537 14967 9571
rect 15393 9537 15427 9571
rect 17417 9537 17451 9571
rect 18521 9537 18555 9571
rect 18705 9537 18739 9571
rect 19073 9537 19107 9571
rect 1409 9469 1443 9503
rect 3341 9469 3375 9503
rect 4905 9469 4939 9503
rect 7757 9469 7791 9503
rect 8033 9469 8067 9503
rect 14749 9469 14783 9503
rect 16129 9469 16163 9503
rect 17141 9469 17175 9503
rect 19441 9469 19475 9503
rect 3985 9401 4019 9435
rect 14289 9401 14323 9435
rect 17785 9401 17819 9435
rect 18429 9401 18463 9435
rect 4445 9333 4479 9367
rect 4997 9333 5031 9367
rect 6009 9333 6043 9367
rect 7573 9333 7607 9367
rect 10977 9333 11011 9367
rect 14381 9333 14415 9367
rect 1593 9129 1627 9163
rect 2513 9129 2547 9163
rect 3433 9129 3467 9163
rect 14473 9129 14507 9163
rect 16681 9129 16715 9163
rect 26709 9129 26743 9163
rect 3065 9061 3099 9095
rect 15546 9061 15580 9095
rect 18582 9061 18616 9095
rect 1409 8993 1443 9027
rect 7481 8993 7515 9027
rect 11437 8993 11471 9027
rect 11529 8993 11563 9027
rect 15301 8993 15335 9027
rect 26525 8993 26559 9027
rect 7573 8925 7607 8959
rect 7757 8925 7791 8959
rect 11621 8925 11655 8959
rect 18337 8925 18371 8959
rect 10793 8857 10827 8891
rect 4629 8789 4663 8823
rect 7113 8789 7147 8823
rect 11069 8789 11103 8823
rect 17969 8789 18003 8823
rect 19717 8789 19751 8823
rect 1593 8585 1627 8619
rect 2053 8585 2087 8619
rect 5181 8585 5215 8619
rect 13553 8585 13587 8619
rect 15025 8585 15059 8619
rect 15301 8585 15335 8619
rect 18337 8585 18371 8619
rect 20545 8585 20579 8619
rect 26617 8585 26651 8619
rect 2697 8517 2731 8551
rect 7113 8517 7147 8551
rect 10333 8517 10367 8551
rect 10701 8517 10735 8551
rect 11805 8517 11839 8551
rect 17417 8517 17451 8551
rect 27353 8517 27387 8551
rect 27721 8517 27755 8551
rect 3157 8449 3191 8483
rect 7849 8449 7883 8483
rect 11437 8449 11471 8483
rect 16221 8449 16255 8483
rect 16773 8449 16807 8483
rect 16957 8449 16991 8483
rect 19165 8449 19199 8483
rect 1409 8381 1443 8415
rect 2421 8381 2455 8415
rect 2513 8381 2547 8415
rect 3801 8381 3835 8415
rect 6561 8381 6595 8415
rect 7665 8381 7699 8415
rect 8217 8381 8251 8415
rect 11161 8381 11195 8415
rect 13737 8381 13771 8415
rect 14013 8381 14047 8415
rect 26433 8381 26467 8415
rect 26985 8381 27019 8415
rect 27537 8381 27571 8415
rect 28089 8381 28123 8415
rect 3709 8313 3743 8347
rect 4046 8313 4080 8347
rect 6285 8313 6319 8347
rect 7573 8313 7607 8347
rect 8585 8313 8619 8347
rect 8769 8313 8803 8347
rect 11253 8313 11287 8347
rect 12265 8313 12299 8347
rect 15853 8313 15887 8347
rect 16681 8313 16715 8347
rect 19073 8313 19107 8347
rect 19432 8313 19466 8347
rect 7205 8245 7239 8279
rect 10793 8245 10827 8279
rect 12449 8245 12483 8279
rect 16313 8245 16347 8279
rect 1593 8041 1627 8075
rect 3893 8041 3927 8075
rect 9965 8041 9999 8075
rect 17877 8041 17911 8075
rect 18429 8041 18463 8075
rect 19165 8041 19199 8075
rect 19993 8041 20027 8075
rect 26709 8041 26743 8075
rect 10517 7973 10551 8007
rect 12909 7973 12943 8007
rect 1409 7905 1443 7939
rect 7021 7905 7055 7939
rect 7369 7905 7403 7939
rect 11253 7905 11287 7939
rect 16681 7905 16715 7939
rect 26525 7905 26559 7939
rect 7113 7837 7147 7871
rect 16773 7837 16807 7871
rect 16865 7837 16899 7871
rect 8493 7701 8527 7735
rect 10793 7701 10827 7735
rect 13461 7701 13495 7735
rect 15945 7701 15979 7735
rect 16313 7701 16347 7735
rect 2053 7497 2087 7531
rect 4721 7497 4755 7531
rect 9045 7497 9079 7531
rect 11805 7497 11839 7531
rect 14749 7497 14783 7531
rect 1593 7429 1627 7463
rect 6653 7429 6687 7463
rect 15761 7429 15795 7463
rect 19993 7429 20027 7463
rect 27353 7429 27387 7463
rect 7297 7361 7331 7395
rect 7481 7361 7515 7395
rect 8953 7361 8987 7395
rect 10149 7361 10183 7395
rect 16313 7361 16347 7395
rect 16405 7361 16439 7395
rect 19533 7361 19567 7395
rect 20637 7361 20671 7395
rect 1409 7293 1443 7327
rect 2421 7293 2455 7327
rect 3341 7293 3375 7327
rect 6285 7293 6319 7327
rect 7205 7293 7239 7327
rect 9229 7293 9263 7327
rect 9965 7293 9999 7327
rect 10425 7293 10459 7327
rect 10681 7293 10715 7327
rect 13369 7293 13403 7327
rect 16957 7293 16991 7327
rect 20361 7293 20395 7327
rect 26433 7293 26467 7327
rect 26985 7293 27019 7327
rect 3249 7225 3283 7259
rect 3608 7225 3642 7259
rect 8309 7225 8343 7259
rect 13614 7225 13648 7259
rect 15393 7225 15427 7259
rect 16221 7225 16255 7259
rect 6837 7157 6871 7191
rect 7849 7157 7883 7191
rect 9597 7157 9631 7191
rect 10057 7157 10091 7191
rect 13277 7157 13311 7191
rect 15853 7157 15887 7191
rect 19901 7157 19935 7191
rect 20453 7157 20487 7191
rect 26617 7157 26651 7191
rect 3433 6953 3467 6987
rect 4445 6953 4479 6987
rect 7021 6953 7055 6987
rect 9137 6953 9171 6987
rect 9965 6953 9999 6987
rect 15945 6953 15979 6987
rect 6285 6885 6319 6919
rect 17386 6885 17420 6919
rect 1409 6817 1443 6851
rect 10609 6817 10643 6851
rect 10701 6817 10735 6851
rect 11621 6817 11655 6851
rect 12173 6817 12207 6851
rect 19993 6817 20027 6851
rect 26525 6817 26559 6851
rect 4537 6749 4571 6783
rect 4721 6749 4755 6783
rect 6377 6749 6411 6783
rect 6561 6749 6595 6783
rect 10793 6749 10827 6783
rect 12265 6749 12299 6783
rect 12449 6749 12483 6783
rect 17141 6749 17175 6783
rect 1593 6681 1627 6715
rect 26709 6681 26743 6715
rect 4077 6613 4111 6647
rect 5917 6613 5951 6647
rect 7573 6613 7607 6647
rect 10241 6613 10275 6647
rect 11253 6613 11287 6647
rect 11805 6613 11839 6647
rect 12909 6613 12943 6647
rect 13277 6613 13311 6647
rect 16313 6613 16347 6647
rect 18521 6613 18555 6647
rect 21649 6613 21683 6647
rect 2329 6409 2363 6443
rect 3801 6409 3835 6443
rect 4629 6409 4663 6443
rect 5917 6409 5951 6443
rect 6285 6409 6319 6443
rect 8953 6409 8987 6443
rect 10149 6409 10183 6443
rect 10517 6409 10551 6443
rect 10701 6409 10735 6443
rect 12173 6409 12207 6443
rect 14841 6409 14875 6443
rect 17141 6409 17175 6443
rect 18245 6409 18279 6443
rect 27353 6409 27387 6443
rect 1593 6341 1627 6375
rect 2053 6341 2087 6375
rect 4169 6341 4203 6375
rect 19993 6341 20027 6375
rect 26617 6341 26651 6375
rect 4537 6273 4571 6307
rect 5273 6273 5307 6307
rect 7573 6273 7607 6307
rect 11253 6273 11287 6307
rect 12725 6273 12759 6307
rect 13461 6273 13495 6307
rect 18889 6273 18923 6307
rect 18981 6273 19015 6307
rect 19809 6273 19843 6307
rect 20453 6273 20487 6307
rect 20637 6273 20671 6307
rect 22109 6273 22143 6307
rect 1409 6205 1443 6239
rect 11069 6205 11103 6239
rect 11161 6205 11195 6239
rect 13185 6205 13219 6239
rect 13277 6205 13311 6239
rect 14565 6205 14599 6239
rect 17877 6205 17911 6239
rect 18797 6205 18831 6239
rect 19533 6205 19567 6239
rect 21925 6205 21959 6239
rect 26433 6205 26467 6239
rect 26985 6205 27019 6239
rect 7818 6137 7852 6171
rect 9873 6137 9907 6171
rect 20361 6137 20395 6171
rect 22017 6137 22051 6171
rect 4997 6069 5031 6103
rect 5089 6069 5123 6103
rect 7481 6069 7515 6103
rect 11897 6069 11931 6103
rect 12817 6069 12851 6103
rect 14381 6069 14415 6103
rect 16773 6069 16807 6103
rect 18429 6069 18463 6103
rect 21373 6069 21407 6103
rect 21557 6069 21591 6103
rect 4353 5865 4387 5899
rect 4997 5865 5031 5899
rect 5457 5865 5491 5899
rect 5917 5865 5951 5899
rect 7021 5865 7055 5899
rect 9505 5865 9539 5899
rect 10333 5865 10367 5899
rect 11161 5865 11195 5899
rect 11713 5865 11747 5899
rect 13277 5865 13311 5899
rect 15761 5865 15795 5899
rect 18521 5865 18555 5899
rect 19625 5865 19659 5899
rect 19717 5865 19751 5899
rect 21649 5865 21683 5899
rect 4721 5797 4755 5831
rect 6929 5797 6963 5831
rect 10701 5797 10735 5831
rect 13185 5797 13219 5831
rect 1409 5729 1443 5763
rect 5825 5729 5859 5763
rect 7389 5729 7423 5763
rect 11621 5729 11655 5763
rect 26525 5729 26559 5763
rect 6009 5661 6043 5695
rect 7481 5661 7515 5695
rect 7573 5661 7607 5695
rect 11805 5661 11839 5695
rect 12357 5661 12391 5695
rect 13461 5661 13495 5695
rect 15853 5661 15887 5695
rect 16037 5661 16071 5695
rect 19809 5661 19843 5695
rect 1593 5593 1627 5627
rect 11253 5593 11287 5627
rect 26709 5593 26743 5627
rect 6561 5525 6595 5559
rect 12817 5525 12851 5559
rect 15393 5525 15427 5559
rect 19257 5525 19291 5559
rect 2421 5321 2455 5355
rect 5181 5321 5215 5355
rect 5825 5321 5859 5355
rect 6653 5321 6687 5355
rect 6837 5321 6871 5355
rect 7849 5321 7883 5355
rect 8401 5321 8435 5355
rect 11345 5321 11379 5355
rect 11713 5321 11747 5355
rect 11989 5321 12023 5355
rect 12909 5321 12943 5355
rect 13645 5321 13679 5355
rect 15945 5321 15979 5355
rect 16589 5321 16623 5355
rect 19717 5321 19751 5355
rect 20177 5321 20211 5355
rect 27353 5321 27387 5355
rect 1593 5253 1627 5287
rect 3157 5253 3191 5287
rect 5549 5253 5583 5287
rect 13185 5253 13219 5287
rect 19441 5253 19475 5287
rect 7297 5185 7331 5219
rect 7389 5185 7423 5219
rect 9321 5185 9355 5219
rect 9965 5185 9999 5219
rect 18889 5185 18923 5219
rect 1409 5117 1443 5151
rect 2513 5117 2547 5151
rect 6285 5117 6319 5151
rect 8769 5117 8803 5151
rect 9781 5117 9815 5151
rect 9873 5117 9907 5151
rect 14565 5117 14599 5151
rect 18705 5117 18739 5151
rect 26433 5117 26467 5151
rect 26985 5117 27019 5151
rect 7205 5049 7239 5083
rect 14473 5049 14507 5083
rect 14832 5049 14866 5083
rect 17877 5049 17911 5083
rect 2053 4981 2087 5015
rect 2697 4981 2731 5015
rect 8585 4981 8619 5015
rect 9413 4981 9447 5015
rect 18337 4981 18371 5015
rect 18797 4981 18831 5015
rect 26617 4981 26651 5015
rect 6009 4777 6043 4811
rect 7113 4777 7147 4811
rect 7389 4777 7423 4811
rect 9505 4777 9539 4811
rect 15945 4777 15979 4811
rect 18797 4777 18831 4811
rect 6469 4709 6503 4743
rect 10946 4709 10980 4743
rect 16396 4709 16430 4743
rect 18337 4709 18371 4743
rect 1409 4641 1443 4675
rect 4077 4641 4111 4675
rect 6377 4641 6411 4675
rect 16129 4641 16163 4675
rect 25329 4641 25363 4675
rect 26525 4641 26559 4675
rect 4353 4573 4387 4607
rect 6561 4573 6595 4607
rect 10701 4573 10735 4607
rect 1593 4437 1627 4471
rect 12081 4437 12115 4471
rect 14565 4437 14599 4471
rect 15577 4437 15611 4471
rect 17509 4437 17543 4471
rect 25513 4437 25547 4471
rect 26709 4437 26743 4471
rect 4077 4233 4111 4267
rect 5733 4233 5767 4267
rect 10793 4233 10827 4267
rect 16221 4233 16255 4267
rect 25329 4233 25363 4267
rect 27353 4233 27387 4267
rect 2421 4165 2455 4199
rect 6377 4165 6411 4199
rect 16497 4165 16531 4199
rect 2053 4097 2087 4131
rect 6101 4097 6135 4131
rect 11069 4097 11103 4131
rect 1409 4029 1443 4063
rect 2513 4029 2547 4063
rect 4629 4029 4663 4063
rect 4721 4029 4755 4063
rect 4997 4029 5031 4063
rect 9781 4029 9815 4063
rect 10425 4029 10459 4063
rect 26433 4029 26467 4063
rect 26985 4029 27019 4063
rect 1593 3893 1627 3927
rect 2697 3893 2731 3927
rect 3157 3893 3191 3927
rect 9965 3893 9999 3927
rect 26617 3893 26651 3927
rect 1961 3689 1995 3723
rect 6745 3689 6779 3723
rect 7389 3689 7423 3723
rect 5610 3621 5644 3655
rect 12694 3621 12728 3655
rect 1409 3553 1443 3587
rect 2513 3553 2547 3587
rect 8217 3553 8251 3587
rect 9965 3553 9999 3587
rect 10221 3553 10255 3587
rect 26525 3553 26559 3587
rect 5365 3485 5399 3519
rect 12449 3485 12483 3519
rect 1593 3349 1627 3383
rect 2697 3349 2731 3383
rect 8401 3349 8435 3383
rect 11345 3349 11379 3383
rect 13829 3349 13863 3383
rect 26709 3349 26743 3383
rect 2053 3145 2087 3179
rect 2513 3145 2547 3179
rect 4537 3145 4571 3179
rect 8677 3145 8711 3179
rect 9229 3145 9263 3179
rect 9689 3145 9723 3179
rect 9965 3145 9999 3179
rect 10793 3145 10827 3179
rect 11897 3145 11931 3179
rect 12633 3145 12667 3179
rect 27353 3145 27387 3179
rect 4813 3077 4847 3111
rect 11437 3077 11471 3111
rect 4169 3009 4203 3043
rect 5825 3009 5859 3043
rect 7297 3009 7331 3043
rect 1409 2941 1443 2975
rect 3341 2941 3375 2975
rect 4629 2941 4663 2975
rect 10149 2941 10183 2975
rect 11253 2941 11287 2975
rect 13185 2941 13219 2975
rect 13737 2941 13771 2975
rect 14289 2941 14323 2975
rect 14841 2941 14875 2975
rect 19073 2941 19107 2975
rect 19625 2941 19659 2975
rect 25329 2941 25363 2975
rect 25881 2941 25915 2975
rect 26433 2941 26467 2975
rect 26985 2941 27019 2975
rect 3617 2873 3651 2907
rect 5457 2873 5491 2907
rect 7205 2873 7239 2907
rect 7542 2873 7576 2907
rect 1593 2805 1627 2839
rect 10333 2805 10367 2839
rect 13001 2805 13035 2839
rect 13369 2805 13403 2839
rect 14473 2805 14507 2839
rect 19257 2805 19291 2839
rect 25513 2805 25547 2839
rect 26617 2805 26651 2839
rect 3525 2601 3559 2635
rect 4905 2601 4939 2635
rect 9137 2601 9171 2635
rect 11161 2601 11195 2635
rect 12449 2601 12483 2635
rect 14013 2601 14047 2635
rect 17325 2601 17359 2635
rect 25881 2601 25915 2635
rect 2973 2533 3007 2567
rect 6745 2533 6779 2567
rect 7174 2533 7208 2567
rect 9505 2533 9539 2567
rect 10026 2533 10060 2567
rect 12878 2533 12912 2567
rect 1409 2465 1443 2499
rect 2145 2465 2179 2499
rect 2697 2465 2731 2499
rect 4077 2465 4111 2499
rect 12081 2465 12115 2499
rect 12633 2465 12667 2499
rect 15485 2465 15519 2499
rect 16037 2465 16071 2499
rect 16773 2465 16807 2499
rect 19073 2465 19107 2499
rect 19625 2465 19659 2499
rect 24409 2465 24443 2499
rect 24961 2465 24995 2499
rect 26893 2465 26927 2499
rect 27445 2465 27479 2499
rect 1593 2397 1627 2431
rect 4261 2397 4295 2431
rect 6377 2397 6411 2431
rect 6929 2397 6963 2431
rect 9781 2397 9815 2431
rect 19257 2329 19291 2363
rect 24593 2329 24627 2363
rect 8309 2261 8343 2295
rect 15669 2261 15703 2295
rect 16957 2261 16991 2295
rect 27077 2261 27111 2295
<< metal1 >>
rect 3142 22176 3148 22228
rect 3200 22216 3206 22228
rect 9398 22216 9404 22228
rect 3200 22188 9404 22216
rect 3200 22176 3206 22188
rect 9398 22176 9404 22188
rect 9456 22176 9462 22228
rect 2958 22108 2964 22160
rect 3016 22148 3022 22160
rect 15654 22148 15660 22160
rect 3016 22120 15660 22148
rect 3016 22108 3022 22120
rect 15654 22108 15660 22120
rect 15712 22108 15718 22160
rect 1104 21786 28888 21808
rect 1104 21734 5982 21786
rect 6034 21734 6046 21786
rect 6098 21734 6110 21786
rect 6162 21734 6174 21786
rect 6226 21734 15982 21786
rect 16034 21734 16046 21786
rect 16098 21734 16110 21786
rect 16162 21734 16174 21786
rect 16226 21734 25982 21786
rect 26034 21734 26046 21786
rect 26098 21734 26110 21786
rect 26162 21734 26174 21786
rect 26226 21734 28888 21786
rect 1104 21712 28888 21734
rect 3878 21632 3884 21684
rect 3936 21672 3942 21684
rect 6914 21672 6920 21684
rect 3936 21644 6920 21672
rect 3936 21632 3942 21644
rect 6914 21632 6920 21644
rect 6972 21632 6978 21684
rect 1104 21242 28888 21264
rect 1104 21190 10982 21242
rect 11034 21190 11046 21242
rect 11098 21190 11110 21242
rect 11162 21190 11174 21242
rect 11226 21190 20982 21242
rect 21034 21190 21046 21242
rect 21098 21190 21110 21242
rect 21162 21190 21174 21242
rect 21226 21190 28888 21242
rect 1104 21168 28888 21190
rect 3510 20816 3516 20868
rect 3568 20856 3574 20868
rect 10778 20856 10784 20868
rect 3568 20828 10784 20856
rect 3568 20816 3574 20828
rect 10778 20816 10784 20828
rect 10836 20816 10842 20868
rect 11514 20816 11520 20868
rect 11572 20856 11578 20868
rect 25774 20856 25780 20868
rect 11572 20828 25780 20856
rect 11572 20816 11578 20828
rect 25774 20816 25780 20828
rect 25832 20816 25838 20868
rect 8938 20748 8944 20800
rect 8996 20788 9002 20800
rect 25406 20788 25412 20800
rect 8996 20760 25412 20788
rect 8996 20748 9002 20760
rect 25406 20748 25412 20760
rect 25464 20748 25470 20800
rect 1104 20698 28888 20720
rect 1104 20646 5982 20698
rect 6034 20646 6046 20698
rect 6098 20646 6110 20698
rect 6162 20646 6174 20698
rect 6226 20646 15982 20698
rect 16034 20646 16046 20698
rect 16098 20646 16110 20698
rect 16162 20646 16174 20698
rect 16226 20646 25982 20698
rect 26034 20646 26046 20698
rect 26098 20646 26110 20698
rect 26162 20646 26174 20698
rect 26226 20646 28888 20698
rect 1104 20624 28888 20646
rect 4893 20587 4951 20593
rect 4893 20553 4905 20587
rect 4939 20584 4951 20587
rect 5166 20584 5172 20596
rect 4939 20556 5172 20584
rect 4939 20553 4951 20556
rect 4893 20547 4951 20553
rect 5166 20544 5172 20556
rect 5224 20544 5230 20596
rect 6730 20544 6736 20596
rect 6788 20584 6794 20596
rect 7009 20587 7067 20593
rect 7009 20584 7021 20587
rect 6788 20556 7021 20584
rect 6788 20544 6794 20556
rect 7009 20553 7021 20556
rect 7055 20553 7067 20587
rect 7009 20547 7067 20553
rect 8113 20587 8171 20593
rect 8113 20553 8125 20587
rect 8159 20584 8171 20587
rect 8202 20584 8208 20596
rect 8159 20556 8208 20584
rect 8159 20553 8171 20556
rect 8113 20547 8171 20553
rect 8202 20544 8208 20556
rect 8260 20544 8266 20596
rect 10137 20587 10195 20593
rect 10137 20553 10149 20587
rect 10183 20584 10195 20587
rect 11330 20584 11336 20596
rect 10183 20556 11336 20584
rect 10183 20553 10195 20556
rect 10137 20547 10195 20553
rect 11330 20544 11336 20556
rect 11388 20544 11394 20596
rect 18230 20584 18236 20596
rect 18191 20556 18236 20584
rect 18230 20544 18236 20556
rect 18288 20544 18294 20596
rect 16666 20516 16672 20528
rect 16627 20488 16672 20516
rect 16666 20476 16672 20488
rect 16724 20476 16730 20528
rect 25774 20516 25780 20528
rect 25735 20488 25780 20516
rect 25774 20476 25780 20488
rect 25832 20476 25838 20528
rect 20533 20451 20591 20457
rect 20533 20448 20545 20451
rect 19996 20420 20545 20448
rect 19996 20392 20024 20420
rect 20533 20417 20545 20420
rect 20579 20417 20591 20451
rect 20533 20411 20591 20417
rect 4709 20383 4767 20389
rect 4709 20349 4721 20383
rect 4755 20380 4767 20383
rect 6825 20383 6883 20389
rect 4755 20352 5396 20380
rect 4755 20349 4767 20352
rect 4709 20343 4767 20349
rect 5368 20256 5396 20352
rect 6825 20349 6837 20383
rect 6871 20349 6883 20383
rect 6825 20343 6883 20349
rect 7929 20383 7987 20389
rect 7929 20349 7941 20383
rect 7975 20380 7987 20383
rect 14093 20383 14151 20389
rect 7975 20352 8616 20380
rect 7975 20349 7987 20352
rect 7929 20343 7987 20349
rect 6840 20312 6868 20343
rect 7466 20312 7472 20324
rect 6840 20284 7472 20312
rect 7466 20272 7472 20284
rect 7524 20272 7530 20324
rect 8588 20256 8616 20352
rect 14093 20349 14105 20383
rect 14139 20380 14151 20383
rect 14737 20383 14795 20389
rect 14737 20380 14749 20383
rect 14139 20352 14749 20380
rect 14139 20349 14151 20352
rect 14093 20343 14151 20349
rect 14737 20349 14749 20352
rect 14783 20380 14795 20383
rect 15381 20383 15439 20389
rect 15381 20380 15393 20383
rect 14783 20352 15393 20380
rect 14783 20349 14795 20352
rect 14737 20343 14795 20349
rect 15381 20349 15393 20352
rect 15427 20380 15439 20383
rect 16485 20383 16543 20389
rect 15427 20352 16068 20380
rect 15427 20349 15439 20352
rect 15381 20343 15439 20349
rect 5350 20244 5356 20256
rect 5311 20216 5356 20244
rect 5350 20204 5356 20216
rect 5408 20204 5414 20256
rect 8570 20244 8576 20256
rect 8531 20216 8576 20244
rect 8570 20204 8576 20216
rect 8628 20204 8634 20256
rect 14274 20244 14280 20256
rect 14235 20216 14280 20244
rect 14274 20204 14280 20216
rect 14332 20204 14338 20256
rect 15562 20244 15568 20256
rect 15523 20216 15568 20244
rect 15562 20204 15568 20216
rect 15620 20204 15626 20256
rect 16040 20253 16068 20352
rect 16485 20349 16497 20383
rect 16531 20380 16543 20383
rect 18049 20383 18107 20389
rect 16531 20352 17080 20380
rect 16531 20349 16543 20352
rect 16485 20343 16543 20349
rect 17052 20256 17080 20352
rect 18049 20349 18061 20383
rect 18095 20380 18107 20383
rect 19978 20380 19984 20392
rect 18095 20352 18736 20380
rect 19939 20352 19984 20380
rect 18095 20349 18107 20352
rect 18049 20343 18107 20349
rect 16025 20247 16083 20253
rect 16025 20213 16037 20247
rect 16071 20244 16083 20247
rect 16390 20244 16396 20256
rect 16071 20216 16396 20244
rect 16071 20213 16083 20216
rect 16025 20207 16083 20213
rect 16390 20204 16396 20216
rect 16448 20204 16454 20256
rect 17034 20244 17040 20256
rect 16995 20216 17040 20244
rect 17034 20204 17040 20216
rect 17092 20204 17098 20256
rect 18708 20253 18736 20352
rect 19978 20340 19984 20352
rect 20036 20340 20042 20392
rect 20162 20340 20168 20392
rect 20220 20380 20226 20392
rect 20622 20380 20628 20392
rect 20220 20352 20628 20380
rect 20220 20340 20226 20352
rect 20622 20340 20628 20352
rect 20680 20340 20686 20392
rect 20806 20340 20812 20392
rect 20864 20380 20870 20392
rect 21085 20383 21143 20389
rect 21085 20380 21097 20383
rect 20864 20352 21097 20380
rect 20864 20340 20870 20352
rect 21085 20349 21097 20352
rect 21131 20380 21143 20383
rect 21637 20383 21695 20389
rect 21637 20380 21649 20383
rect 21131 20352 21649 20380
rect 21131 20349 21143 20352
rect 21085 20343 21143 20349
rect 21637 20349 21649 20352
rect 21683 20349 21695 20383
rect 24210 20380 24216 20392
rect 24171 20352 24216 20380
rect 21637 20343 21695 20349
rect 24210 20340 24216 20352
rect 24268 20380 24274 20392
rect 24765 20383 24823 20389
rect 24765 20380 24777 20383
rect 24268 20352 24777 20380
rect 24268 20340 24274 20352
rect 24765 20349 24777 20352
rect 24811 20349 24823 20383
rect 25590 20380 25596 20392
rect 25551 20352 25596 20380
rect 24765 20343 24823 20349
rect 25590 20340 25596 20352
rect 25648 20380 25654 20392
rect 26145 20383 26203 20389
rect 26145 20380 26157 20383
rect 25648 20352 26157 20380
rect 25648 20340 25654 20352
rect 26145 20349 26157 20352
rect 26191 20349 26203 20383
rect 26145 20343 26203 20349
rect 26697 20383 26755 20389
rect 26697 20349 26709 20383
rect 26743 20380 26755 20383
rect 26743 20352 27292 20380
rect 26743 20349 26755 20352
rect 26697 20343 26755 20349
rect 27264 20256 27292 20352
rect 18693 20247 18751 20253
rect 18693 20213 18705 20247
rect 18739 20244 18751 20247
rect 19150 20244 19156 20256
rect 18739 20216 19156 20244
rect 18739 20213 18751 20216
rect 18693 20207 18751 20213
rect 19150 20204 19156 20216
rect 19208 20204 19214 20256
rect 20162 20244 20168 20256
rect 20123 20216 20168 20244
rect 20162 20204 20168 20216
rect 20220 20204 20226 20256
rect 21266 20244 21272 20256
rect 21227 20216 21272 20244
rect 21266 20204 21272 20216
rect 21324 20204 21330 20256
rect 24394 20244 24400 20256
rect 24355 20216 24400 20244
rect 24394 20204 24400 20216
rect 24452 20204 24458 20256
rect 26878 20244 26884 20256
rect 26839 20216 26884 20244
rect 26878 20204 26884 20216
rect 26936 20204 26942 20256
rect 27246 20244 27252 20256
rect 27207 20216 27252 20244
rect 27246 20204 27252 20216
rect 27304 20204 27310 20256
rect 1104 20154 28888 20176
rect 1104 20102 10982 20154
rect 11034 20102 11046 20154
rect 11098 20102 11110 20154
rect 11162 20102 11174 20154
rect 11226 20102 20982 20154
rect 21034 20102 21046 20154
rect 21098 20102 21110 20154
rect 21162 20102 21174 20154
rect 21226 20102 28888 20154
rect 1104 20080 28888 20102
rect 16574 20040 16580 20052
rect 16535 20012 16580 20040
rect 16574 20000 16580 20012
rect 16632 20000 16638 20052
rect 26694 20040 26700 20052
rect 26655 20012 26700 20040
rect 26694 20000 26700 20012
rect 26752 20000 26758 20052
rect 15286 19904 15292 19916
rect 15247 19876 15292 19904
rect 15286 19864 15292 19876
rect 15344 19864 15350 19916
rect 16393 19907 16451 19913
rect 16393 19873 16405 19907
rect 16439 19904 16451 19907
rect 16482 19904 16488 19916
rect 16439 19876 16488 19904
rect 16439 19873 16451 19876
rect 16393 19867 16451 19873
rect 16482 19864 16488 19876
rect 16540 19864 16546 19916
rect 26510 19904 26516 19916
rect 26471 19876 26516 19904
rect 26510 19864 26516 19876
rect 26568 19864 26574 19916
rect 15470 19768 15476 19780
rect 15431 19740 15476 19768
rect 15470 19728 15476 19740
rect 15528 19728 15534 19780
rect 15378 19660 15384 19712
rect 15436 19700 15442 19712
rect 16574 19700 16580 19712
rect 15436 19672 16580 19700
rect 15436 19660 15442 19672
rect 16574 19660 16580 19672
rect 16632 19660 16638 19712
rect 1104 19610 28888 19632
rect 1104 19558 5982 19610
rect 6034 19558 6046 19610
rect 6098 19558 6110 19610
rect 6162 19558 6174 19610
rect 6226 19558 15982 19610
rect 16034 19558 16046 19610
rect 16098 19558 16110 19610
rect 16162 19558 16174 19610
rect 16226 19558 25982 19610
rect 26034 19558 26046 19610
rect 26098 19558 26110 19610
rect 26162 19558 26174 19610
rect 26226 19558 28888 19610
rect 1104 19536 28888 19558
rect 15286 19388 15292 19440
rect 15344 19428 15350 19440
rect 15381 19431 15439 19437
rect 15381 19428 15393 19431
rect 15344 19400 15393 19428
rect 15344 19388 15350 19400
rect 15381 19397 15393 19400
rect 15427 19428 15439 19431
rect 17034 19428 17040 19440
rect 15427 19400 17040 19428
rect 15427 19397 15439 19400
rect 15381 19391 15439 19397
rect 17034 19388 17040 19400
rect 17092 19388 17098 19440
rect 15562 19320 15568 19372
rect 15620 19360 15626 19372
rect 15746 19360 15752 19372
rect 15620 19332 15752 19360
rect 15620 19320 15626 19332
rect 15746 19320 15752 19332
rect 15804 19320 15810 19372
rect 16482 19360 16488 19372
rect 16395 19332 16488 19360
rect 16482 19320 16488 19332
rect 16540 19360 16546 19372
rect 19150 19360 19156 19372
rect 16540 19332 19156 19360
rect 16540 19320 16546 19332
rect 19150 19320 19156 19332
rect 19208 19320 19214 19372
rect 6914 19252 6920 19304
rect 6972 19252 6978 19304
rect 16942 19252 16948 19304
rect 17000 19292 17006 19304
rect 17126 19292 17132 19304
rect 17000 19264 17132 19292
rect 17000 19252 17006 19264
rect 17126 19252 17132 19264
rect 17184 19252 17190 19304
rect 6932 19224 6960 19252
rect 7190 19224 7196 19236
rect 6932 19196 7196 19224
rect 7190 19184 7196 19196
rect 7248 19184 7254 19236
rect 26510 19156 26516 19168
rect 26471 19128 26516 19156
rect 26510 19116 26516 19128
rect 26568 19116 26574 19168
rect 1104 19066 28888 19088
rect 1104 19014 10982 19066
rect 11034 19014 11046 19066
rect 11098 19014 11110 19066
rect 11162 19014 11174 19066
rect 11226 19014 20982 19066
rect 21034 19014 21046 19066
rect 21098 19014 21110 19066
rect 21162 19014 21174 19066
rect 21226 19014 28888 19066
rect 1104 18992 28888 19014
rect 1104 18522 28888 18544
rect 1104 18470 5982 18522
rect 6034 18470 6046 18522
rect 6098 18470 6110 18522
rect 6162 18470 6174 18522
rect 6226 18470 15982 18522
rect 16034 18470 16046 18522
rect 16098 18470 16110 18522
rect 16162 18470 16174 18522
rect 16226 18470 25982 18522
rect 26034 18470 26046 18522
rect 26098 18470 26110 18522
rect 26162 18470 26174 18522
rect 26226 18470 28888 18522
rect 1104 18448 28888 18470
rect 1104 17978 28888 18000
rect 1104 17926 10982 17978
rect 11034 17926 11046 17978
rect 11098 17926 11110 17978
rect 11162 17926 11174 17978
rect 11226 17926 20982 17978
rect 21034 17926 21046 17978
rect 21098 17926 21110 17978
rect 21162 17926 21174 17978
rect 21226 17926 28888 17978
rect 1104 17904 28888 17926
rect 1104 17434 28888 17456
rect 1104 17382 5982 17434
rect 6034 17382 6046 17434
rect 6098 17382 6110 17434
rect 6162 17382 6174 17434
rect 6226 17382 15982 17434
rect 16034 17382 16046 17434
rect 16098 17382 16110 17434
rect 16162 17382 16174 17434
rect 16226 17382 25982 17434
rect 26034 17382 26046 17434
rect 26098 17382 26110 17434
rect 26162 17382 26174 17434
rect 26226 17382 28888 17434
rect 1104 17360 28888 17382
rect 1104 16890 28888 16912
rect 1104 16838 10982 16890
rect 11034 16838 11046 16890
rect 11098 16838 11110 16890
rect 11162 16838 11174 16890
rect 11226 16838 20982 16890
rect 21034 16838 21046 16890
rect 21098 16838 21110 16890
rect 21162 16838 21174 16890
rect 21226 16838 28888 16890
rect 1104 16816 28888 16838
rect 1104 16346 28888 16368
rect 1104 16294 5982 16346
rect 6034 16294 6046 16346
rect 6098 16294 6110 16346
rect 6162 16294 6174 16346
rect 6226 16294 15982 16346
rect 16034 16294 16046 16346
rect 16098 16294 16110 16346
rect 16162 16294 16174 16346
rect 16226 16294 25982 16346
rect 26034 16294 26046 16346
rect 26098 16294 26110 16346
rect 26162 16294 26174 16346
rect 26226 16294 28888 16346
rect 1104 16272 28888 16294
rect 24854 16192 24860 16244
rect 24912 16232 24918 16244
rect 25866 16232 25872 16244
rect 24912 16204 25872 16232
rect 24912 16192 24918 16204
rect 25866 16192 25872 16204
rect 25924 16192 25930 16244
rect 1104 15802 28888 15824
rect 1104 15750 10982 15802
rect 11034 15750 11046 15802
rect 11098 15750 11110 15802
rect 11162 15750 11174 15802
rect 11226 15750 20982 15802
rect 21034 15750 21046 15802
rect 21098 15750 21110 15802
rect 21162 15750 21174 15802
rect 21226 15750 28888 15802
rect 1104 15728 28888 15750
rect 1104 15258 28888 15280
rect 1104 15206 5982 15258
rect 6034 15206 6046 15258
rect 6098 15206 6110 15258
rect 6162 15206 6174 15258
rect 6226 15206 15982 15258
rect 16034 15206 16046 15258
rect 16098 15206 16110 15258
rect 16162 15206 16174 15258
rect 16226 15206 25982 15258
rect 26034 15206 26046 15258
rect 26098 15206 26110 15258
rect 26162 15206 26174 15258
rect 26226 15206 28888 15258
rect 1104 15184 28888 15206
rect 24946 15104 24952 15156
rect 25004 15144 25010 15156
rect 25774 15144 25780 15156
rect 25004 15116 25780 15144
rect 25004 15104 25010 15116
rect 25774 15104 25780 15116
rect 25832 15104 25838 15156
rect 1104 14714 28888 14736
rect 1104 14662 10982 14714
rect 11034 14662 11046 14714
rect 11098 14662 11110 14714
rect 11162 14662 11174 14714
rect 11226 14662 20982 14714
rect 21034 14662 21046 14714
rect 21098 14662 21110 14714
rect 21162 14662 21174 14714
rect 21226 14662 28888 14714
rect 1104 14640 28888 14662
rect 1104 14170 28888 14192
rect 1104 14118 5982 14170
rect 6034 14118 6046 14170
rect 6098 14118 6110 14170
rect 6162 14118 6174 14170
rect 6226 14118 15982 14170
rect 16034 14118 16046 14170
rect 16098 14118 16110 14170
rect 16162 14118 16174 14170
rect 16226 14118 25982 14170
rect 26034 14118 26046 14170
rect 26098 14118 26110 14170
rect 26162 14118 26174 14170
rect 26226 14118 28888 14170
rect 1104 14096 28888 14118
rect 1104 13626 28888 13648
rect 1104 13574 10982 13626
rect 11034 13574 11046 13626
rect 11098 13574 11110 13626
rect 11162 13574 11174 13626
rect 11226 13574 20982 13626
rect 21034 13574 21046 13626
rect 21098 13574 21110 13626
rect 21162 13574 21174 13626
rect 21226 13574 28888 13626
rect 1104 13552 28888 13574
rect 8573 13379 8631 13385
rect 8573 13345 8585 13379
rect 8619 13376 8631 13379
rect 10045 13379 10103 13385
rect 10045 13376 10057 13379
rect 8619 13348 10057 13376
rect 8619 13345 8631 13348
rect 8573 13339 8631 13345
rect 10045 13345 10057 13348
rect 10091 13376 10103 13379
rect 10410 13376 10416 13388
rect 10091 13348 10416 13376
rect 10091 13345 10103 13348
rect 10045 13339 10103 13345
rect 10410 13336 10416 13348
rect 10468 13336 10474 13388
rect 11606 13385 11612 13388
rect 11600 13376 11612 13385
rect 11567 13348 11612 13376
rect 11600 13339 11612 13348
rect 11606 13336 11612 13339
rect 11664 13336 11670 13388
rect 2038 13268 2044 13320
rect 2096 13308 2102 13320
rect 2501 13311 2559 13317
rect 2501 13308 2513 13311
rect 2096 13280 2513 13308
rect 2096 13268 2102 13280
rect 2501 13277 2513 13280
rect 2547 13277 2559 13311
rect 10134 13308 10140 13320
rect 10095 13280 10140 13308
rect 2501 13271 2559 13277
rect 10134 13268 10140 13280
rect 10192 13268 10198 13320
rect 10226 13268 10232 13320
rect 10284 13308 10290 13320
rect 11330 13308 11336 13320
rect 10284 13280 10329 13308
rect 11291 13280 11336 13308
rect 10284 13268 10290 13280
rect 11330 13268 11336 13280
rect 11388 13268 11394 13320
rect 9677 13243 9735 13249
rect 9677 13209 9689 13243
rect 9723 13240 9735 13243
rect 10962 13240 10968 13252
rect 9723 13212 10968 13240
rect 9723 13209 9735 13212
rect 9677 13203 9735 13209
rect 10962 13200 10968 13212
rect 11020 13240 11026 13252
rect 11057 13243 11115 13249
rect 11057 13240 11069 13243
rect 11020 13212 11069 13240
rect 11020 13200 11026 13212
rect 11057 13209 11069 13212
rect 11103 13209 11115 13243
rect 11057 13203 11115 13209
rect 3053 13175 3111 13181
rect 3053 13141 3065 13175
rect 3099 13172 3111 13175
rect 3142 13172 3148 13184
rect 3099 13144 3148 13172
rect 3099 13141 3111 13144
rect 3053 13135 3111 13141
rect 3142 13132 3148 13144
rect 3200 13132 3206 13184
rect 9122 13172 9128 13184
rect 9083 13144 9128 13172
rect 9122 13132 9128 13144
rect 9180 13132 9186 13184
rect 9490 13132 9496 13184
rect 9548 13172 9554 13184
rect 10689 13175 10747 13181
rect 10689 13172 10701 13175
rect 9548 13144 10701 13172
rect 9548 13132 9554 13144
rect 10689 13141 10701 13144
rect 10735 13172 10747 13175
rect 11146 13172 11152 13184
rect 10735 13144 11152 13172
rect 10735 13141 10747 13144
rect 10689 13135 10747 13141
rect 11146 13132 11152 13144
rect 11204 13132 11210 13184
rect 12710 13172 12716 13184
rect 12671 13144 12716 13172
rect 12710 13132 12716 13144
rect 12768 13132 12774 13184
rect 1104 13082 28888 13104
rect 1104 13030 5982 13082
rect 6034 13030 6046 13082
rect 6098 13030 6110 13082
rect 6162 13030 6174 13082
rect 6226 13030 15982 13082
rect 16034 13030 16046 13082
rect 16098 13030 16110 13082
rect 16162 13030 16174 13082
rect 16226 13030 25982 13082
rect 26034 13030 26046 13082
rect 26098 13030 26110 13082
rect 26162 13030 26174 13082
rect 26226 13030 28888 13082
rect 1104 13008 28888 13030
rect 10410 12968 10416 12980
rect 10371 12940 10416 12968
rect 10410 12928 10416 12940
rect 10468 12928 10474 12980
rect 13814 12968 13820 12980
rect 13775 12940 13820 12968
rect 13814 12928 13820 12940
rect 13872 12968 13878 12980
rect 15105 12971 15163 12977
rect 15105 12968 15117 12971
rect 13872 12940 15117 12968
rect 13872 12928 13878 12940
rect 15105 12937 15117 12940
rect 15151 12937 15163 12971
rect 15105 12931 15163 12937
rect 10042 12900 10048 12912
rect 10003 12872 10048 12900
rect 10042 12860 10048 12872
rect 10100 12860 10106 12912
rect 11606 12900 11612 12912
rect 10980 12872 11612 12900
rect 3142 12832 3148 12844
rect 3103 12804 3148 12832
rect 3142 12792 3148 12804
rect 3200 12832 3206 12844
rect 4065 12835 4123 12841
rect 4065 12832 4077 12835
rect 3200 12804 4077 12832
rect 3200 12792 3206 12804
rect 4065 12801 4077 12804
rect 4111 12832 4123 12835
rect 4111 12804 4384 12832
rect 4111 12801 4123 12804
rect 4065 12795 4123 12801
rect 1394 12764 1400 12776
rect 1355 12736 1400 12764
rect 1394 12724 1400 12736
rect 1452 12724 1458 12776
rect 2961 12767 3019 12773
rect 2961 12764 2973 12767
rect 1964 12736 2973 12764
rect 1394 12588 1400 12640
rect 1452 12628 1458 12640
rect 1581 12631 1639 12637
rect 1581 12628 1593 12631
rect 1452 12600 1593 12628
rect 1452 12588 1458 12600
rect 1581 12597 1593 12600
rect 1627 12597 1639 12631
rect 1581 12591 1639 12597
rect 1762 12588 1768 12640
rect 1820 12628 1826 12640
rect 1964 12637 1992 12736
rect 2961 12733 2973 12736
rect 3007 12764 3019 12767
rect 3970 12764 3976 12776
rect 3007 12736 3976 12764
rect 3007 12733 3019 12736
rect 2961 12727 3019 12733
rect 3970 12724 3976 12736
rect 4028 12724 4034 12776
rect 4246 12764 4252 12776
rect 4207 12736 4252 12764
rect 4246 12724 4252 12736
rect 4304 12724 4310 12776
rect 4356 12764 4384 12804
rect 9122 12792 9128 12844
rect 9180 12832 9186 12844
rect 9585 12835 9643 12841
rect 9585 12832 9597 12835
rect 9180 12804 9597 12832
rect 9180 12792 9186 12804
rect 9585 12801 9597 12804
rect 9631 12832 9643 12835
rect 10226 12832 10232 12844
rect 9631 12804 10232 12832
rect 9631 12801 9643 12804
rect 9585 12795 9643 12801
rect 10226 12792 10232 12804
rect 10284 12832 10290 12844
rect 10502 12832 10508 12844
rect 10284 12804 10508 12832
rect 10284 12792 10290 12804
rect 10502 12792 10508 12804
rect 10560 12832 10566 12844
rect 10980 12832 11008 12872
rect 11606 12860 11612 12872
rect 11664 12860 11670 12912
rect 11146 12832 11152 12844
rect 10560 12804 11008 12832
rect 11107 12804 11152 12832
rect 10560 12792 10566 12804
rect 11146 12792 11152 12804
rect 11204 12832 11210 12844
rect 12161 12835 12219 12841
rect 12161 12832 12173 12835
rect 11204 12804 12173 12832
rect 11204 12792 11210 12804
rect 12161 12801 12173 12804
rect 12207 12832 12219 12835
rect 15120 12832 15148 12931
rect 12207 12804 12572 12832
rect 15120 12804 15424 12832
rect 12207 12801 12219 12804
rect 12161 12795 12219 12801
rect 4505 12767 4563 12773
rect 4505 12764 4517 12767
rect 4356 12736 4517 12764
rect 4505 12733 4517 12736
rect 4551 12733 4563 12767
rect 4505 12727 4563 12733
rect 8941 12767 8999 12773
rect 8941 12733 8953 12767
rect 8987 12764 8999 12767
rect 9398 12764 9404 12776
rect 8987 12736 9404 12764
rect 8987 12733 8999 12736
rect 8941 12727 8999 12733
rect 9398 12724 9404 12736
rect 9456 12724 9462 12776
rect 10962 12764 10968 12776
rect 10923 12736 10968 12764
rect 10962 12724 10968 12736
rect 11020 12724 11026 12776
rect 12434 12764 12440 12776
rect 12395 12736 12440 12764
rect 12434 12724 12440 12736
rect 12492 12724 12498 12776
rect 12544 12764 12572 12804
rect 12710 12773 12716 12776
rect 12704 12764 12716 12773
rect 12544 12736 12716 12764
rect 12704 12727 12716 12736
rect 12710 12724 12716 12727
rect 12768 12724 12774 12776
rect 15194 12764 15200 12776
rect 14752 12736 15200 12764
rect 2409 12699 2467 12705
rect 2409 12665 2421 12699
rect 2455 12696 2467 12699
rect 2866 12696 2872 12708
rect 2455 12668 2872 12696
rect 2455 12665 2467 12668
rect 2409 12659 2467 12665
rect 2866 12656 2872 12668
rect 2924 12696 2930 12708
rect 7466 12696 7472 12708
rect 2924 12668 7472 12696
rect 2924 12656 2930 12668
rect 7466 12656 7472 12668
rect 7524 12656 7530 12708
rect 10686 12696 10692 12708
rect 9048 12668 10692 12696
rect 1949 12631 2007 12637
rect 1949 12628 1961 12631
rect 1820 12600 1961 12628
rect 1820 12588 1826 12600
rect 1949 12597 1961 12600
rect 1995 12597 2007 12631
rect 2498 12628 2504 12640
rect 2459 12600 2504 12628
rect 1949 12591 2007 12597
rect 2498 12588 2504 12600
rect 2556 12588 2562 12640
rect 5534 12588 5540 12640
rect 5592 12628 5598 12640
rect 9048 12637 9076 12668
rect 10686 12656 10692 12668
rect 10744 12696 10750 12708
rect 11057 12699 11115 12705
rect 11057 12696 11069 12699
rect 10744 12668 11069 12696
rect 10744 12656 10750 12668
rect 11057 12665 11069 12668
rect 11103 12665 11115 12699
rect 11057 12659 11115 12665
rect 5629 12631 5687 12637
rect 5629 12628 5641 12631
rect 5592 12600 5641 12628
rect 5592 12588 5598 12600
rect 5629 12597 5641 12600
rect 5675 12597 5687 12631
rect 5629 12591 5687 12597
rect 9033 12631 9091 12637
rect 9033 12597 9045 12631
rect 9079 12597 9091 12631
rect 9033 12591 9091 12597
rect 9306 12588 9312 12640
rect 9364 12628 9370 12640
rect 9493 12631 9551 12637
rect 9493 12628 9505 12631
rect 9364 12600 9505 12628
rect 9364 12588 9370 12600
rect 9493 12597 9505 12600
rect 9539 12597 9551 12631
rect 9493 12591 9551 12597
rect 9674 12588 9680 12640
rect 9732 12628 9738 12640
rect 10597 12631 10655 12637
rect 10597 12628 10609 12631
rect 9732 12600 10609 12628
rect 9732 12588 9738 12600
rect 10597 12597 10609 12600
rect 10643 12597 10655 12631
rect 10597 12591 10655 12597
rect 12434 12588 12440 12640
rect 12492 12628 12498 12640
rect 13906 12628 13912 12640
rect 12492 12600 13912 12628
rect 12492 12588 12498 12600
rect 13906 12588 13912 12600
rect 13964 12628 13970 12640
rect 14752 12637 14780 12736
rect 15194 12724 15200 12736
rect 15252 12764 15258 12776
rect 15289 12767 15347 12773
rect 15289 12764 15301 12767
rect 15252 12736 15301 12764
rect 15252 12724 15258 12736
rect 15289 12733 15301 12736
rect 15335 12733 15347 12767
rect 15396 12764 15424 12804
rect 15545 12767 15603 12773
rect 15545 12764 15557 12767
rect 15396 12736 15557 12764
rect 15289 12727 15347 12733
rect 15545 12733 15557 12736
rect 15591 12733 15603 12767
rect 15545 12727 15603 12733
rect 14737 12631 14795 12637
rect 14737 12628 14749 12631
rect 13964 12600 14749 12628
rect 13964 12588 13970 12600
rect 14737 12597 14749 12600
rect 14783 12597 14795 12631
rect 16666 12628 16672 12640
rect 16627 12600 16672 12628
rect 14737 12591 14795 12597
rect 16666 12588 16672 12600
rect 16724 12588 16730 12640
rect 1104 12538 28888 12560
rect 1104 12486 10982 12538
rect 11034 12486 11046 12538
rect 11098 12486 11110 12538
rect 11162 12486 11174 12538
rect 11226 12486 20982 12538
rect 21034 12486 21046 12538
rect 21098 12486 21110 12538
rect 21162 12486 21174 12538
rect 21226 12486 28888 12538
rect 1104 12464 28888 12486
rect 1486 12384 1492 12436
rect 1544 12424 1550 12436
rect 1581 12427 1639 12433
rect 1581 12424 1593 12427
rect 1544 12396 1593 12424
rect 1544 12384 1550 12396
rect 1581 12393 1593 12396
rect 1627 12393 1639 12427
rect 1581 12387 1639 12393
rect 3050 12384 3056 12436
rect 3108 12424 3114 12436
rect 3108 12396 3740 12424
rect 3108 12384 3114 12396
rect 2038 12248 2044 12300
rect 2096 12288 2102 12300
rect 2777 12291 2835 12297
rect 2777 12288 2789 12291
rect 2096 12260 2789 12288
rect 2096 12248 2102 12260
rect 2777 12257 2789 12260
rect 2823 12257 2835 12291
rect 2777 12251 2835 12257
rect 2869 12291 2927 12297
rect 2869 12257 2881 12291
rect 2915 12288 2927 12291
rect 3712 12288 3740 12396
rect 4062 12384 4068 12436
rect 4120 12424 4126 12436
rect 4338 12424 4344 12436
rect 4120 12396 4344 12424
rect 4120 12384 4126 12396
rect 4338 12384 4344 12396
rect 4396 12384 4402 12436
rect 7929 12427 7987 12433
rect 7929 12393 7941 12427
rect 7975 12424 7987 12427
rect 8389 12427 8447 12433
rect 8389 12424 8401 12427
rect 7975 12396 8401 12424
rect 7975 12393 7987 12396
rect 7929 12387 7987 12393
rect 8389 12393 8401 12396
rect 8435 12424 8447 12427
rect 9582 12424 9588 12436
rect 8435 12396 9588 12424
rect 8435 12393 8447 12396
rect 8389 12387 8447 12393
rect 9582 12384 9588 12396
rect 9640 12384 9646 12436
rect 10686 12384 10692 12436
rect 10744 12424 10750 12436
rect 10965 12427 11023 12433
rect 10965 12424 10977 12427
rect 10744 12396 10977 12424
rect 10744 12384 10750 12396
rect 10965 12393 10977 12396
rect 11011 12393 11023 12427
rect 11330 12424 11336 12436
rect 11291 12396 11336 12424
rect 10965 12387 11023 12393
rect 11330 12384 11336 12396
rect 11388 12424 11394 12436
rect 12434 12424 12440 12436
rect 11388 12396 12440 12424
rect 11388 12384 11394 12396
rect 12434 12384 12440 12396
rect 12492 12384 12498 12436
rect 5534 12316 5540 12368
rect 5592 12356 5598 12368
rect 5690 12359 5748 12365
rect 5690 12356 5702 12359
rect 5592 12328 5702 12356
rect 5592 12316 5598 12328
rect 5690 12325 5702 12328
rect 5736 12325 5748 12359
rect 5690 12319 5748 12325
rect 16666 12316 16672 12368
rect 16724 12356 16730 12368
rect 17402 12356 17408 12368
rect 16724 12328 17408 12356
rect 16724 12316 16730 12328
rect 17402 12316 17408 12328
rect 17460 12356 17466 12368
rect 17558 12359 17616 12365
rect 17558 12356 17570 12359
rect 17460 12328 17570 12356
rect 17460 12316 17466 12328
rect 17558 12325 17570 12328
rect 17604 12325 17616 12359
rect 17558 12319 17616 12325
rect 19426 12316 19432 12368
rect 19484 12356 19490 12368
rect 20070 12356 20076 12368
rect 19484 12328 20076 12356
rect 19484 12316 19490 12328
rect 20070 12316 20076 12328
rect 20128 12316 20134 12368
rect 9674 12288 9680 12300
rect 2915 12260 3280 12288
rect 3712 12260 9680 12288
rect 2915 12257 2927 12260
rect 2869 12251 2927 12257
rect 3252 12232 3280 12260
rect 9674 12248 9680 12260
rect 9732 12248 9738 12300
rect 9858 12248 9864 12300
rect 9916 12288 9922 12300
rect 10321 12291 10379 12297
rect 10321 12288 10333 12291
rect 9916 12260 10333 12288
rect 9916 12248 9922 12260
rect 10321 12257 10333 12260
rect 10367 12257 10379 12291
rect 10321 12251 10379 12257
rect 10410 12248 10416 12300
rect 10468 12288 10474 12300
rect 10468 12260 10513 12288
rect 10468 12248 10474 12260
rect 15194 12248 15200 12300
rect 15252 12288 15258 12300
rect 17310 12288 17316 12300
rect 15252 12260 17316 12288
rect 15252 12248 15258 12260
rect 17310 12248 17316 12260
rect 17368 12248 17374 12300
rect 3050 12220 3056 12232
rect 3011 12192 3056 12220
rect 3050 12180 3056 12192
rect 3108 12180 3114 12232
rect 3234 12180 3240 12232
rect 3292 12180 3298 12232
rect 4246 12180 4252 12232
rect 4304 12220 4310 12232
rect 4341 12223 4399 12229
rect 4341 12220 4353 12223
rect 4304 12192 4353 12220
rect 4304 12180 4310 12192
rect 4341 12189 4353 12192
rect 4387 12220 4399 12223
rect 5166 12220 5172 12232
rect 4387 12192 5172 12220
rect 4387 12189 4399 12192
rect 4341 12183 4399 12189
rect 5166 12180 5172 12192
rect 5224 12220 5230 12232
rect 5445 12223 5503 12229
rect 5445 12220 5457 12223
rect 5224 12192 5457 12220
rect 5224 12180 5230 12192
rect 5445 12189 5457 12192
rect 5491 12189 5503 12223
rect 8478 12220 8484 12232
rect 8439 12192 8484 12220
rect 5445 12183 5503 12189
rect 8478 12180 8484 12192
rect 8536 12180 8542 12232
rect 8570 12180 8576 12232
rect 8628 12220 8634 12232
rect 10502 12220 10508 12232
rect 8628 12192 8673 12220
rect 10463 12192 10508 12220
rect 8628 12180 8634 12192
rect 10502 12180 10508 12192
rect 10560 12180 10566 12232
rect 15289 12223 15347 12229
rect 15289 12189 15301 12223
rect 15335 12220 15347 12223
rect 15746 12220 15752 12232
rect 15335 12192 15752 12220
rect 15335 12189 15347 12192
rect 15289 12183 15347 12189
rect 15746 12180 15752 12192
rect 15804 12180 15810 12232
rect 2225 12155 2283 12161
rect 2225 12121 2237 12155
rect 2271 12152 2283 12155
rect 2682 12152 2688 12164
rect 2271 12124 2688 12152
rect 2271 12121 2283 12124
rect 2225 12115 2283 12121
rect 2682 12112 2688 12124
rect 2740 12112 2746 12164
rect 3142 12112 3148 12164
rect 3200 12152 3206 12164
rect 3510 12152 3516 12164
rect 3200 12124 3516 12152
rect 3200 12112 3206 12124
rect 3510 12112 3516 12124
rect 3568 12112 3574 12164
rect 2406 12084 2412 12096
rect 2367 12056 2412 12084
rect 2406 12044 2412 12056
rect 2464 12044 2470 12096
rect 2498 12044 2504 12096
rect 2556 12084 2562 12096
rect 3421 12087 3479 12093
rect 3421 12084 3433 12087
rect 2556 12056 3433 12084
rect 2556 12044 2562 12056
rect 3421 12053 3433 12056
rect 3467 12053 3479 12087
rect 3786 12084 3792 12096
rect 3747 12056 3792 12084
rect 3421 12047 3479 12053
rect 3786 12044 3792 12056
rect 3844 12044 3850 12096
rect 6822 12084 6828 12096
rect 6783 12056 6828 12084
rect 6822 12044 6828 12056
rect 6880 12044 6886 12096
rect 8018 12084 8024 12096
rect 7979 12056 8024 12084
rect 8018 12044 8024 12056
rect 8076 12044 8082 12096
rect 9122 12084 9128 12096
rect 9083 12056 9128 12084
rect 9122 12044 9128 12056
rect 9180 12084 9186 12096
rect 9306 12084 9312 12096
rect 9180 12056 9312 12084
rect 9180 12044 9186 12056
rect 9306 12044 9312 12056
rect 9364 12044 9370 12096
rect 9493 12087 9551 12093
rect 9493 12053 9505 12087
rect 9539 12084 9551 12087
rect 9582 12084 9588 12096
rect 9539 12056 9588 12084
rect 9539 12053 9551 12056
rect 9493 12047 9551 12053
rect 9582 12044 9588 12056
rect 9640 12044 9646 12096
rect 9950 12084 9956 12096
rect 9911 12056 9956 12084
rect 9950 12044 9956 12056
rect 10008 12044 10014 12096
rect 14274 12084 14280 12096
rect 14235 12056 14280 12084
rect 14274 12044 14280 12056
rect 14332 12044 14338 12096
rect 18690 12084 18696 12096
rect 18651 12056 18696 12084
rect 18690 12044 18696 12056
rect 18748 12044 18754 12096
rect 1104 11994 28888 12016
rect 1104 11942 5982 11994
rect 6034 11942 6046 11994
rect 6098 11942 6110 11994
rect 6162 11942 6174 11994
rect 6226 11942 15982 11994
rect 16034 11942 16046 11994
rect 16098 11942 16110 11994
rect 16162 11942 16174 11994
rect 16226 11942 25982 11994
rect 26034 11942 26046 11994
rect 26098 11942 26110 11994
rect 26162 11942 26174 11994
rect 26226 11942 28888 11994
rect 1104 11920 28888 11942
rect 2038 11880 2044 11892
rect 1999 11852 2044 11880
rect 2038 11840 2044 11852
rect 2096 11840 2102 11892
rect 3050 11880 3056 11892
rect 2700 11852 3056 11880
rect 1673 11815 1731 11821
rect 1673 11781 1685 11815
rect 1719 11812 1731 11815
rect 2700 11812 2728 11852
rect 3050 11840 3056 11852
rect 3108 11880 3114 11892
rect 3602 11880 3608 11892
rect 3108 11852 3608 11880
rect 3108 11840 3114 11852
rect 3602 11840 3608 11852
rect 3660 11840 3666 11892
rect 8113 11883 8171 11889
rect 8113 11849 8125 11883
rect 8159 11880 8171 11883
rect 8570 11880 8576 11892
rect 8159 11852 8576 11880
rect 8159 11849 8171 11852
rect 8113 11843 8171 11849
rect 8570 11840 8576 11852
rect 8628 11840 8634 11892
rect 12342 11840 12348 11892
rect 12400 11880 12406 11892
rect 15473 11883 15531 11889
rect 15473 11880 15485 11883
rect 12400 11852 15485 11880
rect 12400 11840 12406 11852
rect 15473 11849 15485 11852
rect 15519 11880 15531 11883
rect 15565 11883 15623 11889
rect 15565 11880 15577 11883
rect 15519 11852 15577 11880
rect 15519 11849 15531 11852
rect 15473 11843 15531 11849
rect 15565 11849 15577 11852
rect 15611 11849 15623 11883
rect 15565 11843 15623 11849
rect 17310 11840 17316 11892
rect 17368 11880 17374 11892
rect 17681 11883 17739 11889
rect 17681 11880 17693 11883
rect 17368 11852 17693 11880
rect 17368 11840 17374 11852
rect 17681 11849 17693 11852
rect 17727 11849 17739 11883
rect 17681 11843 17739 11849
rect 3786 11812 3792 11824
rect 1719 11784 2728 11812
rect 3528 11784 3792 11812
rect 1719 11781 1731 11784
rect 1673 11775 1731 11781
rect 2498 11704 2504 11756
rect 2556 11744 2562 11756
rect 2593 11747 2651 11753
rect 2593 11744 2605 11747
rect 2556 11716 2605 11744
rect 2556 11704 2562 11716
rect 2593 11713 2605 11716
rect 2639 11713 2651 11747
rect 2593 11707 2651 11713
rect 2682 11704 2688 11756
rect 2740 11744 2746 11756
rect 3234 11744 3240 11756
rect 2740 11716 2785 11744
rect 3195 11716 3240 11744
rect 2740 11704 2746 11716
rect 3234 11704 3240 11716
rect 3292 11704 3298 11756
rect 2222 11636 2228 11688
rect 2280 11676 2286 11688
rect 3528 11676 3556 11784
rect 3786 11772 3792 11784
rect 3844 11772 3850 11824
rect 7377 11815 7435 11821
rect 7377 11781 7389 11815
rect 7423 11812 7435 11815
rect 8478 11812 8484 11824
rect 7423 11784 8484 11812
rect 7423 11781 7435 11784
rect 7377 11775 7435 11781
rect 8478 11772 8484 11784
rect 8536 11772 8542 11824
rect 15749 11815 15807 11821
rect 15749 11812 15761 11815
rect 14568 11784 15761 11812
rect 3605 11747 3663 11753
rect 3605 11713 3617 11747
rect 3651 11744 3663 11747
rect 4249 11747 4307 11753
rect 4249 11744 4261 11747
rect 3651 11716 4261 11744
rect 3651 11713 3663 11716
rect 3605 11707 3663 11713
rect 4249 11713 4261 11716
rect 4295 11744 4307 11747
rect 6822 11744 6828 11756
rect 4295 11716 6828 11744
rect 4295 11713 4307 11716
rect 4249 11707 4307 11713
rect 6822 11704 6828 11716
rect 6880 11704 6886 11756
rect 8662 11704 8668 11756
rect 8720 11744 8726 11756
rect 9033 11747 9091 11753
rect 9033 11744 9045 11747
rect 8720 11716 9045 11744
rect 8720 11704 8726 11716
rect 9033 11713 9045 11716
rect 9079 11744 9091 11747
rect 9490 11744 9496 11756
rect 9079 11716 9496 11744
rect 9079 11713 9091 11716
rect 9033 11707 9091 11713
rect 9490 11704 9496 11716
rect 9548 11704 9554 11756
rect 9582 11704 9588 11756
rect 9640 11744 9646 11756
rect 10502 11744 10508 11756
rect 9640 11716 10508 11744
rect 9640 11704 9646 11716
rect 10502 11704 10508 11716
rect 10560 11744 10566 11756
rect 10597 11747 10655 11753
rect 10597 11744 10609 11747
rect 10560 11716 10609 11744
rect 10560 11704 10566 11716
rect 10597 11713 10609 11716
rect 10643 11713 10655 11747
rect 10597 11707 10655 11713
rect 4157 11679 4215 11685
rect 4157 11676 4169 11679
rect 2280 11648 4169 11676
rect 2280 11636 2286 11648
rect 4157 11645 4169 11648
rect 4203 11645 4215 11679
rect 5534 11676 5540 11688
rect 5495 11648 5540 11676
rect 4157 11639 4215 11645
rect 5534 11636 5540 11648
rect 5592 11636 5598 11688
rect 8849 11679 8907 11685
rect 8849 11645 8861 11679
rect 8895 11676 8907 11679
rect 9122 11676 9128 11688
rect 8895 11648 9128 11676
rect 8895 11645 8907 11648
rect 8849 11639 8907 11645
rect 9122 11636 9128 11648
rect 9180 11676 9186 11688
rect 9950 11676 9956 11688
rect 9180 11648 9956 11676
rect 9180 11636 9186 11648
rect 9950 11636 9956 11648
rect 10008 11636 10014 11688
rect 14274 11636 14280 11688
rect 14332 11676 14338 11688
rect 14568 11685 14596 11784
rect 15749 11781 15761 11784
rect 15795 11781 15807 11815
rect 17402 11812 17408 11824
rect 17363 11784 17408 11812
rect 15749 11775 15807 11781
rect 17402 11772 17408 11784
rect 17460 11772 17466 11824
rect 14737 11747 14795 11753
rect 14737 11713 14749 11747
rect 14783 11713 14795 11747
rect 14737 11707 14795 11713
rect 15289 11747 15347 11753
rect 15289 11713 15301 11747
rect 15335 11744 15347 11747
rect 16390 11744 16396 11756
rect 15335 11716 16396 11744
rect 15335 11713 15347 11716
rect 15289 11707 15347 11713
rect 14553 11679 14611 11685
rect 14553 11676 14565 11679
rect 14332 11648 14565 11676
rect 14332 11636 14338 11648
rect 14553 11645 14565 11648
rect 14599 11645 14611 11679
rect 14553 11639 14611 11645
rect 14752 11676 14780 11707
rect 16390 11704 16396 11716
rect 16448 11704 16454 11756
rect 15194 11676 15200 11688
rect 14752 11648 15200 11676
rect 4065 11611 4123 11617
rect 4065 11608 4077 11611
rect 2148 11580 4077 11608
rect 2148 11549 2176 11580
rect 4065 11577 4077 11580
rect 4111 11608 4123 11611
rect 4709 11611 4767 11617
rect 4709 11608 4721 11611
rect 4111 11580 4721 11608
rect 4111 11577 4123 11580
rect 4065 11571 4123 11577
rect 4709 11577 4721 11580
rect 4755 11577 4767 11611
rect 4709 11571 4767 11577
rect 7745 11611 7803 11617
rect 7745 11577 7757 11611
rect 7791 11608 7803 11611
rect 8941 11611 8999 11617
rect 8941 11608 8953 11611
rect 7791 11580 8953 11608
rect 7791 11577 7803 11580
rect 7745 11571 7803 11577
rect 8941 11577 8953 11580
rect 8987 11608 8999 11611
rect 10413 11611 10471 11617
rect 8987 11580 10088 11608
rect 8987 11577 8999 11580
rect 8941 11571 8999 11577
rect 2133 11543 2191 11549
rect 2133 11509 2145 11543
rect 2179 11509 2191 11543
rect 2498 11540 2504 11552
rect 2459 11512 2504 11540
rect 2133 11503 2191 11509
rect 2498 11500 2504 11512
rect 2556 11500 2562 11552
rect 3694 11540 3700 11552
rect 3655 11512 3700 11540
rect 3694 11500 3700 11512
rect 3752 11500 3758 11552
rect 5902 11540 5908 11552
rect 5863 11512 5908 11540
rect 5902 11500 5908 11512
rect 5960 11500 5966 11552
rect 9858 11540 9864 11552
rect 9819 11512 9864 11540
rect 9858 11500 9864 11512
rect 9916 11500 9922 11552
rect 10060 11549 10088 11580
rect 10413 11577 10425 11611
rect 10459 11608 10471 11611
rect 10594 11608 10600 11620
rect 10459 11580 10600 11608
rect 10459 11577 10471 11580
rect 10413 11571 10471 11577
rect 10594 11568 10600 11580
rect 10652 11608 10658 11620
rect 11425 11611 11483 11617
rect 11425 11608 11437 11611
rect 10652 11580 11437 11608
rect 10652 11568 10658 11580
rect 11425 11577 11437 11580
rect 11471 11577 11483 11611
rect 11425 11571 11483 11577
rect 14093 11611 14151 11617
rect 14093 11577 14105 11611
rect 14139 11608 14151 11611
rect 14752 11608 14780 11648
rect 15194 11636 15200 11648
rect 15252 11636 15258 11688
rect 15746 11636 15752 11688
rect 15804 11676 15810 11688
rect 16117 11679 16175 11685
rect 16117 11676 16129 11679
rect 15804 11648 16129 11676
rect 15804 11636 15810 11648
rect 16117 11645 16129 11648
rect 16163 11645 16175 11679
rect 26418 11676 26424 11688
rect 26379 11648 26424 11676
rect 16117 11639 16175 11645
rect 26418 11636 26424 11648
rect 26476 11676 26482 11688
rect 26973 11679 27031 11685
rect 26973 11676 26985 11679
rect 26476 11648 26985 11676
rect 26476 11636 26482 11648
rect 26973 11645 26985 11648
rect 27019 11645 27031 11679
rect 26973 11639 27031 11645
rect 14139 11580 14780 11608
rect 15473 11611 15531 11617
rect 14139 11577 14151 11580
rect 14093 11571 14151 11577
rect 15473 11577 15485 11611
rect 15519 11608 15531 11611
rect 16206 11608 16212 11620
rect 15519 11580 16212 11608
rect 15519 11577 15531 11580
rect 15473 11571 15531 11577
rect 16206 11568 16212 11580
rect 16264 11568 16270 11620
rect 10045 11543 10103 11549
rect 10045 11509 10057 11543
rect 10091 11509 10103 11543
rect 10045 11503 10103 11509
rect 10505 11543 10563 11549
rect 10505 11509 10517 11543
rect 10551 11540 10563 11543
rect 10686 11540 10692 11552
rect 10551 11512 10692 11540
rect 10551 11509 10563 11512
rect 10505 11503 10563 11509
rect 10686 11500 10692 11512
rect 10744 11540 10750 11552
rect 11057 11543 11115 11549
rect 11057 11540 11069 11543
rect 10744 11512 11069 11540
rect 10744 11500 10750 11512
rect 11057 11509 11069 11512
rect 11103 11509 11115 11543
rect 14182 11540 14188 11552
rect 14143 11512 14188 11540
rect 11057 11503 11115 11509
rect 14182 11500 14188 11512
rect 14240 11500 14246 11552
rect 14642 11500 14648 11552
rect 14700 11540 14706 11552
rect 26602 11540 26608 11552
rect 14700 11512 14745 11540
rect 26563 11512 26608 11540
rect 14700 11500 14706 11512
rect 26602 11500 26608 11512
rect 26660 11500 26666 11552
rect 1104 11450 28888 11472
rect 1104 11398 10982 11450
rect 11034 11398 11046 11450
rect 11098 11398 11110 11450
rect 11162 11398 11174 11450
rect 11226 11398 20982 11450
rect 21034 11398 21046 11450
rect 21098 11398 21110 11450
rect 21162 11398 21174 11450
rect 21226 11398 28888 11450
rect 1104 11376 28888 11398
rect 2222 11336 2228 11348
rect 2183 11308 2228 11336
rect 2222 11296 2228 11308
rect 2280 11296 2286 11348
rect 2498 11296 2504 11348
rect 2556 11336 2562 11348
rect 3605 11339 3663 11345
rect 3605 11336 3617 11339
rect 2556 11308 3617 11336
rect 2556 11296 2562 11308
rect 3605 11305 3617 11308
rect 3651 11305 3663 11339
rect 8662 11336 8668 11348
rect 8623 11308 8668 11336
rect 3605 11299 3663 11305
rect 8662 11296 8668 11308
rect 8720 11296 8726 11348
rect 9033 11339 9091 11345
rect 9033 11305 9045 11339
rect 9079 11336 9091 11339
rect 9122 11336 9128 11348
rect 9079 11308 9128 11336
rect 9079 11305 9091 11308
rect 9033 11299 9091 11305
rect 9122 11296 9128 11308
rect 9180 11296 9186 11348
rect 9493 11339 9551 11345
rect 9493 11305 9505 11339
rect 9539 11336 9551 11339
rect 10410 11336 10416 11348
rect 9539 11308 10416 11336
rect 9539 11305 9551 11308
rect 9493 11299 9551 11305
rect 10410 11296 10416 11308
rect 10468 11296 10474 11348
rect 14277 11339 14335 11345
rect 14277 11305 14289 11339
rect 14323 11336 14335 11339
rect 14642 11336 14648 11348
rect 14323 11308 14648 11336
rect 14323 11305 14335 11308
rect 14277 11299 14335 11305
rect 14642 11296 14648 11308
rect 14700 11336 14706 11348
rect 15289 11339 15347 11345
rect 15289 11336 15301 11339
rect 14700 11308 15301 11336
rect 14700 11296 14706 11308
rect 15289 11305 15301 11308
rect 15335 11305 15347 11339
rect 15654 11336 15660 11348
rect 15615 11308 15660 11336
rect 15289 11299 15347 11305
rect 15654 11296 15660 11308
rect 15712 11296 15718 11348
rect 18417 11339 18475 11345
rect 18417 11305 18429 11339
rect 18463 11336 18475 11339
rect 19242 11336 19248 11348
rect 18463 11308 19248 11336
rect 18463 11305 18475 11308
rect 18417 11299 18475 11305
rect 19242 11296 19248 11308
rect 19300 11296 19306 11348
rect 26694 11336 26700 11348
rect 26655 11308 26700 11336
rect 26694 11296 26700 11308
rect 26752 11296 26758 11348
rect 6822 11228 6828 11280
rect 6880 11277 6886 11280
rect 6880 11271 6944 11277
rect 6880 11237 6898 11271
rect 6932 11237 6944 11271
rect 6880 11231 6944 11237
rect 10137 11271 10195 11277
rect 10137 11237 10149 11271
rect 10183 11268 10195 11271
rect 10502 11268 10508 11280
rect 10183 11240 10508 11268
rect 10183 11237 10195 11240
rect 10137 11231 10195 11237
rect 6880 11228 6886 11231
rect 10502 11228 10508 11240
rect 10560 11228 10566 11280
rect 17402 11228 17408 11280
rect 17460 11268 17466 11280
rect 17460 11240 18644 11268
rect 17460 11228 17466 11240
rect 1765 11203 1823 11209
rect 1765 11169 1777 11203
rect 1811 11200 1823 11203
rect 2498 11200 2504 11212
rect 1811 11172 2504 11200
rect 1811 11169 1823 11172
rect 1765 11163 1823 11169
rect 2498 11160 2504 11172
rect 2556 11200 2562 11212
rect 2593 11203 2651 11209
rect 2593 11200 2605 11203
rect 2556 11172 2605 11200
rect 2556 11160 2562 11172
rect 2593 11169 2605 11172
rect 2639 11169 2651 11203
rect 2593 11163 2651 11169
rect 10781 11203 10839 11209
rect 10781 11169 10793 11203
rect 10827 11200 10839 11203
rect 12158 11200 12164 11212
rect 10827 11172 12164 11200
rect 10827 11169 10839 11172
rect 10781 11163 10839 11169
rect 12158 11160 12164 11172
rect 12216 11160 12222 11212
rect 16298 11200 16304 11212
rect 15764 11172 16304 11200
rect 1946 11092 1952 11144
rect 2004 11132 2010 11144
rect 2685 11135 2743 11141
rect 2685 11132 2697 11135
rect 2004 11104 2697 11132
rect 2004 11092 2010 11104
rect 2685 11101 2697 11104
rect 2731 11101 2743 11135
rect 2685 11095 2743 11101
rect 2777 11135 2835 11141
rect 2777 11101 2789 11135
rect 2823 11101 2835 11135
rect 2777 11095 2835 11101
rect 2314 11024 2320 11076
rect 2372 11064 2378 11076
rect 2792 11064 2820 11095
rect 5166 11092 5172 11144
rect 5224 11132 5230 11144
rect 5902 11132 5908 11144
rect 5224 11104 5908 11132
rect 5224 11092 5230 11104
rect 5902 11092 5908 11104
rect 5960 11132 5966 11144
rect 6641 11135 6699 11141
rect 6641 11132 6653 11135
rect 5960 11104 6653 11132
rect 5960 11092 5966 11104
rect 6641 11101 6653 11104
rect 6687 11101 6699 11135
rect 6641 11095 6699 11101
rect 2372 11036 2820 11064
rect 2372 11024 2378 11036
rect 2700 11008 2728 11036
rect 2130 10996 2136 11008
rect 2091 10968 2136 10996
rect 2130 10956 2136 10968
rect 2188 10956 2194 11008
rect 2682 10956 2688 11008
rect 2740 10956 2746 11008
rect 3329 10999 3387 11005
rect 3329 10965 3341 10999
rect 3375 10996 3387 10999
rect 3602 10996 3608 11008
rect 3375 10968 3608 10996
rect 3375 10965 3387 10968
rect 3329 10959 3387 10965
rect 3602 10956 3608 10968
rect 3660 10956 3666 11008
rect 6656 10996 6684 11095
rect 10042 11092 10048 11144
rect 10100 11132 10106 11144
rect 10410 11132 10416 11144
rect 10100 11104 10416 11132
rect 10100 11092 10106 11104
rect 10410 11092 10416 11104
rect 10468 11132 10474 11144
rect 10873 11135 10931 11141
rect 10873 11132 10885 11135
rect 10468 11104 10885 11132
rect 10468 11092 10474 11104
rect 10873 11101 10885 11104
rect 10919 11101 10931 11135
rect 10873 11095 10931 11101
rect 10965 11135 11023 11141
rect 10965 11101 10977 11135
rect 11011 11101 11023 11135
rect 10965 11095 11023 11101
rect 10318 11024 10324 11076
rect 10376 11064 10382 11076
rect 10980 11064 11008 11095
rect 15470 11092 15476 11144
rect 15528 11132 15534 11144
rect 15764 11141 15792 11172
rect 16298 11160 16304 11172
rect 16356 11160 16362 11212
rect 18616 11144 18644 11240
rect 26510 11200 26516 11212
rect 26471 11172 26516 11200
rect 26510 11160 26516 11172
rect 26568 11160 26574 11212
rect 15749 11135 15807 11141
rect 15749 11132 15761 11135
rect 15528 11104 15761 11132
rect 15528 11092 15534 11104
rect 15749 11101 15761 11104
rect 15795 11101 15807 11135
rect 15749 11095 15807 11101
rect 15933 11135 15991 11141
rect 15933 11101 15945 11135
rect 15979 11132 15991 11135
rect 16390 11132 16396 11144
rect 15979 11104 16396 11132
rect 15979 11101 15991 11104
rect 15933 11095 15991 11101
rect 16390 11092 16396 11104
rect 16448 11092 16454 11144
rect 17954 11092 17960 11144
rect 18012 11132 18018 11144
rect 18509 11135 18567 11141
rect 18509 11132 18521 11135
rect 18012 11104 18521 11132
rect 18012 11092 18018 11104
rect 18509 11101 18521 11104
rect 18555 11101 18567 11135
rect 18509 11095 18567 11101
rect 11425 11067 11483 11073
rect 11425 11064 11437 11067
rect 10376 11036 11437 11064
rect 10376 11024 10382 11036
rect 11425 11033 11437 11036
rect 11471 11033 11483 11067
rect 16850 11064 16856 11076
rect 16763 11036 16856 11064
rect 11425 11027 11483 11033
rect 16850 11024 16856 11036
rect 16908 11064 16914 11076
rect 18049 11067 18107 11073
rect 18049 11064 18061 11067
rect 16908 11036 18061 11064
rect 16908 11024 16914 11036
rect 18049 11033 18061 11036
rect 18095 11033 18107 11067
rect 18524 11064 18552 11095
rect 18598 11092 18604 11144
rect 18656 11132 18662 11144
rect 18656 11104 18749 11132
rect 18656 11092 18662 11104
rect 19058 11064 19064 11076
rect 18524 11036 19064 11064
rect 18049 11027 18107 11033
rect 19058 11024 19064 11036
rect 19116 11024 19122 11076
rect 7374 10996 7380 11008
rect 6656 10968 7380 10996
rect 7374 10956 7380 10968
rect 7432 10956 7438 11008
rect 8021 10999 8079 11005
rect 8021 10965 8033 10999
rect 8067 10996 8079 10999
rect 8110 10996 8116 11008
rect 8067 10968 8116 10996
rect 8067 10965 8079 10968
rect 8021 10959 8079 10965
rect 8110 10956 8116 10968
rect 8168 10956 8174 11008
rect 16390 10996 16396 11008
rect 16351 10968 16396 10996
rect 16390 10956 16396 10968
rect 16448 10956 16454 11008
rect 1104 10906 28888 10928
rect 1104 10854 5982 10906
rect 6034 10854 6046 10906
rect 6098 10854 6110 10906
rect 6162 10854 6174 10906
rect 6226 10854 15982 10906
rect 16034 10854 16046 10906
rect 16098 10854 16110 10906
rect 16162 10854 16174 10906
rect 16226 10854 25982 10906
rect 26034 10854 26046 10906
rect 26098 10854 26110 10906
rect 26162 10854 26174 10906
rect 26226 10854 28888 10906
rect 1104 10832 28888 10854
rect 1578 10792 1584 10804
rect 1539 10764 1584 10792
rect 1578 10752 1584 10764
rect 1636 10752 1642 10804
rect 2498 10792 2504 10804
rect 2459 10764 2504 10792
rect 2498 10752 2504 10764
rect 2556 10752 2562 10804
rect 6914 10752 6920 10804
rect 6972 10792 6978 10804
rect 7009 10795 7067 10801
rect 7009 10792 7021 10795
rect 6972 10764 7021 10792
rect 6972 10752 6978 10764
rect 7009 10761 7021 10764
rect 7055 10761 7067 10795
rect 8110 10792 8116 10804
rect 8071 10764 8116 10792
rect 7009 10755 7067 10761
rect 8110 10752 8116 10764
rect 8168 10752 8174 10804
rect 9582 10792 9588 10804
rect 9543 10764 9588 10792
rect 9582 10752 9588 10764
rect 9640 10752 9646 10804
rect 10686 10792 10692 10804
rect 10647 10764 10692 10792
rect 10686 10752 10692 10764
rect 10744 10752 10750 10804
rect 12158 10792 12164 10804
rect 12119 10764 12164 10792
rect 12158 10752 12164 10764
rect 12216 10752 12222 10804
rect 15194 10752 15200 10804
rect 15252 10792 15258 10804
rect 15289 10795 15347 10801
rect 15289 10792 15301 10795
rect 15252 10764 15301 10792
rect 15252 10752 15258 10764
rect 15289 10761 15301 10764
rect 15335 10761 15347 10795
rect 15289 10755 15347 10761
rect 15654 10752 15660 10804
rect 15712 10792 15718 10804
rect 15841 10795 15899 10801
rect 15841 10792 15853 10795
rect 15712 10764 15853 10792
rect 15712 10752 15718 10764
rect 15841 10761 15853 10764
rect 15887 10761 15899 10795
rect 17862 10792 17868 10804
rect 17823 10764 17868 10792
rect 15841 10755 15899 10761
rect 17862 10752 17868 10764
rect 17920 10752 17926 10804
rect 19153 10795 19211 10801
rect 19153 10761 19165 10795
rect 19199 10792 19211 10795
rect 19242 10792 19248 10804
rect 19199 10764 19248 10792
rect 19199 10761 19211 10764
rect 19153 10755 19211 10761
rect 19242 10752 19248 10764
rect 19300 10752 19306 10804
rect 26510 10752 26516 10804
rect 26568 10792 26574 10804
rect 27341 10795 27399 10801
rect 27341 10792 27353 10795
rect 26568 10764 27353 10792
rect 26568 10752 26574 10764
rect 27341 10761 27353 10764
rect 27387 10761 27399 10795
rect 27341 10755 27399 10761
rect 2041 10727 2099 10733
rect 2041 10693 2053 10727
rect 2087 10724 2099 10727
rect 7929 10727 7987 10733
rect 7929 10724 7941 10727
rect 2087 10696 7941 10724
rect 2087 10693 2099 10696
rect 2041 10687 2099 10693
rect 7929 10693 7941 10696
rect 7975 10693 7987 10727
rect 7929 10687 7987 10693
rect 1397 10591 1455 10597
rect 1397 10557 1409 10591
rect 1443 10588 1455 10591
rect 2056 10588 2084 10687
rect 3145 10659 3203 10665
rect 3145 10625 3157 10659
rect 3191 10656 3203 10659
rect 3602 10656 3608 10668
rect 3191 10628 3608 10656
rect 3191 10625 3203 10628
rect 3145 10619 3203 10625
rect 3602 10616 3608 10628
rect 3660 10616 3666 10668
rect 4709 10659 4767 10665
rect 4709 10625 4721 10659
rect 4755 10656 4767 10659
rect 5442 10656 5448 10668
rect 4755 10628 5448 10656
rect 4755 10625 4767 10628
rect 4709 10619 4767 10625
rect 5442 10616 5448 10628
rect 5500 10616 5506 10668
rect 8128 10656 8156 10752
rect 16301 10727 16359 10733
rect 16301 10693 16313 10727
rect 16347 10724 16359 10727
rect 16390 10724 16396 10736
rect 16347 10696 16396 10724
rect 16347 10693 16359 10696
rect 16301 10687 16359 10693
rect 11241 10659 11299 10665
rect 11241 10656 11253 10659
rect 8128 10628 8340 10656
rect 1443 10560 2084 10588
rect 1443 10557 1455 10560
rect 1397 10551 1455 10557
rect 2498 10548 2504 10600
rect 2556 10588 2562 10600
rect 2556 10560 3648 10588
rect 2556 10548 2562 10560
rect 2130 10480 2136 10532
rect 2188 10520 2194 10532
rect 3620 10529 3648 10560
rect 3878 10548 3884 10600
rect 3936 10588 3942 10600
rect 3973 10591 4031 10597
rect 3973 10588 3985 10591
rect 3936 10560 3985 10588
rect 3936 10548 3942 10560
rect 3973 10557 3985 10560
rect 4019 10588 4031 10591
rect 8205 10591 8263 10597
rect 8205 10588 8217 10591
rect 4019 10560 4568 10588
rect 4019 10557 4031 10560
rect 3973 10551 4031 10557
rect 2961 10523 3019 10529
rect 2961 10520 2973 10523
rect 2188 10492 2973 10520
rect 2188 10480 2194 10492
rect 2961 10489 2973 10492
rect 3007 10489 3019 10523
rect 2961 10483 3019 10489
rect 3605 10523 3663 10529
rect 3605 10489 3617 10523
rect 3651 10520 3663 10523
rect 3651 10492 4476 10520
rect 3651 10489 3663 10492
rect 3605 10483 3663 10489
rect 4448 10464 4476 10492
rect 4540 10464 4568 10560
rect 7392 10560 8217 10588
rect 7392 10464 7420 10560
rect 8205 10557 8217 10560
rect 8251 10557 8263 10591
rect 8312 10588 8340 10628
rect 10336 10628 11253 10656
rect 10336 10600 10364 10628
rect 11241 10625 11253 10628
rect 11287 10625 11299 10659
rect 11241 10619 11299 10625
rect 13817 10659 13875 10665
rect 13817 10625 13829 10659
rect 13863 10656 13875 10659
rect 13863 10628 14044 10656
rect 13863 10625 13875 10628
rect 13817 10619 13875 10625
rect 8461 10591 8519 10597
rect 8461 10588 8473 10591
rect 8312 10560 8473 10588
rect 8205 10551 8263 10557
rect 8461 10557 8473 10560
rect 8507 10588 8519 10591
rect 10318 10588 10324 10600
rect 8507 10560 10324 10588
rect 8507 10557 8519 10560
rect 8461 10551 8519 10557
rect 10318 10548 10324 10560
rect 10376 10548 10382 10600
rect 11882 10588 11888 10600
rect 10980 10560 11888 10588
rect 7466 10480 7472 10532
rect 7524 10520 7530 10532
rect 9582 10520 9588 10532
rect 7524 10492 9588 10520
rect 7524 10480 7530 10492
rect 9582 10480 9588 10492
rect 9640 10480 9646 10532
rect 10229 10523 10287 10529
rect 10229 10489 10241 10523
rect 10275 10520 10287 10523
rect 10410 10520 10416 10532
rect 10275 10492 10416 10520
rect 10275 10489 10287 10492
rect 10229 10483 10287 10489
rect 10410 10480 10416 10492
rect 10468 10480 10474 10532
rect 2409 10455 2467 10461
rect 2409 10421 2421 10455
rect 2455 10452 2467 10455
rect 2869 10455 2927 10461
rect 2869 10452 2881 10455
rect 2455 10424 2881 10452
rect 2455 10421 2467 10424
rect 2409 10415 2467 10421
rect 2869 10421 2881 10424
rect 2915 10452 2927 10455
rect 3786 10452 3792 10464
rect 2915 10424 3792 10452
rect 2915 10421 2927 10424
rect 2869 10415 2927 10421
rect 3786 10412 3792 10424
rect 3844 10412 3850 10464
rect 4062 10452 4068 10464
rect 4023 10424 4068 10452
rect 4062 10412 4068 10424
rect 4120 10412 4126 10464
rect 4430 10452 4436 10464
rect 4391 10424 4436 10452
rect 4430 10412 4436 10424
rect 4488 10412 4494 10464
rect 4522 10412 4528 10464
rect 4580 10452 4586 10464
rect 7374 10452 7380 10464
rect 4580 10424 4625 10452
rect 7335 10424 7380 10452
rect 4580 10412 4586 10424
rect 7374 10412 7380 10424
rect 7432 10412 7438 10464
rect 7929 10455 7987 10461
rect 7929 10421 7941 10455
rect 7975 10452 7987 10455
rect 9490 10452 9496 10464
rect 7975 10424 9496 10452
rect 7975 10421 7987 10424
rect 7929 10415 7987 10421
rect 9490 10412 9496 10424
rect 9548 10412 9554 10464
rect 10502 10452 10508 10464
rect 10463 10424 10508 10452
rect 10502 10412 10508 10424
rect 10560 10452 10566 10464
rect 10980 10452 11008 10560
rect 11882 10548 11888 10560
rect 11940 10548 11946 10600
rect 13906 10588 13912 10600
rect 13867 10560 13912 10588
rect 13906 10548 13912 10560
rect 13964 10548 13970 10600
rect 14016 10588 14044 10628
rect 14176 10591 14234 10597
rect 14176 10588 14188 10591
rect 14016 10560 14188 10588
rect 14176 10557 14188 10560
rect 14222 10588 14234 10591
rect 16316 10588 16344 10687
rect 16390 10684 16396 10696
rect 16448 10724 16454 10736
rect 16448 10696 17080 10724
rect 16448 10684 16454 10696
rect 16850 10656 16856 10668
rect 16811 10628 16856 10656
rect 16850 10616 16856 10628
rect 16908 10616 16914 10668
rect 17052 10665 17080 10696
rect 17037 10659 17095 10665
rect 17037 10625 17049 10659
rect 17083 10656 17095 10659
rect 17310 10656 17316 10668
rect 17083 10628 17316 10656
rect 17083 10625 17095 10628
rect 17037 10619 17095 10625
rect 17310 10616 17316 10628
rect 17368 10616 17374 10668
rect 18598 10656 18604 10668
rect 18559 10628 18604 10656
rect 18598 10616 18604 10628
rect 18656 10656 18662 10668
rect 19429 10659 19487 10665
rect 19429 10656 19441 10659
rect 18656 10628 19441 10656
rect 18656 10616 18662 10628
rect 19429 10625 19441 10628
rect 19475 10656 19487 10659
rect 19797 10659 19855 10665
rect 19797 10656 19809 10659
rect 19475 10628 19809 10656
rect 19475 10625 19487 10628
rect 19429 10619 19487 10625
rect 19797 10625 19809 10628
rect 19843 10625 19855 10659
rect 19797 10619 19855 10625
rect 14222 10560 16344 10588
rect 14222 10557 14234 10560
rect 14176 10551 14234 10557
rect 16574 10548 16580 10600
rect 16632 10588 16638 10600
rect 17497 10591 17555 10597
rect 17497 10588 17509 10591
rect 16632 10560 17509 10588
rect 16632 10548 16638 10560
rect 17497 10557 17509 10560
rect 17543 10588 17555 10591
rect 26418 10588 26424 10600
rect 17543 10560 18552 10588
rect 26379 10560 26424 10588
rect 17543 10557 17555 10560
rect 17497 10551 17555 10557
rect 11057 10523 11115 10529
rect 11057 10489 11069 10523
rect 11103 10520 11115 10523
rect 16761 10523 16819 10529
rect 11103 10492 11836 10520
rect 11103 10489 11115 10492
rect 11057 10483 11115 10489
rect 11808 10464 11836 10492
rect 16761 10489 16773 10523
rect 16807 10520 16819 10523
rect 16807 10492 17908 10520
rect 16807 10489 16819 10492
rect 16761 10483 16819 10489
rect 17880 10464 17908 10492
rect 11149 10455 11207 10461
rect 11149 10452 11161 10455
rect 10560 10424 11161 10452
rect 10560 10412 10566 10424
rect 11149 10421 11161 10424
rect 11195 10421 11207 10455
rect 11790 10452 11796 10464
rect 11751 10424 11796 10452
rect 11149 10415 11207 10421
rect 11790 10412 11796 10424
rect 11848 10412 11854 10464
rect 16390 10452 16396 10464
rect 16351 10424 16396 10452
rect 16390 10412 16396 10424
rect 16448 10412 16454 10464
rect 17862 10412 17868 10464
rect 17920 10452 17926 10464
rect 18049 10455 18107 10461
rect 18049 10452 18061 10455
rect 17920 10424 18061 10452
rect 17920 10412 17926 10424
rect 18049 10421 18061 10424
rect 18095 10421 18107 10455
rect 18414 10452 18420 10464
rect 18375 10424 18420 10452
rect 18049 10415 18107 10421
rect 18414 10412 18420 10424
rect 18472 10412 18478 10464
rect 18524 10461 18552 10560
rect 26418 10548 26424 10560
rect 26476 10588 26482 10600
rect 26973 10591 27031 10597
rect 26973 10588 26985 10591
rect 26476 10560 26985 10588
rect 26476 10548 26482 10560
rect 26973 10557 26985 10560
rect 27019 10557 27031 10591
rect 26973 10551 27031 10557
rect 18509 10455 18567 10461
rect 18509 10421 18521 10455
rect 18555 10452 18567 10455
rect 18874 10452 18880 10464
rect 18555 10424 18880 10452
rect 18555 10421 18567 10424
rect 18509 10415 18567 10421
rect 18874 10412 18880 10424
rect 18932 10412 18938 10464
rect 26602 10452 26608 10464
rect 26563 10424 26608 10452
rect 26602 10412 26608 10424
rect 26660 10412 26666 10464
rect 1104 10362 28888 10384
rect 1104 10310 10982 10362
rect 11034 10310 11046 10362
rect 11098 10310 11110 10362
rect 11162 10310 11174 10362
rect 11226 10310 20982 10362
rect 21034 10310 21046 10362
rect 21098 10310 21110 10362
rect 21162 10310 21174 10362
rect 21226 10310 28888 10362
rect 1104 10288 28888 10310
rect 1946 10248 1952 10260
rect 1907 10220 1952 10248
rect 1946 10208 1952 10220
rect 2004 10208 2010 10260
rect 2130 10208 2136 10260
rect 2188 10248 2194 10260
rect 2409 10251 2467 10257
rect 2409 10248 2421 10251
rect 2188 10220 2421 10248
rect 2188 10208 2194 10220
rect 2409 10217 2421 10220
rect 2455 10217 2467 10251
rect 2409 10211 2467 10217
rect 2590 10208 2596 10260
rect 2648 10248 2654 10260
rect 2869 10251 2927 10257
rect 2869 10248 2881 10251
rect 2648 10220 2881 10248
rect 2648 10208 2654 10220
rect 2869 10217 2881 10220
rect 2915 10217 2927 10251
rect 2869 10211 2927 10217
rect 3326 10208 3332 10260
rect 3384 10248 3390 10260
rect 3513 10251 3571 10257
rect 3513 10248 3525 10251
rect 3384 10220 3525 10248
rect 3384 10208 3390 10220
rect 3513 10217 3525 10220
rect 3559 10248 3571 10251
rect 4062 10248 4068 10260
rect 3559 10220 4068 10248
rect 3559 10217 3571 10220
rect 3513 10211 3571 10217
rect 4062 10208 4068 10220
rect 4120 10208 4126 10260
rect 4430 10208 4436 10260
rect 4488 10248 4494 10260
rect 9582 10248 9588 10260
rect 4488 10220 9588 10248
rect 4488 10208 4494 10220
rect 9582 10208 9588 10220
rect 9640 10208 9646 10260
rect 10318 10248 10324 10260
rect 10279 10220 10324 10248
rect 10318 10208 10324 10220
rect 10376 10208 10382 10260
rect 10505 10251 10563 10257
rect 10505 10217 10517 10251
rect 10551 10248 10563 10251
rect 10594 10248 10600 10260
rect 10551 10220 10600 10248
rect 10551 10217 10563 10220
rect 10505 10211 10563 10217
rect 10594 10208 10600 10220
rect 10652 10208 10658 10260
rect 13906 10248 13912 10260
rect 13867 10220 13912 10248
rect 13906 10208 13912 10220
rect 13964 10208 13970 10260
rect 14182 10208 14188 10260
rect 14240 10248 14246 10260
rect 14369 10251 14427 10257
rect 14369 10248 14381 10251
rect 14240 10220 14381 10248
rect 14240 10208 14246 10220
rect 14369 10217 14381 10220
rect 14415 10217 14427 10251
rect 14369 10211 14427 10217
rect 16390 10208 16396 10260
rect 16448 10248 16454 10260
rect 16577 10251 16635 10257
rect 16577 10248 16589 10251
rect 16448 10220 16589 10248
rect 16448 10208 16454 10220
rect 16577 10217 16589 10220
rect 16623 10217 16635 10251
rect 16577 10211 16635 10217
rect 17221 10251 17279 10257
rect 17221 10217 17233 10251
rect 17267 10248 17279 10251
rect 17862 10248 17868 10260
rect 17267 10220 17868 10248
rect 17267 10217 17279 10220
rect 17221 10211 17279 10217
rect 17862 10208 17868 10220
rect 17920 10208 17926 10260
rect 18322 10248 18328 10260
rect 18248 10220 18328 10248
rect 2314 10180 2320 10192
rect 2275 10152 2320 10180
rect 2314 10140 2320 10152
rect 2372 10140 2378 10192
rect 2958 10140 2964 10192
rect 3016 10180 3022 10192
rect 3142 10180 3148 10192
rect 3016 10152 3148 10180
rect 3016 10140 3022 10152
rect 3142 10140 3148 10152
rect 3200 10140 3206 10192
rect 10336 10180 10364 10208
rect 10336 10152 11008 10180
rect 2777 10115 2835 10121
rect 2777 10081 2789 10115
rect 2823 10112 2835 10115
rect 2866 10112 2872 10124
rect 2823 10084 2872 10112
rect 2823 10081 2835 10084
rect 2777 10075 2835 10081
rect 2866 10072 2872 10084
rect 2924 10072 2930 10124
rect 4154 10072 4160 10124
rect 4212 10112 4218 10124
rect 5166 10112 5172 10124
rect 4212 10084 5172 10112
rect 4212 10072 4218 10084
rect 5166 10072 5172 10084
rect 5224 10072 5230 10124
rect 5442 10121 5448 10124
rect 5436 10112 5448 10121
rect 5403 10084 5448 10112
rect 5436 10075 5448 10084
rect 5442 10072 5448 10075
rect 5500 10072 5506 10124
rect 10870 10112 10876 10124
rect 10831 10084 10876 10112
rect 10870 10072 10876 10084
rect 10928 10072 10934 10124
rect 10980 10112 11008 10152
rect 10980 10084 11100 10112
rect 2958 10044 2964 10056
rect 2919 10016 2964 10044
rect 2958 10004 2964 10016
rect 3016 10044 3022 10056
rect 4249 10047 4307 10053
rect 4249 10044 4261 10047
rect 3016 10016 4261 10044
rect 3016 10004 3022 10016
rect 4249 10013 4261 10016
rect 4295 10013 4307 10047
rect 4249 10007 4307 10013
rect 9674 10004 9680 10056
rect 9732 10044 9738 10056
rect 10502 10044 10508 10056
rect 9732 10016 10508 10044
rect 9732 10004 9738 10016
rect 10502 10004 10508 10016
rect 10560 10044 10566 10056
rect 11072 10053 11100 10084
rect 13814 10072 13820 10124
rect 13872 10112 13878 10124
rect 14737 10115 14795 10121
rect 14737 10112 14749 10115
rect 13872 10084 14749 10112
rect 13872 10072 13878 10084
rect 14737 10081 14749 10084
rect 14783 10112 14795 10115
rect 15102 10112 15108 10124
rect 14783 10084 15108 10112
rect 14783 10081 14795 10084
rect 14737 10075 14795 10081
rect 15102 10072 15108 10084
rect 15160 10072 15166 10124
rect 16298 10072 16304 10124
rect 16356 10112 16362 10124
rect 16485 10115 16543 10121
rect 16485 10112 16497 10115
rect 16356 10084 16497 10112
rect 16356 10072 16362 10084
rect 16485 10081 16497 10084
rect 16531 10081 16543 10115
rect 16485 10075 16543 10081
rect 18138 10072 18144 10124
rect 18196 10112 18202 10124
rect 18248 10121 18276 10220
rect 18322 10208 18328 10220
rect 18380 10208 18386 10260
rect 18233 10115 18291 10121
rect 18233 10112 18245 10115
rect 18196 10084 18245 10112
rect 18196 10072 18202 10084
rect 18233 10081 18245 10084
rect 18279 10081 18291 10115
rect 18233 10075 18291 10081
rect 18322 10072 18328 10124
rect 18380 10112 18386 10124
rect 18380 10084 18425 10112
rect 18380 10072 18386 10084
rect 10965 10047 11023 10053
rect 10965 10044 10977 10047
rect 10560 10016 10977 10044
rect 10560 10004 10566 10016
rect 10965 10013 10977 10016
rect 11011 10013 11023 10047
rect 10965 10007 11023 10013
rect 11057 10047 11115 10053
rect 11057 10013 11069 10047
rect 11103 10044 11115 10047
rect 11238 10044 11244 10056
rect 11103 10016 11244 10044
rect 11103 10013 11115 10016
rect 11057 10007 11115 10013
rect 11238 10004 11244 10016
rect 11296 10004 11302 10056
rect 15194 10004 15200 10056
rect 15252 10044 15258 10056
rect 16669 10047 16727 10053
rect 16669 10044 16681 10047
rect 15252 10016 16681 10044
rect 15252 10004 15258 10016
rect 16669 10013 16681 10016
rect 16715 10013 16727 10047
rect 16669 10007 16727 10013
rect 18509 10047 18567 10053
rect 18509 10013 18521 10047
rect 18555 10044 18567 10047
rect 18598 10044 18604 10056
rect 18555 10016 18604 10044
rect 18555 10013 18567 10016
rect 18509 10007 18567 10013
rect 18598 10004 18604 10016
rect 18656 10004 18662 10056
rect 13906 9936 13912 9988
rect 13964 9976 13970 9988
rect 14550 9976 14556 9988
rect 13964 9948 14556 9976
rect 13964 9936 13970 9948
rect 14550 9936 14556 9948
rect 14608 9936 14614 9988
rect 18414 9976 18420 9988
rect 15304 9948 18420 9976
rect 5534 9868 5540 9920
rect 5592 9908 5598 9920
rect 6549 9911 6607 9917
rect 6549 9908 6561 9911
rect 5592 9880 6561 9908
rect 5592 9868 5598 9880
rect 6549 9877 6561 9880
rect 6595 9877 6607 9911
rect 6549 9871 6607 9877
rect 7374 9868 7380 9920
rect 7432 9908 7438 9920
rect 8205 9911 8263 9917
rect 8205 9908 8217 9911
rect 7432 9880 8217 9908
rect 7432 9868 7438 9880
rect 8205 9877 8217 9880
rect 8251 9877 8263 9911
rect 8205 9871 8263 9877
rect 13170 9868 13176 9920
rect 13228 9908 13234 9920
rect 15304 9908 15332 9948
rect 18414 9936 18420 9948
rect 18472 9976 18478 9988
rect 18877 9979 18935 9985
rect 18877 9976 18889 9979
rect 18472 9948 18889 9976
rect 18472 9936 18478 9948
rect 18877 9945 18889 9948
rect 18923 9976 18935 9979
rect 18966 9976 18972 9988
rect 18923 9948 18972 9976
rect 18923 9945 18935 9948
rect 18877 9939 18935 9945
rect 18966 9936 18972 9948
rect 19024 9936 19030 9988
rect 15470 9908 15476 9920
rect 13228 9880 15332 9908
rect 15431 9880 15476 9908
rect 13228 9868 13234 9880
rect 15470 9868 15476 9880
rect 15528 9868 15534 9920
rect 15654 9868 15660 9920
rect 15712 9908 15718 9920
rect 16117 9911 16175 9917
rect 16117 9908 16129 9911
rect 15712 9880 16129 9908
rect 15712 9868 15718 9880
rect 16117 9877 16129 9880
rect 16163 9877 16175 9911
rect 17862 9908 17868 9920
rect 17823 9880 17868 9908
rect 16117 9871 16175 9877
rect 17862 9868 17868 9880
rect 17920 9868 17926 9920
rect 1104 9818 28888 9840
rect 1104 9766 5982 9818
rect 6034 9766 6046 9818
rect 6098 9766 6110 9818
rect 6162 9766 6174 9818
rect 6226 9766 15982 9818
rect 16034 9766 16046 9818
rect 16098 9766 16110 9818
rect 16162 9766 16174 9818
rect 16226 9766 25982 9818
rect 26034 9766 26046 9818
rect 26098 9766 26110 9818
rect 26162 9766 26174 9818
rect 26226 9766 28888 9818
rect 1104 9744 28888 9766
rect 1946 9664 1952 9716
rect 2004 9704 2010 9716
rect 2866 9704 2872 9716
rect 2004 9676 2728 9704
rect 2779 9676 2872 9704
rect 2004 9664 2010 9676
rect 1578 9636 1584 9648
rect 1539 9608 1584 9636
rect 1578 9596 1584 9608
rect 1636 9596 1642 9648
rect 2501 9639 2559 9645
rect 2501 9605 2513 9639
rect 2547 9636 2559 9639
rect 2590 9636 2596 9648
rect 2547 9608 2596 9636
rect 2547 9605 2559 9608
rect 2501 9599 2559 9605
rect 2590 9596 2596 9608
rect 2648 9596 2654 9648
rect 2700 9636 2728 9676
rect 2866 9664 2872 9676
rect 2924 9704 2930 9716
rect 3878 9704 3884 9716
rect 2924 9676 3884 9704
rect 2924 9664 2930 9676
rect 3878 9664 3884 9676
rect 3936 9664 3942 9716
rect 10502 9704 10508 9716
rect 10463 9676 10508 9704
rect 10502 9664 10508 9676
rect 10560 9664 10566 9716
rect 11238 9704 11244 9716
rect 11199 9676 11244 9704
rect 11238 9664 11244 9676
rect 11296 9664 11302 9716
rect 12250 9664 12256 9716
rect 12308 9704 12314 9716
rect 13170 9704 13176 9716
rect 12308 9676 13176 9704
rect 12308 9664 12314 9676
rect 13170 9664 13176 9676
rect 13228 9664 13234 9716
rect 15654 9704 15660 9716
rect 15120 9676 15660 9704
rect 2961 9639 3019 9645
rect 2961 9636 2973 9639
rect 2700 9608 2973 9636
rect 2961 9605 2973 9608
rect 3007 9605 3019 9639
rect 4525 9639 4583 9645
rect 4525 9636 4537 9639
rect 2961 9599 3019 9605
rect 3436 9608 4537 9636
rect 3436 9580 3464 9608
rect 4525 9605 4537 9608
rect 4571 9605 4583 9639
rect 15120 9636 15148 9676
rect 15654 9664 15660 9676
rect 15712 9664 15718 9716
rect 16390 9664 16396 9716
rect 16448 9704 16454 9716
rect 16485 9707 16543 9713
rect 16485 9704 16497 9707
rect 16448 9676 16497 9704
rect 16448 9664 16454 9676
rect 16485 9673 16497 9676
rect 16531 9673 16543 9707
rect 16485 9667 16543 9673
rect 16942 9664 16948 9716
rect 17000 9704 17006 9716
rect 17218 9704 17224 9716
rect 17000 9676 17224 9704
rect 17000 9664 17006 9676
rect 17218 9664 17224 9676
rect 17276 9664 17282 9716
rect 4525 9599 4583 9605
rect 14844 9608 15148 9636
rect 15841 9639 15899 9645
rect 2041 9571 2099 9577
rect 2041 9537 2053 9571
rect 2087 9568 2099 9571
rect 2682 9568 2688 9580
rect 2087 9540 2688 9568
rect 2087 9537 2099 9540
rect 2041 9531 2099 9537
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9500 1455 9503
rect 2056 9500 2084 9531
rect 2682 9528 2688 9540
rect 2740 9528 2746 9580
rect 3418 9568 3424 9580
rect 3331 9540 3424 9568
rect 3418 9528 3424 9540
rect 3476 9528 3482 9580
rect 3602 9568 3608 9580
rect 3563 9540 3608 9568
rect 3602 9528 3608 9540
rect 3660 9528 3666 9580
rect 5077 9571 5135 9577
rect 5077 9568 5089 9571
rect 3988 9540 5089 9568
rect 3326 9500 3332 9512
rect 1443 9472 2084 9500
rect 3287 9472 3332 9500
rect 1443 9469 1455 9472
rect 1397 9463 1455 9469
rect 3326 9460 3332 9472
rect 3384 9460 3390 9512
rect 2958 9392 2964 9444
rect 3016 9432 3022 9444
rect 3988 9441 4016 9540
rect 5077 9537 5089 9540
rect 5123 9568 5135 9571
rect 5442 9568 5448 9580
rect 5123 9540 5448 9568
rect 5123 9537 5135 9540
rect 5077 9531 5135 9537
rect 5442 9528 5448 9540
rect 5500 9568 5506 9580
rect 5537 9571 5595 9577
rect 5537 9568 5549 9571
rect 5500 9540 5549 9568
rect 5500 9528 5506 9540
rect 5537 9537 5549 9540
rect 5583 9537 5595 9571
rect 5537 9531 5595 9537
rect 14458 9528 14464 9580
rect 14516 9568 14522 9580
rect 14844 9577 14872 9608
rect 15841 9605 15853 9639
rect 15887 9636 15899 9639
rect 16298 9636 16304 9648
rect 15887 9608 16304 9636
rect 15887 9605 15899 9608
rect 15841 9599 15899 9605
rect 16298 9596 16304 9608
rect 16356 9636 16362 9648
rect 18049 9639 18107 9645
rect 18049 9636 18061 9639
rect 16356 9608 18061 9636
rect 16356 9596 16362 9608
rect 18049 9605 18061 9608
rect 18095 9605 18107 9639
rect 18049 9599 18107 9605
rect 14829 9571 14887 9577
rect 14829 9568 14841 9571
rect 14516 9540 14841 9568
rect 14516 9528 14522 9540
rect 14829 9537 14841 9540
rect 14875 9537 14887 9571
rect 14829 9531 14887 9537
rect 14921 9571 14979 9577
rect 14921 9537 14933 9571
rect 14967 9537 14979 9571
rect 14921 9531 14979 9537
rect 4614 9460 4620 9512
rect 4672 9500 4678 9512
rect 4893 9503 4951 9509
rect 4893 9500 4905 9503
rect 4672 9472 4905 9500
rect 4672 9460 4678 9472
rect 4893 9469 4905 9472
rect 4939 9469 4951 9503
rect 4893 9463 4951 9469
rect 7745 9503 7803 9509
rect 7745 9469 7757 9503
rect 7791 9500 7803 9503
rect 8021 9503 8079 9509
rect 8021 9500 8033 9503
rect 7791 9472 8033 9500
rect 7791 9469 7803 9472
rect 7745 9463 7803 9469
rect 8021 9469 8033 9472
rect 8067 9500 8079 9503
rect 8294 9500 8300 9512
rect 8067 9472 8300 9500
rect 8067 9469 8079 9472
rect 8021 9463 8079 9469
rect 8294 9460 8300 9472
rect 8352 9460 8358 9512
rect 14182 9460 14188 9512
rect 14240 9500 14246 9512
rect 14737 9503 14795 9509
rect 14737 9500 14749 9503
rect 14240 9472 14749 9500
rect 14240 9460 14246 9472
rect 14737 9469 14749 9472
rect 14783 9469 14795 9503
rect 14737 9463 14795 9469
rect 14936 9444 14964 9531
rect 15102 9528 15108 9580
rect 15160 9568 15166 9580
rect 15381 9571 15439 9577
rect 15381 9568 15393 9571
rect 15160 9540 15393 9568
rect 15160 9528 15166 9540
rect 15381 9537 15393 9540
rect 15427 9537 15439 9571
rect 17402 9568 17408 9580
rect 17363 9540 17408 9568
rect 15381 9531 15439 9537
rect 17402 9528 17408 9540
rect 17460 9528 17466 9580
rect 17954 9528 17960 9580
rect 18012 9568 18018 9580
rect 18509 9571 18567 9577
rect 18509 9568 18521 9571
rect 18012 9540 18521 9568
rect 18012 9528 18018 9540
rect 18509 9537 18521 9540
rect 18555 9537 18567 9571
rect 18690 9568 18696 9580
rect 18603 9540 18696 9568
rect 18509 9531 18567 9537
rect 15194 9460 15200 9512
rect 15252 9500 15258 9512
rect 16117 9503 16175 9509
rect 16117 9500 16129 9503
rect 15252 9472 16129 9500
rect 15252 9460 15258 9472
rect 16117 9469 16129 9472
rect 16163 9469 16175 9503
rect 16117 9463 16175 9469
rect 17129 9503 17187 9509
rect 17129 9469 17141 9503
rect 17175 9500 17187 9503
rect 17310 9500 17316 9512
rect 17175 9472 17316 9500
rect 17175 9469 17187 9472
rect 17129 9463 17187 9469
rect 17310 9460 17316 9472
rect 17368 9460 17374 9512
rect 18524 9500 18552 9531
rect 18690 9528 18696 9540
rect 18748 9568 18754 9580
rect 19061 9571 19119 9577
rect 19061 9568 19073 9571
rect 18748 9540 19073 9568
rect 18748 9528 18754 9540
rect 19061 9537 19073 9540
rect 19107 9537 19119 9571
rect 19061 9531 19119 9537
rect 19429 9503 19487 9509
rect 19429 9500 19441 9503
rect 18524 9472 19441 9500
rect 19429 9469 19441 9472
rect 19475 9469 19487 9503
rect 19429 9463 19487 9469
rect 3973 9435 4031 9441
rect 3973 9432 3985 9435
rect 3016 9404 3985 9432
rect 3016 9392 3022 9404
rect 3973 9401 3985 9404
rect 4019 9401 4031 9435
rect 3973 9395 4031 9401
rect 14277 9435 14335 9441
rect 14277 9401 14289 9435
rect 14323 9432 14335 9435
rect 14918 9432 14924 9444
rect 14323 9404 14924 9432
rect 14323 9401 14335 9404
rect 14277 9395 14335 9401
rect 14918 9392 14924 9404
rect 14976 9392 14982 9444
rect 17770 9432 17776 9444
rect 17731 9404 17776 9432
rect 17770 9392 17776 9404
rect 17828 9432 17834 9444
rect 18417 9435 18475 9441
rect 18417 9432 18429 9435
rect 17828 9404 18429 9432
rect 17828 9392 17834 9404
rect 18417 9401 18429 9404
rect 18463 9401 18475 9435
rect 18417 9395 18475 9401
rect 4062 9324 4068 9376
rect 4120 9364 4126 9376
rect 4433 9367 4491 9373
rect 4433 9364 4445 9367
rect 4120 9336 4445 9364
rect 4120 9324 4126 9336
rect 4433 9333 4445 9336
rect 4479 9364 4491 9367
rect 4982 9364 4988 9376
rect 4479 9336 4988 9364
rect 4479 9333 4491 9336
rect 4433 9327 4491 9333
rect 4982 9324 4988 9336
rect 5040 9324 5046 9376
rect 5997 9367 6055 9373
rect 5997 9333 6009 9367
rect 6043 9364 6055 9367
rect 7374 9364 7380 9376
rect 6043 9336 7380 9364
rect 6043 9333 6055 9336
rect 5997 9327 6055 9333
rect 7374 9324 7380 9336
rect 7432 9364 7438 9376
rect 7561 9367 7619 9373
rect 7561 9364 7573 9367
rect 7432 9336 7573 9364
rect 7432 9324 7438 9336
rect 7561 9333 7573 9336
rect 7607 9333 7619 9367
rect 7561 9327 7619 9333
rect 10870 9324 10876 9376
rect 10928 9364 10934 9376
rect 10965 9367 11023 9373
rect 10965 9364 10977 9367
rect 10928 9336 10977 9364
rect 10928 9324 10934 9336
rect 10965 9333 10977 9336
rect 11011 9364 11023 9367
rect 11330 9364 11336 9376
rect 11011 9336 11336 9364
rect 11011 9333 11023 9336
rect 10965 9327 11023 9333
rect 11330 9324 11336 9336
rect 11388 9324 11394 9376
rect 14366 9364 14372 9376
rect 14327 9336 14372 9364
rect 14366 9324 14372 9336
rect 14424 9324 14430 9376
rect 1104 9274 28888 9296
rect 1104 9222 10982 9274
rect 11034 9222 11046 9274
rect 11098 9222 11110 9274
rect 11162 9222 11174 9274
rect 11226 9222 20982 9274
rect 21034 9222 21046 9274
rect 21098 9222 21110 9274
rect 21162 9222 21174 9274
rect 21226 9222 28888 9274
rect 1104 9200 28888 9222
rect 1486 9120 1492 9172
rect 1544 9160 1550 9172
rect 1581 9163 1639 9169
rect 1581 9160 1593 9163
rect 1544 9132 1593 9160
rect 1544 9120 1550 9132
rect 1581 9129 1593 9132
rect 1627 9129 1639 9163
rect 1581 9123 1639 9129
rect 2501 9163 2559 9169
rect 2501 9129 2513 9163
rect 2547 9160 2559 9163
rect 2958 9160 2964 9172
rect 2547 9132 2964 9160
rect 2547 9129 2559 9132
rect 2501 9123 2559 9129
rect 2958 9120 2964 9132
rect 3016 9120 3022 9172
rect 3418 9160 3424 9172
rect 3379 9132 3424 9160
rect 3418 9120 3424 9132
rect 3476 9120 3482 9172
rect 14458 9160 14464 9172
rect 14419 9132 14464 9160
rect 14458 9120 14464 9132
rect 14516 9120 14522 9172
rect 16666 9160 16672 9172
rect 16627 9132 16672 9160
rect 16666 9120 16672 9132
rect 16724 9120 16730 9172
rect 26694 9160 26700 9172
rect 26655 9132 26700 9160
rect 26694 9120 26700 9132
rect 26752 9120 26758 9172
rect 3053 9095 3111 9101
rect 3053 9061 3065 9095
rect 3099 9092 3111 9095
rect 3602 9092 3608 9104
rect 3099 9064 3608 9092
rect 3099 9061 3111 9064
rect 3053 9055 3111 9061
rect 3602 9052 3608 9064
rect 3660 9052 3666 9104
rect 15194 9052 15200 9104
rect 15252 9092 15258 9104
rect 15534 9095 15592 9101
rect 15534 9092 15546 9095
rect 15252 9064 15546 9092
rect 15252 9052 15258 9064
rect 15534 9061 15546 9064
rect 15580 9061 15592 9095
rect 16684 9092 16712 9120
rect 18322 9092 18328 9104
rect 16684 9064 18328 9092
rect 15534 9055 15592 9061
rect 18322 9052 18328 9064
rect 18380 9092 18386 9104
rect 18570 9095 18628 9101
rect 18570 9092 18582 9095
rect 18380 9064 18582 9092
rect 18380 9052 18386 9064
rect 18570 9061 18582 9064
rect 18616 9061 18628 9095
rect 18570 9055 18628 9061
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 9024 1455 9027
rect 2406 9024 2412 9036
rect 1443 8996 2412 9024
rect 1443 8993 1455 8996
rect 1397 8987 1455 8993
rect 2406 8984 2412 8996
rect 2464 8984 2470 9036
rect 7190 8984 7196 9036
rect 7248 9024 7254 9036
rect 7469 9027 7527 9033
rect 7469 9024 7481 9027
rect 7248 8996 7481 9024
rect 7248 8984 7254 8996
rect 7469 8993 7481 8996
rect 7515 8993 7527 9027
rect 7469 8987 7527 8993
rect 10318 8984 10324 9036
rect 10376 9024 10382 9036
rect 11422 9024 11428 9036
rect 10376 8996 11428 9024
rect 10376 8984 10382 8996
rect 11422 8984 11428 8996
rect 11480 8984 11486 9036
rect 11514 8984 11520 9036
rect 11572 9024 11578 9036
rect 11572 8996 11617 9024
rect 11572 8984 11578 8996
rect 14550 8984 14556 9036
rect 14608 9024 14614 9036
rect 15010 9024 15016 9036
rect 14608 8996 15016 9024
rect 14608 8984 14614 8996
rect 15010 8984 15016 8996
rect 15068 9024 15074 9036
rect 15289 9027 15347 9033
rect 15289 9024 15301 9027
rect 15068 8996 15301 9024
rect 15068 8984 15074 8996
rect 15289 8993 15301 8996
rect 15335 9024 15347 9027
rect 18414 9024 18420 9036
rect 15335 8996 18420 9024
rect 15335 8993 15347 8996
rect 15289 8987 15347 8993
rect 6546 8916 6552 8968
rect 6604 8956 6610 8968
rect 7558 8956 7564 8968
rect 6604 8928 7564 8956
rect 6604 8916 6610 8928
rect 7558 8916 7564 8928
rect 7616 8916 7622 8968
rect 7745 8959 7803 8965
rect 7745 8925 7757 8959
rect 7791 8956 7803 8959
rect 7834 8956 7840 8968
rect 7791 8928 7840 8956
rect 7791 8925 7803 8928
rect 7745 8919 7803 8925
rect 7834 8916 7840 8928
rect 7892 8916 7898 8968
rect 11606 8956 11612 8968
rect 11567 8928 11612 8956
rect 11606 8916 11612 8928
rect 11664 8916 11670 8968
rect 18340 8965 18368 8996
rect 18414 8984 18420 8996
rect 18472 8984 18478 9036
rect 26510 9024 26516 9036
rect 26471 8996 26516 9024
rect 26510 8984 26516 8996
rect 26568 8984 26574 9036
rect 18325 8959 18383 8965
rect 18325 8925 18337 8959
rect 18371 8925 18383 8959
rect 18325 8919 18383 8925
rect 10502 8848 10508 8900
rect 10560 8888 10566 8900
rect 10781 8891 10839 8897
rect 10781 8888 10793 8891
rect 10560 8860 10793 8888
rect 10560 8848 10566 8860
rect 10781 8857 10793 8860
rect 10827 8888 10839 8891
rect 11624 8888 11652 8916
rect 10827 8860 11652 8888
rect 10827 8857 10839 8860
rect 10781 8851 10839 8857
rect 4614 8820 4620 8832
rect 4575 8792 4620 8820
rect 4614 8780 4620 8792
rect 4672 8780 4678 8832
rect 7098 8820 7104 8832
rect 7059 8792 7104 8820
rect 7098 8780 7104 8792
rect 7156 8780 7162 8832
rect 10870 8780 10876 8832
rect 10928 8820 10934 8832
rect 11057 8823 11115 8829
rect 11057 8820 11069 8823
rect 10928 8792 11069 8820
rect 10928 8780 10934 8792
rect 11057 8789 11069 8792
rect 11103 8789 11115 8823
rect 11057 8783 11115 8789
rect 17957 8823 18015 8829
rect 17957 8789 17969 8823
rect 18003 8820 18015 8823
rect 18138 8820 18144 8832
rect 18003 8792 18144 8820
rect 18003 8789 18015 8792
rect 17957 8783 18015 8789
rect 18138 8780 18144 8792
rect 18196 8820 18202 8832
rect 18598 8820 18604 8832
rect 18196 8792 18604 8820
rect 18196 8780 18202 8792
rect 18598 8780 18604 8792
rect 18656 8780 18662 8832
rect 19518 8780 19524 8832
rect 19576 8820 19582 8832
rect 19705 8823 19763 8829
rect 19705 8820 19717 8823
rect 19576 8792 19717 8820
rect 19576 8780 19582 8792
rect 19705 8789 19717 8792
rect 19751 8789 19763 8823
rect 19705 8783 19763 8789
rect 1104 8730 28888 8752
rect 1104 8678 5982 8730
rect 6034 8678 6046 8730
rect 6098 8678 6110 8730
rect 6162 8678 6174 8730
rect 6226 8678 15982 8730
rect 16034 8678 16046 8730
rect 16098 8678 16110 8730
rect 16162 8678 16174 8730
rect 16226 8678 25982 8730
rect 26034 8678 26046 8730
rect 26098 8678 26110 8730
rect 26162 8678 26174 8730
rect 26226 8678 28888 8730
rect 1104 8656 28888 8678
rect 1394 8576 1400 8628
rect 1452 8616 1458 8628
rect 1581 8619 1639 8625
rect 1581 8616 1593 8619
rect 1452 8588 1593 8616
rect 1452 8576 1458 8588
rect 1581 8585 1593 8588
rect 1627 8585 1639 8619
rect 2038 8616 2044 8628
rect 1999 8588 2044 8616
rect 1581 8579 1639 8585
rect 2038 8576 2044 8588
rect 2096 8576 2102 8628
rect 5169 8619 5227 8625
rect 5169 8585 5181 8619
rect 5215 8616 5227 8619
rect 5442 8616 5448 8628
rect 5215 8588 5448 8616
rect 5215 8585 5227 8588
rect 5169 8579 5227 8585
rect 5442 8576 5448 8588
rect 5500 8576 5506 8628
rect 13541 8619 13599 8625
rect 13541 8585 13553 8619
rect 13587 8616 13599 8619
rect 13722 8616 13728 8628
rect 13587 8588 13728 8616
rect 13587 8585 13599 8588
rect 13541 8579 13599 8585
rect 13722 8576 13728 8588
rect 13780 8576 13786 8628
rect 15010 8616 15016 8628
rect 14971 8588 15016 8616
rect 15010 8576 15016 8588
rect 15068 8576 15074 8628
rect 15194 8576 15200 8628
rect 15252 8616 15258 8628
rect 15289 8619 15347 8625
rect 15289 8616 15301 8619
rect 15252 8588 15301 8616
rect 15252 8576 15258 8588
rect 15289 8585 15301 8588
rect 15335 8585 15347 8619
rect 18322 8616 18328 8628
rect 18283 8588 18328 8616
rect 15289 8579 15347 8585
rect 18322 8576 18328 8588
rect 18380 8576 18386 8628
rect 20533 8619 20591 8625
rect 20533 8616 20545 8619
rect 18432 8588 20545 8616
rect 2682 8548 2688 8560
rect 2643 8520 2688 8548
rect 2682 8508 2688 8520
rect 2740 8508 2746 8560
rect 7101 8551 7159 8557
rect 7101 8517 7113 8551
rect 7147 8548 7159 8551
rect 7190 8548 7196 8560
rect 7147 8520 7196 8548
rect 7147 8517 7159 8520
rect 7101 8511 7159 8517
rect 7190 8508 7196 8520
rect 7248 8508 7254 8560
rect 10318 8548 10324 8560
rect 10279 8520 10324 8548
rect 10318 8508 10324 8520
rect 10376 8508 10382 8560
rect 10689 8551 10747 8557
rect 10689 8517 10701 8551
rect 10735 8548 10747 8551
rect 10778 8548 10784 8560
rect 10735 8520 10784 8548
rect 10735 8517 10747 8520
rect 10689 8511 10747 8517
rect 10778 8508 10784 8520
rect 10836 8548 10842 8560
rect 10836 8520 11192 8548
rect 10836 8508 10842 8520
rect 3142 8480 3148 8492
rect 2516 8452 3148 8480
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8412 1455 8415
rect 2038 8412 2044 8424
rect 1443 8384 2044 8412
rect 1443 8381 1455 8384
rect 1397 8375 1455 8381
rect 2038 8372 2044 8384
rect 2096 8372 2102 8424
rect 2406 8412 2412 8424
rect 2367 8384 2412 8412
rect 2406 8372 2412 8384
rect 2464 8372 2470 8424
rect 2516 8421 2544 8452
rect 3142 8440 3148 8452
rect 3200 8440 3206 8492
rect 7834 8480 7840 8492
rect 7795 8452 7840 8480
rect 7834 8440 7840 8452
rect 7892 8440 7898 8492
rect 2501 8415 2559 8421
rect 2501 8381 2513 8415
rect 2547 8381 2559 8415
rect 2501 8375 2559 8381
rect 3789 8415 3847 8421
rect 3789 8381 3801 8415
rect 3835 8412 3847 8415
rect 3878 8412 3884 8424
rect 3835 8384 3884 8412
rect 3835 8381 3847 8384
rect 3789 8375 3847 8381
rect 3878 8372 3884 8384
rect 3936 8372 3942 8424
rect 6546 8412 6552 8424
rect 6507 8384 6552 8412
rect 6546 8372 6552 8384
rect 6604 8372 6610 8424
rect 7650 8412 7656 8424
rect 7611 8384 7656 8412
rect 7650 8372 7656 8384
rect 7708 8412 7714 8424
rect 8205 8415 8263 8421
rect 8205 8412 8217 8415
rect 7708 8384 8217 8412
rect 7708 8372 7714 8384
rect 8205 8381 8217 8384
rect 8251 8412 8263 8415
rect 8938 8412 8944 8424
rect 8251 8384 8944 8412
rect 8251 8381 8263 8384
rect 8205 8375 8263 8381
rect 8938 8372 8944 8384
rect 8996 8372 9002 8424
rect 11164 8421 11192 8520
rect 11514 8508 11520 8560
rect 11572 8548 11578 8560
rect 11793 8551 11851 8557
rect 11793 8548 11805 8551
rect 11572 8520 11805 8548
rect 11572 8508 11578 8520
rect 11793 8517 11805 8520
rect 11839 8517 11851 8551
rect 17405 8551 17463 8557
rect 17405 8548 17417 8551
rect 11793 8511 11851 8517
rect 16960 8520 17417 8548
rect 11425 8483 11483 8489
rect 11425 8449 11437 8483
rect 11471 8480 11483 8483
rect 11606 8480 11612 8492
rect 11471 8452 11612 8480
rect 11471 8449 11483 8452
rect 11425 8443 11483 8449
rect 11606 8440 11612 8452
rect 11664 8480 11670 8492
rect 11664 8452 12296 8480
rect 11664 8440 11670 8452
rect 11149 8415 11207 8421
rect 11149 8381 11161 8415
rect 11195 8381 11207 8415
rect 11149 8375 11207 8381
rect 12268 8356 12296 8452
rect 15470 8440 15476 8492
rect 15528 8480 15534 8492
rect 16209 8483 16267 8489
rect 16209 8480 16221 8483
rect 15528 8452 16221 8480
rect 15528 8440 15534 8452
rect 16209 8449 16221 8452
rect 16255 8480 16267 8483
rect 16758 8480 16764 8492
rect 16255 8452 16764 8480
rect 16255 8449 16267 8452
rect 16209 8443 16267 8449
rect 16758 8440 16764 8452
rect 16816 8440 16822 8492
rect 16850 8440 16856 8492
rect 16908 8480 16914 8492
rect 16960 8489 16988 8520
rect 17405 8517 17417 8520
rect 17451 8548 17463 8551
rect 18432 8548 18460 8588
rect 20533 8585 20545 8588
rect 20579 8585 20591 8619
rect 26602 8616 26608 8628
rect 26563 8588 26608 8616
rect 20533 8579 20591 8585
rect 26602 8576 26608 8588
rect 26660 8576 26666 8628
rect 17451 8520 18460 8548
rect 17451 8517 17463 8520
rect 17405 8511 17463 8517
rect 26510 8508 26516 8560
rect 26568 8548 26574 8560
rect 27341 8551 27399 8557
rect 27341 8548 27353 8551
rect 26568 8520 27353 8548
rect 26568 8508 26574 8520
rect 27341 8517 27353 8520
rect 27387 8517 27399 8551
rect 27706 8548 27712 8560
rect 27667 8520 27712 8548
rect 27341 8511 27399 8517
rect 27706 8508 27712 8520
rect 27764 8508 27770 8560
rect 16945 8483 17003 8489
rect 16945 8480 16957 8483
rect 16908 8452 16957 8480
rect 16908 8440 16914 8452
rect 16945 8449 16957 8452
rect 16991 8449 17003 8483
rect 16945 8443 17003 8449
rect 18414 8440 18420 8492
rect 18472 8480 18478 8492
rect 19153 8483 19211 8489
rect 19153 8480 19165 8483
rect 18472 8452 19165 8480
rect 18472 8440 18478 8452
rect 19153 8449 19165 8452
rect 19199 8449 19211 8483
rect 19153 8443 19211 8449
rect 12894 8372 12900 8424
rect 12952 8412 12958 8424
rect 13725 8415 13783 8421
rect 13725 8412 13737 8415
rect 12952 8384 13737 8412
rect 12952 8372 12958 8384
rect 13725 8381 13737 8384
rect 13771 8412 13783 8415
rect 14001 8415 14059 8421
rect 14001 8412 14013 8415
rect 13771 8384 14013 8412
rect 13771 8381 13783 8384
rect 13725 8375 13783 8381
rect 14001 8381 14013 8384
rect 14047 8381 14059 8415
rect 26418 8412 26424 8424
rect 26379 8384 26424 8412
rect 14001 8375 14059 8381
rect 26418 8372 26424 8384
rect 26476 8412 26482 8424
rect 26973 8415 27031 8421
rect 26973 8412 26985 8415
rect 26476 8384 26985 8412
rect 26476 8372 26482 8384
rect 26973 8381 26985 8384
rect 27019 8381 27031 8415
rect 27522 8412 27528 8424
rect 27483 8384 27528 8412
rect 26973 8375 27031 8381
rect 27522 8372 27528 8384
rect 27580 8412 27586 8424
rect 28077 8415 28135 8421
rect 28077 8412 28089 8415
rect 27580 8384 28089 8412
rect 27580 8372 27586 8384
rect 28077 8381 28089 8384
rect 28123 8381 28135 8415
rect 28077 8375 28135 8381
rect 3697 8347 3755 8353
rect 3697 8313 3709 8347
rect 3743 8344 3755 8347
rect 4034 8347 4092 8353
rect 4034 8344 4046 8347
rect 3743 8316 4046 8344
rect 3743 8313 3755 8316
rect 3697 8307 3755 8313
rect 4034 8313 4046 8316
rect 4080 8344 4092 8347
rect 6273 8347 6331 8353
rect 4080 8316 4200 8344
rect 4080 8313 4092 8316
rect 4034 8307 4092 8313
rect 1394 8236 1400 8288
rect 1452 8276 1458 8288
rect 1762 8276 1768 8288
rect 1452 8248 1768 8276
rect 1452 8236 1458 8248
rect 1762 8236 1768 8248
rect 1820 8236 1826 8288
rect 4172 8276 4200 8316
rect 6273 8313 6285 8347
rect 6319 8344 6331 8347
rect 6914 8344 6920 8356
rect 6319 8316 6920 8344
rect 6319 8313 6331 8316
rect 6273 8307 6331 8313
rect 6914 8304 6920 8316
rect 6972 8304 6978 8356
rect 7561 8347 7619 8353
rect 7561 8313 7573 8347
rect 7607 8344 7619 8347
rect 8573 8347 8631 8353
rect 8573 8344 8585 8347
rect 7607 8316 8585 8344
rect 7607 8313 7619 8316
rect 7561 8307 7619 8313
rect 8573 8313 8585 8316
rect 8619 8344 8631 8347
rect 8757 8347 8815 8353
rect 8757 8344 8769 8347
rect 8619 8316 8769 8344
rect 8619 8313 8631 8316
rect 8573 8307 8631 8313
rect 8757 8313 8769 8316
rect 8803 8313 8815 8347
rect 8757 8307 8815 8313
rect 10686 8304 10692 8356
rect 10744 8344 10750 8356
rect 11241 8347 11299 8353
rect 11241 8344 11253 8347
rect 10744 8316 11253 8344
rect 10744 8304 10750 8316
rect 11241 8313 11253 8316
rect 11287 8344 11299 8347
rect 11698 8344 11704 8356
rect 11287 8316 11704 8344
rect 11287 8313 11299 8316
rect 11241 8307 11299 8313
rect 11698 8304 11704 8316
rect 11756 8304 11762 8356
rect 12250 8344 12256 8356
rect 12211 8316 12256 8344
rect 12250 8304 12256 8316
rect 12308 8304 12314 8356
rect 15841 8347 15899 8353
rect 15841 8313 15853 8347
rect 15887 8344 15899 8347
rect 16669 8347 16727 8353
rect 16669 8344 16681 8347
rect 15887 8316 16681 8344
rect 15887 8313 15899 8316
rect 15841 8307 15899 8313
rect 16669 8313 16681 8316
rect 16715 8344 16727 8347
rect 17862 8344 17868 8356
rect 16715 8316 17868 8344
rect 16715 8313 16727 8316
rect 16669 8307 16727 8313
rect 17862 8304 17868 8316
rect 17920 8304 17926 8356
rect 19061 8347 19119 8353
rect 19061 8313 19073 8347
rect 19107 8344 19119 8347
rect 19420 8347 19478 8353
rect 19420 8344 19432 8347
rect 19107 8316 19432 8344
rect 19107 8313 19119 8316
rect 19061 8307 19119 8313
rect 19420 8313 19432 8316
rect 19466 8344 19478 8347
rect 19518 8344 19524 8356
rect 19466 8316 19524 8344
rect 19466 8313 19478 8316
rect 19420 8307 19478 8313
rect 19518 8304 19524 8316
rect 19576 8304 19582 8356
rect 4706 8276 4712 8288
rect 4172 8248 4712 8276
rect 4706 8236 4712 8248
rect 4764 8236 4770 8288
rect 7190 8276 7196 8288
rect 7151 8248 7196 8276
rect 7190 8236 7196 8248
rect 7248 8236 7254 8288
rect 10778 8276 10784 8288
rect 10739 8248 10784 8276
rect 10778 8236 10784 8248
rect 10836 8236 10842 8288
rect 11422 8236 11428 8288
rect 11480 8276 11486 8288
rect 12437 8279 12495 8285
rect 12437 8276 12449 8279
rect 11480 8248 12449 8276
rect 11480 8236 11486 8248
rect 12437 8245 12449 8248
rect 12483 8245 12495 8279
rect 12437 8239 12495 8245
rect 16301 8279 16359 8285
rect 16301 8245 16313 8279
rect 16347 8276 16359 8279
rect 16390 8276 16396 8288
rect 16347 8248 16396 8276
rect 16347 8245 16359 8248
rect 16301 8239 16359 8245
rect 16390 8236 16396 8248
rect 16448 8236 16454 8288
rect 20806 8236 20812 8288
rect 20864 8276 20870 8288
rect 21358 8276 21364 8288
rect 20864 8248 21364 8276
rect 20864 8236 20870 8248
rect 21358 8236 21364 8248
rect 21416 8236 21422 8288
rect 1104 8186 28888 8208
rect 1104 8134 10982 8186
rect 11034 8134 11046 8186
rect 11098 8134 11110 8186
rect 11162 8134 11174 8186
rect 11226 8134 20982 8186
rect 21034 8134 21046 8186
rect 21098 8134 21110 8186
rect 21162 8134 21174 8186
rect 21226 8134 28888 8186
rect 1104 8112 28888 8134
rect 1578 8072 1584 8084
rect 1539 8044 1584 8072
rect 1578 8032 1584 8044
rect 1636 8032 1642 8084
rect 3881 8075 3939 8081
rect 3881 8041 3893 8075
rect 3927 8072 3939 8075
rect 4062 8072 4068 8084
rect 3927 8044 4068 8072
rect 3927 8041 3939 8044
rect 3881 8035 3939 8041
rect 4062 8032 4068 8044
rect 4120 8032 4126 8084
rect 9950 8072 9956 8084
rect 9863 8044 9956 8072
rect 9950 8032 9956 8044
rect 10008 8072 10014 8084
rect 10870 8072 10876 8084
rect 10008 8044 10876 8072
rect 10008 8032 10014 8044
rect 10870 8032 10876 8044
rect 10928 8032 10934 8084
rect 17862 8072 17868 8084
rect 17823 8044 17868 8072
rect 17862 8032 17868 8044
rect 17920 8032 17926 8084
rect 18414 8072 18420 8084
rect 18375 8044 18420 8072
rect 18414 8032 18420 8044
rect 18472 8072 18478 8084
rect 19153 8075 19211 8081
rect 19153 8072 19165 8075
rect 18472 8044 19165 8072
rect 18472 8032 18478 8044
rect 19153 8041 19165 8044
rect 19199 8041 19211 8075
rect 19978 8072 19984 8084
rect 19939 8044 19984 8072
rect 19153 8035 19211 8041
rect 19978 8032 19984 8044
rect 20036 8032 20042 8084
rect 26694 8072 26700 8084
rect 26655 8044 26700 8072
rect 26694 8032 26700 8044
rect 26752 8032 26758 8084
rect 10502 8004 10508 8016
rect 10463 7976 10508 8004
rect 10502 7964 10508 7976
rect 10560 7964 10566 8016
rect 11054 7964 11060 8016
rect 11112 8004 11118 8016
rect 12894 8004 12900 8016
rect 11112 7976 12900 8004
rect 11112 7964 11118 7976
rect 12894 7964 12900 7976
rect 12952 7964 12958 8016
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7936 1455 7939
rect 2406 7936 2412 7948
rect 1443 7908 2412 7936
rect 1443 7905 1455 7908
rect 1397 7899 1455 7905
rect 2406 7896 2412 7908
rect 2464 7896 2470 7948
rect 6914 7896 6920 7948
rect 6972 7936 6978 7948
rect 7009 7939 7067 7945
rect 7009 7936 7021 7939
rect 6972 7908 7021 7936
rect 6972 7896 6978 7908
rect 7009 7905 7021 7908
rect 7055 7936 7067 7939
rect 7357 7939 7415 7945
rect 7357 7936 7369 7939
rect 7055 7908 7369 7936
rect 7055 7905 7067 7908
rect 7009 7899 7067 7905
rect 7357 7905 7369 7908
rect 7403 7936 7415 7939
rect 7834 7936 7840 7948
rect 7403 7908 7840 7936
rect 7403 7905 7415 7908
rect 7357 7899 7415 7905
rect 7834 7896 7840 7908
rect 7892 7896 7898 7948
rect 11241 7939 11299 7945
rect 11241 7905 11253 7939
rect 11287 7936 11299 7939
rect 11330 7936 11336 7948
rect 11287 7908 11336 7936
rect 11287 7905 11299 7908
rect 11241 7899 11299 7905
rect 11330 7896 11336 7908
rect 11388 7896 11394 7948
rect 16669 7939 16727 7945
rect 16669 7905 16681 7939
rect 16715 7936 16727 7939
rect 16942 7936 16948 7948
rect 16715 7908 16948 7936
rect 16715 7905 16727 7908
rect 16669 7899 16727 7905
rect 16942 7896 16948 7908
rect 17000 7896 17006 7948
rect 26510 7936 26516 7948
rect 26471 7908 26516 7936
rect 26510 7896 26516 7908
rect 26568 7896 26574 7948
rect 7101 7871 7159 7877
rect 7101 7837 7113 7871
rect 7147 7837 7159 7871
rect 16758 7868 16764 7880
rect 16719 7840 16764 7868
rect 7101 7831 7159 7837
rect 7116 7732 7144 7831
rect 16758 7828 16764 7840
rect 16816 7828 16822 7880
rect 16850 7828 16856 7880
rect 16908 7868 16914 7880
rect 16908 7840 16953 7868
rect 16908 7828 16914 7840
rect 16776 7800 16804 7828
rect 17494 7800 17500 7812
rect 16776 7772 17500 7800
rect 17494 7760 17500 7772
rect 17552 7760 17558 7812
rect 7282 7732 7288 7744
rect 7116 7704 7288 7732
rect 7282 7692 7288 7704
rect 7340 7692 7346 7744
rect 7466 7692 7472 7744
rect 7524 7732 7530 7744
rect 8481 7735 8539 7741
rect 8481 7732 8493 7735
rect 7524 7704 8493 7732
rect 7524 7692 7530 7704
rect 8481 7701 8493 7704
rect 8527 7701 8539 7735
rect 8481 7695 8539 7701
rect 10686 7692 10692 7744
rect 10744 7732 10750 7744
rect 10781 7735 10839 7741
rect 10781 7732 10793 7735
rect 10744 7704 10793 7732
rect 10744 7692 10750 7704
rect 10781 7701 10793 7704
rect 10827 7701 10839 7735
rect 10781 7695 10839 7701
rect 13449 7735 13507 7741
rect 13449 7701 13461 7735
rect 13495 7732 13507 7735
rect 13722 7732 13728 7744
rect 13495 7704 13728 7732
rect 13495 7701 13507 7704
rect 13449 7695 13507 7701
rect 13722 7692 13728 7704
rect 13780 7692 13786 7744
rect 15933 7735 15991 7741
rect 15933 7701 15945 7735
rect 15979 7732 15991 7735
rect 16298 7732 16304 7744
rect 15979 7704 16304 7732
rect 15979 7701 15991 7704
rect 15933 7695 15991 7701
rect 16298 7692 16304 7704
rect 16356 7692 16362 7744
rect 1104 7642 28888 7664
rect 1104 7590 5982 7642
rect 6034 7590 6046 7642
rect 6098 7590 6110 7642
rect 6162 7590 6174 7642
rect 6226 7590 15982 7642
rect 16034 7590 16046 7642
rect 16098 7590 16110 7642
rect 16162 7590 16174 7642
rect 16226 7590 25982 7642
rect 26034 7590 26046 7642
rect 26098 7590 26110 7642
rect 26162 7590 26174 7642
rect 26226 7590 28888 7642
rect 1104 7568 28888 7590
rect 2038 7528 2044 7540
rect 1999 7500 2044 7528
rect 2038 7488 2044 7500
rect 2096 7488 2102 7540
rect 4706 7528 4712 7540
rect 4667 7500 4712 7528
rect 4706 7488 4712 7500
rect 4764 7488 4770 7540
rect 8294 7488 8300 7540
rect 8352 7528 8358 7540
rect 9033 7531 9091 7537
rect 9033 7528 9045 7531
rect 8352 7500 9045 7528
rect 8352 7488 8358 7500
rect 9033 7497 9045 7500
rect 9079 7497 9091 7531
rect 11793 7531 11851 7537
rect 11793 7528 11805 7531
rect 9033 7491 9091 7497
rect 10152 7500 11805 7528
rect 1578 7460 1584 7472
rect 1539 7432 1584 7460
rect 1578 7420 1584 7432
rect 1636 7420 1642 7472
rect 5442 7420 5448 7472
rect 5500 7460 5506 7472
rect 6641 7463 6699 7469
rect 6641 7460 6653 7463
rect 5500 7432 6653 7460
rect 5500 7420 5506 7432
rect 6641 7429 6653 7432
rect 6687 7460 6699 7463
rect 6687 7432 7512 7460
rect 6687 7429 6699 7432
rect 6641 7423 6699 7429
rect 7484 7404 7512 7432
rect 10152 7404 10180 7500
rect 11793 7497 11805 7500
rect 11839 7497 11851 7531
rect 14734 7528 14740 7540
rect 14695 7500 14740 7528
rect 11793 7491 11851 7497
rect 14734 7488 14740 7500
rect 14792 7488 14798 7540
rect 17954 7488 17960 7540
rect 18012 7528 18018 7540
rect 19150 7528 19156 7540
rect 18012 7500 19156 7528
rect 18012 7488 18018 7500
rect 19150 7488 19156 7500
rect 19208 7488 19214 7540
rect 15749 7463 15807 7469
rect 15749 7429 15761 7463
rect 15795 7460 15807 7463
rect 16850 7460 16856 7472
rect 15795 7432 16856 7460
rect 15795 7429 15807 7432
rect 15749 7423 15807 7429
rect 16850 7420 16856 7432
rect 16908 7420 16914 7472
rect 19334 7420 19340 7472
rect 19392 7460 19398 7472
rect 19981 7463 20039 7469
rect 19981 7460 19993 7463
rect 19392 7432 19993 7460
rect 19392 7420 19398 7432
rect 19981 7429 19993 7432
rect 20027 7429 20039 7463
rect 19981 7423 20039 7429
rect 26510 7420 26516 7472
rect 26568 7460 26574 7472
rect 27341 7463 27399 7469
rect 27341 7460 27353 7463
rect 26568 7432 27353 7460
rect 26568 7420 26574 7432
rect 27341 7429 27353 7432
rect 27387 7429 27399 7463
rect 27341 7423 27399 7429
rect 7098 7352 7104 7404
rect 7156 7392 7162 7404
rect 7285 7395 7343 7401
rect 7285 7392 7297 7395
rect 7156 7364 7297 7392
rect 7156 7352 7162 7364
rect 7285 7361 7297 7364
rect 7331 7361 7343 7395
rect 7466 7392 7472 7404
rect 7427 7364 7472 7392
rect 7285 7355 7343 7361
rect 7466 7352 7472 7364
rect 7524 7352 7530 7404
rect 8941 7395 8999 7401
rect 8941 7361 8953 7395
rect 8987 7392 8999 7395
rect 10134 7392 10140 7404
rect 8987 7364 10140 7392
rect 8987 7361 8999 7364
rect 8941 7355 8999 7361
rect 10134 7352 10140 7364
rect 10192 7352 10198 7404
rect 16298 7392 16304 7404
rect 16259 7364 16304 7392
rect 16298 7352 16304 7364
rect 16356 7352 16362 7404
rect 16393 7395 16451 7401
rect 16393 7361 16405 7395
rect 16439 7361 16451 7395
rect 19518 7392 19524 7404
rect 19431 7364 19524 7392
rect 16393 7355 16451 7361
rect 1397 7327 1455 7333
rect 1397 7293 1409 7327
rect 1443 7324 1455 7327
rect 2038 7324 2044 7336
rect 1443 7296 2044 7324
rect 1443 7293 1455 7296
rect 1397 7287 1455 7293
rect 2038 7284 2044 7296
rect 2096 7284 2102 7336
rect 2406 7324 2412 7336
rect 2367 7296 2412 7324
rect 2406 7284 2412 7296
rect 2464 7284 2470 7336
rect 3329 7327 3387 7333
rect 3329 7293 3341 7327
rect 3375 7324 3387 7327
rect 3878 7324 3884 7336
rect 3375 7296 3884 7324
rect 3375 7293 3387 7296
rect 3329 7287 3387 7293
rect 3878 7284 3884 7296
rect 3936 7284 3942 7336
rect 6273 7327 6331 7333
rect 6273 7293 6285 7327
rect 6319 7324 6331 7327
rect 7190 7324 7196 7336
rect 6319 7296 7196 7324
rect 6319 7293 6331 7296
rect 6273 7287 6331 7293
rect 7190 7284 7196 7296
rect 7248 7284 7254 7336
rect 9214 7324 9220 7336
rect 9175 7296 9220 7324
rect 9214 7284 9220 7296
rect 9272 7284 9278 7336
rect 9950 7324 9956 7336
rect 9911 7296 9956 7324
rect 9950 7284 9956 7296
rect 10008 7284 10014 7336
rect 10318 7284 10324 7336
rect 10376 7324 10382 7336
rect 10413 7327 10471 7333
rect 10413 7324 10425 7327
rect 10376 7296 10425 7324
rect 10376 7284 10382 7296
rect 10413 7293 10425 7296
rect 10459 7293 10471 7327
rect 10413 7287 10471 7293
rect 10502 7284 10508 7336
rect 10560 7324 10566 7336
rect 10669 7327 10727 7333
rect 10669 7324 10681 7327
rect 10560 7296 10681 7324
rect 10560 7284 10566 7296
rect 10669 7293 10681 7296
rect 10715 7293 10727 7327
rect 10669 7287 10727 7293
rect 13357 7327 13415 7333
rect 13357 7293 13369 7327
rect 13403 7324 13415 7327
rect 13403 7296 13768 7324
rect 13403 7293 13415 7296
rect 13357 7287 13415 7293
rect 3237 7259 3295 7265
rect 3237 7225 3249 7259
rect 3283 7256 3295 7259
rect 3596 7259 3654 7265
rect 3596 7256 3608 7259
rect 3283 7228 3608 7256
rect 3283 7225 3295 7228
rect 3237 7219 3295 7225
rect 3596 7225 3608 7228
rect 3642 7256 3654 7259
rect 4062 7256 4068 7268
rect 3642 7228 4068 7256
rect 3642 7225 3654 7228
rect 3596 7219 3654 7225
rect 4062 7216 4068 7228
rect 4120 7216 4126 7268
rect 7282 7216 7288 7268
rect 7340 7256 7346 7268
rect 8297 7259 8355 7265
rect 8297 7256 8309 7259
rect 7340 7228 8309 7256
rect 7340 7216 7346 7228
rect 8297 7225 8309 7228
rect 8343 7256 8355 7259
rect 10336 7256 10364 7284
rect 13740 7268 13768 7296
rect 15930 7284 15936 7336
rect 15988 7324 15994 7336
rect 16408 7324 16436 7355
rect 19518 7352 19524 7364
rect 19576 7392 19582 7404
rect 20622 7392 20628 7404
rect 19576 7364 20628 7392
rect 19576 7352 19582 7364
rect 20622 7352 20628 7364
rect 20680 7352 20686 7404
rect 16942 7324 16948 7336
rect 15988 7296 16436 7324
rect 16903 7296 16948 7324
rect 15988 7284 15994 7296
rect 16942 7284 16948 7296
rect 17000 7284 17006 7336
rect 19978 7284 19984 7336
rect 20036 7324 20042 7336
rect 20349 7327 20407 7333
rect 20349 7324 20361 7327
rect 20036 7296 20361 7324
rect 20036 7284 20042 7296
rect 20349 7293 20361 7296
rect 20395 7293 20407 7327
rect 26418 7324 26424 7336
rect 26379 7296 26424 7324
rect 20349 7287 20407 7293
rect 26418 7284 26424 7296
rect 26476 7324 26482 7336
rect 26973 7327 27031 7333
rect 26973 7324 26985 7327
rect 26476 7296 26985 7324
rect 26476 7284 26482 7296
rect 26973 7293 26985 7296
rect 27019 7293 27031 7327
rect 26973 7287 27031 7293
rect 13602 7259 13660 7265
rect 13602 7256 13614 7259
rect 8343 7228 10364 7256
rect 13464 7228 13614 7256
rect 8343 7225 8355 7228
rect 8297 7219 8355 7225
rect 13464 7200 13492 7228
rect 13602 7225 13614 7228
rect 13648 7225 13660 7259
rect 13602 7219 13660 7225
rect 13722 7216 13728 7268
rect 13780 7216 13786 7268
rect 15381 7259 15439 7265
rect 15381 7225 15393 7259
rect 15427 7256 15439 7259
rect 16209 7259 16267 7265
rect 16209 7256 16221 7259
rect 15427 7228 16221 7256
rect 15427 7225 15439 7228
rect 15381 7219 15439 7225
rect 16209 7225 16221 7228
rect 16255 7256 16267 7259
rect 16390 7256 16396 7268
rect 16255 7228 16396 7256
rect 16255 7225 16267 7228
rect 16209 7219 16267 7225
rect 16390 7216 16396 7228
rect 16448 7216 16454 7268
rect 6822 7188 6828 7200
rect 6783 7160 6828 7188
rect 6822 7148 6828 7160
rect 6880 7148 6886 7200
rect 7834 7188 7840 7200
rect 7795 7160 7840 7188
rect 7834 7148 7840 7160
rect 7892 7148 7898 7200
rect 9582 7188 9588 7200
rect 9543 7160 9588 7188
rect 9582 7148 9588 7160
rect 9640 7148 9646 7200
rect 9950 7148 9956 7200
rect 10008 7188 10014 7200
rect 10045 7191 10103 7197
rect 10045 7188 10057 7191
rect 10008 7160 10057 7188
rect 10008 7148 10014 7160
rect 10045 7157 10057 7160
rect 10091 7188 10103 7191
rect 10778 7188 10784 7200
rect 10091 7160 10784 7188
rect 10091 7157 10103 7160
rect 10045 7151 10103 7157
rect 10778 7148 10784 7160
rect 10836 7148 10842 7200
rect 13265 7191 13323 7197
rect 13265 7157 13277 7191
rect 13311 7188 13323 7191
rect 13446 7188 13452 7200
rect 13311 7160 13452 7188
rect 13311 7157 13323 7160
rect 13265 7151 13323 7157
rect 13446 7148 13452 7160
rect 13504 7148 13510 7200
rect 15838 7188 15844 7200
rect 15799 7160 15844 7188
rect 15838 7148 15844 7160
rect 15896 7148 15902 7200
rect 19889 7191 19947 7197
rect 19889 7157 19901 7191
rect 19935 7188 19947 7191
rect 19978 7188 19984 7200
rect 19935 7160 19984 7188
rect 19935 7157 19947 7160
rect 19889 7151 19947 7157
rect 19978 7148 19984 7160
rect 20036 7188 20042 7200
rect 20441 7191 20499 7197
rect 20441 7188 20453 7191
rect 20036 7160 20453 7188
rect 20036 7148 20042 7160
rect 20441 7157 20453 7160
rect 20487 7157 20499 7191
rect 26602 7188 26608 7200
rect 26563 7160 26608 7188
rect 20441 7151 20499 7157
rect 26602 7148 26608 7160
rect 26660 7148 26666 7200
rect 1104 7098 28888 7120
rect 1104 7046 10982 7098
rect 11034 7046 11046 7098
rect 11098 7046 11110 7098
rect 11162 7046 11174 7098
rect 11226 7046 20982 7098
rect 21034 7046 21046 7098
rect 21098 7046 21110 7098
rect 21162 7046 21174 7098
rect 21226 7046 28888 7098
rect 1104 7024 28888 7046
rect 3421 6987 3479 6993
rect 3421 6953 3433 6987
rect 3467 6984 3479 6987
rect 3878 6984 3884 6996
rect 3467 6956 3884 6984
rect 3467 6953 3479 6956
rect 3421 6947 3479 6953
rect 3878 6944 3884 6956
rect 3936 6944 3942 6996
rect 4338 6944 4344 6996
rect 4396 6984 4402 6996
rect 4433 6987 4491 6993
rect 4433 6984 4445 6987
rect 4396 6956 4445 6984
rect 4396 6944 4402 6956
rect 4433 6953 4445 6956
rect 4479 6984 4491 6987
rect 6822 6984 6828 6996
rect 4479 6956 6828 6984
rect 4479 6953 4491 6956
rect 4433 6947 4491 6953
rect 6822 6944 6828 6956
rect 6880 6944 6886 6996
rect 7009 6987 7067 6993
rect 7009 6953 7021 6987
rect 7055 6984 7067 6987
rect 7098 6984 7104 6996
rect 7055 6956 7104 6984
rect 7055 6953 7067 6956
rect 7009 6947 7067 6953
rect 7098 6944 7104 6956
rect 7156 6944 7162 6996
rect 9125 6987 9183 6993
rect 9125 6953 9137 6987
rect 9171 6984 9183 6987
rect 9214 6984 9220 6996
rect 9171 6956 9220 6984
rect 9171 6953 9183 6956
rect 9125 6947 9183 6953
rect 9214 6944 9220 6956
rect 9272 6944 9278 6996
rect 9950 6984 9956 6996
rect 9911 6956 9956 6984
rect 9950 6944 9956 6956
rect 10008 6944 10014 6996
rect 10778 6944 10784 6996
rect 10836 6984 10842 6996
rect 11606 6984 11612 6996
rect 10836 6956 11612 6984
rect 10836 6944 10842 6956
rect 11606 6944 11612 6956
rect 11664 6944 11670 6996
rect 15930 6984 15936 6996
rect 15891 6956 15936 6984
rect 15930 6944 15936 6956
rect 15988 6984 15994 6996
rect 16390 6984 16396 6996
rect 15988 6956 16396 6984
rect 15988 6944 15994 6956
rect 16390 6944 16396 6956
rect 16448 6944 16454 6996
rect 6270 6916 6276 6928
rect 6231 6888 6276 6916
rect 6270 6876 6276 6888
rect 6328 6876 6334 6928
rect 10318 6876 10324 6928
rect 10376 6916 10382 6928
rect 16758 6916 16764 6928
rect 10376 6888 11008 6916
rect 10376 6876 10382 6888
rect 1394 6848 1400 6860
rect 1355 6820 1400 6848
rect 1394 6808 1400 6820
rect 1452 6808 1458 6860
rect 10594 6848 10600 6860
rect 10555 6820 10600 6848
rect 10594 6808 10600 6820
rect 10652 6808 10658 6860
rect 10689 6851 10747 6857
rect 10689 6817 10701 6851
rect 10735 6848 10747 6851
rect 10870 6848 10876 6860
rect 10735 6820 10876 6848
rect 10735 6817 10747 6820
rect 10689 6811 10747 6817
rect 10870 6808 10876 6820
rect 10928 6808 10934 6860
rect 10980 6848 11008 6888
rect 16500 6888 16764 6916
rect 11609 6851 11667 6857
rect 11609 6848 11621 6851
rect 10980 6820 11621 6848
rect 11609 6817 11621 6820
rect 11655 6817 11667 6851
rect 12158 6848 12164 6860
rect 12119 6820 12164 6848
rect 11609 6811 11667 6817
rect 12158 6808 12164 6820
rect 12216 6808 12222 6860
rect 16500 6848 16528 6888
rect 16758 6876 16764 6888
rect 16816 6876 16822 6928
rect 16850 6876 16856 6928
rect 16908 6916 16914 6928
rect 17374 6919 17432 6925
rect 17374 6916 17386 6919
rect 16908 6888 17386 6916
rect 16908 6876 16914 6888
rect 17374 6885 17386 6888
rect 17420 6885 17432 6919
rect 17374 6879 17432 6885
rect 16316 6820 16528 6848
rect 4522 6780 4528 6792
rect 4483 6752 4528 6780
rect 4522 6740 4528 6752
rect 4580 6740 4586 6792
rect 4706 6780 4712 6792
rect 4667 6752 4712 6780
rect 4706 6740 4712 6752
rect 4764 6740 4770 6792
rect 5626 6740 5632 6792
rect 5684 6780 5690 6792
rect 6365 6783 6423 6789
rect 6365 6780 6377 6783
rect 5684 6752 6377 6780
rect 5684 6740 5690 6752
rect 6365 6749 6377 6752
rect 6411 6749 6423 6783
rect 6546 6780 6552 6792
rect 6507 6752 6552 6780
rect 6365 6743 6423 6749
rect 1578 6712 1584 6724
rect 1539 6684 1584 6712
rect 1578 6672 1584 6684
rect 1636 6672 1642 6724
rect 6380 6712 6408 6743
rect 6546 6740 6552 6752
rect 6604 6740 6610 6792
rect 10134 6740 10140 6792
rect 10192 6780 10198 6792
rect 10781 6783 10839 6789
rect 10781 6780 10793 6783
rect 10192 6752 10793 6780
rect 10192 6740 10198 6752
rect 10781 6749 10793 6752
rect 10827 6749 10839 6783
rect 10781 6743 10839 6749
rect 11974 6740 11980 6792
rect 12032 6780 12038 6792
rect 12253 6783 12311 6789
rect 12253 6780 12265 6783
rect 12032 6752 12265 6780
rect 12032 6740 12038 6752
rect 12253 6749 12265 6752
rect 12299 6749 12311 6783
rect 12253 6743 12311 6749
rect 12437 6783 12495 6789
rect 12437 6749 12449 6783
rect 12483 6780 12495 6783
rect 12483 6752 13308 6780
rect 12483 6749 12495 6752
rect 12437 6743 12495 6749
rect 6822 6712 6828 6724
rect 6380 6684 6828 6712
rect 6822 6672 6828 6684
rect 6880 6672 6886 6724
rect 10042 6672 10048 6724
rect 10100 6712 10106 6724
rect 11992 6712 12020 6740
rect 10100 6684 12020 6712
rect 10100 6672 10106 6684
rect 12342 6672 12348 6724
rect 12400 6712 12406 6724
rect 12400 6684 12940 6712
rect 12400 6672 12406 6684
rect 12912 6656 12940 6684
rect 3602 6604 3608 6656
rect 3660 6644 3666 6656
rect 4065 6647 4123 6653
rect 4065 6644 4077 6647
rect 3660 6616 4077 6644
rect 3660 6604 3666 6616
rect 4065 6613 4077 6616
rect 4111 6613 4123 6647
rect 4065 6607 4123 6613
rect 5810 6604 5816 6656
rect 5868 6644 5874 6656
rect 5905 6647 5963 6653
rect 5905 6644 5917 6647
rect 5868 6616 5917 6644
rect 5868 6604 5874 6616
rect 5905 6613 5917 6616
rect 5951 6613 5963 6647
rect 7558 6644 7564 6656
rect 7519 6616 7564 6644
rect 5905 6607 5963 6613
rect 7558 6604 7564 6616
rect 7616 6604 7622 6656
rect 10226 6644 10232 6656
rect 10187 6616 10232 6644
rect 10226 6604 10232 6616
rect 10284 6604 10290 6656
rect 10778 6604 10784 6656
rect 10836 6644 10842 6656
rect 11241 6647 11299 6653
rect 11241 6644 11253 6647
rect 10836 6616 11253 6644
rect 10836 6604 10842 6616
rect 11241 6613 11253 6616
rect 11287 6644 11299 6647
rect 11330 6644 11336 6656
rect 11287 6616 11336 6644
rect 11287 6613 11299 6616
rect 11241 6607 11299 6613
rect 11330 6604 11336 6616
rect 11388 6604 11394 6656
rect 11790 6644 11796 6656
rect 11751 6616 11796 6644
rect 11790 6604 11796 6616
rect 11848 6604 11854 6656
rect 12894 6644 12900 6656
rect 12855 6616 12900 6644
rect 12894 6604 12900 6616
rect 12952 6604 12958 6656
rect 13280 6653 13308 6752
rect 13265 6647 13323 6653
rect 13265 6613 13277 6647
rect 13311 6644 13323 6647
rect 13446 6644 13452 6656
rect 13311 6616 13452 6644
rect 13311 6613 13323 6616
rect 13265 6607 13323 6613
rect 13446 6604 13452 6616
rect 13504 6604 13510 6656
rect 15470 6604 15476 6656
rect 15528 6644 15534 6656
rect 16316 6653 16344 6820
rect 19886 6808 19892 6860
rect 19944 6848 19950 6860
rect 19981 6851 20039 6857
rect 19981 6848 19993 6851
rect 19944 6820 19993 6848
rect 19944 6808 19950 6820
rect 19981 6817 19993 6820
rect 20027 6817 20039 6851
rect 26510 6848 26516 6860
rect 26471 6820 26516 6848
rect 19981 6811 20039 6817
rect 26510 6808 26516 6820
rect 26568 6808 26574 6860
rect 16666 6740 16672 6792
rect 16724 6780 16730 6792
rect 17129 6783 17187 6789
rect 17129 6780 17141 6783
rect 16724 6752 17141 6780
rect 16724 6740 16730 6752
rect 17129 6749 17141 6752
rect 17175 6749 17187 6783
rect 17129 6743 17187 6749
rect 26694 6712 26700 6724
rect 26655 6684 26700 6712
rect 26694 6672 26700 6684
rect 26752 6672 26758 6724
rect 16301 6647 16359 6653
rect 16301 6644 16313 6647
rect 15528 6616 16313 6644
rect 15528 6604 15534 6616
rect 16301 6613 16313 6616
rect 16347 6613 16359 6647
rect 16301 6607 16359 6613
rect 18138 6604 18144 6656
rect 18196 6644 18202 6656
rect 18509 6647 18567 6653
rect 18509 6644 18521 6647
rect 18196 6616 18521 6644
rect 18196 6604 18202 6616
rect 18509 6613 18521 6616
rect 18555 6613 18567 6647
rect 21634 6644 21640 6656
rect 21595 6616 21640 6644
rect 18509 6607 18567 6613
rect 21634 6604 21640 6616
rect 21692 6604 21698 6656
rect 1104 6554 28888 6576
rect 1104 6502 5982 6554
rect 6034 6502 6046 6554
rect 6098 6502 6110 6554
rect 6162 6502 6174 6554
rect 6226 6502 15982 6554
rect 16034 6502 16046 6554
rect 16098 6502 16110 6554
rect 16162 6502 16174 6554
rect 16226 6502 25982 6554
rect 26034 6502 26046 6554
rect 26098 6502 26110 6554
rect 26162 6502 26174 6554
rect 26226 6502 28888 6554
rect 1104 6480 28888 6502
rect 1394 6400 1400 6452
rect 1452 6440 1458 6452
rect 2317 6443 2375 6449
rect 2317 6440 2329 6443
rect 1452 6412 2329 6440
rect 1452 6400 1458 6412
rect 2317 6409 2329 6412
rect 2363 6409 2375 6443
rect 2317 6403 2375 6409
rect 3789 6443 3847 6449
rect 3789 6409 3801 6443
rect 3835 6440 3847 6443
rect 4522 6440 4528 6452
rect 3835 6412 4528 6440
rect 3835 6409 3847 6412
rect 3789 6403 3847 6409
rect 4522 6400 4528 6412
rect 4580 6440 4586 6452
rect 4617 6443 4675 6449
rect 4617 6440 4629 6443
rect 4580 6412 4629 6440
rect 4580 6400 4586 6412
rect 4617 6409 4629 6412
rect 4663 6409 4675 6443
rect 4617 6403 4675 6409
rect 5626 6400 5632 6452
rect 5684 6440 5690 6452
rect 5905 6443 5963 6449
rect 5905 6440 5917 6443
rect 5684 6412 5917 6440
rect 5684 6400 5690 6412
rect 5905 6409 5917 6412
rect 5951 6409 5963 6443
rect 6270 6440 6276 6452
rect 6231 6412 6276 6440
rect 5905 6403 5963 6409
rect 6270 6400 6276 6412
rect 6328 6400 6334 6452
rect 7834 6400 7840 6452
rect 7892 6440 7898 6452
rect 8941 6443 8999 6449
rect 8941 6440 8953 6443
rect 7892 6412 8953 6440
rect 7892 6400 7898 6412
rect 8941 6409 8953 6412
rect 8987 6409 8999 6443
rect 10134 6440 10140 6452
rect 10095 6412 10140 6440
rect 8941 6403 8999 6409
rect 10134 6400 10140 6412
rect 10192 6400 10198 6452
rect 10318 6400 10324 6452
rect 10376 6440 10382 6452
rect 10505 6443 10563 6449
rect 10505 6440 10517 6443
rect 10376 6412 10517 6440
rect 10376 6400 10382 6412
rect 1578 6372 1584 6384
rect 1539 6344 1584 6372
rect 1578 6332 1584 6344
rect 1636 6332 1642 6384
rect 2038 6372 2044 6384
rect 1999 6344 2044 6372
rect 2038 6332 2044 6344
rect 2096 6332 2102 6384
rect 4157 6375 4215 6381
rect 4157 6341 4169 6375
rect 4203 6372 4215 6375
rect 4706 6372 4712 6384
rect 4203 6344 4712 6372
rect 4203 6341 4215 6344
rect 4157 6335 4215 6341
rect 4706 6332 4712 6344
rect 4764 6332 4770 6384
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6236 1455 6239
rect 2056 6236 2084 6332
rect 4246 6264 4252 6316
rect 4304 6304 4310 6316
rect 4525 6307 4583 6313
rect 4525 6304 4537 6307
rect 4304 6276 4537 6304
rect 4304 6264 4310 6276
rect 4525 6273 4537 6276
rect 4571 6304 4583 6307
rect 5261 6307 5319 6313
rect 5261 6304 5273 6307
rect 4571 6276 5273 6304
rect 4571 6273 4583 6276
rect 4525 6267 4583 6273
rect 5261 6273 5273 6276
rect 5307 6304 5319 6307
rect 5442 6304 5448 6316
rect 5307 6276 5448 6304
rect 5307 6273 5319 6276
rect 5261 6267 5319 6273
rect 5442 6264 5448 6276
rect 5500 6264 5506 6316
rect 7558 6304 7564 6316
rect 7519 6276 7564 6304
rect 7558 6264 7564 6276
rect 7616 6264 7622 6316
rect 1443 6208 2084 6236
rect 7576 6236 7604 6264
rect 8202 6236 8208 6248
rect 7576 6208 8208 6236
rect 1443 6205 1455 6208
rect 1397 6199 1455 6205
rect 8202 6196 8208 6208
rect 8260 6196 8266 6248
rect 10428 6236 10456 6412
rect 10505 6409 10517 6412
rect 10551 6409 10563 6443
rect 10505 6403 10563 6409
rect 10594 6400 10600 6452
rect 10652 6440 10658 6452
rect 10689 6443 10747 6449
rect 10689 6440 10701 6443
rect 10652 6412 10701 6440
rect 10652 6400 10658 6412
rect 10689 6409 10701 6412
rect 10735 6409 10747 6443
rect 12158 6440 12164 6452
rect 12119 6412 12164 6440
rect 10689 6403 10747 6409
rect 12158 6400 12164 6412
rect 12216 6400 12222 6452
rect 13814 6400 13820 6452
rect 13872 6440 13878 6452
rect 14829 6443 14887 6449
rect 14829 6440 14841 6443
rect 13872 6412 14841 6440
rect 13872 6400 13878 6412
rect 10502 6264 10508 6316
rect 10560 6304 10566 6316
rect 11241 6307 11299 6313
rect 11241 6304 11253 6307
rect 10560 6276 11253 6304
rect 10560 6264 10566 6276
rect 11241 6273 11253 6276
rect 11287 6273 11299 6307
rect 11241 6267 11299 6273
rect 12713 6307 12771 6313
rect 12713 6273 12725 6307
rect 12759 6304 12771 6307
rect 13446 6304 13452 6316
rect 12759 6276 13308 6304
rect 13407 6276 13452 6304
rect 12759 6273 12771 6276
rect 12713 6267 12771 6273
rect 11054 6236 11060 6248
rect 10428 6208 11060 6236
rect 11054 6196 11060 6208
rect 11112 6196 11118 6248
rect 11149 6239 11207 6245
rect 11149 6205 11161 6239
rect 11195 6236 11207 6239
rect 11330 6236 11336 6248
rect 11195 6208 11336 6236
rect 11195 6205 11207 6208
rect 11149 6199 11207 6205
rect 11330 6196 11336 6208
rect 11388 6236 11394 6248
rect 11790 6236 11796 6248
rect 11388 6208 11796 6236
rect 11388 6196 11394 6208
rect 11790 6196 11796 6208
rect 11848 6196 11854 6248
rect 12894 6196 12900 6248
rect 12952 6236 12958 6248
rect 13280 6245 13308 6276
rect 13446 6264 13452 6276
rect 13504 6264 13510 6316
rect 13173 6239 13231 6245
rect 13173 6236 13185 6239
rect 12952 6208 13185 6236
rect 12952 6196 12958 6208
rect 13173 6205 13185 6208
rect 13219 6205 13231 6239
rect 13173 6199 13231 6205
rect 13265 6239 13323 6245
rect 13265 6205 13277 6239
rect 13311 6236 13323 6239
rect 13354 6236 13360 6248
rect 13311 6208 13360 6236
rect 13311 6205 13323 6208
rect 13265 6199 13323 6205
rect 13354 6196 13360 6208
rect 13412 6196 13418 6248
rect 14568 6245 14596 6412
rect 14829 6409 14841 6412
rect 14875 6409 14887 6443
rect 14829 6403 14887 6409
rect 16850 6400 16856 6452
rect 16908 6440 16914 6452
rect 17129 6443 17187 6449
rect 17129 6440 17141 6443
rect 16908 6412 17141 6440
rect 16908 6400 16914 6412
rect 17129 6409 17141 6412
rect 17175 6440 17187 6443
rect 18233 6443 18291 6449
rect 18233 6440 18245 6443
rect 17175 6412 18245 6440
rect 17175 6409 17187 6412
rect 17129 6403 17187 6409
rect 18233 6409 18245 6412
rect 18279 6440 18291 6443
rect 18966 6440 18972 6452
rect 18279 6412 18972 6440
rect 18279 6409 18291 6412
rect 18233 6403 18291 6409
rect 18966 6400 18972 6412
rect 19024 6400 19030 6452
rect 26510 6400 26516 6452
rect 26568 6440 26574 6452
rect 27341 6443 27399 6449
rect 27341 6440 27353 6443
rect 26568 6412 27353 6440
rect 26568 6400 26574 6412
rect 27341 6409 27353 6412
rect 27387 6409 27399 6443
rect 27341 6403 27399 6409
rect 19981 6375 20039 6381
rect 19981 6372 19993 6375
rect 18892 6344 19993 6372
rect 18506 6264 18512 6316
rect 18564 6304 18570 6316
rect 18892 6313 18920 6344
rect 19981 6341 19993 6344
rect 20027 6341 20039 6375
rect 26602 6372 26608 6384
rect 26563 6344 26608 6372
rect 19981 6335 20039 6341
rect 26602 6332 26608 6344
rect 26660 6332 26666 6384
rect 18877 6307 18935 6313
rect 18877 6304 18889 6307
rect 18564 6276 18889 6304
rect 18564 6264 18570 6276
rect 18877 6273 18889 6276
rect 18923 6273 18935 6307
rect 18877 6267 18935 6273
rect 18966 6264 18972 6316
rect 19024 6304 19030 6316
rect 19794 6304 19800 6316
rect 19024 6276 19069 6304
rect 19755 6276 19800 6304
rect 19024 6264 19030 6276
rect 19794 6264 19800 6276
rect 19852 6304 19858 6316
rect 20441 6307 20499 6313
rect 20441 6304 20453 6307
rect 19852 6276 20453 6304
rect 19852 6264 19858 6276
rect 20441 6273 20453 6276
rect 20487 6273 20499 6307
rect 20622 6304 20628 6316
rect 20535 6276 20628 6304
rect 20441 6267 20499 6273
rect 20622 6264 20628 6276
rect 20680 6304 20686 6316
rect 21634 6304 21640 6316
rect 20680 6276 21640 6304
rect 20680 6264 20686 6276
rect 21634 6264 21640 6276
rect 21692 6304 21698 6316
rect 22097 6307 22155 6313
rect 22097 6304 22109 6307
rect 21692 6276 22109 6304
rect 21692 6264 21698 6276
rect 22097 6273 22109 6276
rect 22143 6273 22155 6307
rect 22097 6267 22155 6273
rect 14553 6239 14611 6245
rect 14553 6205 14565 6239
rect 14599 6205 14611 6239
rect 14553 6199 14611 6205
rect 17865 6239 17923 6245
rect 17865 6205 17877 6239
rect 17911 6236 17923 6239
rect 18785 6239 18843 6245
rect 18785 6236 18797 6239
rect 17911 6208 18797 6236
rect 17911 6205 17923 6208
rect 17865 6199 17923 6205
rect 18785 6205 18797 6208
rect 18831 6236 18843 6239
rect 19242 6236 19248 6248
rect 18831 6208 19248 6236
rect 18831 6205 18843 6208
rect 18785 6199 18843 6205
rect 19242 6196 19248 6208
rect 19300 6196 19306 6248
rect 19521 6239 19579 6245
rect 19521 6205 19533 6239
rect 19567 6236 19579 6239
rect 20640 6236 20668 6264
rect 21910 6236 21916 6248
rect 19567 6208 20668 6236
rect 21871 6208 21916 6236
rect 19567 6205 19579 6208
rect 19521 6199 19579 6205
rect 21910 6196 21916 6208
rect 21968 6196 21974 6248
rect 26418 6236 26424 6248
rect 26379 6208 26424 6236
rect 26418 6196 26424 6208
rect 26476 6236 26482 6248
rect 26973 6239 27031 6245
rect 26973 6236 26985 6239
rect 26476 6208 26985 6236
rect 26476 6196 26482 6208
rect 26973 6205 26985 6208
rect 27019 6205 27031 6239
rect 26973 6199 27031 6205
rect 7806 6171 7864 6177
rect 7806 6168 7818 6171
rect 7484 6140 7818 6168
rect 7484 6112 7512 6140
rect 7806 6137 7818 6140
rect 7852 6137 7864 6171
rect 7806 6131 7864 6137
rect 9861 6171 9919 6177
rect 9861 6137 9873 6171
rect 9907 6168 9919 6171
rect 10870 6168 10876 6180
rect 9907 6140 10876 6168
rect 9907 6137 9919 6140
rect 9861 6131 9919 6137
rect 10870 6128 10876 6140
rect 10928 6128 10934 6180
rect 19886 6128 19892 6180
rect 19944 6168 19950 6180
rect 20349 6171 20407 6177
rect 20349 6168 20361 6171
rect 19944 6140 20361 6168
rect 19944 6128 19950 6140
rect 20349 6137 20361 6140
rect 20395 6137 20407 6171
rect 22005 6171 22063 6177
rect 22005 6168 22017 6171
rect 20349 6131 20407 6137
rect 21376 6140 22017 6168
rect 4982 6100 4988 6112
rect 4943 6072 4988 6100
rect 4982 6060 4988 6072
rect 5040 6060 5046 6112
rect 5074 6060 5080 6112
rect 5132 6100 5138 6112
rect 7466 6100 7472 6112
rect 5132 6072 5177 6100
rect 7427 6072 7472 6100
rect 5132 6060 5138 6072
rect 7466 6060 7472 6072
rect 7524 6060 7530 6112
rect 11882 6100 11888 6112
rect 11843 6072 11888 6100
rect 11882 6060 11888 6072
rect 11940 6060 11946 6112
rect 12802 6100 12808 6112
rect 12763 6072 12808 6100
rect 12802 6060 12808 6072
rect 12860 6060 12866 6112
rect 13722 6060 13728 6112
rect 13780 6100 13786 6112
rect 14369 6103 14427 6109
rect 14369 6100 14381 6103
rect 13780 6072 14381 6100
rect 13780 6060 13786 6072
rect 14369 6069 14381 6072
rect 14415 6100 14427 6103
rect 14550 6100 14556 6112
rect 14415 6072 14556 6100
rect 14415 6069 14427 6072
rect 14369 6063 14427 6069
rect 14550 6060 14556 6072
rect 14608 6060 14614 6112
rect 16666 6060 16672 6112
rect 16724 6100 16730 6112
rect 16761 6103 16819 6109
rect 16761 6100 16773 6103
rect 16724 6072 16773 6100
rect 16724 6060 16730 6072
rect 16761 6069 16773 6072
rect 16807 6069 16819 6103
rect 18414 6100 18420 6112
rect 18375 6072 18420 6100
rect 16761 6063 16819 6069
rect 18414 6060 18420 6072
rect 18472 6060 18478 6112
rect 20806 6060 20812 6112
rect 20864 6100 20870 6112
rect 21376 6109 21404 6140
rect 22005 6137 22017 6140
rect 22051 6137 22063 6171
rect 22005 6131 22063 6137
rect 21361 6103 21419 6109
rect 21361 6100 21373 6103
rect 20864 6072 21373 6100
rect 20864 6060 20870 6072
rect 21361 6069 21373 6072
rect 21407 6069 21419 6103
rect 21542 6100 21548 6112
rect 21503 6072 21548 6100
rect 21361 6063 21419 6069
rect 21542 6060 21548 6072
rect 21600 6060 21606 6112
rect 1104 6010 28888 6032
rect 1104 5958 10982 6010
rect 11034 5958 11046 6010
rect 11098 5958 11110 6010
rect 11162 5958 11174 6010
rect 11226 5958 20982 6010
rect 21034 5958 21046 6010
rect 21098 5958 21110 6010
rect 21162 5958 21174 6010
rect 21226 5958 28888 6010
rect 1104 5936 28888 5958
rect 4338 5896 4344 5908
rect 4299 5868 4344 5896
rect 4338 5856 4344 5868
rect 4396 5856 4402 5908
rect 4982 5896 4988 5908
rect 4943 5868 4988 5896
rect 4982 5856 4988 5868
rect 5040 5896 5046 5908
rect 5445 5899 5503 5905
rect 5445 5896 5457 5899
rect 5040 5868 5457 5896
rect 5040 5856 5046 5868
rect 5445 5865 5457 5868
rect 5491 5865 5503 5899
rect 5445 5859 5503 5865
rect 5534 5856 5540 5908
rect 5592 5896 5598 5908
rect 5810 5896 5816 5908
rect 5592 5868 5816 5896
rect 5592 5856 5598 5868
rect 5810 5856 5816 5868
rect 5868 5896 5874 5908
rect 5905 5899 5963 5905
rect 5905 5896 5917 5899
rect 5868 5868 5917 5896
rect 5868 5856 5874 5868
rect 5905 5865 5917 5868
rect 5951 5865 5963 5899
rect 7006 5896 7012 5908
rect 6967 5868 7012 5896
rect 5905 5859 5963 5865
rect 7006 5856 7012 5868
rect 7064 5856 7070 5908
rect 9493 5899 9551 5905
rect 9493 5865 9505 5899
rect 9539 5896 9551 5899
rect 9582 5896 9588 5908
rect 9539 5868 9588 5896
rect 9539 5865 9551 5868
rect 9493 5859 9551 5865
rect 9582 5856 9588 5868
rect 9640 5856 9646 5908
rect 10321 5899 10379 5905
rect 10321 5865 10333 5899
rect 10367 5896 10379 5899
rect 10594 5896 10600 5908
rect 10367 5868 10600 5896
rect 10367 5865 10379 5868
rect 10321 5859 10379 5865
rect 10594 5856 10600 5868
rect 10652 5856 10658 5908
rect 11149 5899 11207 5905
rect 11149 5865 11161 5899
rect 11195 5896 11207 5899
rect 11330 5896 11336 5908
rect 11195 5868 11336 5896
rect 11195 5865 11207 5868
rect 11149 5859 11207 5865
rect 11330 5856 11336 5868
rect 11388 5856 11394 5908
rect 11698 5896 11704 5908
rect 11611 5868 11704 5896
rect 11698 5856 11704 5868
rect 11756 5896 11762 5908
rect 12802 5896 12808 5908
rect 11756 5868 12808 5896
rect 11756 5856 11762 5868
rect 12802 5856 12808 5868
rect 12860 5856 12866 5908
rect 13262 5896 13268 5908
rect 13223 5868 13268 5896
rect 13262 5856 13268 5868
rect 13320 5856 13326 5908
rect 15749 5899 15807 5905
rect 15749 5865 15761 5899
rect 15795 5896 15807 5899
rect 15838 5896 15844 5908
rect 15795 5868 15844 5896
rect 15795 5865 15807 5868
rect 15749 5859 15807 5865
rect 15838 5856 15844 5868
rect 15896 5896 15902 5908
rect 16574 5896 16580 5908
rect 15896 5868 16580 5896
rect 15896 5856 15902 5868
rect 16574 5856 16580 5868
rect 16632 5856 16638 5908
rect 18506 5896 18512 5908
rect 18467 5868 18512 5896
rect 18506 5856 18512 5868
rect 18564 5856 18570 5908
rect 19610 5896 19616 5908
rect 19571 5868 19616 5896
rect 19610 5856 19616 5868
rect 19668 5856 19674 5908
rect 19705 5899 19763 5905
rect 19705 5865 19717 5899
rect 19751 5896 19763 5899
rect 20162 5896 20168 5908
rect 19751 5868 20168 5896
rect 19751 5865 19763 5868
rect 19705 5859 19763 5865
rect 20162 5856 20168 5868
rect 20220 5896 20226 5908
rect 21542 5896 21548 5908
rect 20220 5868 21548 5896
rect 20220 5856 20226 5868
rect 21542 5856 21548 5868
rect 21600 5856 21606 5908
rect 21637 5899 21695 5905
rect 21637 5865 21649 5899
rect 21683 5896 21695 5899
rect 21910 5896 21916 5908
rect 21683 5868 21916 5896
rect 21683 5865 21695 5868
rect 21637 5859 21695 5865
rect 21910 5856 21916 5868
rect 21968 5856 21974 5908
rect 4709 5831 4767 5837
rect 4709 5797 4721 5831
rect 4755 5828 4767 5831
rect 5074 5828 5080 5840
rect 4755 5800 5080 5828
rect 4755 5797 4767 5800
rect 4709 5791 4767 5797
rect 5074 5788 5080 5800
rect 5132 5788 5138 5840
rect 6917 5831 6975 5837
rect 6917 5797 6929 5831
rect 6963 5828 6975 5831
rect 7190 5828 7196 5840
rect 6963 5800 7196 5828
rect 6963 5797 6975 5800
rect 6917 5791 6975 5797
rect 7190 5788 7196 5800
rect 7248 5828 7254 5840
rect 7742 5828 7748 5840
rect 7248 5800 7748 5828
rect 7248 5788 7254 5800
rect 7742 5788 7748 5800
rect 7800 5788 7806 5840
rect 10502 5788 10508 5840
rect 10560 5828 10566 5840
rect 10689 5831 10747 5837
rect 10689 5828 10701 5831
rect 10560 5800 10701 5828
rect 10560 5788 10566 5800
rect 10689 5797 10701 5800
rect 10735 5797 10747 5831
rect 13170 5828 13176 5840
rect 13131 5800 13176 5828
rect 10689 5791 10747 5797
rect 1397 5763 1455 5769
rect 1397 5729 1409 5763
rect 1443 5760 1455 5763
rect 2406 5760 2412 5772
rect 1443 5732 2412 5760
rect 1443 5729 1455 5732
rect 1397 5723 1455 5729
rect 2406 5720 2412 5732
rect 2464 5720 2470 5772
rect 5810 5760 5816 5772
rect 5771 5732 5816 5760
rect 5810 5720 5816 5732
rect 5868 5720 5874 5772
rect 7374 5760 7380 5772
rect 7335 5732 7380 5760
rect 7374 5720 7380 5732
rect 7432 5720 7438 5772
rect 5997 5695 6055 5701
rect 5997 5661 6009 5695
rect 6043 5661 6055 5695
rect 5997 5655 6055 5661
rect 1578 5624 1584 5636
rect 1539 5596 1584 5624
rect 1578 5584 1584 5596
rect 1636 5584 1642 5636
rect 5810 5584 5816 5636
rect 5868 5624 5874 5636
rect 6012 5624 6040 5655
rect 7098 5652 7104 5704
rect 7156 5692 7162 5704
rect 7469 5695 7527 5701
rect 7469 5692 7481 5695
rect 7156 5664 7481 5692
rect 7156 5652 7162 5664
rect 7469 5661 7481 5664
rect 7515 5661 7527 5695
rect 7469 5655 7527 5661
rect 7561 5695 7619 5701
rect 7561 5661 7573 5695
rect 7607 5661 7619 5695
rect 10704 5692 10732 5791
rect 13170 5788 13176 5800
rect 13228 5788 13234 5840
rect 11609 5763 11667 5769
rect 11609 5729 11621 5763
rect 11655 5760 11667 5763
rect 11974 5760 11980 5772
rect 11655 5732 11980 5760
rect 11655 5729 11667 5732
rect 11609 5723 11667 5729
rect 11974 5720 11980 5732
rect 12032 5720 12038 5772
rect 26510 5760 26516 5772
rect 26471 5732 26516 5760
rect 26510 5720 26516 5732
rect 26568 5720 26574 5772
rect 11330 5692 11336 5704
rect 10704 5664 11336 5692
rect 7561 5655 7619 5661
rect 7576 5624 7604 5655
rect 11330 5652 11336 5664
rect 11388 5692 11394 5704
rect 11793 5695 11851 5701
rect 11793 5692 11805 5695
rect 11388 5664 11805 5692
rect 11388 5652 11394 5664
rect 11793 5661 11805 5664
rect 11839 5661 11851 5695
rect 11793 5655 11851 5661
rect 12345 5695 12403 5701
rect 12345 5661 12357 5695
rect 12391 5692 12403 5695
rect 13446 5692 13452 5704
rect 12391 5664 13452 5692
rect 12391 5661 12403 5664
rect 12345 5655 12403 5661
rect 13446 5652 13452 5664
rect 13504 5652 13510 5704
rect 15838 5692 15844 5704
rect 15799 5664 15844 5692
rect 15838 5652 15844 5664
rect 15896 5652 15902 5704
rect 16025 5695 16083 5701
rect 16025 5661 16037 5695
rect 16071 5692 16083 5695
rect 16298 5692 16304 5704
rect 16071 5664 16304 5692
rect 16071 5661 16083 5664
rect 16025 5655 16083 5661
rect 16298 5652 16304 5664
rect 16356 5652 16362 5704
rect 18966 5652 18972 5704
rect 19024 5692 19030 5704
rect 19702 5692 19708 5704
rect 19024 5664 19708 5692
rect 19024 5652 19030 5664
rect 19702 5652 19708 5664
rect 19760 5692 19766 5704
rect 19797 5695 19855 5701
rect 19797 5692 19809 5695
rect 19760 5664 19809 5692
rect 19760 5652 19766 5664
rect 19797 5661 19809 5664
rect 19843 5661 19855 5695
rect 19797 5655 19855 5661
rect 7834 5624 7840 5636
rect 5868 5596 7840 5624
rect 5868 5584 5874 5596
rect 7834 5584 7840 5596
rect 7892 5584 7898 5636
rect 10870 5584 10876 5636
rect 10928 5624 10934 5636
rect 11241 5627 11299 5633
rect 11241 5624 11253 5627
rect 10928 5596 11253 5624
rect 10928 5584 10934 5596
rect 11241 5593 11253 5596
rect 11287 5593 11299 5627
rect 26694 5624 26700 5636
rect 26655 5596 26700 5624
rect 11241 5587 11299 5593
rect 26694 5584 26700 5596
rect 26752 5584 26758 5636
rect 6546 5556 6552 5568
rect 6507 5528 6552 5556
rect 6546 5516 6552 5528
rect 6604 5516 6610 5568
rect 11974 5516 11980 5568
rect 12032 5556 12038 5568
rect 12805 5559 12863 5565
rect 12805 5556 12817 5559
rect 12032 5528 12817 5556
rect 12032 5516 12038 5528
rect 12805 5525 12817 5528
rect 12851 5525 12863 5559
rect 15378 5556 15384 5568
rect 15339 5528 15384 5556
rect 12805 5519 12863 5525
rect 15378 5516 15384 5528
rect 15436 5516 15442 5568
rect 19242 5556 19248 5568
rect 19203 5528 19248 5556
rect 19242 5516 19248 5528
rect 19300 5516 19306 5568
rect 1104 5466 28888 5488
rect 1104 5414 5982 5466
rect 6034 5414 6046 5466
rect 6098 5414 6110 5466
rect 6162 5414 6174 5466
rect 6226 5414 15982 5466
rect 16034 5414 16046 5466
rect 16098 5414 16110 5466
rect 16162 5414 16174 5466
rect 16226 5414 25982 5466
rect 26034 5414 26046 5466
rect 26098 5414 26110 5466
rect 26162 5414 26174 5466
rect 26226 5414 28888 5466
rect 1104 5392 28888 5414
rect 2406 5352 2412 5364
rect 2367 5324 2412 5352
rect 2406 5312 2412 5324
rect 2464 5312 2470 5364
rect 5169 5355 5227 5361
rect 5169 5321 5181 5355
rect 5215 5352 5227 5355
rect 5442 5352 5448 5364
rect 5215 5324 5448 5352
rect 5215 5321 5227 5324
rect 5169 5315 5227 5321
rect 5442 5312 5448 5324
rect 5500 5312 5506 5364
rect 5810 5352 5816 5364
rect 5771 5324 5816 5352
rect 5810 5312 5816 5324
rect 5868 5312 5874 5364
rect 6638 5352 6644 5364
rect 6599 5324 6644 5352
rect 6638 5312 6644 5324
rect 6696 5312 6702 5364
rect 6825 5355 6883 5361
rect 6825 5321 6837 5355
rect 6871 5352 6883 5355
rect 7374 5352 7380 5364
rect 6871 5324 7380 5352
rect 6871 5321 6883 5324
rect 6825 5315 6883 5321
rect 7374 5312 7380 5324
rect 7432 5312 7438 5364
rect 7834 5352 7840 5364
rect 7795 5324 7840 5352
rect 7834 5312 7840 5324
rect 7892 5312 7898 5364
rect 8294 5312 8300 5364
rect 8352 5352 8358 5364
rect 8389 5355 8447 5361
rect 8389 5352 8401 5355
rect 8352 5324 8401 5352
rect 8352 5312 8358 5324
rect 8389 5321 8401 5324
rect 8435 5321 8447 5355
rect 11330 5352 11336 5364
rect 11291 5324 11336 5352
rect 8389 5315 8447 5321
rect 1581 5287 1639 5293
rect 1581 5253 1593 5287
rect 1627 5284 1639 5287
rect 2774 5284 2780 5296
rect 1627 5256 2780 5284
rect 1627 5253 1639 5256
rect 1581 5247 1639 5253
rect 2774 5244 2780 5256
rect 2832 5244 2838 5296
rect 3142 5284 3148 5296
rect 3103 5256 3148 5284
rect 3142 5244 3148 5256
rect 3200 5244 3206 5296
rect 5537 5287 5595 5293
rect 5537 5253 5549 5287
rect 5583 5284 5595 5287
rect 5718 5284 5724 5296
rect 5583 5256 5724 5284
rect 5583 5253 5595 5256
rect 5537 5247 5595 5253
rect 5718 5244 5724 5256
rect 5776 5244 5782 5296
rect 6656 5216 6684 5312
rect 7285 5219 7343 5225
rect 7285 5216 7297 5219
rect 6656 5188 7297 5216
rect 7285 5185 7297 5188
rect 7331 5185 7343 5219
rect 7285 5179 7343 5185
rect 7377 5219 7435 5225
rect 7377 5185 7389 5219
rect 7423 5216 7435 5219
rect 7466 5216 7472 5228
rect 7423 5188 7472 5216
rect 7423 5185 7435 5188
rect 7377 5179 7435 5185
rect 1397 5151 1455 5157
rect 1397 5117 1409 5151
rect 1443 5148 1455 5151
rect 2501 5151 2559 5157
rect 1443 5120 2084 5148
rect 1443 5117 1455 5120
rect 1397 5111 1455 5117
rect 2056 5024 2084 5120
rect 2501 5117 2513 5151
rect 2547 5117 2559 5151
rect 2501 5111 2559 5117
rect 6273 5151 6331 5157
rect 6273 5117 6285 5151
rect 6319 5148 6331 5151
rect 6546 5148 6552 5160
rect 6319 5120 6552 5148
rect 6319 5117 6331 5120
rect 6273 5111 6331 5117
rect 2516 5080 2544 5111
rect 6546 5108 6552 5120
rect 6604 5148 6610 5160
rect 7392 5148 7420 5179
rect 7466 5176 7472 5188
rect 7524 5176 7530 5228
rect 6604 5120 7420 5148
rect 8404 5148 8432 5315
rect 11330 5312 11336 5324
rect 11388 5312 11394 5364
rect 11698 5352 11704 5364
rect 11659 5324 11704 5352
rect 11698 5312 11704 5324
rect 11756 5312 11762 5364
rect 11974 5352 11980 5364
rect 11935 5324 11980 5352
rect 11974 5312 11980 5324
rect 12032 5312 12038 5364
rect 12897 5355 12955 5361
rect 12897 5321 12909 5355
rect 12943 5352 12955 5355
rect 13262 5352 13268 5364
rect 12943 5324 13268 5352
rect 12943 5321 12955 5324
rect 12897 5315 12955 5321
rect 13262 5312 13268 5324
rect 13320 5312 13326 5364
rect 13446 5312 13452 5364
rect 13504 5352 13510 5364
rect 13633 5355 13691 5361
rect 13633 5352 13645 5355
rect 13504 5324 13645 5352
rect 13504 5312 13510 5324
rect 13633 5321 13645 5324
rect 13679 5352 13691 5355
rect 15933 5355 15991 5361
rect 15933 5352 15945 5355
rect 13679 5324 15945 5352
rect 13679 5321 13691 5324
rect 13633 5315 13691 5321
rect 15933 5321 15945 5324
rect 15979 5321 15991 5355
rect 16574 5352 16580 5364
rect 16535 5324 16580 5352
rect 15933 5315 15991 5321
rect 16574 5312 16580 5324
rect 16632 5312 16638 5364
rect 19702 5352 19708 5364
rect 19663 5324 19708 5352
rect 19702 5312 19708 5324
rect 19760 5312 19766 5364
rect 20162 5352 20168 5364
rect 20123 5324 20168 5352
rect 20162 5312 20168 5324
rect 20220 5312 20226 5364
rect 26510 5312 26516 5364
rect 26568 5352 26574 5364
rect 27341 5355 27399 5361
rect 27341 5352 27353 5355
rect 26568 5324 27353 5352
rect 26568 5312 26574 5324
rect 27341 5321 27353 5324
rect 27387 5321 27399 5355
rect 27341 5315 27399 5321
rect 13170 5284 13176 5296
rect 13131 5256 13176 5284
rect 13170 5244 13176 5256
rect 13228 5244 13234 5296
rect 19429 5287 19487 5293
rect 19429 5253 19441 5287
rect 19475 5284 19487 5287
rect 19610 5284 19616 5296
rect 19475 5256 19616 5284
rect 19475 5253 19487 5256
rect 19429 5247 19487 5253
rect 19610 5244 19616 5256
rect 19668 5244 19674 5296
rect 9309 5219 9367 5225
rect 9309 5185 9321 5219
rect 9355 5216 9367 5219
rect 9950 5216 9956 5228
rect 9355 5188 9956 5216
rect 9355 5185 9367 5188
rect 9309 5179 9367 5185
rect 9950 5176 9956 5188
rect 10008 5176 10014 5228
rect 18138 5176 18144 5228
rect 18196 5216 18202 5228
rect 18877 5219 18935 5225
rect 18877 5216 18889 5219
rect 18196 5188 18889 5216
rect 18196 5176 18202 5188
rect 18877 5185 18889 5188
rect 18923 5185 18935 5219
rect 18877 5179 18935 5185
rect 8757 5151 8815 5157
rect 8757 5148 8769 5151
rect 8404 5120 8769 5148
rect 6604 5108 6610 5120
rect 8757 5117 8769 5120
rect 8803 5117 8815 5151
rect 8757 5111 8815 5117
rect 9674 5108 9680 5160
rect 9732 5148 9738 5160
rect 9769 5151 9827 5157
rect 9769 5148 9781 5151
rect 9732 5120 9781 5148
rect 9732 5108 9738 5120
rect 9769 5117 9781 5120
rect 9815 5117 9827 5151
rect 9769 5111 9827 5117
rect 9861 5151 9919 5157
rect 9861 5117 9873 5151
rect 9907 5148 9919 5151
rect 10226 5148 10232 5160
rect 9907 5120 10232 5148
rect 9907 5117 9919 5120
rect 9861 5111 9919 5117
rect 10226 5108 10232 5120
rect 10284 5108 10290 5160
rect 14550 5148 14556 5160
rect 14511 5120 14556 5148
rect 14550 5108 14556 5120
rect 14608 5108 14614 5160
rect 18693 5151 18751 5157
rect 18693 5117 18705 5151
rect 18739 5148 18751 5151
rect 18782 5148 18788 5160
rect 18739 5120 18788 5148
rect 18739 5117 18751 5120
rect 18693 5111 18751 5117
rect 18782 5108 18788 5120
rect 18840 5148 18846 5160
rect 19242 5148 19248 5160
rect 18840 5120 19248 5148
rect 18840 5108 18846 5120
rect 19242 5108 19248 5120
rect 19300 5108 19306 5160
rect 26418 5148 26424 5160
rect 26379 5120 26424 5148
rect 26418 5108 26424 5120
rect 26476 5148 26482 5160
rect 26973 5151 27031 5157
rect 26973 5148 26985 5151
rect 26476 5120 26985 5148
rect 26476 5108 26482 5120
rect 26973 5117 26985 5120
rect 27019 5117 27031 5151
rect 26973 5111 27031 5117
rect 3142 5080 3148 5092
rect 2516 5052 3148 5080
rect 3142 5040 3148 5052
rect 3200 5040 3206 5092
rect 7190 5080 7196 5092
rect 7151 5052 7196 5080
rect 7190 5040 7196 5052
rect 7248 5040 7254 5092
rect 14461 5083 14519 5089
rect 14461 5049 14473 5083
rect 14507 5080 14519 5083
rect 14820 5083 14878 5089
rect 14820 5080 14832 5083
rect 14507 5052 14832 5080
rect 14507 5049 14519 5052
rect 14461 5043 14519 5049
rect 14820 5049 14832 5052
rect 14866 5080 14878 5083
rect 16298 5080 16304 5092
rect 14866 5052 16304 5080
rect 14866 5049 14878 5052
rect 14820 5043 14878 5049
rect 16298 5040 16304 5052
rect 16356 5040 16362 5092
rect 17865 5083 17923 5089
rect 17865 5049 17877 5083
rect 17911 5080 17923 5083
rect 17911 5052 18460 5080
rect 17911 5049 17923 5052
rect 17865 5043 17923 5049
rect 18432 5024 18460 5052
rect 2038 5012 2044 5024
rect 1999 4984 2044 5012
rect 2038 4972 2044 4984
rect 2096 4972 2102 5024
rect 2682 5012 2688 5024
rect 2643 4984 2688 5012
rect 2682 4972 2688 4984
rect 2740 4972 2746 5024
rect 8294 4972 8300 5024
rect 8352 5012 8358 5024
rect 8573 5015 8631 5021
rect 8573 5012 8585 5015
rect 8352 4984 8585 5012
rect 8352 4972 8358 4984
rect 8573 4981 8585 4984
rect 8619 4981 8631 5015
rect 9398 5012 9404 5024
rect 9359 4984 9404 5012
rect 8573 4975 8631 4981
rect 9398 4972 9404 4984
rect 9456 4972 9462 5024
rect 18322 5012 18328 5024
rect 18283 4984 18328 5012
rect 18322 4972 18328 4984
rect 18380 4972 18386 5024
rect 18414 4972 18420 5024
rect 18472 5012 18478 5024
rect 18785 5015 18843 5021
rect 18785 5012 18797 5015
rect 18472 4984 18797 5012
rect 18472 4972 18478 4984
rect 18785 4981 18797 4984
rect 18831 4981 18843 5015
rect 26602 5012 26608 5024
rect 26563 4984 26608 5012
rect 18785 4975 18843 4981
rect 26602 4972 26608 4984
rect 26660 4972 26666 5024
rect 1104 4922 28888 4944
rect 1104 4870 10982 4922
rect 11034 4870 11046 4922
rect 11098 4870 11110 4922
rect 11162 4870 11174 4922
rect 11226 4870 20982 4922
rect 21034 4870 21046 4922
rect 21098 4870 21110 4922
rect 21162 4870 21174 4922
rect 21226 4870 28888 4922
rect 1104 4848 28888 4870
rect 5997 4811 6055 4817
rect 5997 4777 6009 4811
rect 6043 4808 6055 4811
rect 7098 4808 7104 4820
rect 6043 4780 7104 4808
rect 6043 4777 6055 4780
rect 5997 4771 6055 4777
rect 7098 4768 7104 4780
rect 7156 4768 7162 4820
rect 7374 4808 7380 4820
rect 7335 4780 7380 4808
rect 7374 4768 7380 4780
rect 7432 4768 7438 4820
rect 9493 4811 9551 4817
rect 9493 4777 9505 4811
rect 9539 4808 9551 4811
rect 10226 4808 10232 4820
rect 9539 4780 10232 4808
rect 9539 4777 9551 4780
rect 9493 4771 9551 4777
rect 10226 4768 10232 4780
rect 10284 4768 10290 4820
rect 15930 4808 15936 4820
rect 15891 4780 15936 4808
rect 15930 4768 15936 4780
rect 15988 4768 15994 4820
rect 18782 4808 18788 4820
rect 18743 4780 18788 4808
rect 18782 4768 18788 4780
rect 18840 4768 18846 4820
rect 6454 4740 6460 4752
rect 6415 4712 6460 4740
rect 6454 4700 6460 4712
rect 6512 4700 6518 4752
rect 10134 4700 10140 4752
rect 10192 4740 10198 4752
rect 10778 4740 10784 4752
rect 10192 4712 10784 4740
rect 10192 4700 10198 4712
rect 10778 4700 10784 4712
rect 10836 4740 10842 4752
rect 16390 4749 16396 4752
rect 10934 4743 10992 4749
rect 10934 4740 10946 4743
rect 10836 4712 10946 4740
rect 10836 4700 10842 4712
rect 10934 4709 10946 4712
rect 10980 4709 10992 4743
rect 16384 4740 16396 4749
rect 16351 4712 16396 4740
rect 10934 4703 10992 4709
rect 16384 4703 16396 4712
rect 16448 4740 16454 4752
rect 18138 4740 18144 4752
rect 16448 4712 18144 4740
rect 16390 4700 16396 4703
rect 16448 4700 16454 4712
rect 18138 4700 18144 4712
rect 18196 4740 18202 4752
rect 18325 4743 18383 4749
rect 18325 4740 18337 4743
rect 18196 4712 18337 4740
rect 18196 4700 18202 4712
rect 18325 4709 18337 4712
rect 18371 4709 18383 4743
rect 18325 4703 18383 4709
rect 1397 4675 1455 4681
rect 1397 4641 1409 4675
rect 1443 4672 1455 4675
rect 2406 4672 2412 4684
rect 1443 4644 2412 4672
rect 1443 4641 1455 4644
rect 1397 4635 1455 4641
rect 2406 4632 2412 4644
rect 2464 4632 2470 4684
rect 4062 4672 4068 4684
rect 4023 4644 4068 4672
rect 4062 4632 4068 4644
rect 4120 4632 4126 4684
rect 6362 4672 6368 4684
rect 6323 4644 6368 4672
rect 6362 4632 6368 4644
rect 6420 4632 6426 4684
rect 14550 4632 14556 4684
rect 14608 4672 14614 4684
rect 15838 4672 15844 4684
rect 14608 4644 15844 4672
rect 14608 4632 14614 4644
rect 15838 4632 15844 4644
rect 15896 4672 15902 4684
rect 16117 4675 16175 4681
rect 16117 4672 16129 4675
rect 15896 4644 16129 4672
rect 15896 4632 15902 4644
rect 16117 4641 16129 4644
rect 16163 4672 16175 4675
rect 16666 4672 16672 4684
rect 16163 4644 16672 4672
rect 16163 4641 16175 4644
rect 16117 4635 16175 4641
rect 16666 4632 16672 4644
rect 16724 4632 16730 4684
rect 25314 4672 25320 4684
rect 25275 4644 25320 4672
rect 25314 4632 25320 4644
rect 25372 4632 25378 4684
rect 26513 4675 26571 4681
rect 26513 4641 26525 4675
rect 26559 4672 26571 4675
rect 26786 4672 26792 4684
rect 26559 4644 26792 4672
rect 26559 4641 26571 4644
rect 26513 4635 26571 4641
rect 26786 4632 26792 4644
rect 26844 4632 26850 4684
rect 4341 4607 4399 4613
rect 4341 4573 4353 4607
rect 4387 4604 4399 4607
rect 4522 4604 4528 4616
rect 4387 4576 4528 4604
rect 4387 4573 4399 4576
rect 4341 4567 4399 4573
rect 4522 4564 4528 4576
rect 4580 4564 4586 4616
rect 6546 4564 6552 4616
rect 6604 4604 6610 4616
rect 10686 4604 10692 4616
rect 6604 4576 6649 4604
rect 10647 4576 10692 4604
rect 6604 4564 6610 4576
rect 10686 4564 10692 4576
rect 10744 4564 10750 4616
rect 1578 4468 1584 4480
rect 1539 4440 1584 4468
rect 1578 4428 1584 4440
rect 1636 4428 1642 4480
rect 9950 4428 9956 4480
rect 10008 4468 10014 4480
rect 12069 4471 12127 4477
rect 12069 4468 12081 4471
rect 10008 4440 12081 4468
rect 10008 4428 10014 4440
rect 12069 4437 12081 4440
rect 12115 4468 12127 4471
rect 12434 4468 12440 4480
rect 12115 4440 12440 4468
rect 12115 4437 12127 4440
rect 12069 4431 12127 4437
rect 12434 4428 12440 4440
rect 12492 4428 12498 4480
rect 13814 4428 13820 4480
rect 13872 4468 13878 4480
rect 14550 4468 14556 4480
rect 13872 4440 14556 4468
rect 13872 4428 13878 4440
rect 14550 4428 14556 4440
rect 14608 4428 14614 4480
rect 15565 4471 15623 4477
rect 15565 4437 15577 4471
rect 15611 4468 15623 4471
rect 16298 4468 16304 4480
rect 15611 4440 16304 4468
rect 15611 4437 15623 4440
rect 15565 4431 15623 4437
rect 16298 4428 16304 4440
rect 16356 4468 16362 4480
rect 17497 4471 17555 4477
rect 17497 4468 17509 4471
rect 16356 4440 17509 4468
rect 16356 4428 16362 4440
rect 17497 4437 17509 4440
rect 17543 4437 17555 4471
rect 17497 4431 17555 4437
rect 25501 4471 25559 4477
rect 25501 4437 25513 4471
rect 25547 4468 25559 4471
rect 25774 4468 25780 4480
rect 25547 4440 25780 4468
rect 25547 4437 25559 4440
rect 25501 4431 25559 4437
rect 25774 4428 25780 4440
rect 25832 4428 25838 4480
rect 26694 4468 26700 4480
rect 26655 4440 26700 4468
rect 26694 4428 26700 4440
rect 26752 4428 26758 4480
rect 1104 4378 28888 4400
rect 1104 4326 5982 4378
rect 6034 4326 6046 4378
rect 6098 4326 6110 4378
rect 6162 4326 6174 4378
rect 6226 4326 15982 4378
rect 16034 4326 16046 4378
rect 16098 4326 16110 4378
rect 16162 4326 16174 4378
rect 16226 4326 25982 4378
rect 26034 4326 26046 4378
rect 26098 4326 26110 4378
rect 26162 4326 26174 4378
rect 26226 4326 28888 4378
rect 1104 4304 28888 4326
rect 4062 4264 4068 4276
rect 4023 4236 4068 4264
rect 4062 4224 4068 4236
rect 4120 4224 4126 4276
rect 5721 4267 5779 4273
rect 5721 4233 5733 4267
rect 5767 4264 5779 4267
rect 6546 4264 6552 4276
rect 5767 4236 6552 4264
rect 5767 4233 5779 4236
rect 5721 4227 5779 4233
rect 6546 4224 6552 4236
rect 6604 4224 6610 4276
rect 10778 4264 10784 4276
rect 10739 4236 10784 4264
rect 10778 4224 10784 4236
rect 10836 4224 10842 4276
rect 16209 4267 16267 4273
rect 16209 4233 16221 4267
rect 16255 4264 16267 4267
rect 16390 4264 16396 4276
rect 16255 4236 16396 4264
rect 16255 4233 16267 4236
rect 16209 4227 16267 4233
rect 16390 4224 16396 4236
rect 16448 4224 16454 4276
rect 25314 4264 25320 4276
rect 25275 4236 25320 4264
rect 25314 4224 25320 4236
rect 25372 4224 25378 4276
rect 26786 4224 26792 4276
rect 26844 4264 26850 4276
rect 27341 4267 27399 4273
rect 27341 4264 27353 4267
rect 26844 4236 27353 4264
rect 26844 4224 26850 4236
rect 27341 4233 27353 4236
rect 27387 4233 27399 4267
rect 27341 4227 27399 4233
rect 2406 4196 2412 4208
rect 2367 4168 2412 4196
rect 2406 4156 2412 4168
rect 2464 4156 2470 4208
rect 6362 4196 6368 4208
rect 6323 4168 6368 4196
rect 6362 4156 6368 4168
rect 6420 4156 6426 4208
rect 15838 4156 15844 4208
rect 15896 4196 15902 4208
rect 16485 4199 16543 4205
rect 16485 4196 16497 4199
rect 15896 4168 16497 4196
rect 15896 4156 15902 4168
rect 16485 4165 16497 4168
rect 16531 4165 16543 4199
rect 16485 4159 16543 4165
rect 2041 4131 2099 4137
rect 2041 4128 2053 4131
rect 1412 4100 2053 4128
rect 1412 4069 1440 4100
rect 2041 4097 2053 4100
rect 2087 4128 2099 4131
rect 6089 4131 6147 4137
rect 2087 4100 5764 4128
rect 2087 4097 2099 4100
rect 2041 4091 2099 4097
rect 1397 4063 1455 4069
rect 1397 4029 1409 4063
rect 1443 4029 1455 4063
rect 1397 4023 1455 4029
rect 2501 4063 2559 4069
rect 2501 4029 2513 4063
rect 2547 4060 2559 4063
rect 4614 4060 4620 4072
rect 2547 4032 3188 4060
rect 4575 4032 4620 4060
rect 2547 4029 2559 4032
rect 2501 4023 2559 4029
rect 3160 3936 3188 4032
rect 4614 4020 4620 4032
rect 4672 4060 4678 4072
rect 4709 4063 4767 4069
rect 4709 4060 4721 4063
rect 4672 4032 4721 4060
rect 4672 4020 4678 4032
rect 4709 4029 4721 4032
rect 4755 4029 4767 4063
rect 4709 4023 4767 4029
rect 4985 4063 5043 4069
rect 4985 4029 4997 4063
rect 5031 4060 5043 4063
rect 5626 4060 5632 4072
rect 5031 4032 5632 4060
rect 5031 4029 5043 4032
rect 4985 4023 5043 4029
rect 5626 4020 5632 4032
rect 5684 4020 5690 4072
rect 5736 4060 5764 4100
rect 6089 4097 6101 4131
rect 6135 4128 6147 4131
rect 6454 4128 6460 4140
rect 6135 4100 6460 4128
rect 6135 4097 6147 4100
rect 6089 4091 6147 4097
rect 6454 4088 6460 4100
rect 6512 4088 6518 4140
rect 10686 4088 10692 4140
rect 10744 4128 10750 4140
rect 11057 4131 11115 4137
rect 11057 4128 11069 4131
rect 10744 4100 11069 4128
rect 10744 4088 10750 4100
rect 11057 4097 11069 4100
rect 11103 4097 11115 4131
rect 11057 4091 11115 4097
rect 8110 4060 8116 4072
rect 5736 4032 8116 4060
rect 8110 4020 8116 4032
rect 8168 4020 8174 4072
rect 9769 4063 9827 4069
rect 9769 4029 9781 4063
rect 9815 4060 9827 4063
rect 10413 4063 10471 4069
rect 10413 4060 10425 4063
rect 9815 4032 10425 4060
rect 9815 4029 9827 4032
rect 9769 4023 9827 4029
rect 10413 4029 10425 4032
rect 10459 4060 10471 4063
rect 10870 4060 10876 4072
rect 10459 4032 10876 4060
rect 10459 4029 10471 4032
rect 10413 4023 10471 4029
rect 10870 4020 10876 4032
rect 10928 4020 10934 4072
rect 26418 4060 26424 4072
rect 26379 4032 26424 4060
rect 26418 4020 26424 4032
rect 26476 4060 26482 4072
rect 26973 4063 27031 4069
rect 26973 4060 26985 4063
rect 26476 4032 26985 4060
rect 26476 4020 26482 4032
rect 26973 4029 26985 4032
rect 27019 4029 27031 4063
rect 26973 4023 27031 4029
rect 10778 3992 10784 4004
rect 9968 3964 10784 3992
rect 1578 3924 1584 3936
rect 1539 3896 1584 3924
rect 1578 3884 1584 3896
rect 1636 3884 1642 3936
rect 2685 3927 2743 3933
rect 2685 3893 2697 3927
rect 2731 3924 2743 3927
rect 2866 3924 2872 3936
rect 2731 3896 2872 3924
rect 2731 3893 2743 3896
rect 2685 3887 2743 3893
rect 2866 3884 2872 3896
rect 2924 3884 2930 3936
rect 3142 3924 3148 3936
rect 3103 3896 3148 3924
rect 3142 3884 3148 3896
rect 3200 3884 3206 3936
rect 9968 3933 9996 3964
rect 10778 3952 10784 3964
rect 10836 3952 10842 4004
rect 9953 3927 10011 3933
rect 9953 3893 9965 3927
rect 9999 3893 10011 3927
rect 26602 3924 26608 3936
rect 26563 3896 26608 3924
rect 9953 3887 10011 3893
rect 26602 3884 26608 3896
rect 26660 3884 26666 3936
rect 1104 3834 28888 3856
rect 1104 3782 10982 3834
rect 11034 3782 11046 3834
rect 11098 3782 11110 3834
rect 11162 3782 11174 3834
rect 11226 3782 20982 3834
rect 21034 3782 21046 3834
rect 21098 3782 21110 3834
rect 21162 3782 21174 3834
rect 21226 3782 28888 3834
rect 1104 3760 28888 3782
rect 1946 3720 1952 3732
rect 1907 3692 1952 3720
rect 1946 3680 1952 3692
rect 2004 3680 2010 3732
rect 6546 3680 6552 3732
rect 6604 3720 6610 3732
rect 6733 3723 6791 3729
rect 6733 3720 6745 3723
rect 6604 3692 6745 3720
rect 6604 3680 6610 3692
rect 6733 3689 6745 3692
rect 6779 3689 6791 3723
rect 6733 3683 6791 3689
rect 7282 3680 7288 3732
rect 7340 3720 7346 3732
rect 7377 3723 7435 3729
rect 7377 3720 7389 3723
rect 7340 3692 7389 3720
rect 7340 3680 7346 3692
rect 7377 3689 7389 3692
rect 7423 3720 7435 3723
rect 8202 3720 8208 3732
rect 7423 3692 8208 3720
rect 7423 3689 7435 3692
rect 7377 3683 7435 3689
rect 8202 3680 8208 3692
rect 8260 3680 8266 3732
rect 1397 3587 1455 3593
rect 1397 3553 1409 3587
rect 1443 3584 1455 3587
rect 1964 3584 1992 3680
rect 5534 3612 5540 3664
rect 5592 3661 5598 3664
rect 5592 3655 5656 3661
rect 5592 3621 5610 3655
rect 5644 3621 5656 3655
rect 10686 3652 10692 3664
rect 5592 3615 5656 3621
rect 9968 3624 10692 3652
rect 5592 3612 5598 3615
rect 2498 3584 2504 3596
rect 1443 3556 1992 3584
rect 2459 3556 2504 3584
rect 1443 3553 1455 3556
rect 1397 3547 1455 3553
rect 2498 3544 2504 3556
rect 2556 3544 2562 3596
rect 8205 3587 8263 3593
rect 8205 3553 8217 3587
rect 8251 3584 8263 3587
rect 8662 3584 8668 3596
rect 8251 3556 8668 3584
rect 8251 3553 8263 3556
rect 8205 3547 8263 3553
rect 8662 3544 8668 3556
rect 8720 3544 8726 3596
rect 9674 3544 9680 3596
rect 9732 3584 9738 3596
rect 9968 3593 9996 3624
rect 10686 3612 10692 3624
rect 10744 3612 10750 3664
rect 12434 3612 12440 3664
rect 12492 3652 12498 3664
rect 12682 3655 12740 3661
rect 12682 3652 12694 3655
rect 12492 3624 12694 3652
rect 12492 3612 12498 3624
rect 12682 3621 12694 3624
rect 12728 3621 12740 3655
rect 12682 3615 12740 3621
rect 9953 3587 10011 3593
rect 9953 3584 9965 3587
rect 9732 3556 9965 3584
rect 9732 3544 9738 3556
rect 9953 3553 9965 3556
rect 9999 3553 10011 3587
rect 10209 3587 10267 3593
rect 10209 3584 10221 3587
rect 9953 3547 10011 3553
rect 10060 3556 10221 3584
rect 5350 3516 5356 3528
rect 5311 3488 5356 3516
rect 5350 3476 5356 3488
rect 5408 3476 5414 3528
rect 10060 3516 10088 3556
rect 10209 3553 10221 3556
rect 10255 3553 10267 3587
rect 10209 3547 10267 3553
rect 18138 3544 18144 3596
rect 18196 3584 18202 3596
rect 26513 3587 26571 3593
rect 26513 3584 26525 3587
rect 18196 3556 26525 3584
rect 18196 3544 18202 3556
rect 26513 3553 26525 3556
rect 26559 3584 26571 3587
rect 27338 3584 27344 3596
rect 26559 3556 27344 3584
rect 26559 3553 26571 3556
rect 26513 3547 26571 3553
rect 27338 3544 27344 3556
rect 27396 3544 27402 3596
rect 9968 3488 10088 3516
rect 12437 3519 12495 3525
rect 9968 3460 9996 3488
rect 12437 3485 12449 3519
rect 12483 3485 12495 3519
rect 12437 3479 12495 3485
rect 9950 3408 9956 3460
rect 10008 3408 10014 3460
rect 1578 3380 1584 3392
rect 1539 3352 1584 3380
rect 1578 3340 1584 3352
rect 1636 3340 1642 3392
rect 2682 3380 2688 3392
rect 2643 3352 2688 3380
rect 2682 3340 2688 3352
rect 2740 3340 2746 3392
rect 8389 3383 8447 3389
rect 8389 3349 8401 3383
rect 8435 3380 8447 3383
rect 9766 3380 9772 3392
rect 8435 3352 9772 3380
rect 8435 3349 8447 3352
rect 8389 3343 8447 3349
rect 9766 3340 9772 3352
rect 9824 3340 9830 3392
rect 11330 3380 11336 3392
rect 11291 3352 11336 3380
rect 11330 3340 11336 3352
rect 11388 3340 11394 3392
rect 12452 3380 12480 3479
rect 13722 3448 13728 3460
rect 13648 3420 13728 3448
rect 12618 3380 12624 3392
rect 12452 3352 12624 3380
rect 12618 3340 12624 3352
rect 12676 3380 12682 3392
rect 13648 3380 13676 3420
rect 13722 3408 13728 3420
rect 13780 3408 13786 3460
rect 13814 3380 13820 3392
rect 12676 3352 13676 3380
rect 13775 3352 13820 3380
rect 12676 3340 12682 3352
rect 13814 3340 13820 3352
rect 13872 3340 13878 3392
rect 26694 3380 26700 3392
rect 26655 3352 26700 3380
rect 26694 3340 26700 3352
rect 26752 3340 26758 3392
rect 1104 3290 28888 3312
rect 1104 3238 5982 3290
rect 6034 3238 6046 3290
rect 6098 3238 6110 3290
rect 6162 3238 6174 3290
rect 6226 3238 15982 3290
rect 16034 3238 16046 3290
rect 16098 3238 16110 3290
rect 16162 3238 16174 3290
rect 16226 3238 25982 3290
rect 26034 3238 26046 3290
rect 26098 3238 26110 3290
rect 26162 3238 26174 3290
rect 26226 3238 28888 3290
rect 1104 3216 28888 3238
rect 2038 3176 2044 3188
rect 1999 3148 2044 3176
rect 2038 3136 2044 3148
rect 2096 3136 2102 3188
rect 2498 3176 2504 3188
rect 2459 3148 2504 3176
rect 2498 3136 2504 3148
rect 2556 3136 2562 3188
rect 4525 3179 4583 3185
rect 4525 3145 4537 3179
rect 4571 3176 4583 3179
rect 4706 3176 4712 3188
rect 4571 3148 4712 3176
rect 4571 3145 4583 3148
rect 4525 3139 4583 3145
rect 4706 3136 4712 3148
rect 4764 3136 4770 3188
rect 8662 3176 8668 3188
rect 8623 3148 8668 3176
rect 8662 3136 8668 3148
rect 8720 3176 8726 3188
rect 9217 3179 9275 3185
rect 9217 3176 9229 3179
rect 8720 3148 9229 3176
rect 8720 3136 8726 3148
rect 9217 3145 9229 3148
rect 9263 3145 9275 3179
rect 9674 3176 9680 3188
rect 9635 3148 9680 3176
rect 9217 3139 9275 3145
rect 9674 3136 9680 3148
rect 9732 3136 9738 3188
rect 9950 3176 9956 3188
rect 9911 3148 9956 3176
rect 9950 3136 9956 3148
rect 10008 3136 10014 3188
rect 10781 3179 10839 3185
rect 10781 3145 10793 3179
rect 10827 3176 10839 3179
rect 11330 3176 11336 3188
rect 10827 3148 11336 3176
rect 10827 3145 10839 3148
rect 10781 3139 10839 3145
rect 4062 3068 4068 3120
rect 4120 3108 4126 3120
rect 4801 3111 4859 3117
rect 4801 3108 4813 3111
rect 4120 3080 4813 3108
rect 4120 3068 4126 3080
rect 4801 3077 4813 3080
rect 4847 3077 4859 3111
rect 4801 3071 4859 3077
rect 4154 3040 4160 3052
rect 3344 3012 4160 3040
rect 1397 2975 1455 2981
rect 1397 2941 1409 2975
rect 1443 2972 1455 2975
rect 2038 2972 2044 2984
rect 1443 2944 2044 2972
rect 1443 2941 1455 2944
rect 1397 2935 1455 2941
rect 2038 2932 2044 2944
rect 2096 2932 2102 2984
rect 3344 2981 3372 3012
rect 4154 3000 4160 3012
rect 4212 3000 4218 3052
rect 5350 3000 5356 3052
rect 5408 3040 5414 3052
rect 5813 3043 5871 3049
rect 5813 3040 5825 3043
rect 5408 3012 5825 3040
rect 5408 3000 5414 3012
rect 5813 3009 5825 3012
rect 5859 3040 5871 3043
rect 6914 3040 6920 3052
rect 5859 3012 6920 3040
rect 5859 3009 5871 3012
rect 5813 3003 5871 3009
rect 6914 3000 6920 3012
rect 6972 3040 6978 3052
rect 7282 3040 7288 3052
rect 6972 3012 7288 3040
rect 6972 3000 6978 3012
rect 7282 3000 7288 3012
rect 7340 3000 7346 3052
rect 3329 2975 3387 2981
rect 3329 2941 3341 2975
rect 3375 2941 3387 2975
rect 3329 2935 3387 2941
rect 4617 2975 4675 2981
rect 4617 2941 4629 2975
rect 4663 2972 4675 2975
rect 4706 2972 4712 2984
rect 4663 2944 4712 2972
rect 4663 2941 4675 2944
rect 4617 2935 4675 2941
rect 4706 2932 4712 2944
rect 4764 2932 4770 2984
rect 10137 2975 10195 2981
rect 10137 2941 10149 2975
rect 10183 2972 10195 2975
rect 10796 2972 10824 3139
rect 11330 3136 11336 3148
rect 11388 3136 11394 3188
rect 11882 3176 11888 3188
rect 11843 3148 11888 3176
rect 11882 3136 11888 3148
rect 11940 3136 11946 3188
rect 12434 3136 12440 3188
rect 12492 3176 12498 3188
rect 12621 3179 12679 3185
rect 12621 3176 12633 3179
rect 12492 3148 12633 3176
rect 12492 3136 12498 3148
rect 12621 3145 12633 3148
rect 12667 3145 12679 3179
rect 27338 3176 27344 3188
rect 27299 3148 27344 3176
rect 12621 3139 12679 3145
rect 27338 3136 27344 3148
rect 27396 3136 27402 3188
rect 11425 3111 11483 3117
rect 11425 3077 11437 3111
rect 11471 3108 11483 3111
rect 12802 3108 12808 3120
rect 11471 3080 12808 3108
rect 11471 3077 11483 3080
rect 11425 3071 11483 3077
rect 12802 3068 12808 3080
rect 12860 3068 12866 3120
rect 10183 2944 10824 2972
rect 11241 2975 11299 2981
rect 10183 2941 10195 2944
rect 10137 2935 10195 2941
rect 11241 2941 11253 2975
rect 11287 2972 11299 2975
rect 11882 2972 11888 2984
rect 11287 2944 11888 2972
rect 11287 2941 11299 2944
rect 11241 2935 11299 2941
rect 11882 2932 11888 2944
rect 11940 2932 11946 2984
rect 13170 2972 13176 2984
rect 13131 2944 13176 2972
rect 13170 2932 13176 2944
rect 13228 2972 13234 2984
rect 13725 2975 13783 2981
rect 13725 2972 13737 2975
rect 13228 2944 13737 2972
rect 13228 2932 13234 2944
rect 13725 2941 13737 2944
rect 13771 2941 13783 2975
rect 13725 2935 13783 2941
rect 13998 2932 14004 2984
rect 14056 2972 14062 2984
rect 14277 2975 14335 2981
rect 14277 2972 14289 2975
rect 14056 2944 14289 2972
rect 14056 2932 14062 2944
rect 14277 2941 14289 2944
rect 14323 2972 14335 2975
rect 14829 2975 14887 2981
rect 14829 2972 14841 2975
rect 14323 2944 14841 2972
rect 14323 2941 14335 2944
rect 14277 2935 14335 2941
rect 14829 2941 14841 2944
rect 14875 2941 14887 2975
rect 19058 2972 19064 2984
rect 18971 2944 19064 2972
rect 14829 2935 14887 2941
rect 19058 2932 19064 2944
rect 19116 2972 19122 2984
rect 19613 2975 19671 2981
rect 19613 2972 19625 2975
rect 19116 2944 19625 2972
rect 19116 2932 19122 2944
rect 19613 2941 19625 2944
rect 19659 2941 19671 2975
rect 25314 2972 25320 2984
rect 25275 2944 25320 2972
rect 19613 2935 19671 2941
rect 25314 2932 25320 2944
rect 25372 2972 25378 2984
rect 25869 2975 25927 2981
rect 25869 2972 25881 2975
rect 25372 2944 25881 2972
rect 25372 2932 25378 2944
rect 25869 2941 25881 2944
rect 25915 2941 25927 2975
rect 25869 2935 25927 2941
rect 26326 2932 26332 2984
rect 26384 2972 26390 2984
rect 26421 2975 26479 2981
rect 26421 2972 26433 2975
rect 26384 2944 26433 2972
rect 26384 2932 26390 2944
rect 26421 2941 26433 2944
rect 26467 2972 26479 2975
rect 26973 2975 27031 2981
rect 26973 2972 26985 2975
rect 26467 2944 26985 2972
rect 26467 2941 26479 2944
rect 26421 2935 26479 2941
rect 26973 2941 26985 2944
rect 27019 2941 27031 2975
rect 26973 2935 27031 2941
rect 3510 2864 3516 2916
rect 3568 2904 3574 2916
rect 3605 2907 3663 2913
rect 3605 2904 3617 2907
rect 3568 2876 3617 2904
rect 3568 2864 3574 2876
rect 3605 2873 3617 2876
rect 3651 2873 3663 2907
rect 3605 2867 3663 2873
rect 5445 2907 5503 2913
rect 5445 2873 5457 2907
rect 5491 2904 5503 2907
rect 5534 2904 5540 2916
rect 5491 2876 5540 2904
rect 5491 2873 5503 2876
rect 5445 2867 5503 2873
rect 5534 2864 5540 2876
rect 5592 2904 5598 2916
rect 6638 2904 6644 2916
rect 5592 2876 6644 2904
rect 5592 2864 5598 2876
rect 6638 2864 6644 2876
rect 6696 2864 6702 2916
rect 7098 2864 7104 2916
rect 7156 2904 7162 2916
rect 7193 2907 7251 2913
rect 7193 2904 7205 2907
rect 7156 2876 7205 2904
rect 7156 2864 7162 2876
rect 7193 2873 7205 2876
rect 7239 2904 7251 2907
rect 7530 2907 7588 2913
rect 7530 2904 7542 2907
rect 7239 2876 7542 2904
rect 7239 2873 7251 2876
rect 7193 2867 7251 2873
rect 7530 2873 7542 2876
rect 7576 2873 7588 2907
rect 7530 2867 7588 2873
rect 1578 2836 1584 2848
rect 1539 2808 1584 2836
rect 1578 2796 1584 2808
rect 1636 2796 1642 2848
rect 10321 2839 10379 2845
rect 10321 2805 10333 2839
rect 10367 2836 10379 2839
rect 11698 2836 11704 2848
rect 10367 2808 11704 2836
rect 10367 2805 10379 2808
rect 10321 2799 10379 2805
rect 11698 2796 11704 2808
rect 11756 2796 11762 2848
rect 12618 2796 12624 2848
rect 12676 2836 12682 2848
rect 12989 2839 13047 2845
rect 12989 2836 13001 2839
rect 12676 2808 13001 2836
rect 12676 2796 12682 2808
rect 12989 2805 13001 2808
rect 13035 2805 13047 2839
rect 13354 2836 13360 2848
rect 13315 2808 13360 2836
rect 12989 2799 13047 2805
rect 13354 2796 13360 2808
rect 13412 2796 13418 2848
rect 13906 2796 13912 2848
rect 13964 2836 13970 2848
rect 14461 2839 14519 2845
rect 14461 2836 14473 2839
rect 13964 2808 14473 2836
rect 13964 2796 13970 2808
rect 14461 2805 14473 2808
rect 14507 2805 14519 2839
rect 14461 2799 14519 2805
rect 19150 2796 19156 2848
rect 19208 2836 19214 2848
rect 19245 2839 19303 2845
rect 19245 2836 19257 2839
rect 19208 2808 19257 2836
rect 19208 2796 19214 2808
rect 19245 2805 19257 2808
rect 19291 2805 19303 2839
rect 25498 2836 25504 2848
rect 25459 2808 25504 2836
rect 19245 2799 19303 2805
rect 25498 2796 25504 2808
rect 25556 2796 25562 2848
rect 26602 2836 26608 2848
rect 26563 2808 26608 2836
rect 26602 2796 26608 2808
rect 26660 2796 26666 2848
rect 1104 2746 28888 2768
rect 1104 2694 10982 2746
rect 11034 2694 11046 2746
rect 11098 2694 11110 2746
rect 11162 2694 11174 2746
rect 11226 2694 20982 2746
rect 21034 2694 21046 2746
rect 21098 2694 21110 2746
rect 21162 2694 21174 2746
rect 21226 2694 28888 2746
rect 1104 2672 28888 2694
rect 3513 2635 3571 2641
rect 3513 2601 3525 2635
rect 3559 2632 3571 2635
rect 3602 2632 3608 2644
rect 3559 2604 3608 2632
rect 3559 2601 3571 2604
rect 3513 2595 3571 2601
rect 2958 2564 2964 2576
rect 2919 2536 2964 2564
rect 2958 2524 2964 2536
rect 3016 2524 3022 2576
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2496 1455 2499
rect 1670 2496 1676 2508
rect 1443 2468 1676 2496
rect 1443 2465 1455 2468
rect 1397 2459 1455 2465
rect 1670 2456 1676 2468
rect 1728 2496 1734 2508
rect 2133 2499 2191 2505
rect 2133 2496 2145 2499
rect 1728 2468 2145 2496
rect 1728 2456 1734 2468
rect 2133 2465 2145 2468
rect 2179 2465 2191 2499
rect 2133 2459 2191 2465
rect 2685 2499 2743 2505
rect 2685 2465 2697 2499
rect 2731 2496 2743 2499
rect 3528 2496 3556 2595
rect 3602 2592 3608 2604
rect 3660 2592 3666 2644
rect 4890 2632 4896 2644
rect 4851 2604 4896 2632
rect 4890 2592 4896 2604
rect 4948 2592 4954 2644
rect 8202 2592 8208 2644
rect 8260 2632 8266 2644
rect 9125 2635 9183 2641
rect 9125 2632 9137 2635
rect 8260 2604 9137 2632
rect 8260 2592 8266 2604
rect 9125 2601 9137 2604
rect 9171 2632 9183 2635
rect 9674 2632 9680 2644
rect 9171 2604 9680 2632
rect 9171 2601 9183 2604
rect 9125 2595 9183 2601
rect 9674 2592 9680 2604
rect 9732 2592 9738 2644
rect 10870 2592 10876 2644
rect 10928 2632 10934 2644
rect 11149 2635 11207 2641
rect 11149 2632 11161 2635
rect 10928 2604 11161 2632
rect 10928 2592 10934 2604
rect 11149 2601 11161 2604
rect 11195 2601 11207 2635
rect 12434 2632 12440 2644
rect 12395 2604 12440 2632
rect 11149 2595 11207 2601
rect 12434 2592 12440 2604
rect 12492 2592 12498 2644
rect 13998 2632 14004 2644
rect 13959 2604 14004 2632
rect 13998 2592 14004 2604
rect 14056 2592 14062 2644
rect 17218 2592 17224 2644
rect 17276 2632 17282 2644
rect 17313 2635 17371 2641
rect 17313 2632 17325 2635
rect 17276 2604 17325 2632
rect 17276 2592 17282 2604
rect 17313 2601 17325 2604
rect 17359 2601 17371 2635
rect 25866 2632 25872 2644
rect 25827 2604 25872 2632
rect 17313 2595 17371 2601
rect 25866 2592 25872 2604
rect 25924 2592 25930 2644
rect 2731 2468 3556 2496
rect 4065 2499 4123 2505
rect 2731 2465 2743 2468
rect 2685 2459 2743 2465
rect 4065 2465 4077 2499
rect 4111 2496 4123 2499
rect 4908 2496 4936 2592
rect 6733 2567 6791 2573
rect 6733 2533 6745 2567
rect 6779 2564 6791 2567
rect 7098 2564 7104 2576
rect 6779 2536 7104 2564
rect 6779 2533 6791 2536
rect 6733 2527 6791 2533
rect 7098 2524 7104 2536
rect 7156 2573 7162 2576
rect 7156 2567 7220 2573
rect 7156 2533 7174 2567
rect 7208 2564 7220 2567
rect 9493 2567 9551 2573
rect 9493 2564 9505 2567
rect 7208 2536 9505 2564
rect 7208 2533 7220 2536
rect 7156 2527 7220 2533
rect 9493 2533 9505 2536
rect 9539 2564 9551 2567
rect 9950 2564 9956 2576
rect 9539 2536 9956 2564
rect 9539 2533 9551 2536
rect 9493 2527 9551 2533
rect 7156 2524 7162 2527
rect 9950 2524 9956 2536
rect 10008 2573 10014 2576
rect 10008 2567 10072 2573
rect 10008 2533 10026 2567
rect 10060 2533 10072 2567
rect 12452 2564 12480 2592
rect 12866 2567 12924 2573
rect 12866 2564 12878 2567
rect 12452 2536 12878 2564
rect 10008 2527 10072 2533
rect 12866 2533 12878 2536
rect 12912 2533 12924 2567
rect 12866 2527 12924 2533
rect 10008 2524 10014 2527
rect 4111 2468 4936 2496
rect 12069 2499 12127 2505
rect 4111 2465 4123 2468
rect 4065 2459 4123 2465
rect 12069 2465 12081 2499
rect 12115 2496 12127 2499
rect 12618 2496 12624 2508
rect 12115 2468 12624 2496
rect 12115 2465 12127 2468
rect 12069 2459 12127 2465
rect 12618 2456 12624 2468
rect 12676 2456 12682 2508
rect 15473 2499 15531 2505
rect 15473 2465 15485 2499
rect 15519 2496 15531 2499
rect 15562 2496 15568 2508
rect 15519 2468 15568 2496
rect 15519 2465 15531 2468
rect 15473 2459 15531 2465
rect 15562 2456 15568 2468
rect 15620 2496 15626 2508
rect 16025 2499 16083 2505
rect 16025 2496 16037 2499
rect 15620 2468 16037 2496
rect 15620 2456 15626 2468
rect 16025 2465 16037 2468
rect 16071 2465 16083 2499
rect 16025 2459 16083 2465
rect 16761 2499 16819 2505
rect 16761 2465 16773 2499
rect 16807 2496 16819 2499
rect 17236 2496 17264 2592
rect 16807 2468 17264 2496
rect 16807 2465 16819 2468
rect 16761 2459 16819 2465
rect 18874 2456 18880 2508
rect 18932 2496 18938 2508
rect 19061 2499 19119 2505
rect 19061 2496 19073 2499
rect 18932 2468 19073 2496
rect 18932 2456 18938 2468
rect 19061 2465 19073 2468
rect 19107 2496 19119 2499
rect 19613 2499 19671 2505
rect 19613 2496 19625 2499
rect 19107 2468 19625 2496
rect 19107 2465 19119 2468
rect 19061 2459 19119 2465
rect 19613 2465 19625 2468
rect 19659 2465 19671 2499
rect 24394 2496 24400 2508
rect 24355 2468 24400 2496
rect 19613 2459 19671 2465
rect 24394 2456 24400 2468
rect 24452 2496 24458 2508
rect 24949 2499 25007 2505
rect 24949 2496 24961 2499
rect 24452 2468 24961 2496
rect 24452 2456 24458 2468
rect 24949 2465 24961 2468
rect 24995 2465 25007 2499
rect 26878 2496 26884 2508
rect 26839 2468 26884 2496
rect 24949 2459 25007 2465
rect 26878 2456 26884 2468
rect 26936 2496 26942 2508
rect 27433 2499 27491 2505
rect 27433 2496 27445 2499
rect 26936 2468 27445 2496
rect 26936 2456 26942 2468
rect 27433 2465 27445 2468
rect 27479 2465 27491 2499
rect 27433 2459 27491 2465
rect 1486 2388 1492 2440
rect 1544 2428 1550 2440
rect 1581 2431 1639 2437
rect 1581 2428 1593 2431
rect 1544 2400 1593 2428
rect 1544 2388 1550 2400
rect 1581 2397 1593 2400
rect 1627 2397 1639 2431
rect 1581 2391 1639 2397
rect 4249 2431 4307 2437
rect 4249 2397 4261 2431
rect 4295 2397 4307 2431
rect 4249 2391 4307 2397
rect 6365 2431 6423 2437
rect 6365 2397 6377 2431
rect 6411 2428 6423 2431
rect 6914 2428 6920 2440
rect 6411 2400 6920 2428
rect 6411 2397 6423 2400
rect 6365 2391 6423 2397
rect 2498 2320 2504 2372
rect 2556 2360 2562 2372
rect 4264 2360 4292 2391
rect 6914 2388 6920 2400
rect 6972 2428 6978 2440
rect 6972 2400 7017 2428
rect 6972 2388 6978 2400
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 9769 2431 9827 2437
rect 9769 2428 9781 2431
rect 9732 2400 9781 2428
rect 9732 2388 9738 2400
rect 9769 2397 9781 2400
rect 9815 2397 9827 2431
rect 9769 2391 9827 2397
rect 19242 2360 19248 2372
rect 2556 2332 4292 2360
rect 19203 2332 19248 2360
rect 2556 2320 2562 2332
rect 19242 2320 19248 2332
rect 19300 2320 19306 2372
rect 24581 2363 24639 2369
rect 24581 2329 24593 2363
rect 24627 2360 24639 2363
rect 26326 2360 26332 2372
rect 24627 2332 26332 2360
rect 24627 2329 24639 2332
rect 24581 2323 24639 2329
rect 26326 2320 26332 2332
rect 26384 2320 26390 2372
rect 7650 2252 7656 2304
rect 7708 2292 7714 2304
rect 8294 2292 8300 2304
rect 7708 2264 8300 2292
rect 7708 2252 7714 2264
rect 8294 2252 8300 2264
rect 8352 2252 8358 2304
rect 15654 2292 15660 2304
rect 15615 2264 15660 2292
rect 15654 2252 15660 2264
rect 15712 2252 15718 2304
rect 16945 2295 17003 2301
rect 16945 2261 16957 2295
rect 16991 2292 17003 2295
rect 17862 2292 17868 2304
rect 16991 2264 17868 2292
rect 16991 2261 17003 2264
rect 16945 2255 17003 2261
rect 17862 2252 17868 2264
rect 17920 2252 17926 2304
rect 27062 2292 27068 2304
rect 27023 2264 27068 2292
rect 27062 2252 27068 2264
rect 27120 2252 27126 2304
rect 1104 2202 28888 2224
rect 1104 2150 5982 2202
rect 6034 2150 6046 2202
rect 6098 2150 6110 2202
rect 6162 2150 6174 2202
rect 6226 2150 15982 2202
rect 16034 2150 16046 2202
rect 16098 2150 16110 2202
rect 16162 2150 16174 2202
rect 16226 2150 25982 2202
rect 26034 2150 26046 2202
rect 26098 2150 26110 2202
rect 26162 2150 26174 2202
rect 26226 2150 28888 2202
rect 1104 2128 28888 2150
rect 15930 1980 15936 2032
rect 15988 2020 15994 2032
rect 16482 2020 16488 2032
rect 15988 1992 16488 2020
rect 15988 1980 15994 1992
rect 16482 1980 16488 1992
rect 16540 1980 16546 2032
rect 8662 552 8668 604
rect 8720 592 8726 604
rect 10594 592 10600 604
rect 8720 564 10600 592
rect 8720 552 8726 564
rect 10594 552 10600 564
rect 10652 552 10658 604
<< via1 >>
rect 3148 22176 3200 22228
rect 9404 22176 9456 22228
rect 2964 22108 3016 22160
rect 15660 22108 15712 22160
rect 5982 21734 6034 21786
rect 6046 21734 6098 21786
rect 6110 21734 6162 21786
rect 6174 21734 6226 21786
rect 15982 21734 16034 21786
rect 16046 21734 16098 21786
rect 16110 21734 16162 21786
rect 16174 21734 16226 21786
rect 25982 21734 26034 21786
rect 26046 21734 26098 21786
rect 26110 21734 26162 21786
rect 26174 21734 26226 21786
rect 3884 21632 3936 21684
rect 6920 21632 6972 21684
rect 10982 21190 11034 21242
rect 11046 21190 11098 21242
rect 11110 21190 11162 21242
rect 11174 21190 11226 21242
rect 20982 21190 21034 21242
rect 21046 21190 21098 21242
rect 21110 21190 21162 21242
rect 21174 21190 21226 21242
rect 3516 20816 3568 20868
rect 10784 20816 10836 20868
rect 11520 20816 11572 20868
rect 25780 20816 25832 20868
rect 8944 20748 8996 20800
rect 25412 20748 25464 20800
rect 5982 20646 6034 20698
rect 6046 20646 6098 20698
rect 6110 20646 6162 20698
rect 6174 20646 6226 20698
rect 15982 20646 16034 20698
rect 16046 20646 16098 20698
rect 16110 20646 16162 20698
rect 16174 20646 16226 20698
rect 25982 20646 26034 20698
rect 26046 20646 26098 20698
rect 26110 20646 26162 20698
rect 26174 20646 26226 20698
rect 5172 20544 5224 20596
rect 6736 20544 6788 20596
rect 8208 20544 8260 20596
rect 11336 20544 11388 20596
rect 18236 20587 18288 20596
rect 18236 20553 18245 20587
rect 18245 20553 18279 20587
rect 18279 20553 18288 20587
rect 18236 20544 18288 20553
rect 16672 20519 16724 20528
rect 16672 20485 16681 20519
rect 16681 20485 16715 20519
rect 16715 20485 16724 20519
rect 16672 20476 16724 20485
rect 25780 20519 25832 20528
rect 25780 20485 25789 20519
rect 25789 20485 25823 20519
rect 25823 20485 25832 20519
rect 25780 20476 25832 20485
rect 7472 20315 7524 20324
rect 7472 20281 7481 20315
rect 7481 20281 7515 20315
rect 7515 20281 7524 20315
rect 7472 20272 7524 20281
rect 5356 20247 5408 20256
rect 5356 20213 5365 20247
rect 5365 20213 5399 20247
rect 5399 20213 5408 20247
rect 5356 20204 5408 20213
rect 8576 20247 8628 20256
rect 8576 20213 8585 20247
rect 8585 20213 8619 20247
rect 8619 20213 8628 20247
rect 8576 20204 8628 20213
rect 14280 20247 14332 20256
rect 14280 20213 14289 20247
rect 14289 20213 14323 20247
rect 14323 20213 14332 20247
rect 14280 20204 14332 20213
rect 15568 20247 15620 20256
rect 15568 20213 15577 20247
rect 15577 20213 15611 20247
rect 15611 20213 15620 20247
rect 15568 20204 15620 20213
rect 19984 20383 20036 20392
rect 16396 20204 16448 20256
rect 17040 20247 17092 20256
rect 17040 20213 17049 20247
rect 17049 20213 17083 20247
rect 17083 20213 17092 20247
rect 17040 20204 17092 20213
rect 19984 20349 19993 20383
rect 19993 20349 20027 20383
rect 20027 20349 20036 20383
rect 19984 20340 20036 20349
rect 20168 20340 20220 20392
rect 20628 20340 20680 20392
rect 20812 20340 20864 20392
rect 24216 20383 24268 20392
rect 24216 20349 24225 20383
rect 24225 20349 24259 20383
rect 24259 20349 24268 20383
rect 24216 20340 24268 20349
rect 25596 20383 25648 20392
rect 25596 20349 25605 20383
rect 25605 20349 25639 20383
rect 25639 20349 25648 20383
rect 25596 20340 25648 20349
rect 19156 20204 19208 20256
rect 20168 20247 20220 20256
rect 20168 20213 20177 20247
rect 20177 20213 20211 20247
rect 20211 20213 20220 20247
rect 20168 20204 20220 20213
rect 21272 20247 21324 20256
rect 21272 20213 21281 20247
rect 21281 20213 21315 20247
rect 21315 20213 21324 20247
rect 21272 20204 21324 20213
rect 24400 20247 24452 20256
rect 24400 20213 24409 20247
rect 24409 20213 24443 20247
rect 24443 20213 24452 20247
rect 24400 20204 24452 20213
rect 26884 20247 26936 20256
rect 26884 20213 26893 20247
rect 26893 20213 26927 20247
rect 26927 20213 26936 20247
rect 26884 20204 26936 20213
rect 27252 20247 27304 20256
rect 27252 20213 27261 20247
rect 27261 20213 27295 20247
rect 27295 20213 27304 20247
rect 27252 20204 27304 20213
rect 10982 20102 11034 20154
rect 11046 20102 11098 20154
rect 11110 20102 11162 20154
rect 11174 20102 11226 20154
rect 20982 20102 21034 20154
rect 21046 20102 21098 20154
rect 21110 20102 21162 20154
rect 21174 20102 21226 20154
rect 16580 20043 16632 20052
rect 16580 20009 16589 20043
rect 16589 20009 16623 20043
rect 16623 20009 16632 20043
rect 16580 20000 16632 20009
rect 26700 20043 26752 20052
rect 26700 20009 26709 20043
rect 26709 20009 26743 20043
rect 26743 20009 26752 20043
rect 26700 20000 26752 20009
rect 15292 19907 15344 19916
rect 15292 19873 15301 19907
rect 15301 19873 15335 19907
rect 15335 19873 15344 19907
rect 15292 19864 15344 19873
rect 16488 19864 16540 19916
rect 26516 19907 26568 19916
rect 26516 19873 26525 19907
rect 26525 19873 26559 19907
rect 26559 19873 26568 19907
rect 26516 19864 26568 19873
rect 15476 19771 15528 19780
rect 15476 19737 15485 19771
rect 15485 19737 15519 19771
rect 15519 19737 15528 19771
rect 15476 19728 15528 19737
rect 15384 19660 15436 19712
rect 16580 19660 16632 19712
rect 5982 19558 6034 19610
rect 6046 19558 6098 19610
rect 6110 19558 6162 19610
rect 6174 19558 6226 19610
rect 15982 19558 16034 19610
rect 16046 19558 16098 19610
rect 16110 19558 16162 19610
rect 16174 19558 16226 19610
rect 25982 19558 26034 19610
rect 26046 19558 26098 19610
rect 26110 19558 26162 19610
rect 26174 19558 26226 19610
rect 15292 19388 15344 19440
rect 17040 19388 17092 19440
rect 15568 19320 15620 19372
rect 15752 19320 15804 19372
rect 16488 19363 16540 19372
rect 16488 19329 16497 19363
rect 16497 19329 16531 19363
rect 16531 19329 16540 19363
rect 16488 19320 16540 19329
rect 19156 19320 19208 19372
rect 6920 19252 6972 19304
rect 16948 19252 17000 19304
rect 17132 19252 17184 19304
rect 7196 19184 7248 19236
rect 26516 19159 26568 19168
rect 26516 19125 26525 19159
rect 26525 19125 26559 19159
rect 26559 19125 26568 19159
rect 26516 19116 26568 19125
rect 10982 19014 11034 19066
rect 11046 19014 11098 19066
rect 11110 19014 11162 19066
rect 11174 19014 11226 19066
rect 20982 19014 21034 19066
rect 21046 19014 21098 19066
rect 21110 19014 21162 19066
rect 21174 19014 21226 19066
rect 5982 18470 6034 18522
rect 6046 18470 6098 18522
rect 6110 18470 6162 18522
rect 6174 18470 6226 18522
rect 15982 18470 16034 18522
rect 16046 18470 16098 18522
rect 16110 18470 16162 18522
rect 16174 18470 16226 18522
rect 25982 18470 26034 18522
rect 26046 18470 26098 18522
rect 26110 18470 26162 18522
rect 26174 18470 26226 18522
rect 10982 17926 11034 17978
rect 11046 17926 11098 17978
rect 11110 17926 11162 17978
rect 11174 17926 11226 17978
rect 20982 17926 21034 17978
rect 21046 17926 21098 17978
rect 21110 17926 21162 17978
rect 21174 17926 21226 17978
rect 5982 17382 6034 17434
rect 6046 17382 6098 17434
rect 6110 17382 6162 17434
rect 6174 17382 6226 17434
rect 15982 17382 16034 17434
rect 16046 17382 16098 17434
rect 16110 17382 16162 17434
rect 16174 17382 16226 17434
rect 25982 17382 26034 17434
rect 26046 17382 26098 17434
rect 26110 17382 26162 17434
rect 26174 17382 26226 17434
rect 10982 16838 11034 16890
rect 11046 16838 11098 16890
rect 11110 16838 11162 16890
rect 11174 16838 11226 16890
rect 20982 16838 21034 16890
rect 21046 16838 21098 16890
rect 21110 16838 21162 16890
rect 21174 16838 21226 16890
rect 5982 16294 6034 16346
rect 6046 16294 6098 16346
rect 6110 16294 6162 16346
rect 6174 16294 6226 16346
rect 15982 16294 16034 16346
rect 16046 16294 16098 16346
rect 16110 16294 16162 16346
rect 16174 16294 16226 16346
rect 25982 16294 26034 16346
rect 26046 16294 26098 16346
rect 26110 16294 26162 16346
rect 26174 16294 26226 16346
rect 24860 16192 24912 16244
rect 25872 16192 25924 16244
rect 10982 15750 11034 15802
rect 11046 15750 11098 15802
rect 11110 15750 11162 15802
rect 11174 15750 11226 15802
rect 20982 15750 21034 15802
rect 21046 15750 21098 15802
rect 21110 15750 21162 15802
rect 21174 15750 21226 15802
rect 5982 15206 6034 15258
rect 6046 15206 6098 15258
rect 6110 15206 6162 15258
rect 6174 15206 6226 15258
rect 15982 15206 16034 15258
rect 16046 15206 16098 15258
rect 16110 15206 16162 15258
rect 16174 15206 16226 15258
rect 25982 15206 26034 15258
rect 26046 15206 26098 15258
rect 26110 15206 26162 15258
rect 26174 15206 26226 15258
rect 24952 15104 25004 15156
rect 25780 15104 25832 15156
rect 10982 14662 11034 14714
rect 11046 14662 11098 14714
rect 11110 14662 11162 14714
rect 11174 14662 11226 14714
rect 20982 14662 21034 14714
rect 21046 14662 21098 14714
rect 21110 14662 21162 14714
rect 21174 14662 21226 14714
rect 5982 14118 6034 14170
rect 6046 14118 6098 14170
rect 6110 14118 6162 14170
rect 6174 14118 6226 14170
rect 15982 14118 16034 14170
rect 16046 14118 16098 14170
rect 16110 14118 16162 14170
rect 16174 14118 16226 14170
rect 25982 14118 26034 14170
rect 26046 14118 26098 14170
rect 26110 14118 26162 14170
rect 26174 14118 26226 14170
rect 10982 13574 11034 13626
rect 11046 13574 11098 13626
rect 11110 13574 11162 13626
rect 11174 13574 11226 13626
rect 20982 13574 21034 13626
rect 21046 13574 21098 13626
rect 21110 13574 21162 13626
rect 21174 13574 21226 13626
rect 10416 13336 10468 13388
rect 11612 13379 11664 13388
rect 11612 13345 11646 13379
rect 11646 13345 11664 13379
rect 11612 13336 11664 13345
rect 2044 13268 2096 13320
rect 10140 13311 10192 13320
rect 10140 13277 10149 13311
rect 10149 13277 10183 13311
rect 10183 13277 10192 13311
rect 10140 13268 10192 13277
rect 10232 13311 10284 13320
rect 10232 13277 10241 13311
rect 10241 13277 10275 13311
rect 10275 13277 10284 13311
rect 11336 13311 11388 13320
rect 10232 13268 10284 13277
rect 11336 13277 11345 13311
rect 11345 13277 11379 13311
rect 11379 13277 11388 13311
rect 11336 13268 11388 13277
rect 10968 13200 11020 13252
rect 3148 13132 3200 13184
rect 9128 13175 9180 13184
rect 9128 13141 9137 13175
rect 9137 13141 9171 13175
rect 9171 13141 9180 13175
rect 9128 13132 9180 13141
rect 9496 13132 9548 13184
rect 11152 13132 11204 13184
rect 12716 13175 12768 13184
rect 12716 13141 12725 13175
rect 12725 13141 12759 13175
rect 12759 13141 12768 13175
rect 12716 13132 12768 13141
rect 5982 13030 6034 13082
rect 6046 13030 6098 13082
rect 6110 13030 6162 13082
rect 6174 13030 6226 13082
rect 15982 13030 16034 13082
rect 16046 13030 16098 13082
rect 16110 13030 16162 13082
rect 16174 13030 16226 13082
rect 25982 13030 26034 13082
rect 26046 13030 26098 13082
rect 26110 13030 26162 13082
rect 26174 13030 26226 13082
rect 10416 12971 10468 12980
rect 10416 12937 10425 12971
rect 10425 12937 10459 12971
rect 10459 12937 10468 12971
rect 10416 12928 10468 12937
rect 13820 12971 13872 12980
rect 13820 12937 13829 12971
rect 13829 12937 13863 12971
rect 13863 12937 13872 12971
rect 13820 12928 13872 12937
rect 10048 12903 10100 12912
rect 10048 12869 10057 12903
rect 10057 12869 10091 12903
rect 10091 12869 10100 12903
rect 10048 12860 10100 12869
rect 11612 12903 11664 12912
rect 3148 12835 3200 12844
rect 3148 12801 3157 12835
rect 3157 12801 3191 12835
rect 3191 12801 3200 12835
rect 3148 12792 3200 12801
rect 1400 12767 1452 12776
rect 1400 12733 1409 12767
rect 1409 12733 1443 12767
rect 1443 12733 1452 12767
rect 1400 12724 1452 12733
rect 1400 12588 1452 12640
rect 1768 12588 1820 12640
rect 3976 12724 4028 12776
rect 4252 12767 4304 12776
rect 4252 12733 4261 12767
rect 4261 12733 4295 12767
rect 4295 12733 4304 12767
rect 4252 12724 4304 12733
rect 9128 12792 9180 12844
rect 10232 12792 10284 12844
rect 10508 12792 10560 12844
rect 11612 12869 11621 12903
rect 11621 12869 11655 12903
rect 11655 12869 11664 12903
rect 11612 12860 11664 12869
rect 11152 12835 11204 12844
rect 11152 12801 11161 12835
rect 11161 12801 11195 12835
rect 11195 12801 11204 12835
rect 11152 12792 11204 12801
rect 9404 12767 9456 12776
rect 9404 12733 9413 12767
rect 9413 12733 9447 12767
rect 9447 12733 9456 12767
rect 9404 12724 9456 12733
rect 10968 12767 11020 12776
rect 10968 12733 10977 12767
rect 10977 12733 11011 12767
rect 11011 12733 11020 12767
rect 10968 12724 11020 12733
rect 12440 12767 12492 12776
rect 12440 12733 12449 12767
rect 12449 12733 12483 12767
rect 12483 12733 12492 12767
rect 12440 12724 12492 12733
rect 12716 12767 12768 12776
rect 12716 12733 12750 12767
rect 12750 12733 12768 12767
rect 12716 12724 12768 12733
rect 2872 12699 2924 12708
rect 2872 12665 2881 12699
rect 2881 12665 2915 12699
rect 2915 12665 2924 12699
rect 2872 12656 2924 12665
rect 7472 12656 7524 12708
rect 2504 12631 2556 12640
rect 2504 12597 2513 12631
rect 2513 12597 2547 12631
rect 2547 12597 2556 12631
rect 2504 12588 2556 12597
rect 5540 12588 5592 12640
rect 10692 12656 10744 12708
rect 9312 12588 9364 12640
rect 9680 12588 9732 12640
rect 12440 12588 12492 12640
rect 13912 12588 13964 12640
rect 15200 12724 15252 12776
rect 16672 12631 16724 12640
rect 16672 12597 16681 12631
rect 16681 12597 16715 12631
rect 16715 12597 16724 12631
rect 16672 12588 16724 12597
rect 10982 12486 11034 12538
rect 11046 12486 11098 12538
rect 11110 12486 11162 12538
rect 11174 12486 11226 12538
rect 20982 12486 21034 12538
rect 21046 12486 21098 12538
rect 21110 12486 21162 12538
rect 21174 12486 21226 12538
rect 1492 12384 1544 12436
rect 3056 12384 3108 12436
rect 2044 12248 2096 12300
rect 4068 12384 4120 12436
rect 4344 12384 4396 12436
rect 9588 12384 9640 12436
rect 10692 12384 10744 12436
rect 11336 12427 11388 12436
rect 11336 12393 11345 12427
rect 11345 12393 11379 12427
rect 11379 12393 11388 12427
rect 12440 12427 12492 12436
rect 11336 12384 11388 12393
rect 12440 12393 12449 12427
rect 12449 12393 12483 12427
rect 12483 12393 12492 12427
rect 12440 12384 12492 12393
rect 5540 12316 5592 12368
rect 16672 12316 16724 12368
rect 17408 12316 17460 12368
rect 19432 12316 19484 12368
rect 20076 12316 20128 12368
rect 9680 12248 9732 12300
rect 9864 12248 9916 12300
rect 10416 12291 10468 12300
rect 10416 12257 10425 12291
rect 10425 12257 10459 12291
rect 10459 12257 10468 12291
rect 10416 12248 10468 12257
rect 15200 12248 15252 12300
rect 17316 12291 17368 12300
rect 17316 12257 17325 12291
rect 17325 12257 17359 12291
rect 17359 12257 17368 12291
rect 17316 12248 17368 12257
rect 3056 12223 3108 12232
rect 3056 12189 3065 12223
rect 3065 12189 3099 12223
rect 3099 12189 3108 12223
rect 3056 12180 3108 12189
rect 3240 12180 3292 12232
rect 4252 12180 4304 12232
rect 5172 12180 5224 12232
rect 8484 12223 8536 12232
rect 8484 12189 8493 12223
rect 8493 12189 8527 12223
rect 8527 12189 8536 12223
rect 8484 12180 8536 12189
rect 8576 12223 8628 12232
rect 8576 12189 8585 12223
rect 8585 12189 8619 12223
rect 8619 12189 8628 12223
rect 10508 12223 10560 12232
rect 8576 12180 8628 12189
rect 10508 12189 10517 12223
rect 10517 12189 10551 12223
rect 10551 12189 10560 12223
rect 10508 12180 10560 12189
rect 15752 12223 15804 12232
rect 15752 12189 15761 12223
rect 15761 12189 15795 12223
rect 15795 12189 15804 12223
rect 15752 12180 15804 12189
rect 2688 12112 2740 12164
rect 3148 12112 3200 12164
rect 3516 12112 3568 12164
rect 2412 12087 2464 12096
rect 2412 12053 2421 12087
rect 2421 12053 2455 12087
rect 2455 12053 2464 12087
rect 2412 12044 2464 12053
rect 2504 12044 2556 12096
rect 3792 12087 3844 12096
rect 3792 12053 3801 12087
rect 3801 12053 3835 12087
rect 3835 12053 3844 12087
rect 3792 12044 3844 12053
rect 6828 12087 6880 12096
rect 6828 12053 6837 12087
rect 6837 12053 6871 12087
rect 6871 12053 6880 12087
rect 6828 12044 6880 12053
rect 8024 12087 8076 12096
rect 8024 12053 8033 12087
rect 8033 12053 8067 12087
rect 8067 12053 8076 12087
rect 8024 12044 8076 12053
rect 9128 12087 9180 12096
rect 9128 12053 9137 12087
rect 9137 12053 9171 12087
rect 9171 12053 9180 12087
rect 9128 12044 9180 12053
rect 9312 12044 9364 12096
rect 9588 12044 9640 12096
rect 9956 12087 10008 12096
rect 9956 12053 9965 12087
rect 9965 12053 9999 12087
rect 9999 12053 10008 12087
rect 9956 12044 10008 12053
rect 14280 12087 14332 12096
rect 14280 12053 14289 12087
rect 14289 12053 14323 12087
rect 14323 12053 14332 12087
rect 14280 12044 14332 12053
rect 18696 12087 18748 12096
rect 18696 12053 18705 12087
rect 18705 12053 18739 12087
rect 18739 12053 18748 12087
rect 18696 12044 18748 12053
rect 5982 11942 6034 11994
rect 6046 11942 6098 11994
rect 6110 11942 6162 11994
rect 6174 11942 6226 11994
rect 15982 11942 16034 11994
rect 16046 11942 16098 11994
rect 16110 11942 16162 11994
rect 16174 11942 16226 11994
rect 25982 11942 26034 11994
rect 26046 11942 26098 11994
rect 26110 11942 26162 11994
rect 26174 11942 26226 11994
rect 2044 11883 2096 11892
rect 2044 11849 2053 11883
rect 2053 11849 2087 11883
rect 2087 11849 2096 11883
rect 2044 11840 2096 11849
rect 3056 11840 3108 11892
rect 3608 11840 3660 11892
rect 8576 11840 8628 11892
rect 12348 11840 12400 11892
rect 17316 11840 17368 11892
rect 2504 11704 2556 11756
rect 2688 11747 2740 11756
rect 2688 11713 2697 11747
rect 2697 11713 2731 11747
rect 2731 11713 2740 11747
rect 3240 11747 3292 11756
rect 2688 11704 2740 11713
rect 3240 11713 3249 11747
rect 3249 11713 3283 11747
rect 3283 11713 3292 11747
rect 3240 11704 3292 11713
rect 2228 11636 2280 11688
rect 3792 11772 3844 11824
rect 8484 11815 8536 11824
rect 8484 11781 8493 11815
rect 8493 11781 8527 11815
rect 8527 11781 8536 11815
rect 8484 11772 8536 11781
rect 6828 11704 6880 11756
rect 8668 11704 8720 11756
rect 9496 11704 9548 11756
rect 9588 11747 9640 11756
rect 9588 11713 9597 11747
rect 9597 11713 9631 11747
rect 9631 11713 9640 11747
rect 9588 11704 9640 11713
rect 10508 11704 10560 11756
rect 5540 11679 5592 11688
rect 5540 11645 5549 11679
rect 5549 11645 5583 11679
rect 5583 11645 5592 11679
rect 5540 11636 5592 11645
rect 9128 11636 9180 11688
rect 9956 11636 10008 11688
rect 14280 11636 14332 11688
rect 17408 11815 17460 11824
rect 17408 11781 17417 11815
rect 17417 11781 17451 11815
rect 17451 11781 17460 11815
rect 17408 11772 17460 11781
rect 16396 11747 16448 11756
rect 16396 11713 16405 11747
rect 16405 11713 16439 11747
rect 16439 11713 16448 11747
rect 16396 11704 16448 11713
rect 2504 11543 2556 11552
rect 2504 11509 2513 11543
rect 2513 11509 2547 11543
rect 2547 11509 2556 11543
rect 2504 11500 2556 11509
rect 3700 11543 3752 11552
rect 3700 11509 3709 11543
rect 3709 11509 3743 11543
rect 3743 11509 3752 11543
rect 3700 11500 3752 11509
rect 5908 11543 5960 11552
rect 5908 11509 5917 11543
rect 5917 11509 5951 11543
rect 5951 11509 5960 11543
rect 5908 11500 5960 11509
rect 9864 11543 9916 11552
rect 9864 11509 9873 11543
rect 9873 11509 9907 11543
rect 9907 11509 9916 11543
rect 9864 11500 9916 11509
rect 10600 11568 10652 11620
rect 15200 11636 15252 11688
rect 15752 11636 15804 11688
rect 26424 11679 26476 11688
rect 26424 11645 26433 11679
rect 26433 11645 26467 11679
rect 26467 11645 26476 11679
rect 26424 11636 26476 11645
rect 16212 11611 16264 11620
rect 16212 11577 16221 11611
rect 16221 11577 16255 11611
rect 16255 11577 16264 11611
rect 16212 11568 16264 11577
rect 10692 11500 10744 11552
rect 14188 11543 14240 11552
rect 14188 11509 14197 11543
rect 14197 11509 14231 11543
rect 14231 11509 14240 11543
rect 14188 11500 14240 11509
rect 14648 11543 14700 11552
rect 14648 11509 14657 11543
rect 14657 11509 14691 11543
rect 14691 11509 14700 11543
rect 26608 11543 26660 11552
rect 14648 11500 14700 11509
rect 26608 11509 26617 11543
rect 26617 11509 26651 11543
rect 26651 11509 26660 11543
rect 26608 11500 26660 11509
rect 10982 11398 11034 11450
rect 11046 11398 11098 11450
rect 11110 11398 11162 11450
rect 11174 11398 11226 11450
rect 20982 11398 21034 11450
rect 21046 11398 21098 11450
rect 21110 11398 21162 11450
rect 21174 11398 21226 11450
rect 2228 11339 2280 11348
rect 2228 11305 2237 11339
rect 2237 11305 2271 11339
rect 2271 11305 2280 11339
rect 2228 11296 2280 11305
rect 2504 11296 2556 11348
rect 8668 11339 8720 11348
rect 8668 11305 8677 11339
rect 8677 11305 8711 11339
rect 8711 11305 8720 11339
rect 8668 11296 8720 11305
rect 9128 11296 9180 11348
rect 10416 11339 10468 11348
rect 10416 11305 10425 11339
rect 10425 11305 10459 11339
rect 10459 11305 10468 11339
rect 10416 11296 10468 11305
rect 14648 11296 14700 11348
rect 15660 11339 15712 11348
rect 15660 11305 15669 11339
rect 15669 11305 15703 11339
rect 15703 11305 15712 11339
rect 15660 11296 15712 11305
rect 19248 11296 19300 11348
rect 26700 11339 26752 11348
rect 26700 11305 26709 11339
rect 26709 11305 26743 11339
rect 26743 11305 26752 11339
rect 26700 11296 26752 11305
rect 6828 11228 6880 11280
rect 10508 11228 10560 11280
rect 17408 11228 17460 11280
rect 2504 11160 2556 11212
rect 12164 11160 12216 11212
rect 1952 11092 2004 11144
rect 2320 11024 2372 11076
rect 5172 11092 5224 11144
rect 5908 11092 5960 11144
rect 2136 10999 2188 11008
rect 2136 10965 2145 10999
rect 2145 10965 2179 10999
rect 2179 10965 2188 10999
rect 2136 10956 2188 10965
rect 2688 10956 2740 11008
rect 3608 10956 3660 11008
rect 10048 11092 10100 11144
rect 10416 11092 10468 11144
rect 10324 11024 10376 11076
rect 15476 11092 15528 11144
rect 16304 11160 16356 11212
rect 26516 11203 26568 11212
rect 26516 11169 26525 11203
rect 26525 11169 26559 11203
rect 26559 11169 26568 11203
rect 26516 11160 26568 11169
rect 16396 11092 16448 11144
rect 17960 11092 18012 11144
rect 16856 11067 16908 11076
rect 16856 11033 16865 11067
rect 16865 11033 16899 11067
rect 16899 11033 16908 11067
rect 16856 11024 16908 11033
rect 18604 11135 18656 11144
rect 18604 11101 18613 11135
rect 18613 11101 18647 11135
rect 18647 11101 18656 11135
rect 18604 11092 18656 11101
rect 19064 11024 19116 11076
rect 7380 10956 7432 11008
rect 8116 10956 8168 11008
rect 16396 10999 16448 11008
rect 16396 10965 16405 10999
rect 16405 10965 16439 10999
rect 16439 10965 16448 10999
rect 16396 10956 16448 10965
rect 5982 10854 6034 10906
rect 6046 10854 6098 10906
rect 6110 10854 6162 10906
rect 6174 10854 6226 10906
rect 15982 10854 16034 10906
rect 16046 10854 16098 10906
rect 16110 10854 16162 10906
rect 16174 10854 16226 10906
rect 25982 10854 26034 10906
rect 26046 10854 26098 10906
rect 26110 10854 26162 10906
rect 26174 10854 26226 10906
rect 1584 10795 1636 10804
rect 1584 10761 1593 10795
rect 1593 10761 1627 10795
rect 1627 10761 1636 10795
rect 1584 10752 1636 10761
rect 2504 10795 2556 10804
rect 2504 10761 2513 10795
rect 2513 10761 2547 10795
rect 2547 10761 2556 10795
rect 2504 10752 2556 10761
rect 6920 10752 6972 10804
rect 8116 10795 8168 10804
rect 8116 10761 8125 10795
rect 8125 10761 8159 10795
rect 8159 10761 8168 10795
rect 8116 10752 8168 10761
rect 9588 10795 9640 10804
rect 9588 10761 9597 10795
rect 9597 10761 9631 10795
rect 9631 10761 9640 10795
rect 9588 10752 9640 10761
rect 10692 10795 10744 10804
rect 10692 10761 10701 10795
rect 10701 10761 10735 10795
rect 10735 10761 10744 10795
rect 10692 10752 10744 10761
rect 12164 10795 12216 10804
rect 12164 10761 12173 10795
rect 12173 10761 12207 10795
rect 12207 10761 12216 10795
rect 12164 10752 12216 10761
rect 15200 10752 15252 10804
rect 15660 10752 15712 10804
rect 17868 10795 17920 10804
rect 17868 10761 17877 10795
rect 17877 10761 17911 10795
rect 17911 10761 17920 10795
rect 17868 10752 17920 10761
rect 19248 10752 19300 10804
rect 26516 10752 26568 10804
rect 3608 10616 3660 10668
rect 5448 10616 5500 10668
rect 2504 10548 2556 10600
rect 2136 10480 2188 10532
rect 3884 10548 3936 10600
rect 10324 10548 10376 10600
rect 7472 10480 7524 10532
rect 9588 10480 9640 10532
rect 10416 10480 10468 10532
rect 3792 10412 3844 10464
rect 4068 10455 4120 10464
rect 4068 10421 4077 10455
rect 4077 10421 4111 10455
rect 4111 10421 4120 10455
rect 4068 10412 4120 10421
rect 4436 10455 4488 10464
rect 4436 10421 4445 10455
rect 4445 10421 4479 10455
rect 4479 10421 4488 10455
rect 4436 10412 4488 10421
rect 4528 10455 4580 10464
rect 4528 10421 4537 10455
rect 4537 10421 4571 10455
rect 4571 10421 4580 10455
rect 7380 10455 7432 10464
rect 4528 10412 4580 10421
rect 7380 10421 7389 10455
rect 7389 10421 7423 10455
rect 7423 10421 7432 10455
rect 7380 10412 7432 10421
rect 9496 10412 9548 10464
rect 10508 10455 10560 10464
rect 10508 10421 10517 10455
rect 10517 10421 10551 10455
rect 10551 10421 10560 10455
rect 11888 10548 11940 10600
rect 13912 10591 13964 10600
rect 13912 10557 13921 10591
rect 13921 10557 13955 10591
rect 13955 10557 13964 10591
rect 13912 10548 13964 10557
rect 16396 10684 16448 10736
rect 16856 10659 16908 10668
rect 16856 10625 16865 10659
rect 16865 10625 16899 10659
rect 16899 10625 16908 10659
rect 16856 10616 16908 10625
rect 17316 10616 17368 10668
rect 18604 10659 18656 10668
rect 18604 10625 18613 10659
rect 18613 10625 18647 10659
rect 18647 10625 18656 10659
rect 18604 10616 18656 10625
rect 16580 10548 16632 10600
rect 26424 10591 26476 10600
rect 10508 10412 10560 10421
rect 11796 10455 11848 10464
rect 11796 10421 11805 10455
rect 11805 10421 11839 10455
rect 11839 10421 11848 10455
rect 11796 10412 11848 10421
rect 16396 10455 16448 10464
rect 16396 10421 16405 10455
rect 16405 10421 16439 10455
rect 16439 10421 16448 10455
rect 16396 10412 16448 10421
rect 17868 10412 17920 10464
rect 18420 10455 18472 10464
rect 18420 10421 18429 10455
rect 18429 10421 18463 10455
rect 18463 10421 18472 10455
rect 18420 10412 18472 10421
rect 26424 10557 26433 10591
rect 26433 10557 26467 10591
rect 26467 10557 26476 10591
rect 26424 10548 26476 10557
rect 18880 10412 18932 10464
rect 26608 10455 26660 10464
rect 26608 10421 26617 10455
rect 26617 10421 26651 10455
rect 26651 10421 26660 10455
rect 26608 10412 26660 10421
rect 10982 10310 11034 10362
rect 11046 10310 11098 10362
rect 11110 10310 11162 10362
rect 11174 10310 11226 10362
rect 20982 10310 21034 10362
rect 21046 10310 21098 10362
rect 21110 10310 21162 10362
rect 21174 10310 21226 10362
rect 1952 10251 2004 10260
rect 1952 10217 1961 10251
rect 1961 10217 1995 10251
rect 1995 10217 2004 10251
rect 1952 10208 2004 10217
rect 2136 10208 2188 10260
rect 2596 10208 2648 10260
rect 3332 10208 3384 10260
rect 4068 10208 4120 10260
rect 4436 10208 4488 10260
rect 9588 10208 9640 10260
rect 10324 10251 10376 10260
rect 10324 10217 10333 10251
rect 10333 10217 10367 10251
rect 10367 10217 10376 10251
rect 10324 10208 10376 10217
rect 10600 10208 10652 10260
rect 13912 10251 13964 10260
rect 13912 10217 13921 10251
rect 13921 10217 13955 10251
rect 13955 10217 13964 10251
rect 13912 10208 13964 10217
rect 14188 10208 14240 10260
rect 16396 10208 16448 10260
rect 17868 10208 17920 10260
rect 2320 10183 2372 10192
rect 2320 10149 2329 10183
rect 2329 10149 2363 10183
rect 2363 10149 2372 10183
rect 2320 10140 2372 10149
rect 2964 10140 3016 10192
rect 3148 10140 3200 10192
rect 2872 10072 2924 10124
rect 4160 10072 4212 10124
rect 5172 10115 5224 10124
rect 5172 10081 5181 10115
rect 5181 10081 5215 10115
rect 5215 10081 5224 10115
rect 5172 10072 5224 10081
rect 5448 10115 5500 10124
rect 5448 10081 5482 10115
rect 5482 10081 5500 10115
rect 5448 10072 5500 10081
rect 10876 10115 10928 10124
rect 10876 10081 10885 10115
rect 10885 10081 10919 10115
rect 10919 10081 10928 10115
rect 10876 10072 10928 10081
rect 2964 10047 3016 10056
rect 2964 10013 2973 10047
rect 2973 10013 3007 10047
rect 3007 10013 3016 10047
rect 2964 10004 3016 10013
rect 9680 10004 9732 10056
rect 10508 10004 10560 10056
rect 13820 10072 13872 10124
rect 15108 10072 15160 10124
rect 16304 10072 16356 10124
rect 18144 10072 18196 10124
rect 18328 10208 18380 10260
rect 18328 10115 18380 10124
rect 18328 10081 18337 10115
rect 18337 10081 18371 10115
rect 18371 10081 18380 10115
rect 18328 10072 18380 10081
rect 11244 10004 11296 10056
rect 15200 10004 15252 10056
rect 18604 10004 18656 10056
rect 13912 9936 13964 9988
rect 14556 9979 14608 9988
rect 14556 9945 14565 9979
rect 14565 9945 14599 9979
rect 14599 9945 14608 9979
rect 14556 9936 14608 9945
rect 5540 9868 5592 9920
rect 7380 9868 7432 9920
rect 13176 9868 13228 9920
rect 18420 9936 18472 9988
rect 18972 9936 19024 9988
rect 15476 9911 15528 9920
rect 15476 9877 15485 9911
rect 15485 9877 15519 9911
rect 15519 9877 15528 9911
rect 15476 9868 15528 9877
rect 15660 9868 15712 9920
rect 17868 9911 17920 9920
rect 17868 9877 17877 9911
rect 17877 9877 17911 9911
rect 17911 9877 17920 9911
rect 17868 9868 17920 9877
rect 5982 9766 6034 9818
rect 6046 9766 6098 9818
rect 6110 9766 6162 9818
rect 6174 9766 6226 9818
rect 15982 9766 16034 9818
rect 16046 9766 16098 9818
rect 16110 9766 16162 9818
rect 16174 9766 16226 9818
rect 25982 9766 26034 9818
rect 26046 9766 26098 9818
rect 26110 9766 26162 9818
rect 26174 9766 26226 9818
rect 1952 9664 2004 9716
rect 2872 9707 2924 9716
rect 1584 9639 1636 9648
rect 1584 9605 1593 9639
rect 1593 9605 1627 9639
rect 1627 9605 1636 9639
rect 1584 9596 1636 9605
rect 2596 9596 2648 9648
rect 2872 9673 2881 9707
rect 2881 9673 2915 9707
rect 2915 9673 2924 9707
rect 2872 9664 2924 9673
rect 3884 9664 3936 9716
rect 10508 9707 10560 9716
rect 10508 9673 10517 9707
rect 10517 9673 10551 9707
rect 10551 9673 10560 9707
rect 10508 9664 10560 9673
rect 11244 9707 11296 9716
rect 11244 9673 11253 9707
rect 11253 9673 11287 9707
rect 11287 9673 11296 9707
rect 11244 9664 11296 9673
rect 12256 9664 12308 9716
rect 13176 9664 13228 9716
rect 15660 9664 15712 9716
rect 16396 9664 16448 9716
rect 16948 9664 17000 9716
rect 17224 9664 17276 9716
rect 2688 9528 2740 9580
rect 3424 9571 3476 9580
rect 3424 9537 3433 9571
rect 3433 9537 3467 9571
rect 3467 9537 3476 9571
rect 3424 9528 3476 9537
rect 3608 9571 3660 9580
rect 3608 9537 3617 9571
rect 3617 9537 3651 9571
rect 3651 9537 3660 9571
rect 3608 9528 3660 9537
rect 3332 9503 3384 9512
rect 3332 9469 3341 9503
rect 3341 9469 3375 9503
rect 3375 9469 3384 9503
rect 3332 9460 3384 9469
rect 2964 9392 3016 9444
rect 5448 9528 5500 9580
rect 14464 9528 14516 9580
rect 16304 9596 16356 9648
rect 4620 9460 4672 9512
rect 8300 9460 8352 9512
rect 14188 9460 14240 9512
rect 15108 9528 15160 9580
rect 17408 9571 17460 9580
rect 17408 9537 17417 9571
rect 17417 9537 17451 9571
rect 17451 9537 17460 9571
rect 17408 9528 17460 9537
rect 17960 9528 18012 9580
rect 18696 9571 18748 9580
rect 15200 9460 15252 9512
rect 17316 9460 17368 9512
rect 18696 9537 18705 9571
rect 18705 9537 18739 9571
rect 18739 9537 18748 9571
rect 18696 9528 18748 9537
rect 14924 9392 14976 9444
rect 17776 9435 17828 9444
rect 17776 9401 17785 9435
rect 17785 9401 17819 9435
rect 17819 9401 17828 9435
rect 17776 9392 17828 9401
rect 4068 9324 4120 9376
rect 4988 9367 5040 9376
rect 4988 9333 4997 9367
rect 4997 9333 5031 9367
rect 5031 9333 5040 9367
rect 4988 9324 5040 9333
rect 7380 9324 7432 9376
rect 10876 9324 10928 9376
rect 11336 9324 11388 9376
rect 14372 9367 14424 9376
rect 14372 9333 14381 9367
rect 14381 9333 14415 9367
rect 14415 9333 14424 9367
rect 14372 9324 14424 9333
rect 10982 9222 11034 9274
rect 11046 9222 11098 9274
rect 11110 9222 11162 9274
rect 11174 9222 11226 9274
rect 20982 9222 21034 9274
rect 21046 9222 21098 9274
rect 21110 9222 21162 9274
rect 21174 9222 21226 9274
rect 1492 9120 1544 9172
rect 2964 9120 3016 9172
rect 3424 9163 3476 9172
rect 3424 9129 3433 9163
rect 3433 9129 3467 9163
rect 3467 9129 3476 9163
rect 3424 9120 3476 9129
rect 14464 9163 14516 9172
rect 14464 9129 14473 9163
rect 14473 9129 14507 9163
rect 14507 9129 14516 9163
rect 14464 9120 14516 9129
rect 16672 9163 16724 9172
rect 16672 9129 16681 9163
rect 16681 9129 16715 9163
rect 16715 9129 16724 9163
rect 16672 9120 16724 9129
rect 26700 9163 26752 9172
rect 26700 9129 26709 9163
rect 26709 9129 26743 9163
rect 26743 9129 26752 9163
rect 26700 9120 26752 9129
rect 3608 9052 3660 9104
rect 15200 9052 15252 9104
rect 18328 9052 18380 9104
rect 2412 8984 2464 9036
rect 7196 8984 7248 9036
rect 10324 8984 10376 9036
rect 11428 9027 11480 9036
rect 11428 8993 11437 9027
rect 11437 8993 11471 9027
rect 11471 8993 11480 9027
rect 11428 8984 11480 8993
rect 11520 9027 11572 9036
rect 11520 8993 11529 9027
rect 11529 8993 11563 9027
rect 11563 8993 11572 9027
rect 11520 8984 11572 8993
rect 14556 8984 14608 9036
rect 15016 8984 15068 9036
rect 6552 8916 6604 8968
rect 7564 8959 7616 8968
rect 7564 8925 7573 8959
rect 7573 8925 7607 8959
rect 7607 8925 7616 8959
rect 7564 8916 7616 8925
rect 7840 8916 7892 8968
rect 11612 8959 11664 8968
rect 11612 8925 11621 8959
rect 11621 8925 11655 8959
rect 11655 8925 11664 8959
rect 11612 8916 11664 8925
rect 18420 8984 18472 9036
rect 26516 9027 26568 9036
rect 26516 8993 26525 9027
rect 26525 8993 26559 9027
rect 26559 8993 26568 9027
rect 26516 8984 26568 8993
rect 10508 8848 10560 8900
rect 4620 8823 4672 8832
rect 4620 8789 4629 8823
rect 4629 8789 4663 8823
rect 4663 8789 4672 8823
rect 4620 8780 4672 8789
rect 7104 8823 7156 8832
rect 7104 8789 7113 8823
rect 7113 8789 7147 8823
rect 7147 8789 7156 8823
rect 7104 8780 7156 8789
rect 10876 8780 10928 8832
rect 18144 8780 18196 8832
rect 18604 8780 18656 8832
rect 19524 8780 19576 8832
rect 5982 8678 6034 8730
rect 6046 8678 6098 8730
rect 6110 8678 6162 8730
rect 6174 8678 6226 8730
rect 15982 8678 16034 8730
rect 16046 8678 16098 8730
rect 16110 8678 16162 8730
rect 16174 8678 16226 8730
rect 25982 8678 26034 8730
rect 26046 8678 26098 8730
rect 26110 8678 26162 8730
rect 26174 8678 26226 8730
rect 1400 8576 1452 8628
rect 2044 8619 2096 8628
rect 2044 8585 2053 8619
rect 2053 8585 2087 8619
rect 2087 8585 2096 8619
rect 2044 8576 2096 8585
rect 5448 8576 5500 8628
rect 13728 8576 13780 8628
rect 15016 8619 15068 8628
rect 15016 8585 15025 8619
rect 15025 8585 15059 8619
rect 15059 8585 15068 8619
rect 15016 8576 15068 8585
rect 15200 8576 15252 8628
rect 18328 8619 18380 8628
rect 18328 8585 18337 8619
rect 18337 8585 18371 8619
rect 18371 8585 18380 8619
rect 18328 8576 18380 8585
rect 2688 8551 2740 8560
rect 2688 8517 2697 8551
rect 2697 8517 2731 8551
rect 2731 8517 2740 8551
rect 2688 8508 2740 8517
rect 7196 8508 7248 8560
rect 10324 8551 10376 8560
rect 10324 8517 10333 8551
rect 10333 8517 10367 8551
rect 10367 8517 10376 8551
rect 10324 8508 10376 8517
rect 10784 8508 10836 8560
rect 3148 8483 3200 8492
rect 2044 8372 2096 8424
rect 2412 8415 2464 8424
rect 2412 8381 2421 8415
rect 2421 8381 2455 8415
rect 2455 8381 2464 8415
rect 2412 8372 2464 8381
rect 3148 8449 3157 8483
rect 3157 8449 3191 8483
rect 3191 8449 3200 8483
rect 3148 8440 3200 8449
rect 7840 8483 7892 8492
rect 7840 8449 7849 8483
rect 7849 8449 7883 8483
rect 7883 8449 7892 8483
rect 7840 8440 7892 8449
rect 3884 8372 3936 8424
rect 6552 8415 6604 8424
rect 6552 8381 6561 8415
rect 6561 8381 6595 8415
rect 6595 8381 6604 8415
rect 6552 8372 6604 8381
rect 7656 8415 7708 8424
rect 7656 8381 7665 8415
rect 7665 8381 7699 8415
rect 7699 8381 7708 8415
rect 7656 8372 7708 8381
rect 8944 8372 8996 8424
rect 11520 8508 11572 8560
rect 11612 8440 11664 8492
rect 15476 8440 15528 8492
rect 16764 8483 16816 8492
rect 16764 8449 16773 8483
rect 16773 8449 16807 8483
rect 16807 8449 16816 8483
rect 16764 8440 16816 8449
rect 16856 8440 16908 8492
rect 26608 8619 26660 8628
rect 26608 8585 26617 8619
rect 26617 8585 26651 8619
rect 26651 8585 26660 8619
rect 26608 8576 26660 8585
rect 26516 8508 26568 8560
rect 27712 8551 27764 8560
rect 27712 8517 27721 8551
rect 27721 8517 27755 8551
rect 27755 8517 27764 8551
rect 27712 8508 27764 8517
rect 18420 8440 18472 8492
rect 12900 8372 12952 8424
rect 26424 8415 26476 8424
rect 26424 8381 26433 8415
rect 26433 8381 26467 8415
rect 26467 8381 26476 8415
rect 26424 8372 26476 8381
rect 27528 8415 27580 8424
rect 27528 8381 27537 8415
rect 27537 8381 27571 8415
rect 27571 8381 27580 8415
rect 27528 8372 27580 8381
rect 1400 8236 1452 8288
rect 1768 8236 1820 8288
rect 6920 8304 6972 8356
rect 10692 8304 10744 8356
rect 11704 8304 11756 8356
rect 12256 8347 12308 8356
rect 12256 8313 12265 8347
rect 12265 8313 12299 8347
rect 12299 8313 12308 8347
rect 12256 8304 12308 8313
rect 17868 8304 17920 8356
rect 19524 8304 19576 8356
rect 4712 8236 4764 8288
rect 7196 8279 7248 8288
rect 7196 8245 7205 8279
rect 7205 8245 7239 8279
rect 7239 8245 7248 8279
rect 7196 8236 7248 8245
rect 10784 8279 10836 8288
rect 10784 8245 10793 8279
rect 10793 8245 10827 8279
rect 10827 8245 10836 8279
rect 10784 8236 10836 8245
rect 11428 8236 11480 8288
rect 16396 8236 16448 8288
rect 20812 8236 20864 8288
rect 21364 8236 21416 8288
rect 10982 8134 11034 8186
rect 11046 8134 11098 8186
rect 11110 8134 11162 8186
rect 11174 8134 11226 8186
rect 20982 8134 21034 8186
rect 21046 8134 21098 8186
rect 21110 8134 21162 8186
rect 21174 8134 21226 8186
rect 1584 8075 1636 8084
rect 1584 8041 1593 8075
rect 1593 8041 1627 8075
rect 1627 8041 1636 8075
rect 1584 8032 1636 8041
rect 4068 8032 4120 8084
rect 9956 8075 10008 8084
rect 9956 8041 9965 8075
rect 9965 8041 9999 8075
rect 9999 8041 10008 8075
rect 9956 8032 10008 8041
rect 10876 8032 10928 8084
rect 17868 8075 17920 8084
rect 17868 8041 17877 8075
rect 17877 8041 17911 8075
rect 17911 8041 17920 8075
rect 17868 8032 17920 8041
rect 18420 8075 18472 8084
rect 18420 8041 18429 8075
rect 18429 8041 18463 8075
rect 18463 8041 18472 8075
rect 18420 8032 18472 8041
rect 19984 8075 20036 8084
rect 19984 8041 19993 8075
rect 19993 8041 20027 8075
rect 20027 8041 20036 8075
rect 19984 8032 20036 8041
rect 26700 8075 26752 8084
rect 26700 8041 26709 8075
rect 26709 8041 26743 8075
rect 26743 8041 26752 8075
rect 26700 8032 26752 8041
rect 10508 8007 10560 8016
rect 10508 7973 10517 8007
rect 10517 7973 10551 8007
rect 10551 7973 10560 8007
rect 10508 7964 10560 7973
rect 11060 7964 11112 8016
rect 12900 8007 12952 8016
rect 12900 7973 12909 8007
rect 12909 7973 12943 8007
rect 12943 7973 12952 8007
rect 12900 7964 12952 7973
rect 2412 7896 2464 7948
rect 6920 7896 6972 7948
rect 7840 7896 7892 7948
rect 11336 7896 11388 7948
rect 16948 7896 17000 7948
rect 26516 7939 26568 7948
rect 26516 7905 26525 7939
rect 26525 7905 26559 7939
rect 26559 7905 26568 7939
rect 26516 7896 26568 7905
rect 16764 7871 16816 7880
rect 16764 7837 16773 7871
rect 16773 7837 16807 7871
rect 16807 7837 16816 7871
rect 16764 7828 16816 7837
rect 16856 7871 16908 7880
rect 16856 7837 16865 7871
rect 16865 7837 16899 7871
rect 16899 7837 16908 7871
rect 16856 7828 16908 7837
rect 17500 7760 17552 7812
rect 7288 7692 7340 7744
rect 7472 7692 7524 7744
rect 10692 7692 10744 7744
rect 13728 7692 13780 7744
rect 16304 7735 16356 7744
rect 16304 7701 16313 7735
rect 16313 7701 16347 7735
rect 16347 7701 16356 7735
rect 16304 7692 16356 7701
rect 5982 7590 6034 7642
rect 6046 7590 6098 7642
rect 6110 7590 6162 7642
rect 6174 7590 6226 7642
rect 15982 7590 16034 7642
rect 16046 7590 16098 7642
rect 16110 7590 16162 7642
rect 16174 7590 16226 7642
rect 25982 7590 26034 7642
rect 26046 7590 26098 7642
rect 26110 7590 26162 7642
rect 26174 7590 26226 7642
rect 2044 7531 2096 7540
rect 2044 7497 2053 7531
rect 2053 7497 2087 7531
rect 2087 7497 2096 7531
rect 2044 7488 2096 7497
rect 4712 7531 4764 7540
rect 4712 7497 4721 7531
rect 4721 7497 4755 7531
rect 4755 7497 4764 7531
rect 4712 7488 4764 7497
rect 8300 7488 8352 7540
rect 1584 7463 1636 7472
rect 1584 7429 1593 7463
rect 1593 7429 1627 7463
rect 1627 7429 1636 7463
rect 1584 7420 1636 7429
rect 5448 7420 5500 7472
rect 14740 7531 14792 7540
rect 14740 7497 14749 7531
rect 14749 7497 14783 7531
rect 14783 7497 14792 7531
rect 14740 7488 14792 7497
rect 17960 7488 18012 7540
rect 19156 7488 19208 7540
rect 16856 7420 16908 7472
rect 19340 7420 19392 7472
rect 26516 7420 26568 7472
rect 7104 7352 7156 7404
rect 7472 7395 7524 7404
rect 7472 7361 7481 7395
rect 7481 7361 7515 7395
rect 7515 7361 7524 7395
rect 7472 7352 7524 7361
rect 10140 7395 10192 7404
rect 10140 7361 10149 7395
rect 10149 7361 10183 7395
rect 10183 7361 10192 7395
rect 10140 7352 10192 7361
rect 16304 7395 16356 7404
rect 16304 7361 16313 7395
rect 16313 7361 16347 7395
rect 16347 7361 16356 7395
rect 16304 7352 16356 7361
rect 19524 7395 19576 7404
rect 2044 7284 2096 7336
rect 2412 7327 2464 7336
rect 2412 7293 2421 7327
rect 2421 7293 2455 7327
rect 2455 7293 2464 7327
rect 2412 7284 2464 7293
rect 3884 7284 3936 7336
rect 7196 7327 7248 7336
rect 7196 7293 7205 7327
rect 7205 7293 7239 7327
rect 7239 7293 7248 7327
rect 7196 7284 7248 7293
rect 9220 7327 9272 7336
rect 9220 7293 9229 7327
rect 9229 7293 9263 7327
rect 9263 7293 9272 7327
rect 9220 7284 9272 7293
rect 9956 7327 10008 7336
rect 9956 7293 9965 7327
rect 9965 7293 9999 7327
rect 9999 7293 10008 7327
rect 9956 7284 10008 7293
rect 10324 7284 10376 7336
rect 10508 7284 10560 7336
rect 4068 7216 4120 7268
rect 7288 7216 7340 7268
rect 15936 7284 15988 7336
rect 19524 7361 19533 7395
rect 19533 7361 19567 7395
rect 19567 7361 19576 7395
rect 20628 7395 20680 7404
rect 19524 7352 19576 7361
rect 20628 7361 20637 7395
rect 20637 7361 20671 7395
rect 20671 7361 20680 7395
rect 20628 7352 20680 7361
rect 16948 7327 17000 7336
rect 16948 7293 16957 7327
rect 16957 7293 16991 7327
rect 16991 7293 17000 7327
rect 16948 7284 17000 7293
rect 19984 7284 20036 7336
rect 26424 7327 26476 7336
rect 26424 7293 26433 7327
rect 26433 7293 26467 7327
rect 26467 7293 26476 7327
rect 26424 7284 26476 7293
rect 13728 7216 13780 7268
rect 16396 7216 16448 7268
rect 6828 7191 6880 7200
rect 6828 7157 6837 7191
rect 6837 7157 6871 7191
rect 6871 7157 6880 7191
rect 6828 7148 6880 7157
rect 7840 7191 7892 7200
rect 7840 7157 7849 7191
rect 7849 7157 7883 7191
rect 7883 7157 7892 7191
rect 7840 7148 7892 7157
rect 9588 7191 9640 7200
rect 9588 7157 9597 7191
rect 9597 7157 9631 7191
rect 9631 7157 9640 7191
rect 9588 7148 9640 7157
rect 9956 7148 10008 7200
rect 10784 7148 10836 7200
rect 13452 7148 13504 7200
rect 15844 7191 15896 7200
rect 15844 7157 15853 7191
rect 15853 7157 15887 7191
rect 15887 7157 15896 7191
rect 15844 7148 15896 7157
rect 19984 7148 20036 7200
rect 26608 7191 26660 7200
rect 26608 7157 26617 7191
rect 26617 7157 26651 7191
rect 26651 7157 26660 7191
rect 26608 7148 26660 7157
rect 10982 7046 11034 7098
rect 11046 7046 11098 7098
rect 11110 7046 11162 7098
rect 11174 7046 11226 7098
rect 20982 7046 21034 7098
rect 21046 7046 21098 7098
rect 21110 7046 21162 7098
rect 21174 7046 21226 7098
rect 3884 6944 3936 6996
rect 4344 6944 4396 6996
rect 6828 6944 6880 6996
rect 7104 6944 7156 6996
rect 9220 6944 9272 6996
rect 9956 6987 10008 6996
rect 9956 6953 9965 6987
rect 9965 6953 9999 6987
rect 9999 6953 10008 6987
rect 9956 6944 10008 6953
rect 10784 6944 10836 6996
rect 11612 6944 11664 6996
rect 15936 6987 15988 6996
rect 15936 6953 15945 6987
rect 15945 6953 15979 6987
rect 15979 6953 15988 6987
rect 15936 6944 15988 6953
rect 16396 6944 16448 6996
rect 6276 6919 6328 6928
rect 6276 6885 6285 6919
rect 6285 6885 6319 6919
rect 6319 6885 6328 6919
rect 6276 6876 6328 6885
rect 10324 6876 10376 6928
rect 1400 6851 1452 6860
rect 1400 6817 1409 6851
rect 1409 6817 1443 6851
rect 1443 6817 1452 6851
rect 1400 6808 1452 6817
rect 10600 6851 10652 6860
rect 10600 6817 10609 6851
rect 10609 6817 10643 6851
rect 10643 6817 10652 6851
rect 10600 6808 10652 6817
rect 10876 6808 10928 6860
rect 12164 6851 12216 6860
rect 12164 6817 12173 6851
rect 12173 6817 12207 6851
rect 12207 6817 12216 6851
rect 12164 6808 12216 6817
rect 16764 6876 16816 6928
rect 16856 6876 16908 6928
rect 4528 6783 4580 6792
rect 4528 6749 4537 6783
rect 4537 6749 4571 6783
rect 4571 6749 4580 6783
rect 4528 6740 4580 6749
rect 4712 6783 4764 6792
rect 4712 6749 4721 6783
rect 4721 6749 4755 6783
rect 4755 6749 4764 6783
rect 4712 6740 4764 6749
rect 5632 6740 5684 6792
rect 6552 6783 6604 6792
rect 1584 6715 1636 6724
rect 1584 6681 1593 6715
rect 1593 6681 1627 6715
rect 1627 6681 1636 6715
rect 1584 6672 1636 6681
rect 6552 6749 6561 6783
rect 6561 6749 6595 6783
rect 6595 6749 6604 6783
rect 6552 6740 6604 6749
rect 10140 6740 10192 6792
rect 11980 6740 12032 6792
rect 6828 6672 6880 6724
rect 10048 6672 10100 6724
rect 12348 6672 12400 6724
rect 3608 6604 3660 6656
rect 5816 6604 5868 6656
rect 7564 6647 7616 6656
rect 7564 6613 7573 6647
rect 7573 6613 7607 6647
rect 7607 6613 7616 6647
rect 7564 6604 7616 6613
rect 10232 6647 10284 6656
rect 10232 6613 10241 6647
rect 10241 6613 10275 6647
rect 10275 6613 10284 6647
rect 10232 6604 10284 6613
rect 10784 6604 10836 6656
rect 11336 6604 11388 6656
rect 11796 6647 11848 6656
rect 11796 6613 11805 6647
rect 11805 6613 11839 6647
rect 11839 6613 11848 6647
rect 11796 6604 11848 6613
rect 12900 6647 12952 6656
rect 12900 6613 12909 6647
rect 12909 6613 12943 6647
rect 12943 6613 12952 6647
rect 12900 6604 12952 6613
rect 13452 6604 13504 6656
rect 15476 6604 15528 6656
rect 19892 6808 19944 6860
rect 26516 6851 26568 6860
rect 26516 6817 26525 6851
rect 26525 6817 26559 6851
rect 26559 6817 26568 6851
rect 26516 6808 26568 6817
rect 16672 6740 16724 6792
rect 26700 6715 26752 6724
rect 26700 6681 26709 6715
rect 26709 6681 26743 6715
rect 26743 6681 26752 6715
rect 26700 6672 26752 6681
rect 18144 6604 18196 6656
rect 21640 6647 21692 6656
rect 21640 6613 21649 6647
rect 21649 6613 21683 6647
rect 21683 6613 21692 6647
rect 21640 6604 21692 6613
rect 5982 6502 6034 6554
rect 6046 6502 6098 6554
rect 6110 6502 6162 6554
rect 6174 6502 6226 6554
rect 15982 6502 16034 6554
rect 16046 6502 16098 6554
rect 16110 6502 16162 6554
rect 16174 6502 16226 6554
rect 25982 6502 26034 6554
rect 26046 6502 26098 6554
rect 26110 6502 26162 6554
rect 26174 6502 26226 6554
rect 1400 6400 1452 6452
rect 4528 6400 4580 6452
rect 5632 6400 5684 6452
rect 6276 6443 6328 6452
rect 6276 6409 6285 6443
rect 6285 6409 6319 6443
rect 6319 6409 6328 6443
rect 6276 6400 6328 6409
rect 7840 6400 7892 6452
rect 10140 6443 10192 6452
rect 10140 6409 10149 6443
rect 10149 6409 10183 6443
rect 10183 6409 10192 6443
rect 10140 6400 10192 6409
rect 10324 6400 10376 6452
rect 1584 6375 1636 6384
rect 1584 6341 1593 6375
rect 1593 6341 1627 6375
rect 1627 6341 1636 6375
rect 1584 6332 1636 6341
rect 2044 6375 2096 6384
rect 2044 6341 2053 6375
rect 2053 6341 2087 6375
rect 2087 6341 2096 6375
rect 2044 6332 2096 6341
rect 4712 6332 4764 6384
rect 4252 6264 4304 6316
rect 5448 6264 5500 6316
rect 7564 6307 7616 6316
rect 7564 6273 7573 6307
rect 7573 6273 7607 6307
rect 7607 6273 7616 6307
rect 7564 6264 7616 6273
rect 8208 6196 8260 6248
rect 10600 6400 10652 6452
rect 12164 6443 12216 6452
rect 12164 6409 12173 6443
rect 12173 6409 12207 6443
rect 12207 6409 12216 6443
rect 12164 6400 12216 6409
rect 13820 6400 13872 6452
rect 10508 6264 10560 6316
rect 13452 6307 13504 6316
rect 11060 6239 11112 6248
rect 11060 6205 11069 6239
rect 11069 6205 11103 6239
rect 11103 6205 11112 6239
rect 11060 6196 11112 6205
rect 11336 6196 11388 6248
rect 11796 6196 11848 6248
rect 12900 6196 12952 6248
rect 13452 6273 13461 6307
rect 13461 6273 13495 6307
rect 13495 6273 13504 6307
rect 13452 6264 13504 6273
rect 13360 6196 13412 6248
rect 16856 6400 16908 6452
rect 18972 6400 19024 6452
rect 26516 6400 26568 6452
rect 18512 6264 18564 6316
rect 26608 6375 26660 6384
rect 26608 6341 26617 6375
rect 26617 6341 26651 6375
rect 26651 6341 26660 6375
rect 26608 6332 26660 6341
rect 18972 6307 19024 6316
rect 18972 6273 18981 6307
rect 18981 6273 19015 6307
rect 19015 6273 19024 6307
rect 19800 6307 19852 6316
rect 18972 6264 19024 6273
rect 19800 6273 19809 6307
rect 19809 6273 19843 6307
rect 19843 6273 19852 6307
rect 19800 6264 19852 6273
rect 20628 6307 20680 6316
rect 20628 6273 20637 6307
rect 20637 6273 20671 6307
rect 20671 6273 20680 6307
rect 20628 6264 20680 6273
rect 21640 6264 21692 6316
rect 19248 6196 19300 6248
rect 21916 6239 21968 6248
rect 21916 6205 21925 6239
rect 21925 6205 21959 6239
rect 21959 6205 21968 6239
rect 21916 6196 21968 6205
rect 26424 6239 26476 6248
rect 26424 6205 26433 6239
rect 26433 6205 26467 6239
rect 26467 6205 26476 6239
rect 26424 6196 26476 6205
rect 10876 6128 10928 6180
rect 19892 6128 19944 6180
rect 4988 6103 5040 6112
rect 4988 6069 4997 6103
rect 4997 6069 5031 6103
rect 5031 6069 5040 6103
rect 4988 6060 5040 6069
rect 5080 6103 5132 6112
rect 5080 6069 5089 6103
rect 5089 6069 5123 6103
rect 5123 6069 5132 6103
rect 7472 6103 7524 6112
rect 5080 6060 5132 6069
rect 7472 6069 7481 6103
rect 7481 6069 7515 6103
rect 7515 6069 7524 6103
rect 7472 6060 7524 6069
rect 11888 6103 11940 6112
rect 11888 6069 11897 6103
rect 11897 6069 11931 6103
rect 11931 6069 11940 6103
rect 11888 6060 11940 6069
rect 12808 6103 12860 6112
rect 12808 6069 12817 6103
rect 12817 6069 12851 6103
rect 12851 6069 12860 6103
rect 12808 6060 12860 6069
rect 13728 6060 13780 6112
rect 14556 6060 14608 6112
rect 16672 6060 16724 6112
rect 18420 6103 18472 6112
rect 18420 6069 18429 6103
rect 18429 6069 18463 6103
rect 18463 6069 18472 6103
rect 18420 6060 18472 6069
rect 20812 6060 20864 6112
rect 21548 6103 21600 6112
rect 21548 6069 21557 6103
rect 21557 6069 21591 6103
rect 21591 6069 21600 6103
rect 21548 6060 21600 6069
rect 10982 5958 11034 6010
rect 11046 5958 11098 6010
rect 11110 5958 11162 6010
rect 11174 5958 11226 6010
rect 20982 5958 21034 6010
rect 21046 5958 21098 6010
rect 21110 5958 21162 6010
rect 21174 5958 21226 6010
rect 4344 5899 4396 5908
rect 4344 5865 4353 5899
rect 4353 5865 4387 5899
rect 4387 5865 4396 5899
rect 4344 5856 4396 5865
rect 4988 5899 5040 5908
rect 4988 5865 4997 5899
rect 4997 5865 5031 5899
rect 5031 5865 5040 5899
rect 4988 5856 5040 5865
rect 5540 5856 5592 5908
rect 5816 5856 5868 5908
rect 7012 5899 7064 5908
rect 7012 5865 7021 5899
rect 7021 5865 7055 5899
rect 7055 5865 7064 5899
rect 7012 5856 7064 5865
rect 9588 5856 9640 5908
rect 10600 5856 10652 5908
rect 11336 5856 11388 5908
rect 11704 5899 11756 5908
rect 11704 5865 11713 5899
rect 11713 5865 11747 5899
rect 11747 5865 11756 5899
rect 11704 5856 11756 5865
rect 12808 5856 12860 5908
rect 13268 5899 13320 5908
rect 13268 5865 13277 5899
rect 13277 5865 13311 5899
rect 13311 5865 13320 5899
rect 13268 5856 13320 5865
rect 15844 5856 15896 5908
rect 16580 5856 16632 5908
rect 18512 5899 18564 5908
rect 18512 5865 18521 5899
rect 18521 5865 18555 5899
rect 18555 5865 18564 5899
rect 18512 5856 18564 5865
rect 19616 5899 19668 5908
rect 19616 5865 19625 5899
rect 19625 5865 19659 5899
rect 19659 5865 19668 5899
rect 19616 5856 19668 5865
rect 20168 5856 20220 5908
rect 21548 5856 21600 5908
rect 21916 5856 21968 5908
rect 5080 5788 5132 5840
rect 7196 5788 7248 5840
rect 7748 5788 7800 5840
rect 10508 5788 10560 5840
rect 13176 5831 13228 5840
rect 2412 5720 2464 5772
rect 5816 5763 5868 5772
rect 5816 5729 5825 5763
rect 5825 5729 5859 5763
rect 5859 5729 5868 5763
rect 5816 5720 5868 5729
rect 7380 5763 7432 5772
rect 7380 5729 7389 5763
rect 7389 5729 7423 5763
rect 7423 5729 7432 5763
rect 7380 5720 7432 5729
rect 1584 5627 1636 5636
rect 1584 5593 1593 5627
rect 1593 5593 1627 5627
rect 1627 5593 1636 5627
rect 1584 5584 1636 5593
rect 5816 5584 5868 5636
rect 7104 5652 7156 5704
rect 13176 5797 13185 5831
rect 13185 5797 13219 5831
rect 13219 5797 13228 5831
rect 13176 5788 13228 5797
rect 11980 5720 12032 5772
rect 26516 5763 26568 5772
rect 26516 5729 26525 5763
rect 26525 5729 26559 5763
rect 26559 5729 26568 5763
rect 26516 5720 26568 5729
rect 11336 5652 11388 5704
rect 13452 5695 13504 5704
rect 13452 5661 13461 5695
rect 13461 5661 13495 5695
rect 13495 5661 13504 5695
rect 13452 5652 13504 5661
rect 15844 5695 15896 5704
rect 15844 5661 15853 5695
rect 15853 5661 15887 5695
rect 15887 5661 15896 5695
rect 15844 5652 15896 5661
rect 16304 5652 16356 5704
rect 18972 5652 19024 5704
rect 19708 5652 19760 5704
rect 7840 5584 7892 5636
rect 10876 5584 10928 5636
rect 26700 5627 26752 5636
rect 26700 5593 26709 5627
rect 26709 5593 26743 5627
rect 26743 5593 26752 5627
rect 26700 5584 26752 5593
rect 6552 5559 6604 5568
rect 6552 5525 6561 5559
rect 6561 5525 6595 5559
rect 6595 5525 6604 5559
rect 6552 5516 6604 5525
rect 11980 5516 12032 5568
rect 15384 5559 15436 5568
rect 15384 5525 15393 5559
rect 15393 5525 15427 5559
rect 15427 5525 15436 5559
rect 15384 5516 15436 5525
rect 19248 5559 19300 5568
rect 19248 5525 19257 5559
rect 19257 5525 19291 5559
rect 19291 5525 19300 5559
rect 19248 5516 19300 5525
rect 5982 5414 6034 5466
rect 6046 5414 6098 5466
rect 6110 5414 6162 5466
rect 6174 5414 6226 5466
rect 15982 5414 16034 5466
rect 16046 5414 16098 5466
rect 16110 5414 16162 5466
rect 16174 5414 16226 5466
rect 25982 5414 26034 5466
rect 26046 5414 26098 5466
rect 26110 5414 26162 5466
rect 26174 5414 26226 5466
rect 2412 5355 2464 5364
rect 2412 5321 2421 5355
rect 2421 5321 2455 5355
rect 2455 5321 2464 5355
rect 2412 5312 2464 5321
rect 5448 5312 5500 5364
rect 5816 5355 5868 5364
rect 5816 5321 5825 5355
rect 5825 5321 5859 5355
rect 5859 5321 5868 5355
rect 5816 5312 5868 5321
rect 6644 5355 6696 5364
rect 6644 5321 6653 5355
rect 6653 5321 6687 5355
rect 6687 5321 6696 5355
rect 6644 5312 6696 5321
rect 7380 5312 7432 5364
rect 7840 5355 7892 5364
rect 7840 5321 7849 5355
rect 7849 5321 7883 5355
rect 7883 5321 7892 5355
rect 7840 5312 7892 5321
rect 8300 5312 8352 5364
rect 11336 5355 11388 5364
rect 2780 5244 2832 5296
rect 3148 5287 3200 5296
rect 3148 5253 3157 5287
rect 3157 5253 3191 5287
rect 3191 5253 3200 5287
rect 3148 5244 3200 5253
rect 5724 5244 5776 5296
rect 6552 5108 6604 5160
rect 7472 5176 7524 5228
rect 11336 5321 11345 5355
rect 11345 5321 11379 5355
rect 11379 5321 11388 5355
rect 11336 5312 11388 5321
rect 11704 5355 11756 5364
rect 11704 5321 11713 5355
rect 11713 5321 11747 5355
rect 11747 5321 11756 5355
rect 11704 5312 11756 5321
rect 11980 5355 12032 5364
rect 11980 5321 11989 5355
rect 11989 5321 12023 5355
rect 12023 5321 12032 5355
rect 11980 5312 12032 5321
rect 13268 5312 13320 5364
rect 13452 5312 13504 5364
rect 16580 5355 16632 5364
rect 16580 5321 16589 5355
rect 16589 5321 16623 5355
rect 16623 5321 16632 5355
rect 16580 5312 16632 5321
rect 19708 5355 19760 5364
rect 19708 5321 19717 5355
rect 19717 5321 19751 5355
rect 19751 5321 19760 5355
rect 19708 5312 19760 5321
rect 20168 5355 20220 5364
rect 20168 5321 20177 5355
rect 20177 5321 20211 5355
rect 20211 5321 20220 5355
rect 20168 5312 20220 5321
rect 26516 5312 26568 5364
rect 13176 5287 13228 5296
rect 13176 5253 13185 5287
rect 13185 5253 13219 5287
rect 13219 5253 13228 5287
rect 13176 5244 13228 5253
rect 19616 5244 19668 5296
rect 9956 5219 10008 5228
rect 9956 5185 9965 5219
rect 9965 5185 9999 5219
rect 9999 5185 10008 5219
rect 9956 5176 10008 5185
rect 18144 5176 18196 5228
rect 9680 5108 9732 5160
rect 10232 5108 10284 5160
rect 14556 5151 14608 5160
rect 14556 5117 14565 5151
rect 14565 5117 14599 5151
rect 14599 5117 14608 5151
rect 14556 5108 14608 5117
rect 18788 5108 18840 5160
rect 19248 5108 19300 5160
rect 26424 5151 26476 5160
rect 26424 5117 26433 5151
rect 26433 5117 26467 5151
rect 26467 5117 26476 5151
rect 26424 5108 26476 5117
rect 3148 5040 3200 5092
rect 7196 5083 7248 5092
rect 7196 5049 7205 5083
rect 7205 5049 7239 5083
rect 7239 5049 7248 5083
rect 7196 5040 7248 5049
rect 16304 5040 16356 5092
rect 2044 5015 2096 5024
rect 2044 4981 2053 5015
rect 2053 4981 2087 5015
rect 2087 4981 2096 5015
rect 2044 4972 2096 4981
rect 2688 5015 2740 5024
rect 2688 4981 2697 5015
rect 2697 4981 2731 5015
rect 2731 4981 2740 5015
rect 2688 4972 2740 4981
rect 8300 4972 8352 5024
rect 9404 5015 9456 5024
rect 9404 4981 9413 5015
rect 9413 4981 9447 5015
rect 9447 4981 9456 5015
rect 9404 4972 9456 4981
rect 18328 5015 18380 5024
rect 18328 4981 18337 5015
rect 18337 4981 18371 5015
rect 18371 4981 18380 5015
rect 18328 4972 18380 4981
rect 18420 4972 18472 5024
rect 26608 5015 26660 5024
rect 26608 4981 26617 5015
rect 26617 4981 26651 5015
rect 26651 4981 26660 5015
rect 26608 4972 26660 4981
rect 10982 4870 11034 4922
rect 11046 4870 11098 4922
rect 11110 4870 11162 4922
rect 11174 4870 11226 4922
rect 20982 4870 21034 4922
rect 21046 4870 21098 4922
rect 21110 4870 21162 4922
rect 21174 4870 21226 4922
rect 7104 4811 7156 4820
rect 7104 4777 7113 4811
rect 7113 4777 7147 4811
rect 7147 4777 7156 4811
rect 7104 4768 7156 4777
rect 7380 4811 7432 4820
rect 7380 4777 7389 4811
rect 7389 4777 7423 4811
rect 7423 4777 7432 4811
rect 7380 4768 7432 4777
rect 10232 4768 10284 4820
rect 15936 4811 15988 4820
rect 15936 4777 15945 4811
rect 15945 4777 15979 4811
rect 15979 4777 15988 4811
rect 15936 4768 15988 4777
rect 18788 4811 18840 4820
rect 18788 4777 18797 4811
rect 18797 4777 18831 4811
rect 18831 4777 18840 4811
rect 18788 4768 18840 4777
rect 6460 4743 6512 4752
rect 6460 4709 6469 4743
rect 6469 4709 6503 4743
rect 6503 4709 6512 4743
rect 6460 4700 6512 4709
rect 10140 4700 10192 4752
rect 10784 4700 10836 4752
rect 16396 4743 16448 4752
rect 16396 4709 16430 4743
rect 16430 4709 16448 4743
rect 16396 4700 16448 4709
rect 18144 4700 18196 4752
rect 2412 4632 2464 4684
rect 4068 4675 4120 4684
rect 4068 4641 4077 4675
rect 4077 4641 4111 4675
rect 4111 4641 4120 4675
rect 4068 4632 4120 4641
rect 6368 4675 6420 4684
rect 6368 4641 6377 4675
rect 6377 4641 6411 4675
rect 6411 4641 6420 4675
rect 6368 4632 6420 4641
rect 14556 4632 14608 4684
rect 15844 4632 15896 4684
rect 16672 4632 16724 4684
rect 25320 4675 25372 4684
rect 25320 4641 25329 4675
rect 25329 4641 25363 4675
rect 25363 4641 25372 4675
rect 25320 4632 25372 4641
rect 26792 4632 26844 4684
rect 4528 4564 4580 4616
rect 6552 4607 6604 4616
rect 6552 4573 6561 4607
rect 6561 4573 6595 4607
rect 6595 4573 6604 4607
rect 10692 4607 10744 4616
rect 6552 4564 6604 4573
rect 10692 4573 10701 4607
rect 10701 4573 10735 4607
rect 10735 4573 10744 4607
rect 10692 4564 10744 4573
rect 1584 4471 1636 4480
rect 1584 4437 1593 4471
rect 1593 4437 1627 4471
rect 1627 4437 1636 4471
rect 1584 4428 1636 4437
rect 9956 4428 10008 4480
rect 12440 4428 12492 4480
rect 13820 4428 13872 4480
rect 14556 4471 14608 4480
rect 14556 4437 14565 4471
rect 14565 4437 14599 4471
rect 14599 4437 14608 4471
rect 14556 4428 14608 4437
rect 16304 4428 16356 4480
rect 25780 4428 25832 4480
rect 26700 4471 26752 4480
rect 26700 4437 26709 4471
rect 26709 4437 26743 4471
rect 26743 4437 26752 4471
rect 26700 4428 26752 4437
rect 5982 4326 6034 4378
rect 6046 4326 6098 4378
rect 6110 4326 6162 4378
rect 6174 4326 6226 4378
rect 15982 4326 16034 4378
rect 16046 4326 16098 4378
rect 16110 4326 16162 4378
rect 16174 4326 16226 4378
rect 25982 4326 26034 4378
rect 26046 4326 26098 4378
rect 26110 4326 26162 4378
rect 26174 4326 26226 4378
rect 4068 4267 4120 4276
rect 4068 4233 4077 4267
rect 4077 4233 4111 4267
rect 4111 4233 4120 4267
rect 4068 4224 4120 4233
rect 6552 4224 6604 4276
rect 10784 4267 10836 4276
rect 10784 4233 10793 4267
rect 10793 4233 10827 4267
rect 10827 4233 10836 4267
rect 10784 4224 10836 4233
rect 16396 4224 16448 4276
rect 25320 4267 25372 4276
rect 25320 4233 25329 4267
rect 25329 4233 25363 4267
rect 25363 4233 25372 4267
rect 25320 4224 25372 4233
rect 26792 4224 26844 4276
rect 2412 4199 2464 4208
rect 2412 4165 2421 4199
rect 2421 4165 2455 4199
rect 2455 4165 2464 4199
rect 2412 4156 2464 4165
rect 6368 4199 6420 4208
rect 6368 4165 6377 4199
rect 6377 4165 6411 4199
rect 6411 4165 6420 4199
rect 6368 4156 6420 4165
rect 15844 4156 15896 4208
rect 4620 4063 4672 4072
rect 4620 4029 4629 4063
rect 4629 4029 4663 4063
rect 4663 4029 4672 4063
rect 4620 4020 4672 4029
rect 5632 4020 5684 4072
rect 6460 4088 6512 4140
rect 10692 4088 10744 4140
rect 8116 4020 8168 4072
rect 10876 4020 10928 4072
rect 26424 4063 26476 4072
rect 26424 4029 26433 4063
rect 26433 4029 26467 4063
rect 26467 4029 26476 4063
rect 26424 4020 26476 4029
rect 1584 3927 1636 3936
rect 1584 3893 1593 3927
rect 1593 3893 1627 3927
rect 1627 3893 1636 3927
rect 1584 3884 1636 3893
rect 2872 3884 2924 3936
rect 3148 3927 3200 3936
rect 3148 3893 3157 3927
rect 3157 3893 3191 3927
rect 3191 3893 3200 3927
rect 3148 3884 3200 3893
rect 10784 3952 10836 4004
rect 26608 3927 26660 3936
rect 26608 3893 26617 3927
rect 26617 3893 26651 3927
rect 26651 3893 26660 3927
rect 26608 3884 26660 3893
rect 10982 3782 11034 3834
rect 11046 3782 11098 3834
rect 11110 3782 11162 3834
rect 11174 3782 11226 3834
rect 20982 3782 21034 3834
rect 21046 3782 21098 3834
rect 21110 3782 21162 3834
rect 21174 3782 21226 3834
rect 1952 3723 2004 3732
rect 1952 3689 1961 3723
rect 1961 3689 1995 3723
rect 1995 3689 2004 3723
rect 1952 3680 2004 3689
rect 6552 3680 6604 3732
rect 7288 3680 7340 3732
rect 8208 3680 8260 3732
rect 5540 3612 5592 3664
rect 2504 3587 2556 3596
rect 2504 3553 2513 3587
rect 2513 3553 2547 3587
rect 2547 3553 2556 3587
rect 2504 3544 2556 3553
rect 8668 3544 8720 3596
rect 9680 3544 9732 3596
rect 10692 3612 10744 3664
rect 12440 3612 12492 3664
rect 5356 3519 5408 3528
rect 5356 3485 5365 3519
rect 5365 3485 5399 3519
rect 5399 3485 5408 3519
rect 5356 3476 5408 3485
rect 18144 3544 18196 3596
rect 27344 3544 27396 3596
rect 9956 3408 10008 3460
rect 1584 3383 1636 3392
rect 1584 3349 1593 3383
rect 1593 3349 1627 3383
rect 1627 3349 1636 3383
rect 1584 3340 1636 3349
rect 2688 3383 2740 3392
rect 2688 3349 2697 3383
rect 2697 3349 2731 3383
rect 2731 3349 2740 3383
rect 2688 3340 2740 3349
rect 9772 3340 9824 3392
rect 11336 3383 11388 3392
rect 11336 3349 11345 3383
rect 11345 3349 11379 3383
rect 11379 3349 11388 3383
rect 11336 3340 11388 3349
rect 12624 3340 12676 3392
rect 13728 3408 13780 3460
rect 13820 3383 13872 3392
rect 13820 3349 13829 3383
rect 13829 3349 13863 3383
rect 13863 3349 13872 3383
rect 13820 3340 13872 3349
rect 26700 3383 26752 3392
rect 26700 3349 26709 3383
rect 26709 3349 26743 3383
rect 26743 3349 26752 3383
rect 26700 3340 26752 3349
rect 5982 3238 6034 3290
rect 6046 3238 6098 3290
rect 6110 3238 6162 3290
rect 6174 3238 6226 3290
rect 15982 3238 16034 3290
rect 16046 3238 16098 3290
rect 16110 3238 16162 3290
rect 16174 3238 16226 3290
rect 25982 3238 26034 3290
rect 26046 3238 26098 3290
rect 26110 3238 26162 3290
rect 26174 3238 26226 3290
rect 2044 3179 2096 3188
rect 2044 3145 2053 3179
rect 2053 3145 2087 3179
rect 2087 3145 2096 3179
rect 2044 3136 2096 3145
rect 2504 3179 2556 3188
rect 2504 3145 2513 3179
rect 2513 3145 2547 3179
rect 2547 3145 2556 3179
rect 2504 3136 2556 3145
rect 4712 3136 4764 3188
rect 8668 3179 8720 3188
rect 8668 3145 8677 3179
rect 8677 3145 8711 3179
rect 8711 3145 8720 3179
rect 8668 3136 8720 3145
rect 9680 3179 9732 3188
rect 9680 3145 9689 3179
rect 9689 3145 9723 3179
rect 9723 3145 9732 3179
rect 9680 3136 9732 3145
rect 9956 3179 10008 3188
rect 9956 3145 9965 3179
rect 9965 3145 9999 3179
rect 9999 3145 10008 3179
rect 9956 3136 10008 3145
rect 4068 3068 4120 3120
rect 4160 3043 4212 3052
rect 2044 2932 2096 2984
rect 4160 3009 4169 3043
rect 4169 3009 4203 3043
rect 4203 3009 4212 3043
rect 4160 3000 4212 3009
rect 5356 3000 5408 3052
rect 6920 3000 6972 3052
rect 7288 3043 7340 3052
rect 7288 3009 7297 3043
rect 7297 3009 7331 3043
rect 7331 3009 7340 3043
rect 7288 3000 7340 3009
rect 4712 2932 4764 2984
rect 11336 3136 11388 3188
rect 11888 3179 11940 3188
rect 11888 3145 11897 3179
rect 11897 3145 11931 3179
rect 11931 3145 11940 3179
rect 11888 3136 11940 3145
rect 12440 3136 12492 3188
rect 27344 3179 27396 3188
rect 27344 3145 27353 3179
rect 27353 3145 27387 3179
rect 27387 3145 27396 3179
rect 27344 3136 27396 3145
rect 12808 3068 12860 3120
rect 11888 2932 11940 2984
rect 13176 2975 13228 2984
rect 13176 2941 13185 2975
rect 13185 2941 13219 2975
rect 13219 2941 13228 2975
rect 13176 2932 13228 2941
rect 14004 2932 14056 2984
rect 19064 2975 19116 2984
rect 19064 2941 19073 2975
rect 19073 2941 19107 2975
rect 19107 2941 19116 2975
rect 19064 2932 19116 2941
rect 25320 2975 25372 2984
rect 25320 2941 25329 2975
rect 25329 2941 25363 2975
rect 25363 2941 25372 2975
rect 25320 2932 25372 2941
rect 26332 2932 26384 2984
rect 3516 2864 3568 2916
rect 5540 2864 5592 2916
rect 6644 2864 6696 2916
rect 7104 2864 7156 2916
rect 1584 2839 1636 2848
rect 1584 2805 1593 2839
rect 1593 2805 1627 2839
rect 1627 2805 1636 2839
rect 1584 2796 1636 2805
rect 11704 2796 11756 2848
rect 12624 2796 12676 2848
rect 13360 2839 13412 2848
rect 13360 2805 13369 2839
rect 13369 2805 13403 2839
rect 13403 2805 13412 2839
rect 13360 2796 13412 2805
rect 13912 2796 13964 2848
rect 19156 2796 19208 2848
rect 25504 2839 25556 2848
rect 25504 2805 25513 2839
rect 25513 2805 25547 2839
rect 25547 2805 25556 2839
rect 25504 2796 25556 2805
rect 26608 2839 26660 2848
rect 26608 2805 26617 2839
rect 26617 2805 26651 2839
rect 26651 2805 26660 2839
rect 26608 2796 26660 2805
rect 10982 2694 11034 2746
rect 11046 2694 11098 2746
rect 11110 2694 11162 2746
rect 11174 2694 11226 2746
rect 20982 2694 21034 2746
rect 21046 2694 21098 2746
rect 21110 2694 21162 2746
rect 21174 2694 21226 2746
rect 2964 2567 3016 2576
rect 2964 2533 2973 2567
rect 2973 2533 3007 2567
rect 3007 2533 3016 2567
rect 2964 2524 3016 2533
rect 1676 2456 1728 2508
rect 3608 2592 3660 2644
rect 4896 2635 4948 2644
rect 4896 2601 4905 2635
rect 4905 2601 4939 2635
rect 4939 2601 4948 2635
rect 4896 2592 4948 2601
rect 8208 2592 8260 2644
rect 9680 2592 9732 2644
rect 10876 2592 10928 2644
rect 12440 2635 12492 2644
rect 12440 2601 12449 2635
rect 12449 2601 12483 2635
rect 12483 2601 12492 2635
rect 12440 2592 12492 2601
rect 14004 2635 14056 2644
rect 14004 2601 14013 2635
rect 14013 2601 14047 2635
rect 14047 2601 14056 2635
rect 14004 2592 14056 2601
rect 17224 2592 17276 2644
rect 25872 2635 25924 2644
rect 25872 2601 25881 2635
rect 25881 2601 25915 2635
rect 25915 2601 25924 2635
rect 25872 2592 25924 2601
rect 7104 2524 7156 2576
rect 9956 2524 10008 2576
rect 12624 2499 12676 2508
rect 12624 2465 12633 2499
rect 12633 2465 12667 2499
rect 12667 2465 12676 2499
rect 12624 2456 12676 2465
rect 15568 2456 15620 2508
rect 18880 2456 18932 2508
rect 24400 2499 24452 2508
rect 24400 2465 24409 2499
rect 24409 2465 24443 2499
rect 24443 2465 24452 2499
rect 24400 2456 24452 2465
rect 26884 2499 26936 2508
rect 26884 2465 26893 2499
rect 26893 2465 26927 2499
rect 26927 2465 26936 2499
rect 26884 2456 26936 2465
rect 1492 2388 1544 2440
rect 6920 2431 6972 2440
rect 2504 2320 2556 2372
rect 6920 2397 6929 2431
rect 6929 2397 6963 2431
rect 6963 2397 6972 2431
rect 6920 2388 6972 2397
rect 9680 2388 9732 2440
rect 19248 2363 19300 2372
rect 19248 2329 19257 2363
rect 19257 2329 19291 2363
rect 19291 2329 19300 2363
rect 19248 2320 19300 2329
rect 26332 2320 26384 2372
rect 7656 2252 7708 2304
rect 8300 2295 8352 2304
rect 8300 2261 8309 2295
rect 8309 2261 8343 2295
rect 8343 2261 8352 2295
rect 8300 2252 8352 2261
rect 15660 2295 15712 2304
rect 15660 2261 15669 2295
rect 15669 2261 15703 2295
rect 15703 2261 15712 2295
rect 15660 2252 15712 2261
rect 17868 2252 17920 2304
rect 27068 2295 27120 2304
rect 27068 2261 27077 2295
rect 27077 2261 27111 2295
rect 27111 2261 27120 2295
rect 27068 2252 27120 2261
rect 5982 2150 6034 2202
rect 6046 2150 6098 2202
rect 6110 2150 6162 2202
rect 6174 2150 6226 2202
rect 15982 2150 16034 2202
rect 16046 2150 16098 2202
rect 16110 2150 16162 2202
rect 16174 2150 16226 2202
rect 25982 2150 26034 2202
rect 26046 2150 26098 2202
rect 26110 2150 26162 2202
rect 26174 2150 26226 2202
rect 15936 1980 15988 2032
rect 16488 1980 16540 2032
rect 8668 552 8720 604
rect 10600 552 10652 604
<< metal2 >>
rect 754 23520 810 24000
rect 2226 23520 2282 24000
rect 2962 23624 3018 23633
rect 2962 23559 3018 23568
rect 768 20233 796 23520
rect 754 20224 810 20233
rect 754 20159 810 20168
rect 2240 19825 2268 23520
rect 2870 22400 2926 22409
rect 2870 22335 2926 22344
rect 2226 19816 2282 19825
rect 2226 19751 2282 19760
rect 2778 15328 2834 15337
rect 2778 15263 2834 15272
rect 2044 13320 2096 13326
rect 2044 13262 2096 13268
rect 1398 12880 1454 12889
rect 1398 12815 1454 12824
rect 1412 12782 1440 12815
rect 1400 12776 1452 12782
rect 1452 12724 1532 12730
rect 1400 12718 1532 12724
rect 1412 12702 1532 12718
rect 1400 12640 1452 12646
rect 1400 12582 1452 12588
rect 1412 11121 1440 12582
rect 1504 12442 1532 12702
rect 1768 12640 1820 12646
rect 1768 12582 1820 12588
rect 1492 12436 1544 12442
rect 1492 12378 1544 12384
rect 1582 11656 1638 11665
rect 1582 11591 1638 11600
rect 1398 11112 1454 11121
rect 1398 11047 1454 11056
rect 1596 10810 1624 11591
rect 1584 10804 1636 10810
rect 1584 10746 1636 10752
rect 1582 10432 1638 10441
rect 1582 10367 1638 10376
rect 1490 9888 1546 9897
rect 1490 9823 1546 9832
rect 1398 9344 1454 9353
rect 1398 9279 1454 9288
rect 1412 8634 1440 9279
rect 1504 9178 1532 9823
rect 1596 9654 1624 10367
rect 1674 9752 1730 9761
rect 1674 9687 1730 9696
rect 1584 9648 1636 9654
rect 1584 9590 1636 9596
rect 1492 9172 1544 9178
rect 1492 9114 1544 9120
rect 1582 8664 1638 8673
rect 1400 8628 1452 8634
rect 1582 8599 1638 8608
rect 1400 8570 1452 8576
rect 1400 8288 1452 8294
rect 1400 8230 1452 8236
rect 1412 6866 1440 8230
rect 1596 8090 1624 8599
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 1584 7472 1636 7478
rect 1582 7440 1584 7449
rect 1636 7440 1638 7449
rect 1582 7375 1638 7384
rect 1582 6896 1638 6905
rect 1400 6860 1452 6866
rect 1582 6831 1638 6840
rect 1400 6802 1452 6808
rect 1412 6458 1440 6802
rect 1596 6730 1624 6831
rect 1584 6724 1636 6730
rect 1584 6666 1636 6672
rect 1400 6452 1452 6458
rect 1400 6394 1452 6400
rect 1584 6384 1636 6390
rect 1582 6352 1584 6361
rect 1636 6352 1638 6361
rect 1582 6287 1638 6296
rect 1582 5672 1638 5681
rect 1582 5607 1584 5616
rect 1636 5607 1638 5616
rect 1584 5578 1636 5584
rect 1584 4480 1636 4486
rect 1582 4448 1584 4457
rect 1636 4448 1638 4457
rect 1582 4383 1638 4392
rect 1584 3936 1636 3942
rect 1582 3904 1584 3913
rect 1636 3904 1638 3913
rect 1582 3839 1638 3848
rect 1584 3392 1636 3398
rect 1582 3360 1584 3369
rect 1636 3360 1638 3369
rect 1582 3295 1638 3304
rect 1584 2848 1636 2854
rect 570 2816 626 2825
rect 492 2774 570 2802
rect 492 480 520 2774
rect 1584 2790 1636 2796
rect 570 2751 626 2760
rect 1596 2689 1624 2790
rect 1582 2680 1638 2689
rect 1582 2615 1638 2624
rect 1688 2514 1716 9687
rect 1780 8294 1808 12582
rect 2056 12306 2084 13262
rect 2504 12640 2556 12646
rect 2504 12582 2556 12588
rect 2044 12300 2096 12306
rect 2044 12242 2096 12248
rect 2056 11898 2084 12242
rect 2516 12102 2544 12582
rect 2792 12322 2820 15263
rect 2884 12714 2912 22335
rect 2976 22166 3004 23559
rect 3698 23520 3754 24000
rect 5170 23520 5226 24000
rect 6734 23520 6790 24000
rect 8206 23520 8262 24000
rect 9678 23520 9734 24000
rect 11242 23520 11298 24000
rect 12714 23520 12770 24000
rect 14186 23520 14242 24000
rect 15750 23520 15806 24000
rect 17222 23520 17278 24000
rect 18694 23520 18750 24000
rect 20166 23520 20222 24000
rect 21730 23520 21786 24000
rect 23202 23520 23258 24000
rect 24674 23520 24730 24000
rect 25686 23624 25742 23633
rect 25686 23559 25742 23568
rect 3146 23080 3202 23089
rect 3146 23015 3202 23024
rect 3160 22234 3188 23015
rect 3148 22228 3200 22234
rect 3148 22170 3200 22176
rect 2964 22160 3016 22166
rect 2964 22102 3016 22108
rect 3514 21312 3570 21321
rect 3514 21247 3570 21256
rect 3528 20874 3556 21247
rect 3516 20868 3568 20874
rect 3516 20810 3568 20816
rect 3238 20632 3294 20641
rect 3238 20567 3294 20576
rect 2962 14648 3018 14657
rect 2962 14583 3018 14592
rect 2872 12708 2924 12714
rect 2872 12650 2924 12656
rect 2608 12294 2820 12322
rect 2412 12096 2464 12102
rect 2412 12038 2464 12044
rect 2504 12096 2556 12102
rect 2504 12038 2556 12044
rect 2044 11892 2096 11898
rect 2044 11834 2096 11840
rect 2228 11688 2280 11694
rect 2228 11630 2280 11636
rect 2424 11642 2452 12038
rect 2516 11762 2544 12038
rect 2504 11756 2556 11762
rect 2504 11698 2556 11704
rect 2240 11354 2268 11630
rect 2424 11614 2544 11642
rect 2516 11558 2544 11614
rect 2504 11552 2556 11558
rect 2504 11494 2556 11500
rect 2516 11354 2544 11494
rect 2228 11348 2280 11354
rect 2228 11290 2280 11296
rect 2504 11348 2556 11354
rect 2504 11290 2556 11296
rect 2504 11212 2556 11218
rect 2504 11154 2556 11160
rect 1952 11144 2004 11150
rect 1952 11086 2004 11092
rect 1964 10266 1992 11086
rect 2320 11076 2372 11082
rect 2320 11018 2372 11024
rect 2136 11008 2188 11014
rect 2136 10950 2188 10956
rect 2148 10538 2176 10950
rect 2136 10532 2188 10538
rect 2136 10474 2188 10480
rect 2148 10266 2176 10474
rect 1952 10260 2004 10266
rect 1952 10202 2004 10208
rect 2136 10260 2188 10266
rect 2136 10202 2188 10208
rect 1964 9722 1992 10202
rect 2332 10198 2360 11018
rect 2516 10810 2544 11154
rect 2504 10804 2556 10810
rect 2504 10746 2556 10752
rect 2504 10600 2556 10606
rect 2504 10542 2556 10548
rect 2320 10192 2372 10198
rect 2320 10134 2372 10140
rect 2042 10024 2098 10033
rect 2042 9959 2098 9968
rect 1952 9716 2004 9722
rect 1952 9658 2004 9664
rect 2056 9058 2084 9959
rect 1964 9030 2084 9058
rect 2412 9036 2464 9042
rect 1768 8288 1820 8294
rect 1768 8230 1820 8236
rect 1964 3738 1992 9030
rect 2412 8978 2464 8984
rect 2042 8936 2098 8945
rect 2042 8871 2098 8880
rect 2056 8634 2084 8871
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 2056 8430 2084 8570
rect 2424 8430 2452 8978
rect 2044 8424 2096 8430
rect 2412 8424 2464 8430
rect 2044 8366 2096 8372
rect 2410 8392 2412 8401
rect 2464 8392 2466 8401
rect 2410 8327 2466 8336
rect 2042 8256 2098 8265
rect 2042 8191 2098 8200
rect 2056 7546 2084 8191
rect 2412 7948 2464 7954
rect 2412 7890 2464 7896
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 2056 7342 2084 7482
rect 2424 7342 2452 7890
rect 2044 7336 2096 7342
rect 2412 7336 2464 7342
rect 2044 7278 2096 7284
rect 2410 7304 2412 7313
rect 2464 7304 2466 7313
rect 2410 7239 2466 7248
rect 2042 6896 2098 6905
rect 2042 6831 2098 6840
rect 2056 6390 2084 6831
rect 2044 6384 2096 6390
rect 2044 6326 2096 6332
rect 2410 5944 2466 5953
rect 2410 5879 2466 5888
rect 2424 5778 2452 5879
rect 2412 5772 2464 5778
rect 2412 5714 2464 5720
rect 2424 5370 2452 5714
rect 2412 5364 2464 5370
rect 2412 5306 2464 5312
rect 2044 5024 2096 5030
rect 2044 4966 2096 4972
rect 2056 4865 2084 4966
rect 2042 4856 2098 4865
rect 2042 4791 2098 4800
rect 2412 4684 2464 4690
rect 2412 4626 2464 4632
rect 2424 4214 2452 4626
rect 2412 4208 2464 4214
rect 2410 4176 2412 4185
rect 2464 4176 2466 4185
rect 2410 4111 2466 4120
rect 1952 3732 2004 3738
rect 1952 3674 2004 3680
rect 2516 3602 2544 10542
rect 2608 10266 2636 12294
rect 2688 12164 2740 12170
rect 2688 12106 2740 12112
rect 2700 11762 2728 12106
rect 2778 11792 2834 11801
rect 2688 11756 2740 11762
rect 2778 11727 2834 11736
rect 2688 11698 2740 11704
rect 2700 11665 2728 11698
rect 2686 11656 2742 11665
rect 2686 11591 2742 11600
rect 2700 11014 2728 11591
rect 2688 11008 2740 11014
rect 2688 10950 2740 10956
rect 2596 10260 2648 10266
rect 2596 10202 2648 10208
rect 2608 9654 2636 10202
rect 2596 9648 2648 9654
rect 2594 9616 2596 9625
rect 2648 9616 2650 9625
rect 2792 9602 2820 11727
rect 2976 10198 3004 14583
rect 3054 13424 3110 13433
rect 3054 13359 3110 13368
rect 3068 12442 3096 13359
rect 3148 13184 3200 13190
rect 3148 13126 3200 13132
rect 3160 12850 3188 13126
rect 3148 12844 3200 12850
rect 3148 12786 3200 12792
rect 3056 12436 3108 12442
rect 3056 12378 3108 12384
rect 3160 12322 3188 12786
rect 3252 12356 3280 20567
rect 3606 20088 3662 20097
rect 3606 20023 3662 20032
rect 3330 19408 3386 19417
rect 3330 19343 3386 19352
rect 3344 12481 3372 19343
rect 3514 17096 3570 17105
rect 3514 17031 3570 17040
rect 3422 16416 3478 16425
rect 3422 16351 3478 16360
rect 3330 12472 3386 12481
rect 3330 12407 3386 12416
rect 3252 12328 3372 12356
rect 3068 12294 3188 12322
rect 3068 12238 3096 12294
rect 3056 12232 3108 12238
rect 3056 12174 3108 12180
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 3068 11898 3096 12174
rect 3148 12164 3200 12170
rect 3148 12106 3200 12112
rect 3056 11892 3108 11898
rect 3056 11834 3108 11840
rect 3160 11778 3188 12106
rect 3252 11801 3280 12174
rect 3068 11750 3188 11778
rect 3238 11792 3294 11801
rect 2964 10192 3016 10198
rect 2964 10134 3016 10140
rect 2872 10124 2924 10130
rect 2872 10066 2924 10072
rect 2884 10033 2912 10066
rect 2964 10056 3016 10062
rect 2870 10024 2926 10033
rect 2964 9998 3016 10004
rect 2870 9959 2926 9968
rect 2884 9722 2912 9959
rect 2872 9716 2924 9722
rect 2872 9658 2924 9664
rect 2700 9586 2820 9602
rect 2594 9551 2650 9560
rect 2688 9580 2820 9586
rect 2740 9574 2820 9580
rect 2688 9522 2740 9528
rect 2976 9450 3004 9998
rect 2964 9444 3016 9450
rect 2964 9386 3016 9392
rect 2976 9178 3004 9386
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 2688 8560 2740 8566
rect 2688 8502 2740 8508
rect 2700 8129 2728 8502
rect 2686 8120 2742 8129
rect 2686 8055 2742 8064
rect 3068 6769 3096 11750
rect 3238 11727 3240 11736
rect 3292 11727 3294 11736
rect 3240 11698 3292 11704
rect 3344 11370 3372 12328
rect 3252 11342 3372 11370
rect 3146 11112 3202 11121
rect 3146 11047 3202 11056
rect 3160 10441 3188 11047
rect 3146 10432 3202 10441
rect 3146 10367 3202 10376
rect 3148 10192 3200 10198
rect 3148 10134 3200 10140
rect 3160 8650 3188 10134
rect 3252 9058 3280 11342
rect 3436 10305 3464 16351
rect 3528 12170 3556 17031
rect 3516 12164 3568 12170
rect 3516 12106 3568 12112
rect 3620 12050 3648 20023
rect 3712 19961 3740 23520
rect 3882 21856 3938 21865
rect 3882 21791 3938 21800
rect 3896 21690 3924 21791
rect 3884 21684 3936 21690
rect 3884 21626 3936 21632
rect 5184 20602 5212 23520
rect 5956 21788 6252 21808
rect 6012 21786 6036 21788
rect 6092 21786 6116 21788
rect 6172 21786 6196 21788
rect 6034 21734 6036 21786
rect 6098 21734 6110 21786
rect 6172 21734 6174 21786
rect 6012 21732 6036 21734
rect 6092 21732 6116 21734
rect 6172 21732 6196 21734
rect 5956 21712 6252 21732
rect 5956 20700 6252 20720
rect 6012 20698 6036 20700
rect 6092 20698 6116 20700
rect 6172 20698 6196 20700
rect 6034 20646 6036 20698
rect 6098 20646 6110 20698
rect 6172 20646 6174 20698
rect 6012 20644 6036 20646
rect 6092 20644 6116 20646
rect 6172 20644 6196 20646
rect 5956 20624 6252 20644
rect 6748 20602 6776 23520
rect 6920 21684 6972 21690
rect 6920 21626 6972 21632
rect 5172 20596 5224 20602
rect 5172 20538 5224 20544
rect 6736 20596 6788 20602
rect 6736 20538 6788 20544
rect 5356 20256 5408 20262
rect 5356 20198 5408 20204
rect 3698 19952 3754 19961
rect 3698 19887 3754 19896
rect 5368 19417 5396 20198
rect 5956 19612 6252 19632
rect 6012 19610 6036 19612
rect 6092 19610 6116 19612
rect 6172 19610 6196 19612
rect 6034 19558 6036 19610
rect 6098 19558 6110 19610
rect 6172 19558 6174 19610
rect 6012 19556 6036 19558
rect 6092 19556 6116 19558
rect 6172 19556 6196 19558
rect 5956 19536 6252 19556
rect 5354 19408 5410 19417
rect 5354 19343 5410 19352
rect 6932 19310 6960 21626
rect 8220 20602 8248 23520
rect 9404 22228 9456 22234
rect 9404 22170 9456 22176
rect 8944 20800 8996 20806
rect 8944 20742 8996 20748
rect 8208 20596 8260 20602
rect 8208 20538 8260 20544
rect 7470 20360 7526 20369
rect 7470 20295 7472 20304
rect 7524 20295 7526 20304
rect 7472 20266 7524 20272
rect 8576 20256 8628 20262
rect 7562 20224 7618 20233
rect 8576 20198 8628 20204
rect 7562 20159 7618 20168
rect 7576 19689 7604 20159
rect 7562 19680 7618 19689
rect 7562 19615 7618 19624
rect 6920 19304 6972 19310
rect 6920 19246 6972 19252
rect 7196 19236 7248 19242
rect 7196 19178 7248 19184
rect 3698 18864 3754 18873
rect 3698 18799 3754 18808
rect 3528 12022 3648 12050
rect 3422 10296 3478 10305
rect 3332 10260 3384 10266
rect 3422 10231 3478 10240
rect 3332 10202 3384 10208
rect 3344 9518 3372 10202
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 3332 9512 3384 9518
rect 3332 9454 3384 9460
rect 3436 9178 3464 9522
rect 3528 9489 3556 12022
rect 3608 11892 3660 11898
rect 3608 11834 3660 11840
rect 3620 11014 3648 11834
rect 3712 11642 3740 18799
rect 5956 18524 6252 18544
rect 6012 18522 6036 18524
rect 6092 18522 6116 18524
rect 6172 18522 6196 18524
rect 6034 18470 6036 18522
rect 6098 18470 6110 18522
rect 6172 18470 6174 18522
rect 6012 18468 6036 18470
rect 6092 18468 6116 18470
rect 6172 18468 6196 18470
rect 5956 18448 6252 18468
rect 5722 18320 5778 18329
rect 5722 18255 5778 18264
rect 3790 17640 3846 17649
rect 3790 17575 3846 17584
rect 3804 12481 3832 17575
rect 3882 14104 3938 14113
rect 3882 14039 3938 14048
rect 3790 12472 3846 12481
rect 3790 12407 3846 12416
rect 3792 12096 3844 12102
rect 3792 12038 3844 12044
rect 3804 11830 3832 12038
rect 3792 11824 3844 11830
rect 3792 11766 3844 11772
rect 3712 11614 3832 11642
rect 3700 11552 3752 11558
rect 3700 11494 3752 11500
rect 3608 11008 3660 11014
rect 3608 10950 3660 10956
rect 3620 10674 3648 10950
rect 3608 10668 3660 10674
rect 3608 10610 3660 10616
rect 3620 9897 3648 10610
rect 3606 9888 3662 9897
rect 3606 9823 3662 9832
rect 3620 9586 3648 9823
rect 3712 9761 3740 11494
rect 3804 10470 3832 11614
rect 3896 10606 3924 14039
rect 3974 12880 4030 12889
rect 3974 12815 4030 12824
rect 3988 12782 4016 12815
rect 3976 12776 4028 12782
rect 4252 12776 4304 12782
rect 3976 12718 4028 12724
rect 4066 12744 4122 12753
rect 4252 12718 4304 12724
rect 4066 12679 4122 12688
rect 4080 12594 4108 12679
rect 4080 12566 4200 12594
rect 4066 12472 4122 12481
rect 4066 12407 4068 12416
rect 4120 12407 4122 12416
rect 4068 12378 4120 12384
rect 4172 12186 4200 12566
rect 4264 12238 4292 12718
rect 5540 12640 5592 12646
rect 5540 12582 5592 12588
rect 4344 12436 4396 12442
rect 4344 12378 4396 12384
rect 3988 12158 4200 12186
rect 4252 12232 4304 12238
rect 4356 12209 4384 12378
rect 5552 12374 5580 12582
rect 5540 12368 5592 12374
rect 5540 12310 5592 12316
rect 5172 12232 5224 12238
rect 4252 12174 4304 12180
rect 4342 12200 4398 12209
rect 3884 10600 3936 10606
rect 3884 10542 3936 10548
rect 3792 10464 3844 10470
rect 3792 10406 3844 10412
rect 3698 9752 3754 9761
rect 3698 9687 3754 9696
rect 3608 9580 3660 9586
rect 3608 9522 3660 9528
rect 3514 9480 3570 9489
rect 3514 9415 3570 9424
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3620 9110 3648 9522
rect 3608 9104 3660 9110
rect 3252 9030 3464 9058
rect 3608 9046 3660 9052
rect 3160 8622 3372 8650
rect 3146 8528 3202 8537
rect 3146 8463 3148 8472
rect 3200 8463 3202 8472
rect 3148 8434 3200 8440
rect 3054 6760 3110 6769
rect 3054 6695 3110 6704
rect 3344 6633 3372 8622
rect 3436 7857 3464 9030
rect 3804 8129 3832 10406
rect 3988 10146 4016 12158
rect 5172 12174 5224 12180
rect 4342 12135 4398 12144
rect 5184 11150 5212 12174
rect 5552 11694 5580 12310
rect 5540 11688 5592 11694
rect 5538 11656 5540 11665
rect 5592 11656 5594 11665
rect 5538 11591 5594 11600
rect 5172 11144 5224 11150
rect 5172 11086 5224 11092
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 4436 10464 4488 10470
rect 4436 10406 4488 10412
rect 4528 10464 4580 10470
rect 4528 10406 4580 10412
rect 4080 10266 4108 10406
rect 4448 10266 4476 10406
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 4436 10260 4488 10266
rect 4436 10202 4488 10208
rect 4540 10169 4568 10406
rect 4526 10160 4582 10169
rect 3988 10118 4108 10146
rect 3882 9752 3938 9761
rect 3882 9687 3884 9696
rect 3936 9687 3938 9696
rect 3884 9658 3936 9664
rect 4080 9382 4108 10118
rect 4160 10124 4212 10130
rect 5184 10130 5212 11086
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 5460 10130 5488 10610
rect 4526 10095 4582 10104
rect 5172 10124 5224 10130
rect 4160 10066 4212 10072
rect 5172 10066 5224 10072
rect 5448 10124 5500 10130
rect 5448 10066 5500 10072
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 3884 8424 3936 8430
rect 4172 8378 4200 10066
rect 5460 9586 5488 10066
rect 5540 9920 5592 9926
rect 5538 9888 5540 9897
rect 5592 9888 5594 9897
rect 5538 9823 5594 9832
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4632 8838 4660 9454
rect 4988 9376 5040 9382
rect 4988 9318 5040 9324
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 3936 8372 4200 8378
rect 3884 8366 4200 8372
rect 3896 8350 4200 8366
rect 3790 8120 3846 8129
rect 3790 8055 3846 8064
rect 3422 7848 3478 7857
rect 3422 7783 3478 7792
rect 3896 7342 3924 8350
rect 4080 8090 4108 8350
rect 4068 8084 4120 8090
rect 4068 8026 4120 8032
rect 3884 7336 3936 7342
rect 3884 7278 3936 7284
rect 3896 7002 3924 7278
rect 4068 7268 4120 7274
rect 4068 7210 4120 7216
rect 4080 7154 4108 7210
rect 4080 7126 4292 7154
rect 3884 6996 3936 7002
rect 3884 6938 3936 6944
rect 3608 6656 3660 6662
rect 3330 6624 3386 6633
rect 3608 6598 3660 6604
rect 3330 6559 3386 6568
rect 2780 5296 2832 5302
rect 3148 5296 3200 5302
rect 2780 5238 2832 5244
rect 3146 5264 3148 5273
rect 3200 5264 3202 5273
rect 2686 5128 2742 5137
rect 2686 5063 2742 5072
rect 2700 5030 2728 5063
rect 2688 5024 2740 5030
rect 2688 4966 2740 4972
rect 2504 3596 2556 3602
rect 2504 3538 2556 3544
rect 2042 3496 2098 3505
rect 2042 3431 2098 3440
rect 2056 3194 2084 3431
rect 2516 3194 2544 3538
rect 2688 3392 2740 3398
rect 2688 3334 2740 3340
rect 2044 3188 2096 3194
rect 2044 3130 2096 3136
rect 2504 3188 2556 3194
rect 2504 3130 2556 3136
rect 2056 2990 2084 3130
rect 2044 2984 2096 2990
rect 2044 2926 2096 2932
rect 1676 2508 1728 2514
rect 1676 2450 1728 2456
rect 1492 2440 1544 2446
rect 1492 2382 1544 2388
rect 1504 480 1532 2382
rect 2504 2372 2556 2378
rect 2504 2314 2556 2320
rect 2516 480 2544 2314
rect 2700 2145 2728 3334
rect 2686 2136 2742 2145
rect 2686 2071 2742 2080
rect 478 0 534 480
rect 1490 0 1546 480
rect 2502 0 2558 480
rect 2792 377 2820 5238
rect 3146 5199 3202 5208
rect 3160 5098 3188 5199
rect 3148 5092 3200 5098
rect 3148 5034 3200 5040
rect 2872 3936 2924 3942
rect 3148 3936 3200 3942
rect 2872 3878 2924 3884
rect 3146 3904 3148 3913
rect 3200 3904 3202 3913
rect 2884 1465 2912 3878
rect 3146 3839 3202 3848
rect 3516 2916 3568 2922
rect 3516 2858 3568 2864
rect 2962 2816 3018 2825
rect 2962 2751 3018 2760
rect 2976 2582 3004 2751
rect 2964 2576 3016 2582
rect 2964 2518 3016 2524
rect 2870 1456 2926 1465
rect 2870 1391 2926 1400
rect 3528 480 3556 2858
rect 3620 2650 3648 6598
rect 4264 6322 4292 7126
rect 4344 6996 4396 7002
rect 4344 6938 4396 6944
rect 4252 6316 4304 6322
rect 4252 6258 4304 6264
rect 4356 5914 4384 6938
rect 4528 6792 4580 6798
rect 4528 6734 4580 6740
rect 4540 6458 4568 6734
rect 4528 6452 4580 6458
rect 4528 6394 4580 6400
rect 4632 6361 4660 8774
rect 4712 8288 4764 8294
rect 4712 8230 4764 8236
rect 4724 7546 4752 8230
rect 4712 7540 4764 7546
rect 4712 7482 4764 7488
rect 4724 6798 4752 7482
rect 5000 7449 5028 9318
rect 5460 8634 5488 9522
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5448 7472 5500 7478
rect 4986 7440 5042 7449
rect 5448 7414 5500 7420
rect 4986 7375 5042 7384
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 4724 6390 4752 6734
rect 4712 6384 4764 6390
rect 4618 6352 4674 6361
rect 4712 6326 4764 6332
rect 5460 6322 5488 7414
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 5644 6633 5672 6734
rect 5630 6624 5686 6633
rect 5630 6559 5686 6568
rect 5644 6458 5672 6559
rect 5632 6452 5684 6458
rect 5632 6394 5684 6400
rect 4618 6287 4674 6296
rect 5448 6316 5500 6322
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 4066 5128 4122 5137
rect 4066 5063 4122 5072
rect 4080 4690 4108 5063
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 4080 4282 4108 4626
rect 4528 4616 4580 4622
rect 4528 4558 4580 4564
rect 4068 4276 4120 4282
rect 4068 4218 4120 4224
rect 4068 3120 4120 3126
rect 4068 3062 4120 3068
rect 4158 3088 4214 3097
rect 3608 2644 3660 2650
rect 3608 2586 3660 2592
rect 4080 921 4108 3062
rect 4158 3023 4160 3032
rect 4212 3023 4214 3032
rect 4160 2994 4212 3000
rect 4066 912 4122 921
rect 4066 847 4122 856
rect 4540 480 4568 4558
rect 4632 4162 4660 6287
rect 5448 6258 5500 6264
rect 4988 6112 5040 6118
rect 5080 6112 5132 6118
rect 4988 6054 5040 6060
rect 5078 6080 5080 6089
rect 5132 6080 5134 6089
rect 5000 5914 5028 6054
rect 5078 6015 5134 6024
rect 4988 5908 5040 5914
rect 4988 5850 5040 5856
rect 5092 5846 5120 6015
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5080 5840 5132 5846
rect 5080 5782 5132 5788
rect 5448 5364 5500 5370
rect 5552 5352 5580 5850
rect 5500 5324 5580 5352
rect 5736 5794 5764 18255
rect 5956 17436 6252 17456
rect 6012 17434 6036 17436
rect 6092 17434 6116 17436
rect 6172 17434 6196 17436
rect 6034 17382 6036 17434
rect 6098 17382 6110 17434
rect 6172 17382 6174 17434
rect 6012 17380 6036 17382
rect 6092 17380 6116 17382
rect 6172 17380 6196 17382
rect 5956 17360 6252 17380
rect 5956 16348 6252 16368
rect 6012 16346 6036 16348
rect 6092 16346 6116 16348
rect 6172 16346 6196 16348
rect 6034 16294 6036 16346
rect 6098 16294 6110 16346
rect 6172 16294 6174 16346
rect 6012 16292 6036 16294
rect 6092 16292 6116 16294
rect 6172 16292 6196 16294
rect 5956 16272 6252 16292
rect 5956 15260 6252 15280
rect 6012 15258 6036 15260
rect 6092 15258 6116 15260
rect 6172 15258 6196 15260
rect 6034 15206 6036 15258
rect 6098 15206 6110 15258
rect 6172 15206 6174 15258
rect 6012 15204 6036 15206
rect 6092 15204 6116 15206
rect 6172 15204 6196 15206
rect 5956 15184 6252 15204
rect 5956 14172 6252 14192
rect 6012 14170 6036 14172
rect 6092 14170 6116 14172
rect 6172 14170 6196 14172
rect 6034 14118 6036 14170
rect 6098 14118 6110 14170
rect 6172 14118 6174 14170
rect 6012 14116 6036 14118
rect 6092 14116 6116 14118
rect 6172 14116 6196 14118
rect 5956 14096 6252 14116
rect 5956 13084 6252 13104
rect 6012 13082 6036 13084
rect 6092 13082 6116 13084
rect 6172 13082 6196 13084
rect 6034 13030 6036 13082
rect 6098 13030 6110 13082
rect 6172 13030 6174 13082
rect 6012 13028 6036 13030
rect 6092 13028 6116 13030
rect 6172 13028 6196 13030
rect 5956 13008 6252 13028
rect 6828 12096 6880 12102
rect 6828 12038 6880 12044
rect 5956 11996 6252 12016
rect 6012 11994 6036 11996
rect 6092 11994 6116 11996
rect 6172 11994 6196 11996
rect 6034 11942 6036 11994
rect 6098 11942 6110 11994
rect 6172 11942 6174 11994
rect 6012 11940 6036 11942
rect 6092 11940 6116 11942
rect 6172 11940 6196 11942
rect 5956 11920 6252 11940
rect 6840 11762 6868 12038
rect 6828 11756 6880 11762
rect 6828 11698 6880 11704
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 5920 11150 5948 11494
rect 6840 11286 6868 11698
rect 6828 11280 6880 11286
rect 6828 11222 6880 11228
rect 5908 11144 5960 11150
rect 5908 11086 5960 11092
rect 6840 11064 6868 11222
rect 6840 11036 6960 11064
rect 5956 10908 6252 10928
rect 6012 10906 6036 10908
rect 6092 10906 6116 10908
rect 6172 10906 6196 10908
rect 6034 10854 6036 10906
rect 6098 10854 6110 10906
rect 6172 10854 6174 10906
rect 6012 10852 6036 10854
rect 6092 10852 6116 10854
rect 6172 10852 6196 10854
rect 5956 10832 6252 10852
rect 6932 10810 6960 11036
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 6458 10432 6514 10441
rect 6458 10367 6514 10376
rect 5956 9820 6252 9840
rect 6012 9818 6036 9820
rect 6092 9818 6116 9820
rect 6172 9818 6196 9820
rect 6034 9766 6036 9818
rect 6098 9766 6110 9818
rect 6172 9766 6174 9818
rect 6012 9764 6036 9766
rect 6092 9764 6116 9766
rect 6172 9764 6196 9766
rect 5956 9744 6252 9764
rect 5956 8732 6252 8752
rect 6012 8730 6036 8732
rect 6092 8730 6116 8732
rect 6172 8730 6196 8732
rect 6034 8678 6036 8730
rect 6098 8678 6110 8730
rect 6172 8678 6174 8730
rect 6012 8676 6036 8678
rect 6092 8676 6116 8678
rect 6172 8676 6196 8678
rect 5956 8656 6252 8676
rect 6366 8120 6422 8129
rect 6366 8055 6422 8064
rect 6274 7984 6330 7993
rect 6274 7919 6330 7928
rect 5956 7644 6252 7664
rect 6012 7642 6036 7644
rect 6092 7642 6116 7644
rect 6172 7642 6196 7644
rect 6034 7590 6036 7642
rect 6098 7590 6110 7642
rect 6172 7590 6174 7642
rect 6012 7588 6036 7590
rect 6092 7588 6116 7590
rect 6172 7588 6196 7590
rect 5956 7568 6252 7588
rect 6288 6934 6316 7919
rect 6380 7721 6408 8055
rect 6366 7712 6422 7721
rect 6366 7647 6422 7656
rect 6366 7032 6422 7041
rect 6366 6967 6422 6976
rect 6276 6928 6328 6934
rect 6276 6870 6328 6876
rect 5816 6656 5868 6662
rect 5816 6598 5868 6604
rect 5828 5914 5856 6598
rect 5956 6556 6252 6576
rect 6012 6554 6036 6556
rect 6092 6554 6116 6556
rect 6172 6554 6196 6556
rect 6034 6502 6036 6554
rect 6098 6502 6110 6554
rect 6172 6502 6174 6554
rect 6012 6500 6036 6502
rect 6092 6500 6116 6502
rect 6172 6500 6196 6502
rect 5956 6480 6252 6500
rect 6288 6458 6316 6870
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 5816 5908 5868 5914
rect 5816 5850 5868 5856
rect 5814 5808 5870 5817
rect 5736 5766 5814 5794
rect 5448 5306 5500 5312
rect 5736 5302 5764 5766
rect 5814 5743 5816 5752
rect 5868 5743 5870 5752
rect 5816 5714 5868 5720
rect 5816 5636 5868 5642
rect 5816 5578 5868 5584
rect 5828 5370 5856 5578
rect 5956 5468 6252 5488
rect 6012 5466 6036 5468
rect 6092 5466 6116 5468
rect 6172 5466 6196 5468
rect 6034 5414 6036 5466
rect 6098 5414 6110 5466
rect 6172 5414 6174 5466
rect 6012 5412 6036 5414
rect 6092 5412 6116 5414
rect 6172 5412 6196 5414
rect 5956 5392 6252 5412
rect 5816 5364 5868 5370
rect 5816 5306 5868 5312
rect 5724 5296 5776 5302
rect 5724 5238 5776 5244
rect 5956 4380 6252 4400
rect 6012 4378 6036 4380
rect 6092 4378 6116 4380
rect 6172 4378 6196 4380
rect 6034 4326 6036 4378
rect 6098 4326 6110 4378
rect 6172 4326 6174 4378
rect 6012 4324 6036 4326
rect 6092 4324 6116 4326
rect 6172 4324 6196 4326
rect 5956 4304 6252 4324
rect 4632 4134 4752 4162
rect 4620 4072 4672 4078
rect 4618 4040 4620 4049
rect 4672 4040 4674 4049
rect 4618 3975 4674 3984
rect 4724 3194 4752 4134
rect 5632 4072 5684 4078
rect 5632 4014 5684 4020
rect 5540 3664 5592 3670
rect 5540 3606 5592 3612
rect 5356 3528 5408 3534
rect 5356 3470 5408 3476
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 4724 2990 4752 3130
rect 5368 3058 5396 3470
rect 5356 3052 5408 3058
rect 5356 2994 5408 3000
rect 4712 2984 4764 2990
rect 4712 2926 4764 2932
rect 5552 2922 5580 3606
rect 5540 2916 5592 2922
rect 5540 2858 5592 2864
rect 4894 2680 4950 2689
rect 4894 2615 4896 2624
rect 4948 2615 4950 2624
rect 4896 2586 4948 2592
rect 5644 480 5672 4014
rect 6288 3505 6316 6394
rect 6380 4865 6408 6967
rect 6366 4856 6422 4865
rect 6366 4791 6422 4800
rect 6380 4690 6408 4791
rect 6472 4758 6500 10367
rect 7208 9042 7236 19178
rect 8588 18737 8616 20198
rect 8574 18728 8630 18737
rect 8574 18663 8630 18672
rect 8574 13016 8630 13025
rect 8574 12951 8630 12960
rect 7472 12708 7524 12714
rect 7472 12650 7524 12656
rect 7380 11008 7432 11014
rect 7380 10950 7432 10956
rect 7392 10470 7420 10950
rect 7484 10538 7512 12650
rect 8588 12238 8616 12951
rect 8484 12232 8536 12238
rect 8484 12174 8536 12180
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 7472 10532 7524 10538
rect 7472 10474 7524 10480
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 7392 9926 7420 10406
rect 7380 9920 7432 9926
rect 7380 9862 7432 9868
rect 7392 9382 7420 9862
rect 7746 9616 7802 9625
rect 7746 9551 7802 9560
rect 7380 9376 7432 9382
rect 7380 9318 7432 9324
rect 7196 9036 7248 9042
rect 7196 8978 7248 8984
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6564 8430 6592 8910
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 6552 8424 6604 8430
rect 6552 8366 6604 8372
rect 6564 6905 6592 8366
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6932 7954 6960 8298
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 7116 7410 7144 8774
rect 7208 8566 7236 8978
rect 7196 8560 7248 8566
rect 7194 8528 7196 8537
rect 7248 8528 7250 8537
rect 7194 8463 7250 8472
rect 7392 8412 7420 9318
rect 7562 9072 7618 9081
rect 7562 9007 7618 9016
rect 7576 8974 7604 9007
rect 7564 8968 7616 8974
rect 7564 8910 7616 8916
rect 7300 8384 7420 8412
rect 7656 8424 7708 8430
rect 7654 8392 7656 8401
rect 7708 8392 7710 8401
rect 7196 8288 7248 8294
rect 7196 8230 7248 8236
rect 7104 7404 7156 7410
rect 7104 7346 7156 7352
rect 6828 7200 6880 7206
rect 6828 7142 6880 7148
rect 6840 7002 6868 7142
rect 7116 7002 7144 7346
rect 7208 7342 7236 8230
rect 7300 7750 7328 8384
rect 7654 8327 7710 8336
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 7472 7744 7524 7750
rect 7472 7686 7524 7692
rect 7196 7336 7248 7342
rect 7196 7278 7248 7284
rect 7300 7274 7328 7686
rect 7484 7410 7512 7686
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 7288 7268 7340 7274
rect 7288 7210 7340 7216
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 7104 6996 7156 7002
rect 7104 6938 7156 6944
rect 6550 6896 6606 6905
rect 6550 6831 6606 6840
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 6564 5574 6592 6734
rect 6828 6724 6880 6730
rect 6828 6666 6880 6672
rect 6840 6361 6868 6666
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 6826 6352 6882 6361
rect 7576 6322 7604 6598
rect 6826 6287 6882 6296
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7472 6112 7524 6118
rect 7010 6080 7066 6089
rect 7472 6054 7524 6060
rect 7010 6015 7066 6024
rect 7024 5914 7052 6015
rect 7012 5908 7064 5914
rect 7012 5850 7064 5856
rect 7196 5840 7248 5846
rect 7196 5782 7248 5788
rect 7104 5704 7156 5710
rect 7104 5646 7156 5652
rect 6552 5568 6604 5574
rect 6552 5510 6604 5516
rect 6564 5166 6592 5510
rect 6642 5400 6698 5409
rect 6642 5335 6644 5344
rect 6696 5335 6698 5344
rect 6644 5306 6696 5312
rect 6552 5160 6604 5166
rect 6552 5102 6604 5108
rect 6460 4752 6512 4758
rect 6460 4694 6512 4700
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 6380 4214 6408 4626
rect 6368 4208 6420 4214
rect 6368 4150 6420 4156
rect 6472 4146 6500 4694
rect 6564 4622 6592 5102
rect 7116 4826 7144 5646
rect 7208 5098 7236 5782
rect 7380 5772 7432 5778
rect 7380 5714 7432 5720
rect 7392 5370 7420 5714
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 7196 5092 7248 5098
rect 7196 5034 7248 5040
rect 7104 4820 7156 4826
rect 7104 4762 7156 4768
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 6564 4282 6592 4558
rect 6552 4276 6604 4282
rect 6552 4218 6604 4224
rect 6460 4140 6512 4146
rect 6460 4082 6512 4088
rect 6564 3738 6592 4218
rect 7208 3913 7236 5034
rect 7392 4826 7420 5306
rect 7484 5234 7512 6054
rect 7760 5846 7788 9551
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 7852 8498 7880 8910
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 7852 7954 7880 8434
rect 7840 7948 7892 7954
rect 7840 7890 7892 7896
rect 7852 7206 7880 7890
rect 7840 7200 7892 7206
rect 7840 7142 7892 7148
rect 7852 6458 7880 7142
rect 7840 6452 7892 6458
rect 7840 6394 7892 6400
rect 7748 5840 7800 5846
rect 7748 5782 7800 5788
rect 7852 5642 7880 6394
rect 7840 5636 7892 5642
rect 7840 5578 7892 5584
rect 7852 5370 7880 5578
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7380 4820 7432 4826
rect 7380 4762 7432 4768
rect 7194 3904 7250 3913
rect 7194 3839 7250 3848
rect 6552 3732 6604 3738
rect 6552 3674 6604 3680
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 6274 3496 6330 3505
rect 6274 3431 6330 3440
rect 5956 3292 6252 3312
rect 6012 3290 6036 3292
rect 6092 3290 6116 3292
rect 6172 3290 6196 3292
rect 6034 3238 6036 3290
rect 6098 3238 6110 3290
rect 6172 3238 6174 3290
rect 6012 3236 6036 3238
rect 6092 3236 6116 3238
rect 6172 3236 6196 3238
rect 5956 3216 6252 3236
rect 7300 3058 7328 3674
rect 6920 3052 6972 3058
rect 6920 2994 6972 3000
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 6644 2916 6696 2922
rect 6644 2858 6696 2864
rect 5956 2204 6252 2224
rect 6012 2202 6036 2204
rect 6092 2202 6116 2204
rect 6172 2202 6196 2204
rect 6034 2150 6036 2202
rect 6098 2150 6110 2202
rect 6172 2150 6174 2202
rect 6012 2148 6036 2150
rect 6092 2148 6116 2150
rect 6172 2148 6196 2150
rect 5956 2128 6252 2148
rect 6656 480 6684 2858
rect 6932 2446 6960 2994
rect 7104 2916 7156 2922
rect 7104 2858 7156 2864
rect 7116 2582 7144 2858
rect 8036 2689 8064 12038
rect 8496 11830 8524 12174
rect 8588 11898 8616 12174
rect 8576 11892 8628 11898
rect 8576 11834 8628 11840
rect 8484 11824 8536 11830
rect 8484 11766 8536 11772
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 8680 11354 8708 11698
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 8128 10810 8156 10950
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 8300 9512 8352 9518
rect 8300 9454 8352 9460
rect 8312 7546 8340 9454
rect 8956 8430 8984 20742
rect 9310 13288 9366 13297
rect 9310 13223 9366 13232
rect 9128 13184 9180 13190
rect 9128 13126 9180 13132
rect 9140 12850 9168 13126
rect 9128 12844 9180 12850
rect 9128 12786 9180 12792
rect 9324 12646 9352 13223
rect 9416 12782 9444 22170
rect 9692 20505 9720 23520
rect 11256 21434 11284 23520
rect 11256 21406 11376 21434
rect 10956 21244 11252 21264
rect 11012 21242 11036 21244
rect 11092 21242 11116 21244
rect 11172 21242 11196 21244
rect 11034 21190 11036 21242
rect 11098 21190 11110 21242
rect 11172 21190 11174 21242
rect 11012 21188 11036 21190
rect 11092 21188 11116 21190
rect 11172 21188 11196 21190
rect 10956 21168 11252 21188
rect 10784 20868 10836 20874
rect 10784 20810 10836 20816
rect 9678 20496 9734 20505
rect 9678 20431 9734 20440
rect 9954 15872 10010 15881
rect 9954 15807 10010 15816
rect 9496 13184 9548 13190
rect 9496 13126 9548 13132
rect 9404 12776 9456 12782
rect 9404 12718 9456 12724
rect 9312 12640 9364 12646
rect 9312 12582 9364 12588
rect 9324 12102 9352 12582
rect 9128 12096 9180 12102
rect 9128 12038 9180 12044
rect 9312 12096 9364 12102
rect 9312 12038 9364 12044
rect 9140 11914 9168 12038
rect 9048 11886 9168 11914
rect 8944 8424 8996 8430
rect 8944 8366 8996 8372
rect 9048 8265 9076 11886
rect 9416 11801 9444 12718
rect 9402 11792 9458 11801
rect 9508 11762 9536 13126
rect 9968 12764 9996 15807
rect 10138 13424 10194 13433
rect 10138 13359 10194 13368
rect 10416 13388 10468 13394
rect 10152 13326 10180 13359
rect 10416 13330 10468 13336
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 10232 13320 10284 13326
rect 10232 13262 10284 13268
rect 10152 13002 10180 13262
rect 10060 12974 10180 13002
rect 10060 12918 10088 12974
rect 10048 12912 10100 12918
rect 10046 12880 10048 12889
rect 10100 12880 10102 12889
rect 10244 12850 10272 13262
rect 10428 12986 10456 13330
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10046 12815 10102 12824
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 10508 12844 10560 12850
rect 10508 12786 10560 12792
rect 9968 12736 10088 12764
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9692 12458 9720 12582
rect 9600 12442 9720 12458
rect 9588 12436 9720 12442
rect 9640 12430 9720 12436
rect 9588 12378 9640 12384
rect 9600 12347 9628 12378
rect 9862 12336 9918 12345
rect 9680 12300 9732 12306
rect 9862 12271 9864 12280
rect 9680 12242 9732 12248
rect 9916 12271 9918 12280
rect 9864 12242 9916 12248
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 9600 11762 9628 12038
rect 9402 11727 9458 11736
rect 9496 11756 9548 11762
rect 9496 11698 9548 11704
rect 9588 11756 9640 11762
rect 9588 11698 9640 11704
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 9140 11354 9168 11630
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 9600 10810 9628 11698
rect 9588 10804 9640 10810
rect 9588 10746 9640 10752
rect 9494 10704 9550 10713
rect 9494 10639 9550 10648
rect 9508 10470 9536 10639
rect 9586 10568 9642 10577
rect 9586 10503 9588 10512
rect 9640 10503 9642 10512
rect 9588 10474 9640 10480
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9588 10260 9640 10266
rect 9588 10202 9640 10208
rect 9600 9897 9628 10202
rect 9692 10062 9720 12242
rect 9876 11558 9904 12242
rect 9956 12096 10008 12102
rect 9956 12038 10008 12044
rect 9968 11694 9996 12038
rect 9956 11688 10008 11694
rect 9956 11630 10008 11636
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9586 9888 9642 9897
rect 9586 9823 9642 9832
rect 9034 8256 9090 8265
rect 9034 8191 9090 8200
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 8208 6248 8260 6254
rect 8208 6190 8260 6196
rect 8220 5012 8248 6190
rect 8312 5370 8340 7482
rect 9218 7440 9274 7449
rect 9218 7375 9274 7384
rect 9232 7342 9260 7375
rect 9220 7336 9272 7342
rect 9220 7278 9272 7284
rect 9232 7002 9260 7278
rect 9588 7200 9640 7206
rect 9588 7142 9640 7148
rect 9220 6996 9272 7002
rect 9220 6938 9272 6944
rect 9600 5914 9628 7142
rect 9588 5908 9640 5914
rect 9588 5850 9640 5856
rect 9600 5658 9628 5850
rect 9692 5794 9720 9998
rect 9876 6905 9904 11494
rect 10060 11150 10088 12736
rect 10416 12300 10468 12306
rect 10416 12242 10468 12248
rect 10230 12200 10286 12209
rect 10230 12135 10286 12144
rect 10048 11144 10100 11150
rect 10048 11086 10100 11092
rect 10046 9344 10102 9353
rect 10046 9279 10102 9288
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 9968 7342 9996 8026
rect 9956 7336 10008 7342
rect 9956 7278 10008 7284
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 9968 7002 9996 7142
rect 9956 6996 10008 7002
rect 9956 6938 10008 6944
rect 9862 6896 9918 6905
rect 9862 6831 9918 6840
rect 10060 6730 10088 9279
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 10152 6798 10180 7346
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10244 6746 10272 12135
rect 10428 11354 10456 12242
rect 10520 12238 10548 12786
rect 10692 12708 10744 12714
rect 10692 12650 10744 12656
rect 10704 12442 10732 12650
rect 10692 12436 10744 12442
rect 10692 12378 10744 12384
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 10520 11762 10548 12174
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10416 11348 10468 11354
rect 10416 11290 10468 11296
rect 10520 11286 10548 11698
rect 10600 11620 10652 11626
rect 10600 11562 10652 11568
rect 10508 11280 10560 11286
rect 10508 11222 10560 11228
rect 10416 11144 10468 11150
rect 10416 11086 10468 11092
rect 10324 11076 10376 11082
rect 10324 11018 10376 11024
rect 10336 10606 10364 11018
rect 10324 10600 10376 10606
rect 10324 10542 10376 10548
rect 10336 10266 10364 10542
rect 10428 10538 10456 11086
rect 10416 10532 10468 10538
rect 10416 10474 10468 10480
rect 10324 10260 10376 10266
rect 10324 10202 10376 10208
rect 10324 9036 10376 9042
rect 10324 8978 10376 8984
rect 10336 8566 10364 8978
rect 10324 8560 10376 8566
rect 10324 8502 10376 8508
rect 10324 7336 10376 7342
rect 10324 7278 10376 7284
rect 10336 6934 10364 7278
rect 10324 6928 10376 6934
rect 10324 6870 10376 6876
rect 10048 6724 10100 6730
rect 10048 6666 10100 6672
rect 10152 6458 10180 6734
rect 10244 6718 10364 6746
rect 10232 6656 10284 6662
rect 10232 6598 10284 6604
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 9692 5766 9812 5794
rect 9600 5630 9720 5658
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 9692 5166 9720 5630
rect 9784 5409 9812 5766
rect 9770 5400 9826 5409
rect 9770 5335 9826 5344
rect 9956 5228 10008 5234
rect 9956 5170 10008 5176
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 8300 5024 8352 5030
rect 8220 4984 8300 5012
rect 8116 4072 8168 4078
rect 8116 4014 8168 4020
rect 8128 3641 8156 4014
rect 8220 3738 8248 4984
rect 8300 4966 8352 4972
rect 9404 5024 9456 5030
rect 9404 4966 9456 4972
rect 9416 4049 9444 4966
rect 9968 4486 9996 5170
rect 10152 4758 10180 6394
rect 10244 5166 10272 6598
rect 10336 6458 10364 6718
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 10232 5160 10284 5166
rect 10232 5102 10284 5108
rect 10244 4826 10272 5102
rect 10232 4820 10284 4826
rect 10232 4762 10284 4768
rect 10140 4752 10192 4758
rect 10140 4694 10192 4700
rect 9956 4480 10008 4486
rect 9956 4422 10008 4428
rect 9402 4040 9458 4049
rect 9402 3975 9458 3984
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 8114 3632 8170 3641
rect 8114 3567 8170 3576
rect 8022 2680 8078 2689
rect 8220 2650 8248 3674
rect 8668 3596 8720 3602
rect 8668 3538 8720 3544
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 8680 3194 8708 3538
rect 9692 3194 9720 3538
rect 9968 3466 9996 4422
rect 10428 4049 10456 10474
rect 10508 10464 10560 10470
rect 10506 10432 10508 10441
rect 10560 10432 10562 10441
rect 10506 10367 10562 10376
rect 10612 10266 10640 11562
rect 10692 11552 10744 11558
rect 10692 11494 10744 11500
rect 10704 10810 10732 11494
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 10600 10260 10652 10266
rect 10600 10202 10652 10208
rect 10508 10056 10560 10062
rect 10508 9998 10560 10004
rect 10520 9722 10548 9998
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10508 8900 10560 8906
rect 10508 8842 10560 8848
rect 10520 8022 10548 8842
rect 10796 8566 10824 20810
rect 11348 20602 11376 21406
rect 11520 20868 11572 20874
rect 11520 20810 11572 20816
rect 11336 20596 11388 20602
rect 11336 20538 11388 20544
rect 10956 20156 11252 20176
rect 11012 20154 11036 20156
rect 11092 20154 11116 20156
rect 11172 20154 11196 20156
rect 11034 20102 11036 20154
rect 11098 20102 11110 20154
rect 11172 20102 11174 20154
rect 11012 20100 11036 20102
rect 11092 20100 11116 20102
rect 11172 20100 11196 20102
rect 10956 20080 11252 20100
rect 10956 19068 11252 19088
rect 11012 19066 11036 19068
rect 11092 19066 11116 19068
rect 11172 19066 11196 19068
rect 11034 19014 11036 19066
rect 11098 19014 11110 19066
rect 11172 19014 11174 19066
rect 11012 19012 11036 19014
rect 11092 19012 11116 19014
rect 11172 19012 11196 19014
rect 10956 18992 11252 19012
rect 10956 17980 11252 18000
rect 11012 17978 11036 17980
rect 11092 17978 11116 17980
rect 11172 17978 11196 17980
rect 11034 17926 11036 17978
rect 11098 17926 11110 17978
rect 11172 17926 11174 17978
rect 11012 17924 11036 17926
rect 11092 17924 11116 17926
rect 11172 17924 11196 17926
rect 10956 17904 11252 17924
rect 10956 16892 11252 16912
rect 11012 16890 11036 16892
rect 11092 16890 11116 16892
rect 11172 16890 11196 16892
rect 11034 16838 11036 16890
rect 11098 16838 11110 16890
rect 11172 16838 11174 16890
rect 11012 16836 11036 16838
rect 11092 16836 11116 16838
rect 11172 16836 11196 16838
rect 10956 16816 11252 16836
rect 10956 15804 11252 15824
rect 11012 15802 11036 15804
rect 11092 15802 11116 15804
rect 11172 15802 11196 15804
rect 11034 15750 11036 15802
rect 11098 15750 11110 15802
rect 11172 15750 11174 15802
rect 11012 15748 11036 15750
rect 11092 15748 11116 15750
rect 11172 15748 11196 15750
rect 10956 15728 11252 15748
rect 10956 14716 11252 14736
rect 11012 14714 11036 14716
rect 11092 14714 11116 14716
rect 11172 14714 11196 14716
rect 11034 14662 11036 14714
rect 11098 14662 11110 14714
rect 11172 14662 11174 14714
rect 11012 14660 11036 14662
rect 11092 14660 11116 14662
rect 11172 14660 11196 14662
rect 10956 14640 11252 14660
rect 10956 13628 11252 13648
rect 11012 13626 11036 13628
rect 11092 13626 11116 13628
rect 11172 13626 11196 13628
rect 11034 13574 11036 13626
rect 11098 13574 11110 13626
rect 11172 13574 11174 13626
rect 11012 13572 11036 13574
rect 11092 13572 11116 13574
rect 11172 13572 11196 13574
rect 10956 13552 11252 13572
rect 11336 13320 11388 13326
rect 11336 13262 11388 13268
rect 10968 13252 11020 13258
rect 10968 13194 11020 13200
rect 10980 12782 11008 13194
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 11164 12850 11192 13126
rect 11152 12844 11204 12850
rect 11152 12786 11204 12792
rect 10968 12776 11020 12782
rect 10968 12718 11020 12724
rect 10956 12540 11252 12560
rect 11012 12538 11036 12540
rect 11092 12538 11116 12540
rect 11172 12538 11196 12540
rect 11034 12486 11036 12538
rect 11098 12486 11110 12538
rect 11172 12486 11174 12538
rect 11012 12484 11036 12486
rect 11092 12484 11116 12486
rect 11172 12484 11196 12486
rect 10956 12464 11252 12484
rect 11348 12442 11376 13262
rect 11336 12436 11388 12442
rect 11336 12378 11388 12384
rect 10956 11452 11252 11472
rect 11012 11450 11036 11452
rect 11092 11450 11116 11452
rect 11172 11450 11196 11452
rect 11034 11398 11036 11450
rect 11098 11398 11110 11450
rect 11172 11398 11174 11450
rect 11012 11396 11036 11398
rect 11092 11396 11116 11398
rect 11172 11396 11196 11398
rect 10956 11376 11252 11396
rect 10956 10364 11252 10384
rect 11012 10362 11036 10364
rect 11092 10362 11116 10364
rect 11172 10362 11196 10364
rect 11034 10310 11036 10362
rect 11098 10310 11110 10362
rect 11172 10310 11174 10362
rect 11012 10308 11036 10310
rect 11092 10308 11116 10310
rect 11172 10308 11196 10310
rect 10956 10288 11252 10308
rect 10876 10124 10928 10130
rect 10876 10066 10928 10072
rect 10888 9625 10916 10066
rect 11244 10056 11296 10062
rect 11244 9998 11296 10004
rect 11256 9722 11284 9998
rect 11244 9716 11296 9722
rect 11244 9658 11296 9664
rect 10874 9616 10930 9625
rect 10874 9551 10930 9560
rect 10888 9382 10916 9551
rect 10876 9376 10928 9382
rect 11336 9376 11388 9382
rect 10876 9318 10928 9324
rect 11334 9344 11336 9353
rect 11388 9344 11390 9353
rect 10956 9276 11252 9296
rect 11334 9279 11390 9288
rect 11012 9274 11036 9276
rect 11092 9274 11116 9276
rect 11172 9274 11196 9276
rect 11034 9222 11036 9274
rect 11098 9222 11110 9274
rect 11172 9222 11174 9274
rect 11012 9220 11036 9222
rect 11092 9220 11116 9222
rect 11172 9220 11196 9222
rect 10956 9200 11252 9220
rect 11532 9042 11560 20810
rect 12728 20233 12756 23520
rect 12714 20224 12770 20233
rect 12714 20159 12770 20168
rect 14200 20097 14228 23520
rect 15660 22160 15712 22166
rect 15660 22102 15712 22108
rect 15382 20360 15438 20369
rect 15382 20295 15438 20304
rect 15566 20360 15622 20369
rect 15566 20295 15622 20304
rect 14280 20256 14332 20262
rect 14280 20198 14332 20204
rect 14186 20088 14242 20097
rect 14186 20023 14242 20032
rect 14292 19689 14320 20198
rect 15292 19916 15344 19922
rect 15292 19858 15344 19864
rect 14278 19680 14334 19689
rect 14278 19615 14334 19624
rect 15304 19446 15332 19858
rect 15396 19718 15424 20295
rect 15580 20262 15608 20295
rect 15568 20256 15620 20262
rect 15568 20198 15620 20204
rect 15474 19816 15530 19825
rect 15474 19751 15476 19760
rect 15528 19751 15530 19760
rect 15476 19722 15528 19728
rect 15384 19712 15436 19718
rect 15384 19654 15436 19660
rect 15292 19440 15344 19446
rect 15292 19382 15344 19388
rect 15568 19372 15620 19378
rect 15568 19314 15620 19320
rect 11702 17096 11758 17105
rect 11702 17031 11758 17040
rect 11612 13388 11664 13394
rect 11612 13330 11664 13336
rect 11624 12918 11652 13330
rect 11612 12912 11664 12918
rect 11612 12854 11664 12860
rect 11428 9036 11480 9042
rect 11428 8978 11480 8984
rect 11520 9036 11572 9042
rect 11520 8978 11572 8984
rect 10876 8832 10928 8838
rect 10876 8774 10928 8780
rect 10784 8560 10836 8566
rect 10782 8528 10784 8537
rect 10836 8528 10838 8537
rect 10782 8463 10838 8472
rect 10692 8356 10744 8362
rect 10692 8298 10744 8304
rect 10508 8016 10560 8022
rect 10508 7958 10560 7964
rect 10520 7342 10548 7958
rect 10704 7750 10732 8298
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 10692 7744 10744 7750
rect 10692 7686 10744 7692
rect 10508 7336 10560 7342
rect 10508 7278 10560 7284
rect 10520 6322 10548 7278
rect 10600 6860 10652 6866
rect 10600 6802 10652 6808
rect 10612 6458 10640 6802
rect 10600 6452 10652 6458
rect 10600 6394 10652 6400
rect 10508 6316 10560 6322
rect 10508 6258 10560 6264
rect 10520 5846 10548 6258
rect 10612 5914 10640 6394
rect 10704 5953 10732 7686
rect 10796 7206 10824 8230
rect 10888 8090 10916 8774
rect 11440 8294 11468 8978
rect 11532 8945 11560 8978
rect 11612 8968 11664 8974
rect 11518 8936 11574 8945
rect 11612 8910 11664 8916
rect 11518 8871 11574 8880
rect 11532 8566 11560 8871
rect 11520 8560 11572 8566
rect 11520 8502 11572 8508
rect 11624 8498 11652 8910
rect 11612 8492 11664 8498
rect 11612 8434 11664 8440
rect 11716 8362 11744 17031
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 12728 12782 12756 13126
rect 13818 13016 13874 13025
rect 13818 12951 13820 12960
rect 13872 12951 13874 12960
rect 13820 12922 13872 12928
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12716 12776 12768 12782
rect 12716 12718 12768 12724
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 12452 12646 12480 12718
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 12452 12442 12480 12582
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 12162 12200 12218 12209
rect 12162 12135 12218 12144
rect 12176 11218 12204 12135
rect 12348 11892 12400 11898
rect 12348 11834 12400 11840
rect 12164 11212 12216 11218
rect 12164 11154 12216 11160
rect 12176 10810 12204 11154
rect 12164 10804 12216 10810
rect 12084 10764 12164 10792
rect 11888 10600 11940 10606
rect 11888 10542 11940 10548
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11704 8356 11756 8362
rect 11704 8298 11756 8304
rect 11428 8288 11480 8294
rect 11428 8230 11480 8236
rect 10956 8188 11252 8208
rect 11012 8186 11036 8188
rect 11092 8186 11116 8188
rect 11172 8186 11196 8188
rect 11034 8134 11036 8186
rect 11098 8134 11110 8186
rect 11172 8134 11174 8186
rect 11012 8132 11036 8134
rect 11092 8132 11116 8134
rect 11172 8132 11196 8134
rect 10956 8112 11252 8132
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 11060 8016 11112 8022
rect 11808 7993 11836 10406
rect 11060 7958 11112 7964
rect 11610 7984 11666 7993
rect 11072 7449 11100 7958
rect 11336 7948 11388 7954
rect 11610 7919 11666 7928
rect 11794 7984 11850 7993
rect 11794 7919 11850 7928
rect 11336 7890 11388 7896
rect 11242 7712 11298 7721
rect 11242 7647 11298 7656
rect 11256 7449 11284 7647
rect 11058 7440 11114 7449
rect 11058 7375 11114 7384
rect 11242 7440 11298 7449
rect 11242 7375 11298 7384
rect 10784 7200 10836 7206
rect 10784 7142 10836 7148
rect 10956 7100 11252 7120
rect 11012 7098 11036 7100
rect 11092 7098 11116 7100
rect 11172 7098 11196 7100
rect 11034 7046 11036 7098
rect 11098 7046 11110 7098
rect 11172 7046 11174 7098
rect 11012 7044 11036 7046
rect 11092 7044 11116 7046
rect 11172 7044 11196 7046
rect 10782 7032 10838 7041
rect 10956 7024 11252 7044
rect 10782 6967 10784 6976
rect 10836 6967 10838 6976
rect 10784 6938 10836 6944
rect 10876 6860 10928 6866
rect 10876 6802 10928 6808
rect 10784 6656 10836 6662
rect 10784 6598 10836 6604
rect 10690 5944 10746 5953
rect 10600 5908 10652 5914
rect 10690 5879 10746 5888
rect 10600 5850 10652 5856
rect 10508 5840 10560 5846
rect 10796 5794 10824 6598
rect 10888 6186 10916 6802
rect 11348 6662 11376 7890
rect 11624 7002 11652 7919
rect 11612 6996 11664 7002
rect 11612 6938 11664 6944
rect 11336 6656 11388 6662
rect 11336 6598 11388 6604
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11426 6352 11482 6361
rect 11426 6287 11482 6296
rect 11060 6248 11112 6254
rect 11058 6216 11060 6225
rect 11336 6248 11388 6254
rect 11112 6216 11114 6225
rect 10876 6180 10928 6186
rect 11336 6190 11388 6196
rect 11058 6151 11114 6160
rect 10876 6122 10928 6128
rect 10508 5782 10560 5788
rect 10612 5766 10824 5794
rect 10414 4040 10470 4049
rect 10414 3975 10470 3984
rect 9956 3460 10008 3466
rect 9956 3402 10008 3408
rect 9772 3392 9824 3398
rect 9772 3334 9824 3340
rect 8668 3188 8720 3194
rect 8668 3130 8720 3136
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 8298 2952 8354 2961
rect 8298 2887 8354 2896
rect 8022 2615 8078 2624
rect 8208 2644 8260 2650
rect 8208 2586 8260 2592
rect 7104 2576 7156 2582
rect 7104 2518 7156 2524
rect 6920 2440 6972 2446
rect 6920 2382 6972 2388
rect 8312 2310 8340 2887
rect 9692 2650 9720 3130
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 9692 2446 9720 2586
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 7656 2304 7708 2310
rect 7656 2246 7708 2252
rect 8300 2304 8352 2310
rect 8300 2246 8352 2252
rect 7668 480 7696 2246
rect 8668 604 8720 610
rect 8668 546 8720 552
rect 8680 480 8708 546
rect 9784 480 9812 3334
rect 9968 3194 9996 3402
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 9968 2582 9996 3130
rect 9956 2576 10008 2582
rect 9956 2518 10008 2524
rect 10612 610 10640 5766
rect 10888 5642 10916 6122
rect 10956 6012 11252 6032
rect 11012 6010 11036 6012
rect 11092 6010 11116 6012
rect 11172 6010 11196 6012
rect 11034 5958 11036 6010
rect 11098 5958 11110 6010
rect 11172 5958 11174 6010
rect 11012 5956 11036 5958
rect 11092 5956 11116 5958
rect 11172 5956 11196 5958
rect 10956 5936 11252 5956
rect 11348 5914 11376 6190
rect 11440 6089 11468 6287
rect 11808 6254 11836 6598
rect 11900 6361 11928 10542
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 11886 6352 11942 6361
rect 11886 6287 11942 6296
rect 11796 6248 11848 6254
rect 11796 6190 11848 6196
rect 11888 6112 11940 6118
rect 11426 6080 11482 6089
rect 11992 6100 12020 6734
rect 11940 6072 12020 6100
rect 11888 6054 11940 6060
rect 11426 6015 11482 6024
rect 11336 5908 11388 5914
rect 11336 5850 11388 5856
rect 11704 5908 11756 5914
rect 11704 5850 11756 5856
rect 11336 5704 11388 5710
rect 11336 5646 11388 5652
rect 10876 5636 10928 5642
rect 10876 5578 10928 5584
rect 11348 5370 11376 5646
rect 11716 5370 11744 5850
rect 11336 5364 11388 5370
rect 11336 5306 11388 5312
rect 11704 5364 11756 5370
rect 11704 5306 11756 5312
rect 10956 4924 11252 4944
rect 11012 4922 11036 4924
rect 11092 4922 11116 4924
rect 11172 4922 11196 4924
rect 11034 4870 11036 4922
rect 11098 4870 11110 4922
rect 11172 4870 11174 4922
rect 11012 4868 11036 4870
rect 11092 4868 11116 4870
rect 11172 4868 11196 4870
rect 10956 4848 11252 4868
rect 10784 4752 10836 4758
rect 10784 4694 10836 4700
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 10704 4146 10732 4558
rect 10796 4282 10824 4694
rect 10784 4276 10836 4282
rect 10784 4218 10836 4224
rect 10692 4140 10744 4146
rect 10692 4082 10744 4088
rect 10704 3670 10732 4082
rect 10876 4072 10928 4078
rect 10876 4014 10928 4020
rect 10784 4004 10836 4010
rect 10784 3946 10836 3952
rect 10692 3664 10744 3670
rect 10692 3606 10744 3612
rect 10600 604 10652 610
rect 10600 546 10652 552
rect 10796 480 10824 3946
rect 10888 2650 10916 4014
rect 10956 3836 11252 3856
rect 11012 3834 11036 3836
rect 11092 3834 11116 3836
rect 11172 3834 11196 3836
rect 11034 3782 11036 3834
rect 11098 3782 11110 3834
rect 11172 3782 11174 3834
rect 11012 3780 11036 3782
rect 11092 3780 11116 3782
rect 11172 3780 11196 3782
rect 10956 3760 11252 3780
rect 11900 3505 11928 6054
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 11992 5574 12020 5714
rect 11980 5568 12032 5574
rect 11980 5510 12032 5516
rect 11992 5370 12020 5510
rect 11980 5364 12032 5370
rect 11980 5306 12032 5312
rect 12084 3641 12112 10764
rect 12164 10746 12216 10752
rect 12360 10713 12388 11834
rect 12346 10704 12402 10713
rect 12346 10639 12402 10648
rect 13924 10606 13952 12582
rect 15212 12306 15240 12718
rect 15200 12300 15252 12306
rect 15200 12242 15252 12248
rect 14280 12096 14332 12102
rect 14280 12038 14332 12044
rect 14292 11694 14320 12038
rect 14280 11688 14332 11694
rect 14280 11630 14332 11636
rect 15200 11688 15252 11694
rect 15200 11630 15252 11636
rect 14188 11552 14240 11558
rect 14188 11494 14240 11500
rect 14648 11552 14700 11558
rect 14648 11494 14700 11500
rect 13912 10600 13964 10606
rect 13912 10542 13964 10548
rect 12162 10296 12218 10305
rect 13924 10266 13952 10542
rect 14200 10266 14228 11494
rect 14660 11354 14688 11494
rect 14648 11348 14700 11354
rect 14648 11290 14700 11296
rect 15212 10810 15240 11630
rect 15476 11144 15528 11150
rect 15476 11086 15528 11092
rect 15200 10804 15252 10810
rect 15200 10746 15252 10752
rect 12162 10231 12218 10240
rect 13912 10260 13964 10266
rect 12176 9761 12204 10231
rect 13912 10202 13964 10208
rect 14188 10260 14240 10266
rect 14188 10202 14240 10208
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 13266 10024 13322 10033
rect 13266 9959 13322 9968
rect 13176 9920 13228 9926
rect 12254 9888 12310 9897
rect 13176 9862 13228 9868
rect 12254 9823 12310 9832
rect 12162 9752 12218 9761
rect 12268 9722 12296 9823
rect 13188 9722 13216 9862
rect 12162 9687 12218 9696
rect 12256 9716 12308 9722
rect 12176 6866 12204 9687
rect 12256 9658 12308 9664
rect 13176 9716 13228 9722
rect 13176 9658 13228 9664
rect 12900 8424 12952 8430
rect 12900 8366 12952 8372
rect 12256 8356 12308 8362
rect 12256 8298 12308 8304
rect 12268 8129 12296 8298
rect 12254 8120 12310 8129
rect 12254 8055 12310 8064
rect 12912 8022 12940 8366
rect 12900 8016 12952 8022
rect 12900 7958 12952 7964
rect 12164 6860 12216 6866
rect 12164 6802 12216 6808
rect 12176 6458 12204 6802
rect 12348 6724 12400 6730
rect 12348 6666 12400 6672
rect 12360 6497 12388 6666
rect 12900 6656 12952 6662
rect 12900 6598 12952 6604
rect 12346 6488 12402 6497
rect 12164 6452 12216 6458
rect 12346 6423 12402 6432
rect 12164 6394 12216 6400
rect 12912 6254 12940 6598
rect 12900 6248 12952 6254
rect 12900 6190 12952 6196
rect 12808 6112 12860 6118
rect 12808 6054 12860 6060
rect 12820 5914 12848 6054
rect 12912 5953 12940 6190
rect 12898 5944 12954 5953
rect 12808 5908 12860 5914
rect 12898 5879 12954 5888
rect 12808 5850 12860 5856
rect 13188 5846 13216 9658
rect 13280 5914 13308 9959
rect 13832 8650 13860 10066
rect 13924 9994 13952 10202
rect 13912 9988 13964 9994
rect 13912 9930 13964 9936
rect 14200 9518 14228 10202
rect 15108 10124 15160 10130
rect 15108 10066 15160 10072
rect 14556 9988 14608 9994
rect 14556 9930 14608 9936
rect 14464 9580 14516 9586
rect 14464 9522 14516 9528
rect 14188 9512 14240 9518
rect 14188 9454 14240 9460
rect 14372 9376 14424 9382
rect 14372 9318 14424 9324
rect 13740 8634 13860 8650
rect 13728 8628 13860 8634
rect 13780 8622 13860 8628
rect 13728 8570 13780 8576
rect 13728 7744 13780 7750
rect 13728 7686 13780 7692
rect 13358 7576 13414 7585
rect 13358 7511 13414 7520
rect 13372 7041 13400 7511
rect 13740 7274 13768 7686
rect 13728 7268 13780 7274
rect 13728 7210 13780 7216
rect 13452 7200 13504 7206
rect 13452 7142 13504 7148
rect 13358 7032 13414 7041
rect 13358 6967 13414 6976
rect 13372 6254 13400 6967
rect 13464 6662 13492 7142
rect 13452 6656 13504 6662
rect 13452 6598 13504 6604
rect 13464 6322 13492 6598
rect 13452 6316 13504 6322
rect 13452 6258 13504 6264
rect 13360 6248 13412 6254
rect 13360 6190 13412 6196
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 13176 5840 13228 5846
rect 13176 5782 13228 5788
rect 13188 5302 13216 5782
rect 13280 5370 13308 5850
rect 13464 5710 13492 6258
rect 13740 6118 13768 7210
rect 13832 6458 13860 8622
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 13728 6112 13780 6118
rect 13728 6054 13780 6060
rect 13452 5704 13504 5710
rect 13452 5646 13504 5652
rect 13464 5370 13492 5646
rect 13268 5364 13320 5370
rect 13268 5306 13320 5312
rect 13452 5364 13504 5370
rect 13452 5306 13504 5312
rect 13176 5296 13228 5302
rect 13176 5238 13228 5244
rect 12440 4480 12492 4486
rect 13820 4480 13872 4486
rect 12440 4422 12492 4428
rect 13740 4428 13820 4434
rect 13740 4422 13872 4428
rect 12452 3670 12480 4422
rect 13740 4406 13860 4422
rect 12440 3664 12492 3670
rect 12070 3632 12126 3641
rect 12440 3606 12492 3612
rect 12070 3567 12126 3576
rect 11886 3496 11942 3505
rect 11886 3431 11942 3440
rect 11336 3392 11388 3398
rect 11336 3334 11388 3340
rect 11348 3194 11376 3334
rect 11886 3224 11942 3233
rect 11336 3188 11388 3194
rect 12452 3194 12480 3606
rect 13740 3466 13768 4406
rect 13728 3460 13780 3466
rect 13728 3402 13780 3408
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 13820 3392 13872 3398
rect 13820 3334 13872 3340
rect 11886 3159 11888 3168
rect 11336 3130 11388 3136
rect 11940 3159 11942 3168
rect 12440 3188 12492 3194
rect 11888 3130 11940 3136
rect 12440 3130 12492 3136
rect 11900 2990 11928 3130
rect 11888 2984 11940 2990
rect 11888 2926 11940 2932
rect 11704 2848 11756 2854
rect 11704 2790 11756 2796
rect 10956 2748 11252 2768
rect 11012 2746 11036 2748
rect 11092 2746 11116 2748
rect 11172 2746 11196 2748
rect 11034 2694 11036 2746
rect 11098 2694 11110 2746
rect 11172 2694 11174 2746
rect 11012 2692 11036 2694
rect 11092 2692 11116 2694
rect 11172 2692 11196 2694
rect 10956 2672 11252 2692
rect 10876 2644 10928 2650
rect 10876 2586 10928 2592
rect 11716 1442 11744 2790
rect 12452 2650 12480 3130
rect 12636 2854 12664 3334
rect 13832 3233 13860 3334
rect 13818 3224 13874 3233
rect 13818 3159 13874 3168
rect 12808 3120 12860 3126
rect 14384 3097 14412 9318
rect 14476 9178 14504 9522
rect 14464 9172 14516 9178
rect 14464 9114 14516 9120
rect 14568 9042 14596 9930
rect 15120 9586 15148 10066
rect 15212 10062 15240 10746
rect 15200 10056 15252 10062
rect 15200 9998 15252 10004
rect 15108 9580 15160 9586
rect 15108 9522 15160 9528
rect 15212 9518 15240 9998
rect 15488 9926 15516 11086
rect 15476 9920 15528 9926
rect 15476 9862 15528 9868
rect 15200 9512 15252 9518
rect 15200 9454 15252 9460
rect 14924 9444 14976 9450
rect 14924 9386 14976 9392
rect 14936 9217 14964 9386
rect 14922 9208 14978 9217
rect 14922 9143 14978 9152
rect 15212 9110 15240 9454
rect 15200 9104 15252 9110
rect 15200 9046 15252 9052
rect 14556 9036 14608 9042
rect 14556 8978 14608 8984
rect 15016 9036 15068 9042
rect 15016 8978 15068 8984
rect 15028 8634 15056 8978
rect 15212 8634 15240 9046
rect 15488 8673 15516 9862
rect 15474 8664 15530 8673
rect 15016 8628 15068 8634
rect 15016 8570 15068 8576
rect 15200 8628 15252 8634
rect 15474 8599 15530 8608
rect 15200 8570 15252 8576
rect 15476 8492 15528 8498
rect 15476 8434 15528 8440
rect 14738 8120 14794 8129
rect 14738 8055 14794 8064
rect 14752 7546 14780 8055
rect 14740 7540 14792 7546
rect 14740 7482 14792 7488
rect 15488 7313 15516 8434
rect 15474 7304 15530 7313
rect 15474 7239 15530 7248
rect 15476 6656 15528 6662
rect 15476 6598 15528 6604
rect 14556 6112 14608 6118
rect 14556 6054 14608 6060
rect 14568 5166 14596 6054
rect 15384 5568 15436 5574
rect 15384 5510 15436 5516
rect 14556 5160 14608 5166
rect 15396 5137 15424 5510
rect 15488 5273 15516 6598
rect 15474 5264 15530 5273
rect 15474 5199 15530 5208
rect 14556 5102 14608 5108
rect 15382 5128 15438 5137
rect 14568 4690 14596 5102
rect 15382 5063 15438 5072
rect 14556 4684 14608 4690
rect 14556 4626 14608 4632
rect 14568 4486 14596 4626
rect 14556 4480 14608 4486
rect 14556 4422 14608 4428
rect 12808 3062 12860 3068
rect 14370 3088 14426 3097
rect 12624 2848 12676 2854
rect 12624 2790 12676 2796
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 12636 2514 12664 2790
rect 12624 2508 12676 2514
rect 12624 2450 12676 2456
rect 11716 1414 11836 1442
rect 11808 480 11836 1414
rect 12820 480 12848 3062
rect 14370 3023 14426 3032
rect 13176 2984 13228 2990
rect 13174 2952 13176 2961
rect 14004 2984 14056 2990
rect 13228 2952 13230 2961
rect 14004 2926 14056 2932
rect 13174 2887 13230 2896
rect 13360 2848 13412 2854
rect 13358 2816 13360 2825
rect 13912 2848 13964 2854
rect 13412 2816 13414 2825
rect 13912 2790 13964 2796
rect 13358 2751 13414 2760
rect 13924 480 13952 2790
rect 14016 2650 14044 2926
rect 14922 2816 14978 2825
rect 14922 2751 14978 2760
rect 14004 2644 14056 2650
rect 14004 2586 14056 2592
rect 14936 480 14964 2751
rect 15580 2514 15608 19314
rect 15672 11354 15700 22102
rect 15764 19378 15792 23520
rect 17236 23474 17264 23520
rect 18708 23474 18736 23520
rect 17236 23446 17356 23474
rect 17328 22114 17356 23446
rect 17144 22086 17356 22114
rect 18156 23446 18736 23474
rect 15956 21788 16252 21808
rect 16012 21786 16036 21788
rect 16092 21786 16116 21788
rect 16172 21786 16196 21788
rect 16034 21734 16036 21786
rect 16098 21734 16110 21786
rect 16172 21734 16174 21786
rect 16012 21732 16036 21734
rect 16092 21732 16116 21734
rect 16172 21732 16196 21734
rect 15956 21712 16252 21732
rect 15956 20700 16252 20720
rect 16012 20698 16036 20700
rect 16092 20698 16116 20700
rect 16172 20698 16196 20700
rect 16034 20646 16036 20698
rect 16098 20646 16110 20698
rect 16172 20646 16174 20698
rect 16012 20644 16036 20646
rect 16092 20644 16116 20646
rect 16172 20644 16196 20646
rect 15956 20624 16252 20644
rect 16672 20528 16724 20534
rect 16302 20496 16358 20505
rect 16302 20431 16358 20440
rect 16670 20496 16672 20505
rect 16724 20496 16726 20505
rect 16670 20431 16726 20440
rect 16316 19825 16344 20431
rect 16396 20256 16448 20262
rect 16396 20198 16448 20204
rect 17040 20256 17092 20262
rect 17040 20198 17092 20204
rect 16302 19816 16358 19825
rect 16302 19751 16358 19760
rect 15956 19612 16252 19632
rect 16012 19610 16036 19612
rect 16092 19610 16116 19612
rect 16172 19610 16196 19612
rect 16034 19558 16036 19610
rect 16098 19558 16110 19610
rect 16172 19558 16174 19610
rect 16012 19556 16036 19558
rect 16092 19556 16116 19558
rect 16172 19556 16196 19558
rect 15956 19536 16252 19556
rect 15752 19372 15804 19378
rect 15752 19314 15804 19320
rect 15956 18524 16252 18544
rect 16012 18522 16036 18524
rect 16092 18522 16116 18524
rect 16172 18522 16196 18524
rect 16034 18470 16036 18522
rect 16098 18470 16110 18522
rect 16172 18470 16174 18522
rect 16012 18468 16036 18470
rect 16092 18468 16116 18470
rect 16172 18468 16196 18470
rect 15956 18448 16252 18468
rect 15956 17436 16252 17456
rect 16012 17434 16036 17436
rect 16092 17434 16116 17436
rect 16172 17434 16196 17436
rect 16034 17382 16036 17434
rect 16098 17382 16110 17434
rect 16172 17382 16174 17434
rect 16012 17380 16036 17382
rect 16092 17380 16116 17382
rect 16172 17380 16196 17382
rect 15956 17360 16252 17380
rect 15956 16348 16252 16368
rect 16012 16346 16036 16348
rect 16092 16346 16116 16348
rect 16172 16346 16196 16348
rect 16034 16294 16036 16346
rect 16098 16294 16110 16346
rect 16172 16294 16174 16346
rect 16012 16292 16036 16294
rect 16092 16292 16116 16294
rect 16172 16292 16196 16294
rect 15956 16272 16252 16292
rect 15956 15260 16252 15280
rect 16012 15258 16036 15260
rect 16092 15258 16116 15260
rect 16172 15258 16196 15260
rect 16034 15206 16036 15258
rect 16098 15206 16110 15258
rect 16172 15206 16174 15258
rect 16012 15204 16036 15206
rect 16092 15204 16116 15206
rect 16172 15204 16196 15206
rect 15956 15184 16252 15204
rect 16302 14512 16358 14521
rect 16408 14498 16436 20198
rect 16580 20052 16632 20058
rect 16580 19994 16632 20000
rect 16592 19961 16620 19994
rect 16578 19952 16634 19961
rect 16488 19916 16540 19922
rect 16578 19887 16634 19896
rect 16488 19858 16540 19864
rect 16500 19378 16528 19858
rect 16580 19712 16632 19718
rect 16578 19680 16580 19689
rect 16632 19680 16634 19689
rect 16578 19615 16634 19624
rect 17052 19446 17080 20198
rect 17040 19440 17092 19446
rect 17040 19382 17092 19388
rect 16488 19372 16540 19378
rect 16488 19314 16540 19320
rect 16948 19304 17000 19310
rect 16948 19246 17000 19252
rect 16408 14470 16620 14498
rect 16302 14447 16358 14456
rect 15956 14172 16252 14192
rect 16012 14170 16036 14172
rect 16092 14170 16116 14172
rect 16172 14170 16196 14172
rect 16034 14118 16036 14170
rect 16098 14118 16110 14170
rect 16172 14118 16174 14170
rect 16012 14116 16036 14118
rect 16092 14116 16116 14118
rect 16172 14116 16196 14118
rect 15956 14096 16252 14116
rect 15956 13084 16252 13104
rect 16012 13082 16036 13084
rect 16092 13082 16116 13084
rect 16172 13082 16196 13084
rect 16034 13030 16036 13082
rect 16098 13030 16110 13082
rect 16172 13030 16174 13082
rect 16012 13028 16036 13030
rect 16092 13028 16116 13030
rect 16172 13028 16196 13030
rect 15956 13008 16252 13028
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 15764 11694 15792 12174
rect 15956 11996 16252 12016
rect 16012 11994 16036 11996
rect 16092 11994 16116 11996
rect 16172 11994 16196 11996
rect 16034 11942 16036 11994
rect 16098 11942 16110 11994
rect 16172 11942 16174 11994
rect 16012 11940 16036 11942
rect 16092 11940 16116 11942
rect 16172 11940 16196 11942
rect 15956 11920 16252 11940
rect 15752 11688 15804 11694
rect 15752 11630 15804 11636
rect 16212 11620 16264 11626
rect 16212 11562 16264 11568
rect 15660 11348 15712 11354
rect 15660 11290 15712 11296
rect 15672 10810 15700 11290
rect 16224 11121 16252 11562
rect 16316 11218 16344 14447
rect 16592 12356 16620 14470
rect 16672 12640 16724 12646
rect 16672 12582 16724 12588
rect 16684 12374 16712 12582
rect 16500 12328 16620 12356
rect 16672 12368 16724 12374
rect 16396 11756 16448 11762
rect 16396 11698 16448 11704
rect 16304 11212 16356 11218
rect 16304 11154 16356 11160
rect 16408 11150 16436 11698
rect 16396 11144 16448 11150
rect 16210 11112 16266 11121
rect 16396 11086 16448 11092
rect 16210 11047 16266 11056
rect 16408 11014 16436 11086
rect 16396 11008 16448 11014
rect 16396 10950 16448 10956
rect 15956 10908 16252 10928
rect 16012 10906 16036 10908
rect 16092 10906 16116 10908
rect 16172 10906 16196 10908
rect 16034 10854 16036 10906
rect 16098 10854 16110 10906
rect 16172 10854 16174 10906
rect 16012 10852 16036 10854
rect 16092 10852 16116 10854
rect 16172 10852 16196 10854
rect 15956 10832 16252 10852
rect 15660 10804 15712 10810
rect 15660 10746 15712 10752
rect 15672 10713 15700 10746
rect 16408 10742 16436 10950
rect 16396 10736 16448 10742
rect 15658 10704 15714 10713
rect 16396 10678 16448 10684
rect 15658 10639 15714 10648
rect 16396 10464 16448 10470
rect 16396 10406 16448 10412
rect 16408 10266 16436 10406
rect 16396 10260 16448 10266
rect 16396 10202 16448 10208
rect 16304 10124 16356 10130
rect 16304 10066 16356 10072
rect 15660 9920 15712 9926
rect 15660 9862 15712 9868
rect 15672 9722 15700 9862
rect 15956 9820 16252 9840
rect 16012 9818 16036 9820
rect 16092 9818 16116 9820
rect 16172 9818 16196 9820
rect 16034 9766 16036 9818
rect 16098 9766 16110 9818
rect 16172 9766 16174 9818
rect 16012 9764 16036 9766
rect 16092 9764 16116 9766
rect 16172 9764 16196 9766
rect 15956 9744 16252 9764
rect 15660 9716 15712 9722
rect 15660 9658 15712 9664
rect 16316 9654 16344 10066
rect 16408 9722 16436 10202
rect 16396 9716 16448 9722
rect 16396 9658 16448 9664
rect 16304 9648 16356 9654
rect 16304 9590 16356 9596
rect 15956 8732 16252 8752
rect 16012 8730 16036 8732
rect 16092 8730 16116 8732
rect 16172 8730 16196 8732
rect 16034 8678 16036 8730
rect 16098 8678 16110 8730
rect 16172 8678 16174 8730
rect 16012 8676 16036 8678
rect 16092 8676 16116 8678
rect 16172 8676 16196 8678
rect 15956 8656 16252 8676
rect 16396 8288 16448 8294
rect 16396 8230 16448 8236
rect 16304 7744 16356 7750
rect 16304 7686 16356 7692
rect 15956 7644 16252 7664
rect 16012 7642 16036 7644
rect 16092 7642 16116 7644
rect 16172 7642 16196 7644
rect 16034 7590 16036 7642
rect 16098 7590 16110 7642
rect 16172 7590 16174 7642
rect 16012 7588 16036 7590
rect 16092 7588 16116 7590
rect 16172 7588 16196 7590
rect 15956 7568 16252 7588
rect 16316 7410 16344 7686
rect 16304 7404 16356 7410
rect 16304 7346 16356 7352
rect 15936 7336 15988 7342
rect 15936 7278 15988 7284
rect 15844 7200 15896 7206
rect 15844 7142 15896 7148
rect 15856 5914 15884 7142
rect 15948 7002 15976 7278
rect 16408 7274 16436 8230
rect 16396 7268 16448 7274
rect 16396 7210 16448 7216
rect 15936 6996 15988 7002
rect 15936 6938 15988 6944
rect 16396 6996 16448 7002
rect 16396 6938 16448 6944
rect 15956 6556 16252 6576
rect 16012 6554 16036 6556
rect 16092 6554 16116 6556
rect 16172 6554 16196 6556
rect 16034 6502 16036 6554
rect 16098 6502 16110 6554
rect 16172 6502 16174 6554
rect 16012 6500 16036 6502
rect 16092 6500 16116 6502
rect 16172 6500 16196 6502
rect 15956 6480 16252 6500
rect 15844 5908 15896 5914
rect 15844 5850 15896 5856
rect 15844 5704 15896 5710
rect 15844 5646 15896 5652
rect 16304 5704 16356 5710
rect 16304 5646 16356 5652
rect 15856 4842 15884 5646
rect 15956 5468 16252 5488
rect 16012 5466 16036 5468
rect 16092 5466 16116 5468
rect 16172 5466 16196 5468
rect 16034 5414 16036 5466
rect 16098 5414 16110 5466
rect 16172 5414 16174 5466
rect 16012 5412 16036 5414
rect 16092 5412 16116 5414
rect 16172 5412 16196 5414
rect 15956 5392 16252 5412
rect 16316 5098 16344 5646
rect 16304 5092 16356 5098
rect 16304 5034 16356 5040
rect 15934 4856 15990 4865
rect 15856 4814 15934 4842
rect 15934 4791 15936 4800
rect 15988 4791 15990 4800
rect 15936 4762 15988 4768
rect 15844 4684 15896 4690
rect 15844 4626 15896 4632
rect 15856 4214 15884 4626
rect 16316 4486 16344 5034
rect 16408 4758 16436 6938
rect 16396 4752 16448 4758
rect 16396 4694 16448 4700
rect 16304 4480 16356 4486
rect 16304 4422 16356 4428
rect 15956 4380 16252 4400
rect 16012 4378 16036 4380
rect 16092 4378 16116 4380
rect 16172 4378 16196 4380
rect 16034 4326 16036 4378
rect 16098 4326 16110 4378
rect 16172 4326 16174 4378
rect 16012 4324 16036 4326
rect 16092 4324 16116 4326
rect 16172 4324 16196 4326
rect 15956 4304 16252 4324
rect 16408 4282 16436 4694
rect 16396 4276 16448 4282
rect 16396 4218 16448 4224
rect 15844 4208 15896 4214
rect 15844 4150 15896 4156
rect 15956 3292 16252 3312
rect 16012 3290 16036 3292
rect 16092 3290 16116 3292
rect 16172 3290 16196 3292
rect 16034 3238 16036 3290
rect 16098 3238 16110 3290
rect 16172 3238 16174 3290
rect 16012 3236 16036 3238
rect 16092 3236 16116 3238
rect 16172 3236 16196 3238
rect 15956 3216 16252 3236
rect 15568 2508 15620 2514
rect 15568 2450 15620 2456
rect 15660 2304 15712 2310
rect 15660 2246 15712 2252
rect 15672 2009 15700 2246
rect 15956 2204 16252 2224
rect 16012 2202 16036 2204
rect 16092 2202 16116 2204
rect 16172 2202 16196 2204
rect 16034 2150 16036 2202
rect 16098 2150 16110 2202
rect 16172 2150 16174 2202
rect 16012 2148 16036 2150
rect 16092 2148 16116 2150
rect 16172 2148 16196 2150
rect 15956 2128 16252 2148
rect 16500 2038 16528 12328
rect 16672 12310 16724 12316
rect 16856 11076 16908 11082
rect 16856 11018 16908 11024
rect 16868 10674 16896 11018
rect 16856 10668 16908 10674
rect 16856 10610 16908 10616
rect 16580 10600 16632 10606
rect 16580 10542 16632 10548
rect 16592 10033 16620 10542
rect 16578 10024 16634 10033
rect 16578 9959 16634 9968
rect 16960 9722 16988 19246
rect 16948 9716 17000 9722
rect 16948 9658 17000 9664
rect 16670 9208 16726 9217
rect 16670 9143 16672 9152
rect 16724 9143 16726 9152
rect 16672 9114 16724 9120
rect 16762 8664 16818 8673
rect 16762 8599 16818 8608
rect 16776 8498 16804 8599
rect 16764 8492 16816 8498
rect 16764 8434 16816 8440
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 16868 7886 16896 8434
rect 16948 7948 17000 7954
rect 16948 7890 17000 7896
rect 16764 7880 16816 7886
rect 16764 7822 16816 7828
rect 16856 7880 16908 7886
rect 16960 7857 16988 7890
rect 16856 7822 16908 7828
rect 16946 7848 17002 7857
rect 16776 6934 16804 7822
rect 16868 7478 16896 7822
rect 16946 7783 17002 7792
rect 16856 7472 16908 7478
rect 16856 7414 16908 7420
rect 16868 6934 16896 7414
rect 16960 7342 16988 7783
rect 16948 7336 17000 7342
rect 16946 7304 16948 7313
rect 17000 7304 17002 7313
rect 16946 7239 17002 7248
rect 16764 6928 16816 6934
rect 16764 6870 16816 6876
rect 16856 6928 16908 6934
rect 16856 6870 16908 6876
rect 16672 6792 16724 6798
rect 16672 6734 16724 6740
rect 16684 6118 16712 6734
rect 16868 6458 16896 6870
rect 16856 6452 16908 6458
rect 16856 6394 16908 6400
rect 16672 6112 16724 6118
rect 16672 6054 16724 6060
rect 16580 5908 16632 5914
rect 16580 5850 16632 5856
rect 16592 5370 16620 5850
rect 16580 5364 16632 5370
rect 16580 5306 16632 5312
rect 16684 4690 16712 6054
rect 16672 4684 16724 4690
rect 16672 4626 16724 4632
rect 17052 2802 17080 19382
rect 17144 19310 17172 22086
rect 18050 19544 18106 19553
rect 18050 19479 18106 19488
rect 17132 19304 17184 19310
rect 17132 19246 17184 19252
rect 17498 15328 17554 15337
rect 17498 15263 17554 15272
rect 17408 12368 17460 12374
rect 17408 12310 17460 12316
rect 17316 12300 17368 12306
rect 17316 12242 17368 12248
rect 17328 11898 17356 12242
rect 17316 11892 17368 11898
rect 17316 11834 17368 11840
rect 17420 11830 17448 12310
rect 17408 11824 17460 11830
rect 17408 11766 17460 11772
rect 17420 11286 17448 11766
rect 17408 11280 17460 11286
rect 17408 11222 17460 11228
rect 17130 10976 17186 10985
rect 17130 10911 17186 10920
rect 17144 10305 17172 10911
rect 17314 10840 17370 10849
rect 17314 10775 17370 10784
rect 17328 10674 17356 10775
rect 17316 10668 17368 10674
rect 17316 10610 17368 10616
rect 17130 10296 17186 10305
rect 17420 10282 17448 11222
rect 17130 10231 17186 10240
rect 17328 10254 17448 10282
rect 17224 9716 17276 9722
rect 17224 9658 17276 9664
rect 17052 2774 17172 2802
rect 17144 2666 17172 2774
rect 16960 2638 17172 2666
rect 17236 2650 17264 9658
rect 17328 9518 17356 10254
rect 17406 10160 17462 10169
rect 17406 10095 17462 10104
rect 17420 9586 17448 10095
rect 17408 9580 17460 9586
rect 17408 9522 17460 9528
rect 17316 9512 17368 9518
rect 17316 9454 17368 9460
rect 17512 7818 17540 15263
rect 17960 11144 18012 11150
rect 17960 11086 18012 11092
rect 17868 10804 17920 10810
rect 17972 10792 18000 11086
rect 17920 10764 18000 10792
rect 17868 10746 17920 10752
rect 17868 10464 17920 10470
rect 17868 10406 17920 10412
rect 17880 10266 17908 10406
rect 17868 10260 17920 10266
rect 17868 10202 17920 10208
rect 17868 9920 17920 9926
rect 17868 9862 17920 9868
rect 17880 9602 17908 9862
rect 17880 9586 18000 9602
rect 17880 9580 18012 9586
rect 17880 9574 17960 9580
rect 17960 9522 18012 9528
rect 17774 9480 17830 9489
rect 17774 9415 17776 9424
rect 17828 9415 17830 9424
rect 17776 9386 17828 9392
rect 17868 8356 17920 8362
rect 17868 8298 17920 8304
rect 17880 8090 17908 8298
rect 17868 8084 17920 8090
rect 17868 8026 17920 8032
rect 17500 7812 17552 7818
rect 17500 7754 17552 7760
rect 17960 7540 18012 7546
rect 17960 7482 18012 7488
rect 17224 2644 17276 2650
rect 15936 2032 15988 2038
rect 15658 2000 15714 2009
rect 15936 1974 15988 1980
rect 16488 2032 16540 2038
rect 16488 1974 16540 1980
rect 15658 1935 15714 1944
rect 15948 480 15976 1974
rect 16960 480 16988 2638
rect 17224 2586 17276 2592
rect 17868 2304 17920 2310
rect 17868 2246 17920 2252
rect 17880 1465 17908 2246
rect 17972 2122 18000 7482
rect 18064 2258 18092 19479
rect 18156 14498 18184 23446
rect 18234 20632 18290 20641
rect 18234 20567 18236 20576
rect 18288 20567 18290 20576
rect 18236 20538 18288 20544
rect 20180 20398 20208 23520
rect 20956 21244 21252 21264
rect 21012 21242 21036 21244
rect 21092 21242 21116 21244
rect 21172 21242 21196 21244
rect 21034 21190 21036 21242
rect 21098 21190 21110 21242
rect 21172 21190 21174 21242
rect 21012 21188 21036 21190
rect 21092 21188 21116 21190
rect 21172 21188 21196 21190
rect 20956 21168 21252 21188
rect 19984 20392 20036 20398
rect 19984 20334 20036 20340
rect 20168 20392 20220 20398
rect 20168 20334 20220 20340
rect 20628 20392 20680 20398
rect 20628 20334 20680 20340
rect 20812 20392 20864 20398
rect 21744 20369 21772 23520
rect 23216 20505 23244 23520
rect 24688 20641 24716 23520
rect 25502 22400 25558 22409
rect 25502 22335 25558 22344
rect 25410 21584 25466 21593
rect 25410 21519 25466 21528
rect 25424 20806 25452 21519
rect 25412 20800 25464 20806
rect 25412 20742 25464 20748
rect 24674 20632 24730 20641
rect 24674 20567 24730 20576
rect 23202 20496 23258 20505
rect 23202 20431 23258 20440
rect 24216 20392 24268 20398
rect 20812 20334 20864 20340
rect 21730 20360 21786 20369
rect 19156 20256 19208 20262
rect 19996 20233 20024 20334
rect 20168 20256 20220 20262
rect 19156 20198 19208 20204
rect 19982 20224 20038 20233
rect 19168 19378 19196 20198
rect 20168 20198 20220 20204
rect 19982 20159 20038 20168
rect 19522 19680 19578 19689
rect 19522 19615 19578 19624
rect 19156 19372 19208 19378
rect 19156 19314 19208 19320
rect 18156 14470 18276 14498
rect 18144 10124 18196 10130
rect 18144 10066 18196 10072
rect 18156 8838 18184 10066
rect 18144 8832 18196 8838
rect 18144 8774 18196 8780
rect 18144 6656 18196 6662
rect 18144 6598 18196 6604
rect 18156 5234 18184 6598
rect 18144 5228 18196 5234
rect 18144 5170 18196 5176
rect 18156 4758 18184 5170
rect 18144 4752 18196 4758
rect 18144 4694 18196 4700
rect 18142 3598 18198 3607
rect 18142 3533 18198 3542
rect 18248 2553 18276 14470
rect 18326 13832 18382 13841
rect 18326 13767 18382 13776
rect 18340 10266 18368 13767
rect 18696 12096 18748 12102
rect 18696 12038 18748 12044
rect 18604 11144 18656 11150
rect 18604 11086 18656 11092
rect 18616 10674 18644 11086
rect 18708 10849 18736 12038
rect 19064 11076 19116 11082
rect 19064 11018 19116 11024
rect 18694 10840 18750 10849
rect 18694 10775 18750 10784
rect 18604 10668 18656 10674
rect 18604 10610 18656 10616
rect 18420 10464 18472 10470
rect 18420 10406 18472 10412
rect 18328 10260 18380 10266
rect 18328 10202 18380 10208
rect 18326 10160 18382 10169
rect 18326 10095 18328 10104
rect 18380 10095 18382 10104
rect 18328 10066 18380 10072
rect 18432 9994 18460 10406
rect 18616 10062 18644 10610
rect 18604 10056 18656 10062
rect 18604 9998 18656 10004
rect 18420 9988 18472 9994
rect 18420 9930 18472 9936
rect 18708 9586 18736 10775
rect 18880 10464 18932 10470
rect 18880 10406 18932 10412
rect 18696 9580 18748 9586
rect 18696 9522 18748 9528
rect 18328 9104 18380 9110
rect 18328 9046 18380 9052
rect 18340 8634 18368 9046
rect 18420 9036 18472 9042
rect 18420 8978 18472 8984
rect 18328 8628 18380 8634
rect 18328 8570 18380 8576
rect 18432 8498 18460 8978
rect 18604 8832 18656 8838
rect 18604 8774 18656 8780
rect 18420 8492 18472 8498
rect 18420 8434 18472 8440
rect 18432 8090 18460 8434
rect 18420 8084 18472 8090
rect 18420 8026 18472 8032
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 18420 6112 18472 6118
rect 18420 6054 18472 6060
rect 18432 5030 18460 6054
rect 18524 5914 18552 6258
rect 18512 5908 18564 5914
rect 18512 5850 18564 5856
rect 18328 5024 18380 5030
rect 18328 4966 18380 4972
rect 18420 5024 18472 5030
rect 18420 4966 18472 4972
rect 18340 4865 18368 4966
rect 18326 4856 18382 4865
rect 18326 4791 18382 4800
rect 18616 4185 18644 8774
rect 18788 5160 18840 5166
rect 18788 5102 18840 5108
rect 18800 4826 18828 5102
rect 18788 4820 18840 4826
rect 18788 4762 18840 4768
rect 18602 4176 18658 4185
rect 18602 4111 18658 4120
rect 18234 2544 18290 2553
rect 18892 2514 18920 10406
rect 18970 10024 19026 10033
rect 18970 9959 18972 9968
rect 19024 9959 19026 9968
rect 18972 9930 19024 9936
rect 19076 7041 19104 11018
rect 19168 7546 19196 19314
rect 19536 14498 19564 19615
rect 19444 14470 19564 14498
rect 19246 12880 19302 12889
rect 19246 12815 19302 12824
rect 19260 11354 19288 12815
rect 19444 12374 19472 14470
rect 20180 12481 20208 20198
rect 20640 14498 20668 20334
rect 20824 20097 20852 20334
rect 24216 20334 24268 20340
rect 24398 20360 24454 20369
rect 21730 20295 21786 20304
rect 21272 20256 21324 20262
rect 21272 20198 21324 20204
rect 20956 20156 21252 20176
rect 21012 20154 21036 20156
rect 21092 20154 21116 20156
rect 21172 20154 21196 20156
rect 21034 20102 21036 20154
rect 21098 20102 21110 20154
rect 21172 20102 21174 20154
rect 21012 20100 21036 20102
rect 21092 20100 21116 20102
rect 21172 20100 21196 20102
rect 20810 20088 20866 20097
rect 20956 20080 21252 20100
rect 20810 20023 20866 20032
rect 20956 19068 21252 19088
rect 21012 19066 21036 19068
rect 21092 19066 21116 19068
rect 21172 19066 21196 19068
rect 21034 19014 21036 19066
rect 21098 19014 21110 19066
rect 21172 19014 21174 19066
rect 21012 19012 21036 19014
rect 21092 19012 21116 19014
rect 21172 19012 21196 19014
rect 20956 18992 21252 19012
rect 20718 18728 20774 18737
rect 20718 18663 20774 18672
rect 20548 14470 20668 14498
rect 20166 12472 20222 12481
rect 20166 12407 20222 12416
rect 19432 12368 19484 12374
rect 19432 12310 19484 12316
rect 20076 12368 20128 12374
rect 20076 12310 20128 12316
rect 20258 12336 20314 12345
rect 19248 11348 19300 11354
rect 19248 11290 19300 11296
rect 19260 10810 19288 11290
rect 19248 10804 19300 10810
rect 19248 10746 19300 10752
rect 19156 7540 19208 7546
rect 19156 7482 19208 7488
rect 19062 7032 19118 7041
rect 19062 6967 19118 6976
rect 18972 6452 19024 6458
rect 18972 6394 19024 6400
rect 18984 6322 19012 6394
rect 18972 6316 19024 6322
rect 18972 6258 19024 6264
rect 18984 5710 19012 6258
rect 18972 5704 19024 5710
rect 18972 5646 19024 5652
rect 19076 2990 19104 6967
rect 19260 6440 19288 10746
rect 19982 9344 20038 9353
rect 19982 9279 20038 9288
rect 19524 8832 19576 8838
rect 19524 8774 19576 8780
rect 19536 8362 19564 8774
rect 19996 8401 20024 9279
rect 19982 8392 20038 8401
rect 19524 8356 19576 8362
rect 19982 8327 20038 8336
rect 19524 8298 19576 8304
rect 19340 7472 19392 7478
rect 19340 7414 19392 7420
rect 19168 6412 19288 6440
rect 19168 5953 19196 6412
rect 19352 6338 19380 7414
rect 19536 7410 19564 8298
rect 19996 8090 20024 8327
rect 19984 8084 20036 8090
rect 19984 8026 20036 8032
rect 19890 7984 19946 7993
rect 19890 7919 19946 7928
rect 19524 7404 19576 7410
rect 19524 7346 19576 7352
rect 19904 6866 19932 7919
rect 19996 7342 20024 8026
rect 19984 7336 20036 7342
rect 19984 7278 20036 7284
rect 19984 7200 20036 7206
rect 19984 7142 20036 7148
rect 19892 6860 19944 6866
rect 19892 6802 19944 6808
rect 19614 6760 19670 6769
rect 19614 6695 19670 6704
rect 19260 6310 19380 6338
rect 19260 6254 19288 6310
rect 19248 6248 19300 6254
rect 19248 6190 19300 6196
rect 19154 5944 19210 5953
rect 19628 5914 19656 6695
rect 19798 6352 19854 6361
rect 19798 6287 19800 6296
rect 19852 6287 19854 6296
rect 19800 6258 19852 6264
rect 19904 6186 19932 6802
rect 19892 6180 19944 6186
rect 19892 6122 19944 6128
rect 19154 5879 19210 5888
rect 19616 5908 19668 5914
rect 19616 5850 19668 5856
rect 19248 5568 19300 5574
rect 19248 5510 19300 5516
rect 19260 5166 19288 5510
rect 19628 5302 19656 5850
rect 19708 5704 19760 5710
rect 19708 5646 19760 5652
rect 19720 5370 19748 5646
rect 19708 5364 19760 5370
rect 19708 5306 19760 5312
rect 19616 5296 19668 5302
rect 19996 5273 20024 7142
rect 19616 5238 19668 5244
rect 19982 5264 20038 5273
rect 19248 5160 19300 5166
rect 19628 5137 19656 5238
rect 19982 5199 20038 5208
rect 19248 5102 19300 5108
rect 19614 5128 19670 5137
rect 19614 5063 19670 5072
rect 19064 2984 19116 2990
rect 19064 2926 19116 2932
rect 19156 2848 19208 2854
rect 19156 2790 19208 2796
rect 18234 2479 18290 2488
rect 18880 2508 18932 2514
rect 18880 2450 18932 2456
rect 18064 2230 19104 2258
rect 17972 2094 18092 2122
rect 17866 1456 17922 1465
rect 17866 1391 17922 1400
rect 18064 480 18092 2094
rect 19076 480 19104 2230
rect 19168 921 19196 2790
rect 19246 2408 19302 2417
rect 19246 2343 19248 2352
rect 19300 2343 19302 2352
rect 19248 2314 19300 2320
rect 19154 912 19210 921
rect 19154 847 19210 856
rect 20088 480 20116 12310
rect 20258 12271 20314 12280
rect 20168 5908 20220 5914
rect 20168 5850 20220 5856
rect 20180 5370 20208 5850
rect 20168 5364 20220 5370
rect 20168 5306 20220 5312
rect 20272 2961 20300 12271
rect 20548 3097 20576 14470
rect 20628 7404 20680 7410
rect 20628 7346 20680 7352
rect 20640 6322 20668 7346
rect 20628 6316 20680 6322
rect 20628 6258 20680 6264
rect 20534 3088 20590 3097
rect 20534 3023 20590 3032
rect 20258 2952 20314 2961
rect 20258 2887 20314 2896
rect 20732 2530 20760 18663
rect 20956 17980 21252 18000
rect 21012 17978 21036 17980
rect 21092 17978 21116 17980
rect 21172 17978 21196 17980
rect 21034 17926 21036 17978
rect 21098 17926 21110 17978
rect 21172 17926 21174 17978
rect 21012 17924 21036 17926
rect 21092 17924 21116 17926
rect 21172 17924 21196 17926
rect 20956 17904 21252 17924
rect 20956 16892 21252 16912
rect 21012 16890 21036 16892
rect 21092 16890 21116 16892
rect 21172 16890 21196 16892
rect 21034 16838 21036 16890
rect 21098 16838 21110 16890
rect 21172 16838 21174 16890
rect 21012 16836 21036 16838
rect 21092 16836 21116 16838
rect 21172 16836 21196 16838
rect 20956 16816 21252 16836
rect 20956 15804 21252 15824
rect 21012 15802 21036 15804
rect 21092 15802 21116 15804
rect 21172 15802 21196 15804
rect 21034 15750 21036 15802
rect 21098 15750 21110 15802
rect 21172 15750 21174 15802
rect 21012 15748 21036 15750
rect 21092 15748 21116 15750
rect 21172 15748 21196 15750
rect 20956 15728 21252 15748
rect 20956 14716 21252 14736
rect 21012 14714 21036 14716
rect 21092 14714 21116 14716
rect 21172 14714 21196 14716
rect 21034 14662 21036 14714
rect 21098 14662 21110 14714
rect 21172 14662 21174 14714
rect 21012 14660 21036 14662
rect 21092 14660 21116 14662
rect 21172 14660 21196 14662
rect 20956 14640 21252 14660
rect 20956 13628 21252 13648
rect 21012 13626 21036 13628
rect 21092 13626 21116 13628
rect 21172 13626 21196 13628
rect 21034 13574 21036 13626
rect 21098 13574 21110 13626
rect 21172 13574 21174 13626
rect 21012 13572 21036 13574
rect 21092 13572 21116 13574
rect 21172 13572 21196 13574
rect 20956 13552 21252 13572
rect 20956 12540 21252 12560
rect 21012 12538 21036 12540
rect 21092 12538 21116 12540
rect 21172 12538 21196 12540
rect 21034 12486 21036 12538
rect 21098 12486 21110 12538
rect 21172 12486 21174 12538
rect 21012 12484 21036 12486
rect 21092 12484 21116 12486
rect 21172 12484 21196 12486
rect 20956 12464 21252 12484
rect 20956 11452 21252 11472
rect 21012 11450 21036 11452
rect 21092 11450 21116 11452
rect 21172 11450 21196 11452
rect 21034 11398 21036 11450
rect 21098 11398 21110 11450
rect 21172 11398 21174 11450
rect 21012 11396 21036 11398
rect 21092 11396 21116 11398
rect 21172 11396 21196 11398
rect 20956 11376 21252 11396
rect 20956 10364 21252 10384
rect 21012 10362 21036 10364
rect 21092 10362 21116 10364
rect 21172 10362 21196 10364
rect 21034 10310 21036 10362
rect 21098 10310 21110 10362
rect 21172 10310 21174 10362
rect 21012 10308 21036 10310
rect 21092 10308 21116 10310
rect 21172 10308 21196 10310
rect 20956 10288 21252 10308
rect 20956 9276 21252 9296
rect 21012 9274 21036 9276
rect 21092 9274 21116 9276
rect 21172 9274 21196 9276
rect 21034 9222 21036 9274
rect 21098 9222 21110 9274
rect 21172 9222 21174 9274
rect 21012 9220 21036 9222
rect 21092 9220 21116 9222
rect 21172 9220 21196 9222
rect 20956 9200 21252 9220
rect 20812 8288 20864 8294
rect 20810 8256 20812 8265
rect 20864 8256 20866 8265
rect 20810 8191 20866 8200
rect 20956 8188 21252 8208
rect 21012 8186 21036 8188
rect 21092 8186 21116 8188
rect 21172 8186 21196 8188
rect 21034 8134 21036 8186
rect 21098 8134 21110 8186
rect 21172 8134 21174 8186
rect 21012 8132 21036 8134
rect 21092 8132 21116 8134
rect 21172 8132 21196 8134
rect 20956 8112 21252 8132
rect 20956 7100 21252 7120
rect 21012 7098 21036 7100
rect 21092 7098 21116 7100
rect 21172 7098 21196 7100
rect 21034 7046 21036 7098
rect 21098 7046 21110 7098
rect 21172 7046 21174 7098
rect 21012 7044 21036 7046
rect 21092 7044 21116 7046
rect 21172 7044 21196 7046
rect 20956 7024 21252 7044
rect 20824 6118 20852 6149
rect 20812 6112 20864 6118
rect 20810 6080 20812 6089
rect 20864 6080 20866 6089
rect 20810 6015 20866 6024
rect 20824 5681 20852 6015
rect 20956 6012 21252 6032
rect 21012 6010 21036 6012
rect 21092 6010 21116 6012
rect 21172 6010 21196 6012
rect 21034 5958 21036 6010
rect 21098 5958 21110 6010
rect 21172 5958 21174 6010
rect 21012 5956 21036 5958
rect 21092 5956 21116 5958
rect 21172 5956 21196 5958
rect 20956 5936 21252 5956
rect 20810 5672 20866 5681
rect 20810 5607 20866 5616
rect 20956 4924 21252 4944
rect 21012 4922 21036 4924
rect 21092 4922 21116 4924
rect 21172 4922 21196 4924
rect 21034 4870 21036 4922
rect 21098 4870 21110 4922
rect 21172 4870 21174 4922
rect 21012 4868 21036 4870
rect 21092 4868 21116 4870
rect 21172 4868 21196 4870
rect 20956 4848 21252 4868
rect 20956 3836 21252 3856
rect 21012 3834 21036 3836
rect 21092 3834 21116 3836
rect 21172 3834 21196 3836
rect 21034 3782 21036 3834
rect 21098 3782 21110 3834
rect 21172 3782 21174 3834
rect 21012 3780 21036 3782
rect 21092 3780 21116 3782
rect 21172 3780 21196 3782
rect 20956 3760 21252 3780
rect 21284 3641 21312 20198
rect 24228 19553 24256 20334
rect 24398 20295 24454 20304
rect 24412 20262 24440 20295
rect 24400 20256 24452 20262
rect 24400 20198 24452 20204
rect 24950 20224 25006 20233
rect 24950 20159 25006 20168
rect 24214 19544 24270 19553
rect 24214 19479 24270 19488
rect 24860 16244 24912 16250
rect 24860 16186 24912 16192
rect 24872 14770 24900 16186
rect 24964 15162 24992 20159
rect 25410 19952 25466 19961
rect 25410 19887 25466 19896
rect 25226 19408 25282 19417
rect 25226 19343 25282 19352
rect 25134 18864 25190 18873
rect 25134 18799 25190 18808
rect 25042 15872 25098 15881
rect 25042 15807 25098 15816
rect 24952 15156 25004 15162
rect 24952 15098 25004 15104
rect 24780 14742 24900 14770
rect 24780 13433 24808 14742
rect 24858 14648 24914 14657
rect 24858 14583 24914 14592
rect 24766 13424 24822 13433
rect 24766 13359 24822 13368
rect 21364 8288 21416 8294
rect 21362 8256 21364 8265
rect 24872 8265 24900 14583
rect 24950 13968 25006 13977
rect 24950 13903 25006 13912
rect 24964 10033 24992 13903
rect 25056 12209 25084 15807
rect 25148 12753 25176 18799
rect 25240 13025 25268 19343
rect 25318 15464 25374 15473
rect 25318 15399 25374 15408
rect 25226 13016 25282 13025
rect 25226 12951 25282 12960
rect 25134 12744 25190 12753
rect 25134 12679 25190 12688
rect 25042 12200 25098 12209
rect 25042 12135 25098 12144
rect 25332 10985 25360 15399
rect 25424 14521 25452 19887
rect 25410 14512 25466 14521
rect 25410 14447 25466 14456
rect 25410 13424 25466 13433
rect 25410 13359 25466 13368
rect 25318 10976 25374 10985
rect 25318 10911 25374 10920
rect 24950 10024 25006 10033
rect 24950 9959 25006 9968
rect 25424 8401 25452 13359
rect 25516 11665 25544 22335
rect 25596 20392 25648 20398
rect 25596 20334 25648 20340
rect 25608 19689 25636 20334
rect 25594 19680 25650 19689
rect 25594 19615 25650 19624
rect 25594 18320 25650 18329
rect 25594 18255 25650 18264
rect 25502 11656 25558 11665
rect 25502 11591 25558 11600
rect 25608 9081 25636 18255
rect 25700 11121 25728 23559
rect 26238 23520 26294 24000
rect 27710 23520 27766 24000
rect 29182 23520 29238 24000
rect 26252 23474 26280 23520
rect 26252 23446 26464 23474
rect 25870 23080 25926 23089
rect 25870 23015 25926 23024
rect 25778 21312 25834 21321
rect 25778 21247 25834 21256
rect 25792 20874 25820 21247
rect 25780 20868 25832 20874
rect 25780 20810 25832 20816
rect 25780 20528 25832 20534
rect 25778 20496 25780 20505
rect 25832 20496 25834 20505
rect 25778 20431 25834 20440
rect 25778 17096 25834 17105
rect 25778 17031 25834 17040
rect 25792 15337 25820 17031
rect 25884 16250 25912 23015
rect 25956 21788 26252 21808
rect 26012 21786 26036 21788
rect 26092 21786 26116 21788
rect 26172 21786 26196 21788
rect 26034 21734 26036 21786
rect 26098 21734 26110 21786
rect 26172 21734 26174 21786
rect 26012 21732 26036 21734
rect 26092 21732 26116 21734
rect 26172 21732 26196 21734
rect 25956 21712 26252 21732
rect 25956 20700 26252 20720
rect 26012 20698 26036 20700
rect 26092 20698 26116 20700
rect 26172 20698 26196 20700
rect 26034 20646 26036 20698
rect 26098 20646 26110 20698
rect 26172 20646 26174 20698
rect 26012 20644 26036 20646
rect 26092 20644 26116 20646
rect 26172 20644 26196 20646
rect 25956 20624 26252 20644
rect 26436 20369 26464 23446
rect 27724 20505 27752 23520
rect 27710 20496 27766 20505
rect 27710 20431 27766 20440
rect 26422 20360 26478 20369
rect 26422 20295 26478 20304
rect 26884 20256 26936 20262
rect 26884 20198 26936 20204
rect 27252 20256 27304 20262
rect 27252 20198 27304 20204
rect 26698 20088 26754 20097
rect 26698 20023 26700 20032
rect 26752 20023 26754 20032
rect 26700 19994 26752 20000
rect 26516 19916 26568 19922
rect 26516 19858 26568 19864
rect 25956 19612 26252 19632
rect 26012 19610 26036 19612
rect 26092 19610 26116 19612
rect 26172 19610 26196 19612
rect 26034 19558 26036 19610
rect 26098 19558 26110 19610
rect 26172 19558 26174 19610
rect 26012 19556 26036 19558
rect 26092 19556 26116 19558
rect 26172 19556 26196 19558
rect 25956 19536 26252 19556
rect 26528 19174 26556 19858
rect 26896 19825 26924 20198
rect 26882 19816 26938 19825
rect 26882 19751 26938 19760
rect 26516 19168 26568 19174
rect 26516 19110 26568 19116
rect 26528 18737 26556 19110
rect 26514 18728 26570 18737
rect 26514 18663 26570 18672
rect 25956 18524 26252 18544
rect 26012 18522 26036 18524
rect 26092 18522 26116 18524
rect 26172 18522 26196 18524
rect 26034 18470 26036 18522
rect 26098 18470 26110 18522
rect 26172 18470 26174 18522
rect 26012 18468 26036 18470
rect 26092 18468 26116 18470
rect 26172 18468 26196 18470
rect 25956 18448 26252 18468
rect 25956 17436 26252 17456
rect 26012 17434 26036 17436
rect 26092 17434 26116 17436
rect 26172 17434 26196 17436
rect 26034 17382 26036 17434
rect 26098 17382 26110 17434
rect 26172 17382 26174 17434
rect 26012 17380 26036 17382
rect 26092 17380 26116 17382
rect 26172 17380 26196 17382
rect 25956 17360 26252 17380
rect 25956 16348 26252 16368
rect 26012 16346 26036 16348
rect 26092 16346 26116 16348
rect 26172 16346 26196 16348
rect 26034 16294 26036 16346
rect 26098 16294 26110 16346
rect 26172 16294 26174 16346
rect 26012 16292 26036 16294
rect 26092 16292 26116 16294
rect 26172 16292 26196 16294
rect 25956 16272 26252 16292
rect 25872 16244 25924 16250
rect 25872 16186 25924 16192
rect 25870 16144 25926 16153
rect 25870 16079 25926 16088
rect 25778 15328 25834 15337
rect 25778 15263 25834 15272
rect 25780 15156 25832 15162
rect 25780 15098 25832 15104
rect 25686 11112 25742 11121
rect 25686 11047 25742 11056
rect 25594 9072 25650 9081
rect 25594 9007 25650 9016
rect 25792 8673 25820 15098
rect 25884 13841 25912 16079
rect 25956 15260 26252 15280
rect 26012 15258 26036 15260
rect 26092 15258 26116 15260
rect 26172 15258 26196 15260
rect 26034 15206 26036 15258
rect 26098 15206 26110 15258
rect 26172 15206 26174 15258
rect 26012 15204 26036 15206
rect 26092 15204 26116 15206
rect 26172 15204 26196 15206
rect 25956 15184 26252 15204
rect 25956 14172 26252 14192
rect 26012 14170 26036 14172
rect 26092 14170 26116 14172
rect 26172 14170 26196 14172
rect 26034 14118 26036 14170
rect 26098 14118 26110 14170
rect 26172 14118 26174 14170
rect 26012 14116 26036 14118
rect 26092 14116 26116 14118
rect 26172 14116 26196 14118
rect 25956 14096 26252 14116
rect 25870 13832 25926 13841
rect 25870 13767 25926 13776
rect 25956 13084 26252 13104
rect 26012 13082 26036 13084
rect 26092 13082 26116 13084
rect 26172 13082 26196 13084
rect 26034 13030 26036 13082
rect 26098 13030 26110 13082
rect 26172 13030 26174 13082
rect 26012 13028 26036 13030
rect 26092 13028 26116 13030
rect 26172 13028 26196 13030
rect 25956 13008 26252 13028
rect 25870 12336 25926 12345
rect 25870 12271 25926 12280
rect 25778 8664 25834 8673
rect 25778 8599 25834 8608
rect 25410 8392 25466 8401
rect 25410 8327 25466 8336
rect 21416 8256 21418 8265
rect 21362 8191 21418 8200
rect 21914 8256 21970 8265
rect 21914 8191 21970 8200
rect 24858 8256 24914 8265
rect 24858 8191 24914 8200
rect 21640 6656 21692 6662
rect 21640 6598 21692 6604
rect 21652 6322 21680 6598
rect 21640 6316 21692 6322
rect 21640 6258 21692 6264
rect 21928 6254 21956 8191
rect 25884 7993 25912 12271
rect 25956 11996 26252 12016
rect 26012 11994 26036 11996
rect 26092 11994 26116 11996
rect 26172 11994 26196 11996
rect 26034 11942 26036 11994
rect 26098 11942 26110 11994
rect 26172 11942 26174 11994
rect 26012 11940 26036 11942
rect 26092 11940 26116 11942
rect 26172 11940 26196 11942
rect 25956 11920 26252 11940
rect 26422 11792 26478 11801
rect 26422 11727 26478 11736
rect 26436 11694 26464 11727
rect 26424 11688 26476 11694
rect 26424 11630 26476 11636
rect 26698 11656 26754 11665
rect 26698 11591 26754 11600
rect 26608 11552 26660 11558
rect 26608 11494 26660 11500
rect 26516 11212 26568 11218
rect 26516 11154 26568 11160
rect 25956 10908 26252 10928
rect 26012 10906 26036 10908
rect 26092 10906 26116 10908
rect 26172 10906 26196 10908
rect 26034 10854 26036 10906
rect 26098 10854 26110 10906
rect 26172 10854 26174 10906
rect 26012 10852 26036 10854
rect 26092 10852 26116 10854
rect 26172 10852 26196 10854
rect 25956 10832 26252 10852
rect 26528 10810 26556 11154
rect 26620 11121 26648 11494
rect 26712 11354 26740 11591
rect 26700 11348 26752 11354
rect 26700 11290 26752 11296
rect 26606 11112 26662 11121
rect 26606 11047 26662 11056
rect 26516 10804 26568 10810
rect 26516 10746 26568 10752
rect 26528 10713 26556 10746
rect 26514 10704 26570 10713
rect 26514 10639 26570 10648
rect 26424 10600 26476 10606
rect 26422 10568 26424 10577
rect 26476 10568 26478 10577
rect 26422 10503 26478 10512
rect 26608 10464 26660 10470
rect 26606 10432 26608 10441
rect 26660 10432 26662 10441
rect 26606 10367 26662 10376
rect 26790 10160 26846 10169
rect 26790 10095 26846 10104
rect 26698 9888 26754 9897
rect 25956 9820 26252 9840
rect 26698 9823 26754 9832
rect 26012 9818 26036 9820
rect 26092 9818 26116 9820
rect 26172 9818 26196 9820
rect 26034 9766 26036 9818
rect 26098 9766 26110 9818
rect 26172 9766 26174 9818
rect 26012 9764 26036 9766
rect 26092 9764 26116 9766
rect 26172 9764 26196 9766
rect 25956 9744 26252 9764
rect 26606 9344 26662 9353
rect 26606 9279 26662 9288
rect 26516 9036 26568 9042
rect 26516 8978 26568 8984
rect 26528 8945 26556 8978
rect 26514 8936 26570 8945
rect 26514 8871 26570 8880
rect 25956 8732 26252 8752
rect 26012 8730 26036 8732
rect 26092 8730 26116 8732
rect 26172 8730 26196 8732
rect 26034 8678 26036 8730
rect 26098 8678 26110 8730
rect 26172 8678 26174 8730
rect 26012 8676 26036 8678
rect 26092 8676 26116 8678
rect 26172 8676 26196 8678
rect 25956 8656 26252 8676
rect 26528 8566 26556 8871
rect 26620 8634 26648 9279
rect 26712 9178 26740 9823
rect 26700 9172 26752 9178
rect 26700 9114 26752 9120
rect 26698 8664 26754 8673
rect 26608 8628 26660 8634
rect 26698 8599 26754 8608
rect 26608 8570 26660 8576
rect 26516 8560 26568 8566
rect 26422 8528 26478 8537
rect 26516 8502 26568 8508
rect 26422 8463 26478 8472
rect 26436 8430 26464 8463
rect 26424 8424 26476 8430
rect 26424 8366 26476 8372
rect 26712 8090 26740 8599
rect 26700 8084 26752 8090
rect 26700 8026 26752 8032
rect 25870 7984 25926 7993
rect 25870 7919 25926 7928
rect 26516 7948 26568 7954
rect 26516 7890 26568 7896
rect 25956 7644 26252 7664
rect 26012 7642 26036 7644
rect 26092 7642 26116 7644
rect 26172 7642 26196 7644
rect 26034 7590 26036 7642
rect 26098 7590 26110 7642
rect 26172 7590 26174 7642
rect 26012 7588 26036 7590
rect 26092 7588 26116 7590
rect 26172 7588 26196 7590
rect 25956 7568 26252 7588
rect 26528 7478 26556 7890
rect 26516 7472 26568 7478
rect 26422 7440 26478 7449
rect 26516 7414 26568 7420
rect 26698 7440 26754 7449
rect 26422 7375 26478 7384
rect 26436 7342 26464 7375
rect 26424 7336 26476 7342
rect 26528 7313 26556 7414
rect 26698 7375 26754 7384
rect 26424 7278 26476 7284
rect 26514 7304 26570 7313
rect 26514 7239 26570 7248
rect 26608 7200 26660 7206
rect 26608 7142 26660 7148
rect 26620 7041 26648 7142
rect 26606 7032 26662 7041
rect 26606 6967 26662 6976
rect 26514 6896 26570 6905
rect 26514 6831 26516 6840
rect 26568 6831 26570 6840
rect 26516 6802 26568 6808
rect 25956 6556 26252 6576
rect 26012 6554 26036 6556
rect 26092 6554 26116 6556
rect 26172 6554 26196 6556
rect 26034 6502 26036 6554
rect 26098 6502 26110 6554
rect 26172 6502 26174 6554
rect 26012 6500 26036 6502
rect 26092 6500 26116 6502
rect 26172 6500 26196 6502
rect 25956 6480 26252 6500
rect 26528 6458 26556 6802
rect 26712 6730 26740 7375
rect 26700 6724 26752 6730
rect 26700 6666 26752 6672
rect 26516 6452 26568 6458
rect 26516 6394 26568 6400
rect 26608 6384 26660 6390
rect 26330 6352 26386 6361
rect 26330 6287 26386 6296
rect 26606 6352 26608 6361
rect 26660 6352 26662 6361
rect 26606 6287 26662 6296
rect 21916 6248 21968 6254
rect 21916 6190 21968 6196
rect 21548 6112 21600 6118
rect 21548 6054 21600 6060
rect 21560 5914 21588 6054
rect 21928 5914 21956 6190
rect 21548 5908 21600 5914
rect 21548 5850 21600 5856
rect 21916 5908 21968 5914
rect 21916 5850 21968 5856
rect 25318 5672 25374 5681
rect 25318 5607 25374 5616
rect 25332 4690 25360 5607
rect 25956 5468 26252 5488
rect 26012 5466 26036 5468
rect 26092 5466 26116 5468
rect 26172 5466 26196 5468
rect 26034 5414 26036 5466
rect 26098 5414 26110 5466
rect 26172 5414 26174 5466
rect 26012 5412 26036 5414
rect 26092 5412 26116 5414
rect 26172 5412 26196 5414
rect 25956 5392 26252 5412
rect 25320 4684 25372 4690
rect 25320 4626 25372 4632
rect 25332 4282 25360 4626
rect 25780 4480 25832 4486
rect 25780 4422 25832 4428
rect 25320 4276 25372 4282
rect 25320 4218 25372 4224
rect 21270 3632 21326 3641
rect 21270 3567 21326 3576
rect 23202 3632 23258 3641
rect 23202 3567 23258 3576
rect 22190 2952 22246 2961
rect 22190 2887 22246 2896
rect 20956 2748 21252 2768
rect 21012 2746 21036 2748
rect 21092 2746 21116 2748
rect 21172 2746 21196 2748
rect 21034 2694 21036 2746
rect 21098 2694 21110 2746
rect 21172 2694 21174 2746
rect 21012 2692 21036 2694
rect 21092 2692 21116 2694
rect 21172 2692 21196 2694
rect 20956 2672 21252 2692
rect 20732 2502 21128 2530
rect 21100 480 21128 2502
rect 22204 480 22232 2887
rect 23216 480 23244 3567
rect 25318 3088 25374 3097
rect 25318 3023 25374 3032
rect 25332 2990 25360 3023
rect 25320 2984 25372 2990
rect 25320 2926 25372 2932
rect 25502 2952 25558 2961
rect 25502 2887 25558 2896
rect 25516 2854 25544 2887
rect 25504 2848 25556 2854
rect 25504 2790 25556 2796
rect 25792 2689 25820 4422
rect 25956 4380 26252 4400
rect 26012 4378 26036 4380
rect 26092 4378 26116 4380
rect 26172 4378 26196 4380
rect 26034 4326 26036 4378
rect 26098 4326 26110 4378
rect 26172 4326 26174 4378
rect 26012 4324 26036 4326
rect 26092 4324 26116 4326
rect 26172 4324 26196 4326
rect 25956 4304 26252 4324
rect 25956 3292 26252 3312
rect 26012 3290 26036 3292
rect 26092 3290 26116 3292
rect 26172 3290 26196 3292
rect 26034 3238 26036 3290
rect 26098 3238 26110 3290
rect 26172 3238 26174 3290
rect 26012 3236 26036 3238
rect 26092 3236 26116 3238
rect 26172 3236 26196 3238
rect 25956 3216 26252 3236
rect 26344 2990 26372 6287
rect 26424 6248 26476 6254
rect 26424 6190 26476 6196
rect 26514 6216 26570 6225
rect 26436 5817 26464 6190
rect 26514 6151 26570 6160
rect 26422 5808 26478 5817
rect 26528 5778 26556 6151
rect 26422 5743 26478 5752
rect 26516 5772 26568 5778
rect 26516 5714 26568 5720
rect 26528 5370 26556 5714
rect 26698 5672 26754 5681
rect 26698 5607 26700 5616
rect 26752 5607 26754 5616
rect 26700 5578 26752 5584
rect 26516 5364 26568 5370
rect 26516 5306 26568 5312
rect 26424 5160 26476 5166
rect 26422 5128 26424 5137
rect 26476 5128 26478 5137
rect 26422 5063 26478 5072
rect 26606 5128 26662 5137
rect 26606 5063 26662 5072
rect 26620 5030 26648 5063
rect 26608 5024 26660 5030
rect 26608 4966 26660 4972
rect 26804 4690 26832 10095
rect 27264 6769 27292 20198
rect 29196 20097 29224 23520
rect 29182 20088 29238 20097
rect 29182 20023 29238 20032
rect 27526 9480 27582 9489
rect 27526 9415 27582 9424
rect 27540 8430 27568 9415
rect 27712 8560 27764 8566
rect 27712 8502 27764 8508
rect 27528 8424 27580 8430
rect 27724 8401 27752 8502
rect 27528 8366 27580 8372
rect 27710 8392 27766 8401
rect 27710 8327 27766 8336
rect 27250 6760 27306 6769
rect 27250 6695 27306 6704
rect 28354 6760 28410 6769
rect 28354 6695 28410 6704
rect 26882 5264 26938 5273
rect 26882 5199 26938 5208
rect 26792 4684 26844 4690
rect 26792 4626 26844 4632
rect 26700 4480 26752 4486
rect 26698 4448 26700 4457
rect 26752 4448 26754 4457
rect 26698 4383 26754 4392
rect 26804 4282 26832 4626
rect 26792 4276 26844 4282
rect 26792 4218 26844 4224
rect 26424 4072 26476 4078
rect 26422 4040 26424 4049
rect 26476 4040 26478 4049
rect 26422 3975 26478 3984
rect 26608 3936 26660 3942
rect 26606 3904 26608 3913
rect 26660 3904 26662 3913
rect 26606 3839 26662 3848
rect 26700 3392 26752 3398
rect 26698 3360 26700 3369
rect 26752 3360 26754 3369
rect 26698 3295 26754 3304
rect 26332 2984 26384 2990
rect 26332 2926 26384 2932
rect 26608 2848 26660 2854
rect 25870 2816 25926 2825
rect 26608 2790 26660 2796
rect 25870 2751 25926 2760
rect 25778 2680 25834 2689
rect 25884 2650 25912 2751
rect 25778 2615 25834 2624
rect 25872 2644 25924 2650
rect 25872 2586 25924 2592
rect 24398 2544 24454 2553
rect 24398 2479 24400 2488
rect 24452 2479 24454 2488
rect 24400 2450 24452 2456
rect 26332 2372 26384 2378
rect 26332 2314 26384 2320
rect 25956 2204 26252 2224
rect 26012 2202 26036 2204
rect 26092 2202 26116 2204
rect 26172 2202 26196 2204
rect 26034 2150 26036 2202
rect 26098 2150 26110 2202
rect 26172 2150 26174 2202
rect 26012 2148 26036 2150
rect 26092 2148 26116 2150
rect 26172 2148 26196 2150
rect 25956 2128 26252 2148
rect 24214 2000 24270 2009
rect 24214 1935 24270 1944
rect 24228 480 24256 1935
rect 25226 1456 25282 1465
rect 25226 1391 25282 1400
rect 25240 480 25268 1391
rect 26344 480 26372 2314
rect 2778 368 2834 377
rect 2778 303 2834 312
rect 3514 0 3570 480
rect 4526 0 4582 480
rect 5630 0 5686 480
rect 6642 0 6698 480
rect 7654 0 7710 480
rect 8666 0 8722 480
rect 9770 0 9826 480
rect 10782 0 10838 480
rect 11794 0 11850 480
rect 12806 0 12862 480
rect 13910 0 13966 480
rect 14922 0 14978 480
rect 15934 0 15990 480
rect 16946 0 17002 480
rect 18050 0 18106 480
rect 19062 0 19118 480
rect 20074 0 20130 480
rect 21086 0 21142 480
rect 22190 0 22246 480
rect 23202 0 23258 480
rect 24214 0 24270 480
rect 25226 0 25282 480
rect 26330 0 26386 480
rect 26620 377 26648 2790
rect 26896 2514 26924 5199
rect 27344 3596 27396 3602
rect 27344 3538 27396 3544
rect 27356 3194 27384 3538
rect 27344 3188 27396 3194
rect 27344 3130 27396 3136
rect 27342 2952 27398 2961
rect 27342 2887 27398 2896
rect 26884 2508 26936 2514
rect 26884 2450 26936 2456
rect 27068 2304 27120 2310
rect 27068 2246 27120 2252
rect 27080 1465 27108 2246
rect 27066 1456 27122 1465
rect 27066 1391 27122 1400
rect 27356 480 27384 2887
rect 28368 480 28396 6695
rect 29366 2816 29422 2825
rect 29366 2751 29422 2760
rect 29380 480 29408 2751
rect 26606 368 26662 377
rect 26606 303 26662 312
rect 27342 0 27398 480
rect 28354 0 28410 480
rect 29366 0 29422 480
<< via2 >>
rect 2962 23568 3018 23624
rect 754 20168 810 20224
rect 2870 22344 2926 22400
rect 2226 19760 2282 19816
rect 2778 15272 2834 15328
rect 1398 12824 1454 12880
rect 1582 11600 1638 11656
rect 1398 11056 1454 11112
rect 1582 10376 1638 10432
rect 1490 9832 1546 9888
rect 1398 9288 1454 9344
rect 1674 9696 1730 9752
rect 1582 8608 1638 8664
rect 1582 7420 1584 7440
rect 1584 7420 1636 7440
rect 1636 7420 1638 7440
rect 1582 7384 1638 7420
rect 1582 6840 1638 6896
rect 1582 6332 1584 6352
rect 1584 6332 1636 6352
rect 1636 6332 1638 6352
rect 1582 6296 1638 6332
rect 1582 5636 1638 5672
rect 1582 5616 1584 5636
rect 1584 5616 1636 5636
rect 1636 5616 1638 5636
rect 1582 4428 1584 4448
rect 1584 4428 1636 4448
rect 1636 4428 1638 4448
rect 1582 4392 1638 4428
rect 1582 3884 1584 3904
rect 1584 3884 1636 3904
rect 1636 3884 1638 3904
rect 1582 3848 1638 3884
rect 1582 3340 1584 3360
rect 1584 3340 1636 3360
rect 1636 3340 1638 3360
rect 1582 3304 1638 3340
rect 570 2760 626 2816
rect 1582 2624 1638 2680
rect 25686 23568 25742 23624
rect 3146 23024 3202 23080
rect 3514 21256 3570 21312
rect 3238 20576 3294 20632
rect 2962 14592 3018 14648
rect 2042 9968 2098 10024
rect 2042 8880 2098 8936
rect 2410 8372 2412 8392
rect 2412 8372 2464 8392
rect 2464 8372 2466 8392
rect 2410 8336 2466 8372
rect 2042 8200 2098 8256
rect 2410 7284 2412 7304
rect 2412 7284 2464 7304
rect 2464 7284 2466 7304
rect 2410 7248 2466 7284
rect 2042 6840 2098 6896
rect 2410 5888 2466 5944
rect 2042 4800 2098 4856
rect 2410 4156 2412 4176
rect 2412 4156 2464 4176
rect 2464 4156 2466 4176
rect 2410 4120 2466 4156
rect 2778 11736 2834 11792
rect 2686 11600 2742 11656
rect 2594 9596 2596 9616
rect 2596 9596 2648 9616
rect 2648 9596 2650 9616
rect 3054 13368 3110 13424
rect 3606 20032 3662 20088
rect 3330 19352 3386 19408
rect 3514 17040 3570 17096
rect 3422 16360 3478 16416
rect 3330 12416 3386 12472
rect 3238 11756 3294 11792
rect 2870 9968 2926 10024
rect 2594 9560 2650 9596
rect 2686 8064 2742 8120
rect 3238 11736 3240 11756
rect 3240 11736 3292 11756
rect 3292 11736 3294 11756
rect 3146 11056 3202 11112
rect 3146 10376 3202 10432
rect 3882 21800 3938 21856
rect 5956 21786 6012 21788
rect 6036 21786 6092 21788
rect 6116 21786 6172 21788
rect 6196 21786 6252 21788
rect 5956 21734 5982 21786
rect 5982 21734 6012 21786
rect 6036 21734 6046 21786
rect 6046 21734 6092 21786
rect 6116 21734 6162 21786
rect 6162 21734 6172 21786
rect 6196 21734 6226 21786
rect 6226 21734 6252 21786
rect 5956 21732 6012 21734
rect 6036 21732 6092 21734
rect 6116 21732 6172 21734
rect 6196 21732 6252 21734
rect 5956 20698 6012 20700
rect 6036 20698 6092 20700
rect 6116 20698 6172 20700
rect 6196 20698 6252 20700
rect 5956 20646 5982 20698
rect 5982 20646 6012 20698
rect 6036 20646 6046 20698
rect 6046 20646 6092 20698
rect 6116 20646 6162 20698
rect 6162 20646 6172 20698
rect 6196 20646 6226 20698
rect 6226 20646 6252 20698
rect 5956 20644 6012 20646
rect 6036 20644 6092 20646
rect 6116 20644 6172 20646
rect 6196 20644 6252 20646
rect 3698 19896 3754 19952
rect 5956 19610 6012 19612
rect 6036 19610 6092 19612
rect 6116 19610 6172 19612
rect 6196 19610 6252 19612
rect 5956 19558 5982 19610
rect 5982 19558 6012 19610
rect 6036 19558 6046 19610
rect 6046 19558 6092 19610
rect 6116 19558 6162 19610
rect 6162 19558 6172 19610
rect 6196 19558 6226 19610
rect 6226 19558 6252 19610
rect 5956 19556 6012 19558
rect 6036 19556 6092 19558
rect 6116 19556 6172 19558
rect 6196 19556 6252 19558
rect 5354 19352 5410 19408
rect 7470 20324 7526 20360
rect 7470 20304 7472 20324
rect 7472 20304 7524 20324
rect 7524 20304 7526 20324
rect 7562 20168 7618 20224
rect 7562 19624 7618 19680
rect 3698 18808 3754 18864
rect 3422 10240 3478 10296
rect 5956 18522 6012 18524
rect 6036 18522 6092 18524
rect 6116 18522 6172 18524
rect 6196 18522 6252 18524
rect 5956 18470 5982 18522
rect 5982 18470 6012 18522
rect 6036 18470 6046 18522
rect 6046 18470 6092 18522
rect 6116 18470 6162 18522
rect 6162 18470 6172 18522
rect 6196 18470 6226 18522
rect 6226 18470 6252 18522
rect 5956 18468 6012 18470
rect 6036 18468 6092 18470
rect 6116 18468 6172 18470
rect 6196 18468 6252 18470
rect 5722 18264 5778 18320
rect 3790 17584 3846 17640
rect 3882 14048 3938 14104
rect 3790 12416 3846 12472
rect 3606 9832 3662 9888
rect 3974 12824 4030 12880
rect 4066 12688 4122 12744
rect 4066 12436 4122 12472
rect 4066 12416 4068 12436
rect 4068 12416 4120 12436
rect 4120 12416 4122 12436
rect 3698 9696 3754 9752
rect 3514 9424 3570 9480
rect 3146 8492 3202 8528
rect 3146 8472 3148 8492
rect 3148 8472 3200 8492
rect 3200 8472 3202 8492
rect 3054 6704 3110 6760
rect 4342 12144 4398 12200
rect 5538 11636 5540 11656
rect 5540 11636 5592 11656
rect 5592 11636 5594 11656
rect 5538 11600 5594 11636
rect 3882 9716 3938 9752
rect 3882 9696 3884 9716
rect 3884 9696 3936 9716
rect 3936 9696 3938 9716
rect 4526 10104 4582 10160
rect 5538 9868 5540 9888
rect 5540 9868 5592 9888
rect 5592 9868 5594 9888
rect 5538 9832 5594 9868
rect 3790 8064 3846 8120
rect 3422 7792 3478 7848
rect 3330 6568 3386 6624
rect 3146 5244 3148 5264
rect 3148 5244 3200 5264
rect 3200 5244 3202 5264
rect 2686 5072 2742 5128
rect 2042 3440 2098 3496
rect 2686 2080 2742 2136
rect 3146 5208 3202 5244
rect 3146 3884 3148 3904
rect 3148 3884 3200 3904
rect 3200 3884 3202 3904
rect 3146 3848 3202 3884
rect 2962 2760 3018 2816
rect 2870 1400 2926 1456
rect 4986 7384 5042 7440
rect 4618 6296 4674 6352
rect 5630 6568 5686 6624
rect 4066 5072 4122 5128
rect 4158 3052 4214 3088
rect 4158 3032 4160 3052
rect 4160 3032 4212 3052
rect 4212 3032 4214 3052
rect 4066 856 4122 912
rect 5078 6060 5080 6080
rect 5080 6060 5132 6080
rect 5132 6060 5134 6080
rect 5078 6024 5134 6060
rect 5956 17434 6012 17436
rect 6036 17434 6092 17436
rect 6116 17434 6172 17436
rect 6196 17434 6252 17436
rect 5956 17382 5982 17434
rect 5982 17382 6012 17434
rect 6036 17382 6046 17434
rect 6046 17382 6092 17434
rect 6116 17382 6162 17434
rect 6162 17382 6172 17434
rect 6196 17382 6226 17434
rect 6226 17382 6252 17434
rect 5956 17380 6012 17382
rect 6036 17380 6092 17382
rect 6116 17380 6172 17382
rect 6196 17380 6252 17382
rect 5956 16346 6012 16348
rect 6036 16346 6092 16348
rect 6116 16346 6172 16348
rect 6196 16346 6252 16348
rect 5956 16294 5982 16346
rect 5982 16294 6012 16346
rect 6036 16294 6046 16346
rect 6046 16294 6092 16346
rect 6116 16294 6162 16346
rect 6162 16294 6172 16346
rect 6196 16294 6226 16346
rect 6226 16294 6252 16346
rect 5956 16292 6012 16294
rect 6036 16292 6092 16294
rect 6116 16292 6172 16294
rect 6196 16292 6252 16294
rect 5956 15258 6012 15260
rect 6036 15258 6092 15260
rect 6116 15258 6172 15260
rect 6196 15258 6252 15260
rect 5956 15206 5982 15258
rect 5982 15206 6012 15258
rect 6036 15206 6046 15258
rect 6046 15206 6092 15258
rect 6116 15206 6162 15258
rect 6162 15206 6172 15258
rect 6196 15206 6226 15258
rect 6226 15206 6252 15258
rect 5956 15204 6012 15206
rect 6036 15204 6092 15206
rect 6116 15204 6172 15206
rect 6196 15204 6252 15206
rect 5956 14170 6012 14172
rect 6036 14170 6092 14172
rect 6116 14170 6172 14172
rect 6196 14170 6252 14172
rect 5956 14118 5982 14170
rect 5982 14118 6012 14170
rect 6036 14118 6046 14170
rect 6046 14118 6092 14170
rect 6116 14118 6162 14170
rect 6162 14118 6172 14170
rect 6196 14118 6226 14170
rect 6226 14118 6252 14170
rect 5956 14116 6012 14118
rect 6036 14116 6092 14118
rect 6116 14116 6172 14118
rect 6196 14116 6252 14118
rect 5956 13082 6012 13084
rect 6036 13082 6092 13084
rect 6116 13082 6172 13084
rect 6196 13082 6252 13084
rect 5956 13030 5982 13082
rect 5982 13030 6012 13082
rect 6036 13030 6046 13082
rect 6046 13030 6092 13082
rect 6116 13030 6162 13082
rect 6162 13030 6172 13082
rect 6196 13030 6226 13082
rect 6226 13030 6252 13082
rect 5956 13028 6012 13030
rect 6036 13028 6092 13030
rect 6116 13028 6172 13030
rect 6196 13028 6252 13030
rect 5956 11994 6012 11996
rect 6036 11994 6092 11996
rect 6116 11994 6172 11996
rect 6196 11994 6252 11996
rect 5956 11942 5982 11994
rect 5982 11942 6012 11994
rect 6036 11942 6046 11994
rect 6046 11942 6092 11994
rect 6116 11942 6162 11994
rect 6162 11942 6172 11994
rect 6196 11942 6226 11994
rect 6226 11942 6252 11994
rect 5956 11940 6012 11942
rect 6036 11940 6092 11942
rect 6116 11940 6172 11942
rect 6196 11940 6252 11942
rect 5956 10906 6012 10908
rect 6036 10906 6092 10908
rect 6116 10906 6172 10908
rect 6196 10906 6252 10908
rect 5956 10854 5982 10906
rect 5982 10854 6012 10906
rect 6036 10854 6046 10906
rect 6046 10854 6092 10906
rect 6116 10854 6162 10906
rect 6162 10854 6172 10906
rect 6196 10854 6226 10906
rect 6226 10854 6252 10906
rect 5956 10852 6012 10854
rect 6036 10852 6092 10854
rect 6116 10852 6172 10854
rect 6196 10852 6252 10854
rect 6458 10376 6514 10432
rect 5956 9818 6012 9820
rect 6036 9818 6092 9820
rect 6116 9818 6172 9820
rect 6196 9818 6252 9820
rect 5956 9766 5982 9818
rect 5982 9766 6012 9818
rect 6036 9766 6046 9818
rect 6046 9766 6092 9818
rect 6116 9766 6162 9818
rect 6162 9766 6172 9818
rect 6196 9766 6226 9818
rect 6226 9766 6252 9818
rect 5956 9764 6012 9766
rect 6036 9764 6092 9766
rect 6116 9764 6172 9766
rect 6196 9764 6252 9766
rect 5956 8730 6012 8732
rect 6036 8730 6092 8732
rect 6116 8730 6172 8732
rect 6196 8730 6252 8732
rect 5956 8678 5982 8730
rect 5982 8678 6012 8730
rect 6036 8678 6046 8730
rect 6046 8678 6092 8730
rect 6116 8678 6162 8730
rect 6162 8678 6172 8730
rect 6196 8678 6226 8730
rect 6226 8678 6252 8730
rect 5956 8676 6012 8678
rect 6036 8676 6092 8678
rect 6116 8676 6172 8678
rect 6196 8676 6252 8678
rect 6366 8064 6422 8120
rect 6274 7928 6330 7984
rect 5956 7642 6012 7644
rect 6036 7642 6092 7644
rect 6116 7642 6172 7644
rect 6196 7642 6252 7644
rect 5956 7590 5982 7642
rect 5982 7590 6012 7642
rect 6036 7590 6046 7642
rect 6046 7590 6092 7642
rect 6116 7590 6162 7642
rect 6162 7590 6172 7642
rect 6196 7590 6226 7642
rect 6226 7590 6252 7642
rect 5956 7588 6012 7590
rect 6036 7588 6092 7590
rect 6116 7588 6172 7590
rect 6196 7588 6252 7590
rect 6366 7656 6422 7712
rect 6366 6976 6422 7032
rect 5956 6554 6012 6556
rect 6036 6554 6092 6556
rect 6116 6554 6172 6556
rect 6196 6554 6252 6556
rect 5956 6502 5982 6554
rect 5982 6502 6012 6554
rect 6036 6502 6046 6554
rect 6046 6502 6092 6554
rect 6116 6502 6162 6554
rect 6162 6502 6172 6554
rect 6196 6502 6226 6554
rect 6226 6502 6252 6554
rect 5956 6500 6012 6502
rect 6036 6500 6092 6502
rect 6116 6500 6172 6502
rect 6196 6500 6252 6502
rect 5814 5772 5870 5808
rect 5814 5752 5816 5772
rect 5816 5752 5868 5772
rect 5868 5752 5870 5772
rect 5956 5466 6012 5468
rect 6036 5466 6092 5468
rect 6116 5466 6172 5468
rect 6196 5466 6252 5468
rect 5956 5414 5982 5466
rect 5982 5414 6012 5466
rect 6036 5414 6046 5466
rect 6046 5414 6092 5466
rect 6116 5414 6162 5466
rect 6162 5414 6172 5466
rect 6196 5414 6226 5466
rect 6226 5414 6252 5466
rect 5956 5412 6012 5414
rect 6036 5412 6092 5414
rect 6116 5412 6172 5414
rect 6196 5412 6252 5414
rect 5956 4378 6012 4380
rect 6036 4378 6092 4380
rect 6116 4378 6172 4380
rect 6196 4378 6252 4380
rect 5956 4326 5982 4378
rect 5982 4326 6012 4378
rect 6036 4326 6046 4378
rect 6046 4326 6092 4378
rect 6116 4326 6162 4378
rect 6162 4326 6172 4378
rect 6196 4326 6226 4378
rect 6226 4326 6252 4378
rect 5956 4324 6012 4326
rect 6036 4324 6092 4326
rect 6116 4324 6172 4326
rect 6196 4324 6252 4326
rect 4618 4020 4620 4040
rect 4620 4020 4672 4040
rect 4672 4020 4674 4040
rect 4618 3984 4674 4020
rect 4894 2644 4950 2680
rect 4894 2624 4896 2644
rect 4896 2624 4948 2644
rect 4948 2624 4950 2644
rect 6366 4800 6422 4856
rect 8574 18672 8630 18728
rect 8574 12960 8630 13016
rect 7746 9560 7802 9616
rect 7194 8508 7196 8528
rect 7196 8508 7248 8528
rect 7248 8508 7250 8528
rect 7194 8472 7250 8508
rect 7562 9016 7618 9072
rect 7654 8372 7656 8392
rect 7656 8372 7708 8392
rect 7708 8372 7710 8392
rect 7654 8336 7710 8372
rect 6550 6840 6606 6896
rect 6826 6296 6882 6352
rect 7010 6024 7066 6080
rect 6642 5364 6698 5400
rect 6642 5344 6644 5364
rect 6644 5344 6696 5364
rect 6696 5344 6698 5364
rect 7194 3848 7250 3904
rect 6274 3440 6330 3496
rect 5956 3290 6012 3292
rect 6036 3290 6092 3292
rect 6116 3290 6172 3292
rect 6196 3290 6252 3292
rect 5956 3238 5982 3290
rect 5982 3238 6012 3290
rect 6036 3238 6046 3290
rect 6046 3238 6092 3290
rect 6116 3238 6162 3290
rect 6162 3238 6172 3290
rect 6196 3238 6226 3290
rect 6226 3238 6252 3290
rect 5956 3236 6012 3238
rect 6036 3236 6092 3238
rect 6116 3236 6172 3238
rect 6196 3236 6252 3238
rect 5956 2202 6012 2204
rect 6036 2202 6092 2204
rect 6116 2202 6172 2204
rect 6196 2202 6252 2204
rect 5956 2150 5982 2202
rect 5982 2150 6012 2202
rect 6036 2150 6046 2202
rect 6046 2150 6092 2202
rect 6116 2150 6162 2202
rect 6162 2150 6172 2202
rect 6196 2150 6226 2202
rect 6226 2150 6252 2202
rect 5956 2148 6012 2150
rect 6036 2148 6092 2150
rect 6116 2148 6172 2150
rect 6196 2148 6252 2150
rect 9310 13232 9366 13288
rect 10956 21242 11012 21244
rect 11036 21242 11092 21244
rect 11116 21242 11172 21244
rect 11196 21242 11252 21244
rect 10956 21190 10982 21242
rect 10982 21190 11012 21242
rect 11036 21190 11046 21242
rect 11046 21190 11092 21242
rect 11116 21190 11162 21242
rect 11162 21190 11172 21242
rect 11196 21190 11226 21242
rect 11226 21190 11252 21242
rect 10956 21188 11012 21190
rect 11036 21188 11092 21190
rect 11116 21188 11172 21190
rect 11196 21188 11252 21190
rect 9678 20440 9734 20496
rect 9954 15816 10010 15872
rect 9402 11736 9458 11792
rect 10138 13368 10194 13424
rect 10046 12860 10048 12880
rect 10048 12860 10100 12880
rect 10100 12860 10102 12880
rect 10046 12824 10102 12860
rect 9862 12300 9918 12336
rect 9862 12280 9864 12300
rect 9864 12280 9916 12300
rect 9916 12280 9918 12300
rect 9494 10648 9550 10704
rect 9586 10532 9642 10568
rect 9586 10512 9588 10532
rect 9588 10512 9640 10532
rect 9640 10512 9642 10532
rect 9586 9832 9642 9888
rect 9034 8200 9090 8256
rect 9218 7384 9274 7440
rect 10230 12144 10286 12200
rect 10046 9288 10102 9344
rect 9862 6840 9918 6896
rect 9770 5344 9826 5400
rect 9402 3984 9458 4040
rect 8114 3576 8170 3632
rect 8022 2624 8078 2680
rect 10506 10412 10508 10432
rect 10508 10412 10560 10432
rect 10560 10412 10562 10432
rect 10506 10376 10562 10412
rect 10956 20154 11012 20156
rect 11036 20154 11092 20156
rect 11116 20154 11172 20156
rect 11196 20154 11252 20156
rect 10956 20102 10982 20154
rect 10982 20102 11012 20154
rect 11036 20102 11046 20154
rect 11046 20102 11092 20154
rect 11116 20102 11162 20154
rect 11162 20102 11172 20154
rect 11196 20102 11226 20154
rect 11226 20102 11252 20154
rect 10956 20100 11012 20102
rect 11036 20100 11092 20102
rect 11116 20100 11172 20102
rect 11196 20100 11252 20102
rect 10956 19066 11012 19068
rect 11036 19066 11092 19068
rect 11116 19066 11172 19068
rect 11196 19066 11252 19068
rect 10956 19014 10982 19066
rect 10982 19014 11012 19066
rect 11036 19014 11046 19066
rect 11046 19014 11092 19066
rect 11116 19014 11162 19066
rect 11162 19014 11172 19066
rect 11196 19014 11226 19066
rect 11226 19014 11252 19066
rect 10956 19012 11012 19014
rect 11036 19012 11092 19014
rect 11116 19012 11172 19014
rect 11196 19012 11252 19014
rect 10956 17978 11012 17980
rect 11036 17978 11092 17980
rect 11116 17978 11172 17980
rect 11196 17978 11252 17980
rect 10956 17926 10982 17978
rect 10982 17926 11012 17978
rect 11036 17926 11046 17978
rect 11046 17926 11092 17978
rect 11116 17926 11162 17978
rect 11162 17926 11172 17978
rect 11196 17926 11226 17978
rect 11226 17926 11252 17978
rect 10956 17924 11012 17926
rect 11036 17924 11092 17926
rect 11116 17924 11172 17926
rect 11196 17924 11252 17926
rect 10956 16890 11012 16892
rect 11036 16890 11092 16892
rect 11116 16890 11172 16892
rect 11196 16890 11252 16892
rect 10956 16838 10982 16890
rect 10982 16838 11012 16890
rect 11036 16838 11046 16890
rect 11046 16838 11092 16890
rect 11116 16838 11162 16890
rect 11162 16838 11172 16890
rect 11196 16838 11226 16890
rect 11226 16838 11252 16890
rect 10956 16836 11012 16838
rect 11036 16836 11092 16838
rect 11116 16836 11172 16838
rect 11196 16836 11252 16838
rect 10956 15802 11012 15804
rect 11036 15802 11092 15804
rect 11116 15802 11172 15804
rect 11196 15802 11252 15804
rect 10956 15750 10982 15802
rect 10982 15750 11012 15802
rect 11036 15750 11046 15802
rect 11046 15750 11092 15802
rect 11116 15750 11162 15802
rect 11162 15750 11172 15802
rect 11196 15750 11226 15802
rect 11226 15750 11252 15802
rect 10956 15748 11012 15750
rect 11036 15748 11092 15750
rect 11116 15748 11172 15750
rect 11196 15748 11252 15750
rect 10956 14714 11012 14716
rect 11036 14714 11092 14716
rect 11116 14714 11172 14716
rect 11196 14714 11252 14716
rect 10956 14662 10982 14714
rect 10982 14662 11012 14714
rect 11036 14662 11046 14714
rect 11046 14662 11092 14714
rect 11116 14662 11162 14714
rect 11162 14662 11172 14714
rect 11196 14662 11226 14714
rect 11226 14662 11252 14714
rect 10956 14660 11012 14662
rect 11036 14660 11092 14662
rect 11116 14660 11172 14662
rect 11196 14660 11252 14662
rect 10956 13626 11012 13628
rect 11036 13626 11092 13628
rect 11116 13626 11172 13628
rect 11196 13626 11252 13628
rect 10956 13574 10982 13626
rect 10982 13574 11012 13626
rect 11036 13574 11046 13626
rect 11046 13574 11092 13626
rect 11116 13574 11162 13626
rect 11162 13574 11172 13626
rect 11196 13574 11226 13626
rect 11226 13574 11252 13626
rect 10956 13572 11012 13574
rect 11036 13572 11092 13574
rect 11116 13572 11172 13574
rect 11196 13572 11252 13574
rect 10956 12538 11012 12540
rect 11036 12538 11092 12540
rect 11116 12538 11172 12540
rect 11196 12538 11252 12540
rect 10956 12486 10982 12538
rect 10982 12486 11012 12538
rect 11036 12486 11046 12538
rect 11046 12486 11092 12538
rect 11116 12486 11162 12538
rect 11162 12486 11172 12538
rect 11196 12486 11226 12538
rect 11226 12486 11252 12538
rect 10956 12484 11012 12486
rect 11036 12484 11092 12486
rect 11116 12484 11172 12486
rect 11196 12484 11252 12486
rect 10956 11450 11012 11452
rect 11036 11450 11092 11452
rect 11116 11450 11172 11452
rect 11196 11450 11252 11452
rect 10956 11398 10982 11450
rect 10982 11398 11012 11450
rect 11036 11398 11046 11450
rect 11046 11398 11092 11450
rect 11116 11398 11162 11450
rect 11162 11398 11172 11450
rect 11196 11398 11226 11450
rect 11226 11398 11252 11450
rect 10956 11396 11012 11398
rect 11036 11396 11092 11398
rect 11116 11396 11172 11398
rect 11196 11396 11252 11398
rect 10956 10362 11012 10364
rect 11036 10362 11092 10364
rect 11116 10362 11172 10364
rect 11196 10362 11252 10364
rect 10956 10310 10982 10362
rect 10982 10310 11012 10362
rect 11036 10310 11046 10362
rect 11046 10310 11092 10362
rect 11116 10310 11162 10362
rect 11162 10310 11172 10362
rect 11196 10310 11226 10362
rect 11226 10310 11252 10362
rect 10956 10308 11012 10310
rect 11036 10308 11092 10310
rect 11116 10308 11172 10310
rect 11196 10308 11252 10310
rect 10874 9560 10930 9616
rect 11334 9324 11336 9344
rect 11336 9324 11388 9344
rect 11388 9324 11390 9344
rect 11334 9288 11390 9324
rect 10956 9274 11012 9276
rect 11036 9274 11092 9276
rect 11116 9274 11172 9276
rect 11196 9274 11252 9276
rect 10956 9222 10982 9274
rect 10982 9222 11012 9274
rect 11036 9222 11046 9274
rect 11046 9222 11092 9274
rect 11116 9222 11162 9274
rect 11162 9222 11172 9274
rect 11196 9222 11226 9274
rect 11226 9222 11252 9274
rect 10956 9220 11012 9222
rect 11036 9220 11092 9222
rect 11116 9220 11172 9222
rect 11196 9220 11252 9222
rect 12714 20168 12770 20224
rect 15382 20304 15438 20360
rect 15566 20304 15622 20360
rect 14186 20032 14242 20088
rect 14278 19624 14334 19680
rect 15474 19780 15530 19816
rect 15474 19760 15476 19780
rect 15476 19760 15528 19780
rect 15528 19760 15530 19780
rect 11702 17040 11758 17096
rect 10782 8508 10784 8528
rect 10784 8508 10836 8528
rect 10836 8508 10838 8528
rect 10782 8472 10838 8508
rect 11518 8880 11574 8936
rect 13818 12980 13874 13016
rect 13818 12960 13820 12980
rect 13820 12960 13872 12980
rect 13872 12960 13874 12980
rect 12162 12144 12218 12200
rect 10956 8186 11012 8188
rect 11036 8186 11092 8188
rect 11116 8186 11172 8188
rect 11196 8186 11252 8188
rect 10956 8134 10982 8186
rect 10982 8134 11012 8186
rect 11036 8134 11046 8186
rect 11046 8134 11092 8186
rect 11116 8134 11162 8186
rect 11162 8134 11172 8186
rect 11196 8134 11226 8186
rect 11226 8134 11252 8186
rect 10956 8132 11012 8134
rect 11036 8132 11092 8134
rect 11116 8132 11172 8134
rect 11196 8132 11252 8134
rect 11610 7928 11666 7984
rect 11794 7928 11850 7984
rect 11242 7656 11298 7712
rect 11058 7384 11114 7440
rect 11242 7384 11298 7440
rect 10956 7098 11012 7100
rect 11036 7098 11092 7100
rect 11116 7098 11172 7100
rect 11196 7098 11252 7100
rect 10956 7046 10982 7098
rect 10982 7046 11012 7098
rect 11036 7046 11046 7098
rect 11046 7046 11092 7098
rect 11116 7046 11162 7098
rect 11162 7046 11172 7098
rect 11196 7046 11226 7098
rect 11226 7046 11252 7098
rect 10956 7044 11012 7046
rect 11036 7044 11092 7046
rect 11116 7044 11172 7046
rect 11196 7044 11252 7046
rect 10782 6996 10838 7032
rect 10782 6976 10784 6996
rect 10784 6976 10836 6996
rect 10836 6976 10838 6996
rect 10690 5888 10746 5944
rect 11426 6296 11482 6352
rect 11058 6196 11060 6216
rect 11060 6196 11112 6216
rect 11112 6196 11114 6216
rect 11058 6160 11114 6196
rect 10414 3984 10470 4040
rect 8298 2896 8354 2952
rect 10956 6010 11012 6012
rect 11036 6010 11092 6012
rect 11116 6010 11172 6012
rect 11196 6010 11252 6012
rect 10956 5958 10982 6010
rect 10982 5958 11012 6010
rect 11036 5958 11046 6010
rect 11046 5958 11092 6010
rect 11116 5958 11162 6010
rect 11162 5958 11172 6010
rect 11196 5958 11226 6010
rect 11226 5958 11252 6010
rect 10956 5956 11012 5958
rect 11036 5956 11092 5958
rect 11116 5956 11172 5958
rect 11196 5956 11252 5958
rect 11886 6296 11942 6352
rect 11426 6024 11482 6080
rect 10956 4922 11012 4924
rect 11036 4922 11092 4924
rect 11116 4922 11172 4924
rect 11196 4922 11252 4924
rect 10956 4870 10982 4922
rect 10982 4870 11012 4922
rect 11036 4870 11046 4922
rect 11046 4870 11092 4922
rect 11116 4870 11162 4922
rect 11162 4870 11172 4922
rect 11196 4870 11226 4922
rect 11226 4870 11252 4922
rect 10956 4868 11012 4870
rect 11036 4868 11092 4870
rect 11116 4868 11172 4870
rect 11196 4868 11252 4870
rect 10956 3834 11012 3836
rect 11036 3834 11092 3836
rect 11116 3834 11172 3836
rect 11196 3834 11252 3836
rect 10956 3782 10982 3834
rect 10982 3782 11012 3834
rect 11036 3782 11046 3834
rect 11046 3782 11092 3834
rect 11116 3782 11162 3834
rect 11162 3782 11172 3834
rect 11196 3782 11226 3834
rect 11226 3782 11252 3834
rect 10956 3780 11012 3782
rect 11036 3780 11092 3782
rect 11116 3780 11172 3782
rect 11196 3780 11252 3782
rect 12346 10648 12402 10704
rect 12162 10240 12218 10296
rect 13266 9968 13322 10024
rect 12254 9832 12310 9888
rect 12162 9696 12218 9752
rect 12254 8064 12310 8120
rect 12346 6432 12402 6488
rect 12898 5888 12954 5944
rect 13358 7520 13414 7576
rect 13358 6976 13414 7032
rect 12070 3576 12126 3632
rect 11886 3440 11942 3496
rect 11886 3188 11942 3224
rect 11886 3168 11888 3188
rect 11888 3168 11940 3188
rect 11940 3168 11942 3188
rect 10956 2746 11012 2748
rect 11036 2746 11092 2748
rect 11116 2746 11172 2748
rect 11196 2746 11252 2748
rect 10956 2694 10982 2746
rect 10982 2694 11012 2746
rect 11036 2694 11046 2746
rect 11046 2694 11092 2746
rect 11116 2694 11162 2746
rect 11162 2694 11172 2746
rect 11196 2694 11226 2746
rect 11226 2694 11252 2746
rect 10956 2692 11012 2694
rect 11036 2692 11092 2694
rect 11116 2692 11172 2694
rect 11196 2692 11252 2694
rect 13818 3168 13874 3224
rect 14922 9152 14978 9208
rect 15474 8608 15530 8664
rect 14738 8064 14794 8120
rect 15474 7248 15530 7304
rect 15474 5208 15530 5264
rect 15382 5072 15438 5128
rect 14370 3032 14426 3088
rect 13174 2932 13176 2952
rect 13176 2932 13228 2952
rect 13228 2932 13230 2952
rect 13174 2896 13230 2932
rect 13358 2796 13360 2816
rect 13360 2796 13412 2816
rect 13412 2796 13414 2816
rect 13358 2760 13414 2796
rect 14922 2760 14978 2816
rect 15956 21786 16012 21788
rect 16036 21786 16092 21788
rect 16116 21786 16172 21788
rect 16196 21786 16252 21788
rect 15956 21734 15982 21786
rect 15982 21734 16012 21786
rect 16036 21734 16046 21786
rect 16046 21734 16092 21786
rect 16116 21734 16162 21786
rect 16162 21734 16172 21786
rect 16196 21734 16226 21786
rect 16226 21734 16252 21786
rect 15956 21732 16012 21734
rect 16036 21732 16092 21734
rect 16116 21732 16172 21734
rect 16196 21732 16252 21734
rect 15956 20698 16012 20700
rect 16036 20698 16092 20700
rect 16116 20698 16172 20700
rect 16196 20698 16252 20700
rect 15956 20646 15982 20698
rect 15982 20646 16012 20698
rect 16036 20646 16046 20698
rect 16046 20646 16092 20698
rect 16116 20646 16162 20698
rect 16162 20646 16172 20698
rect 16196 20646 16226 20698
rect 16226 20646 16252 20698
rect 15956 20644 16012 20646
rect 16036 20644 16092 20646
rect 16116 20644 16172 20646
rect 16196 20644 16252 20646
rect 16302 20440 16358 20496
rect 16670 20476 16672 20496
rect 16672 20476 16724 20496
rect 16724 20476 16726 20496
rect 16670 20440 16726 20476
rect 16302 19760 16358 19816
rect 15956 19610 16012 19612
rect 16036 19610 16092 19612
rect 16116 19610 16172 19612
rect 16196 19610 16252 19612
rect 15956 19558 15982 19610
rect 15982 19558 16012 19610
rect 16036 19558 16046 19610
rect 16046 19558 16092 19610
rect 16116 19558 16162 19610
rect 16162 19558 16172 19610
rect 16196 19558 16226 19610
rect 16226 19558 16252 19610
rect 15956 19556 16012 19558
rect 16036 19556 16092 19558
rect 16116 19556 16172 19558
rect 16196 19556 16252 19558
rect 15956 18522 16012 18524
rect 16036 18522 16092 18524
rect 16116 18522 16172 18524
rect 16196 18522 16252 18524
rect 15956 18470 15982 18522
rect 15982 18470 16012 18522
rect 16036 18470 16046 18522
rect 16046 18470 16092 18522
rect 16116 18470 16162 18522
rect 16162 18470 16172 18522
rect 16196 18470 16226 18522
rect 16226 18470 16252 18522
rect 15956 18468 16012 18470
rect 16036 18468 16092 18470
rect 16116 18468 16172 18470
rect 16196 18468 16252 18470
rect 15956 17434 16012 17436
rect 16036 17434 16092 17436
rect 16116 17434 16172 17436
rect 16196 17434 16252 17436
rect 15956 17382 15982 17434
rect 15982 17382 16012 17434
rect 16036 17382 16046 17434
rect 16046 17382 16092 17434
rect 16116 17382 16162 17434
rect 16162 17382 16172 17434
rect 16196 17382 16226 17434
rect 16226 17382 16252 17434
rect 15956 17380 16012 17382
rect 16036 17380 16092 17382
rect 16116 17380 16172 17382
rect 16196 17380 16252 17382
rect 15956 16346 16012 16348
rect 16036 16346 16092 16348
rect 16116 16346 16172 16348
rect 16196 16346 16252 16348
rect 15956 16294 15982 16346
rect 15982 16294 16012 16346
rect 16036 16294 16046 16346
rect 16046 16294 16092 16346
rect 16116 16294 16162 16346
rect 16162 16294 16172 16346
rect 16196 16294 16226 16346
rect 16226 16294 16252 16346
rect 15956 16292 16012 16294
rect 16036 16292 16092 16294
rect 16116 16292 16172 16294
rect 16196 16292 16252 16294
rect 15956 15258 16012 15260
rect 16036 15258 16092 15260
rect 16116 15258 16172 15260
rect 16196 15258 16252 15260
rect 15956 15206 15982 15258
rect 15982 15206 16012 15258
rect 16036 15206 16046 15258
rect 16046 15206 16092 15258
rect 16116 15206 16162 15258
rect 16162 15206 16172 15258
rect 16196 15206 16226 15258
rect 16226 15206 16252 15258
rect 15956 15204 16012 15206
rect 16036 15204 16092 15206
rect 16116 15204 16172 15206
rect 16196 15204 16252 15206
rect 16302 14456 16358 14512
rect 16578 19896 16634 19952
rect 16578 19660 16580 19680
rect 16580 19660 16632 19680
rect 16632 19660 16634 19680
rect 16578 19624 16634 19660
rect 15956 14170 16012 14172
rect 16036 14170 16092 14172
rect 16116 14170 16172 14172
rect 16196 14170 16252 14172
rect 15956 14118 15982 14170
rect 15982 14118 16012 14170
rect 16036 14118 16046 14170
rect 16046 14118 16092 14170
rect 16116 14118 16162 14170
rect 16162 14118 16172 14170
rect 16196 14118 16226 14170
rect 16226 14118 16252 14170
rect 15956 14116 16012 14118
rect 16036 14116 16092 14118
rect 16116 14116 16172 14118
rect 16196 14116 16252 14118
rect 15956 13082 16012 13084
rect 16036 13082 16092 13084
rect 16116 13082 16172 13084
rect 16196 13082 16252 13084
rect 15956 13030 15982 13082
rect 15982 13030 16012 13082
rect 16036 13030 16046 13082
rect 16046 13030 16092 13082
rect 16116 13030 16162 13082
rect 16162 13030 16172 13082
rect 16196 13030 16226 13082
rect 16226 13030 16252 13082
rect 15956 13028 16012 13030
rect 16036 13028 16092 13030
rect 16116 13028 16172 13030
rect 16196 13028 16252 13030
rect 15956 11994 16012 11996
rect 16036 11994 16092 11996
rect 16116 11994 16172 11996
rect 16196 11994 16252 11996
rect 15956 11942 15982 11994
rect 15982 11942 16012 11994
rect 16036 11942 16046 11994
rect 16046 11942 16092 11994
rect 16116 11942 16162 11994
rect 16162 11942 16172 11994
rect 16196 11942 16226 11994
rect 16226 11942 16252 11994
rect 15956 11940 16012 11942
rect 16036 11940 16092 11942
rect 16116 11940 16172 11942
rect 16196 11940 16252 11942
rect 16210 11056 16266 11112
rect 15956 10906 16012 10908
rect 16036 10906 16092 10908
rect 16116 10906 16172 10908
rect 16196 10906 16252 10908
rect 15956 10854 15982 10906
rect 15982 10854 16012 10906
rect 16036 10854 16046 10906
rect 16046 10854 16092 10906
rect 16116 10854 16162 10906
rect 16162 10854 16172 10906
rect 16196 10854 16226 10906
rect 16226 10854 16252 10906
rect 15956 10852 16012 10854
rect 16036 10852 16092 10854
rect 16116 10852 16172 10854
rect 16196 10852 16252 10854
rect 15658 10648 15714 10704
rect 15956 9818 16012 9820
rect 16036 9818 16092 9820
rect 16116 9818 16172 9820
rect 16196 9818 16252 9820
rect 15956 9766 15982 9818
rect 15982 9766 16012 9818
rect 16036 9766 16046 9818
rect 16046 9766 16092 9818
rect 16116 9766 16162 9818
rect 16162 9766 16172 9818
rect 16196 9766 16226 9818
rect 16226 9766 16252 9818
rect 15956 9764 16012 9766
rect 16036 9764 16092 9766
rect 16116 9764 16172 9766
rect 16196 9764 16252 9766
rect 15956 8730 16012 8732
rect 16036 8730 16092 8732
rect 16116 8730 16172 8732
rect 16196 8730 16252 8732
rect 15956 8678 15982 8730
rect 15982 8678 16012 8730
rect 16036 8678 16046 8730
rect 16046 8678 16092 8730
rect 16116 8678 16162 8730
rect 16162 8678 16172 8730
rect 16196 8678 16226 8730
rect 16226 8678 16252 8730
rect 15956 8676 16012 8678
rect 16036 8676 16092 8678
rect 16116 8676 16172 8678
rect 16196 8676 16252 8678
rect 15956 7642 16012 7644
rect 16036 7642 16092 7644
rect 16116 7642 16172 7644
rect 16196 7642 16252 7644
rect 15956 7590 15982 7642
rect 15982 7590 16012 7642
rect 16036 7590 16046 7642
rect 16046 7590 16092 7642
rect 16116 7590 16162 7642
rect 16162 7590 16172 7642
rect 16196 7590 16226 7642
rect 16226 7590 16252 7642
rect 15956 7588 16012 7590
rect 16036 7588 16092 7590
rect 16116 7588 16172 7590
rect 16196 7588 16252 7590
rect 15956 6554 16012 6556
rect 16036 6554 16092 6556
rect 16116 6554 16172 6556
rect 16196 6554 16252 6556
rect 15956 6502 15982 6554
rect 15982 6502 16012 6554
rect 16036 6502 16046 6554
rect 16046 6502 16092 6554
rect 16116 6502 16162 6554
rect 16162 6502 16172 6554
rect 16196 6502 16226 6554
rect 16226 6502 16252 6554
rect 15956 6500 16012 6502
rect 16036 6500 16092 6502
rect 16116 6500 16172 6502
rect 16196 6500 16252 6502
rect 15956 5466 16012 5468
rect 16036 5466 16092 5468
rect 16116 5466 16172 5468
rect 16196 5466 16252 5468
rect 15956 5414 15982 5466
rect 15982 5414 16012 5466
rect 16036 5414 16046 5466
rect 16046 5414 16092 5466
rect 16116 5414 16162 5466
rect 16162 5414 16172 5466
rect 16196 5414 16226 5466
rect 16226 5414 16252 5466
rect 15956 5412 16012 5414
rect 16036 5412 16092 5414
rect 16116 5412 16172 5414
rect 16196 5412 16252 5414
rect 15934 4820 15990 4856
rect 15934 4800 15936 4820
rect 15936 4800 15988 4820
rect 15988 4800 15990 4820
rect 15956 4378 16012 4380
rect 16036 4378 16092 4380
rect 16116 4378 16172 4380
rect 16196 4378 16252 4380
rect 15956 4326 15982 4378
rect 15982 4326 16012 4378
rect 16036 4326 16046 4378
rect 16046 4326 16092 4378
rect 16116 4326 16162 4378
rect 16162 4326 16172 4378
rect 16196 4326 16226 4378
rect 16226 4326 16252 4378
rect 15956 4324 16012 4326
rect 16036 4324 16092 4326
rect 16116 4324 16172 4326
rect 16196 4324 16252 4326
rect 15956 3290 16012 3292
rect 16036 3290 16092 3292
rect 16116 3290 16172 3292
rect 16196 3290 16252 3292
rect 15956 3238 15982 3290
rect 15982 3238 16012 3290
rect 16036 3238 16046 3290
rect 16046 3238 16092 3290
rect 16116 3238 16162 3290
rect 16162 3238 16172 3290
rect 16196 3238 16226 3290
rect 16226 3238 16252 3290
rect 15956 3236 16012 3238
rect 16036 3236 16092 3238
rect 16116 3236 16172 3238
rect 16196 3236 16252 3238
rect 15956 2202 16012 2204
rect 16036 2202 16092 2204
rect 16116 2202 16172 2204
rect 16196 2202 16252 2204
rect 15956 2150 15982 2202
rect 15982 2150 16012 2202
rect 16036 2150 16046 2202
rect 16046 2150 16092 2202
rect 16116 2150 16162 2202
rect 16162 2150 16172 2202
rect 16196 2150 16226 2202
rect 16226 2150 16252 2202
rect 15956 2148 16012 2150
rect 16036 2148 16092 2150
rect 16116 2148 16172 2150
rect 16196 2148 16252 2150
rect 16578 9968 16634 10024
rect 16670 9172 16726 9208
rect 16670 9152 16672 9172
rect 16672 9152 16724 9172
rect 16724 9152 16726 9172
rect 16762 8608 16818 8664
rect 16946 7792 17002 7848
rect 16946 7284 16948 7304
rect 16948 7284 17000 7304
rect 17000 7284 17002 7304
rect 16946 7248 17002 7284
rect 18050 19488 18106 19544
rect 17498 15272 17554 15328
rect 17130 10920 17186 10976
rect 17314 10784 17370 10840
rect 17130 10240 17186 10296
rect 17406 10104 17462 10160
rect 17774 9444 17830 9480
rect 17774 9424 17776 9444
rect 17776 9424 17828 9444
rect 17828 9424 17830 9444
rect 15658 1944 15714 2000
rect 18234 20596 18290 20632
rect 18234 20576 18236 20596
rect 18236 20576 18288 20596
rect 18288 20576 18290 20596
rect 20956 21242 21012 21244
rect 21036 21242 21092 21244
rect 21116 21242 21172 21244
rect 21196 21242 21252 21244
rect 20956 21190 20982 21242
rect 20982 21190 21012 21242
rect 21036 21190 21046 21242
rect 21046 21190 21092 21242
rect 21116 21190 21162 21242
rect 21162 21190 21172 21242
rect 21196 21190 21226 21242
rect 21226 21190 21252 21242
rect 20956 21188 21012 21190
rect 21036 21188 21092 21190
rect 21116 21188 21172 21190
rect 21196 21188 21252 21190
rect 25502 22344 25558 22400
rect 25410 21528 25466 21584
rect 24674 20576 24730 20632
rect 23202 20440 23258 20496
rect 19982 20168 20038 20224
rect 19522 19624 19578 19680
rect 18142 3596 18198 3598
rect 18142 3544 18144 3596
rect 18144 3544 18196 3596
rect 18196 3544 18198 3596
rect 18142 3542 18198 3544
rect 18326 13776 18382 13832
rect 18694 10784 18750 10840
rect 18326 10124 18382 10160
rect 18326 10104 18328 10124
rect 18328 10104 18380 10124
rect 18380 10104 18382 10124
rect 18326 4800 18382 4856
rect 18602 4120 18658 4176
rect 18234 2488 18290 2544
rect 18970 9988 19026 10024
rect 18970 9968 18972 9988
rect 18972 9968 19024 9988
rect 19024 9968 19026 9988
rect 19246 12824 19302 12880
rect 21730 20304 21786 20360
rect 20956 20154 21012 20156
rect 21036 20154 21092 20156
rect 21116 20154 21172 20156
rect 21196 20154 21252 20156
rect 20956 20102 20982 20154
rect 20982 20102 21012 20154
rect 21036 20102 21046 20154
rect 21046 20102 21092 20154
rect 21116 20102 21162 20154
rect 21162 20102 21172 20154
rect 21196 20102 21226 20154
rect 21226 20102 21252 20154
rect 20956 20100 21012 20102
rect 21036 20100 21092 20102
rect 21116 20100 21172 20102
rect 21196 20100 21252 20102
rect 20810 20032 20866 20088
rect 20956 19066 21012 19068
rect 21036 19066 21092 19068
rect 21116 19066 21172 19068
rect 21196 19066 21252 19068
rect 20956 19014 20982 19066
rect 20982 19014 21012 19066
rect 21036 19014 21046 19066
rect 21046 19014 21092 19066
rect 21116 19014 21162 19066
rect 21162 19014 21172 19066
rect 21196 19014 21226 19066
rect 21226 19014 21252 19066
rect 20956 19012 21012 19014
rect 21036 19012 21092 19014
rect 21116 19012 21172 19014
rect 21196 19012 21252 19014
rect 20718 18672 20774 18728
rect 20166 12416 20222 12472
rect 19062 6976 19118 7032
rect 19982 9288 20038 9344
rect 19982 8336 20038 8392
rect 19890 7928 19946 7984
rect 19614 6704 19670 6760
rect 19154 5888 19210 5944
rect 19798 6316 19854 6352
rect 19798 6296 19800 6316
rect 19800 6296 19852 6316
rect 19852 6296 19854 6316
rect 19982 5208 20038 5264
rect 19614 5072 19670 5128
rect 17866 1400 17922 1456
rect 19246 2372 19302 2408
rect 19246 2352 19248 2372
rect 19248 2352 19300 2372
rect 19300 2352 19302 2372
rect 19154 856 19210 912
rect 20258 12280 20314 12336
rect 20534 3032 20590 3088
rect 20258 2896 20314 2952
rect 20956 17978 21012 17980
rect 21036 17978 21092 17980
rect 21116 17978 21172 17980
rect 21196 17978 21252 17980
rect 20956 17926 20982 17978
rect 20982 17926 21012 17978
rect 21036 17926 21046 17978
rect 21046 17926 21092 17978
rect 21116 17926 21162 17978
rect 21162 17926 21172 17978
rect 21196 17926 21226 17978
rect 21226 17926 21252 17978
rect 20956 17924 21012 17926
rect 21036 17924 21092 17926
rect 21116 17924 21172 17926
rect 21196 17924 21252 17926
rect 20956 16890 21012 16892
rect 21036 16890 21092 16892
rect 21116 16890 21172 16892
rect 21196 16890 21252 16892
rect 20956 16838 20982 16890
rect 20982 16838 21012 16890
rect 21036 16838 21046 16890
rect 21046 16838 21092 16890
rect 21116 16838 21162 16890
rect 21162 16838 21172 16890
rect 21196 16838 21226 16890
rect 21226 16838 21252 16890
rect 20956 16836 21012 16838
rect 21036 16836 21092 16838
rect 21116 16836 21172 16838
rect 21196 16836 21252 16838
rect 20956 15802 21012 15804
rect 21036 15802 21092 15804
rect 21116 15802 21172 15804
rect 21196 15802 21252 15804
rect 20956 15750 20982 15802
rect 20982 15750 21012 15802
rect 21036 15750 21046 15802
rect 21046 15750 21092 15802
rect 21116 15750 21162 15802
rect 21162 15750 21172 15802
rect 21196 15750 21226 15802
rect 21226 15750 21252 15802
rect 20956 15748 21012 15750
rect 21036 15748 21092 15750
rect 21116 15748 21172 15750
rect 21196 15748 21252 15750
rect 20956 14714 21012 14716
rect 21036 14714 21092 14716
rect 21116 14714 21172 14716
rect 21196 14714 21252 14716
rect 20956 14662 20982 14714
rect 20982 14662 21012 14714
rect 21036 14662 21046 14714
rect 21046 14662 21092 14714
rect 21116 14662 21162 14714
rect 21162 14662 21172 14714
rect 21196 14662 21226 14714
rect 21226 14662 21252 14714
rect 20956 14660 21012 14662
rect 21036 14660 21092 14662
rect 21116 14660 21172 14662
rect 21196 14660 21252 14662
rect 20956 13626 21012 13628
rect 21036 13626 21092 13628
rect 21116 13626 21172 13628
rect 21196 13626 21252 13628
rect 20956 13574 20982 13626
rect 20982 13574 21012 13626
rect 21036 13574 21046 13626
rect 21046 13574 21092 13626
rect 21116 13574 21162 13626
rect 21162 13574 21172 13626
rect 21196 13574 21226 13626
rect 21226 13574 21252 13626
rect 20956 13572 21012 13574
rect 21036 13572 21092 13574
rect 21116 13572 21172 13574
rect 21196 13572 21252 13574
rect 20956 12538 21012 12540
rect 21036 12538 21092 12540
rect 21116 12538 21172 12540
rect 21196 12538 21252 12540
rect 20956 12486 20982 12538
rect 20982 12486 21012 12538
rect 21036 12486 21046 12538
rect 21046 12486 21092 12538
rect 21116 12486 21162 12538
rect 21162 12486 21172 12538
rect 21196 12486 21226 12538
rect 21226 12486 21252 12538
rect 20956 12484 21012 12486
rect 21036 12484 21092 12486
rect 21116 12484 21172 12486
rect 21196 12484 21252 12486
rect 20956 11450 21012 11452
rect 21036 11450 21092 11452
rect 21116 11450 21172 11452
rect 21196 11450 21252 11452
rect 20956 11398 20982 11450
rect 20982 11398 21012 11450
rect 21036 11398 21046 11450
rect 21046 11398 21092 11450
rect 21116 11398 21162 11450
rect 21162 11398 21172 11450
rect 21196 11398 21226 11450
rect 21226 11398 21252 11450
rect 20956 11396 21012 11398
rect 21036 11396 21092 11398
rect 21116 11396 21172 11398
rect 21196 11396 21252 11398
rect 20956 10362 21012 10364
rect 21036 10362 21092 10364
rect 21116 10362 21172 10364
rect 21196 10362 21252 10364
rect 20956 10310 20982 10362
rect 20982 10310 21012 10362
rect 21036 10310 21046 10362
rect 21046 10310 21092 10362
rect 21116 10310 21162 10362
rect 21162 10310 21172 10362
rect 21196 10310 21226 10362
rect 21226 10310 21252 10362
rect 20956 10308 21012 10310
rect 21036 10308 21092 10310
rect 21116 10308 21172 10310
rect 21196 10308 21252 10310
rect 20956 9274 21012 9276
rect 21036 9274 21092 9276
rect 21116 9274 21172 9276
rect 21196 9274 21252 9276
rect 20956 9222 20982 9274
rect 20982 9222 21012 9274
rect 21036 9222 21046 9274
rect 21046 9222 21092 9274
rect 21116 9222 21162 9274
rect 21162 9222 21172 9274
rect 21196 9222 21226 9274
rect 21226 9222 21252 9274
rect 20956 9220 21012 9222
rect 21036 9220 21092 9222
rect 21116 9220 21172 9222
rect 21196 9220 21252 9222
rect 20810 8236 20812 8256
rect 20812 8236 20864 8256
rect 20864 8236 20866 8256
rect 20810 8200 20866 8236
rect 20956 8186 21012 8188
rect 21036 8186 21092 8188
rect 21116 8186 21172 8188
rect 21196 8186 21252 8188
rect 20956 8134 20982 8186
rect 20982 8134 21012 8186
rect 21036 8134 21046 8186
rect 21046 8134 21092 8186
rect 21116 8134 21162 8186
rect 21162 8134 21172 8186
rect 21196 8134 21226 8186
rect 21226 8134 21252 8186
rect 20956 8132 21012 8134
rect 21036 8132 21092 8134
rect 21116 8132 21172 8134
rect 21196 8132 21252 8134
rect 20956 7098 21012 7100
rect 21036 7098 21092 7100
rect 21116 7098 21172 7100
rect 21196 7098 21252 7100
rect 20956 7046 20982 7098
rect 20982 7046 21012 7098
rect 21036 7046 21046 7098
rect 21046 7046 21092 7098
rect 21116 7046 21162 7098
rect 21162 7046 21172 7098
rect 21196 7046 21226 7098
rect 21226 7046 21252 7098
rect 20956 7044 21012 7046
rect 21036 7044 21092 7046
rect 21116 7044 21172 7046
rect 21196 7044 21252 7046
rect 20810 6060 20812 6080
rect 20812 6060 20864 6080
rect 20864 6060 20866 6080
rect 20810 6024 20866 6060
rect 20956 6010 21012 6012
rect 21036 6010 21092 6012
rect 21116 6010 21172 6012
rect 21196 6010 21252 6012
rect 20956 5958 20982 6010
rect 20982 5958 21012 6010
rect 21036 5958 21046 6010
rect 21046 5958 21092 6010
rect 21116 5958 21162 6010
rect 21162 5958 21172 6010
rect 21196 5958 21226 6010
rect 21226 5958 21252 6010
rect 20956 5956 21012 5958
rect 21036 5956 21092 5958
rect 21116 5956 21172 5958
rect 21196 5956 21252 5958
rect 20810 5616 20866 5672
rect 20956 4922 21012 4924
rect 21036 4922 21092 4924
rect 21116 4922 21172 4924
rect 21196 4922 21252 4924
rect 20956 4870 20982 4922
rect 20982 4870 21012 4922
rect 21036 4870 21046 4922
rect 21046 4870 21092 4922
rect 21116 4870 21162 4922
rect 21162 4870 21172 4922
rect 21196 4870 21226 4922
rect 21226 4870 21252 4922
rect 20956 4868 21012 4870
rect 21036 4868 21092 4870
rect 21116 4868 21172 4870
rect 21196 4868 21252 4870
rect 20956 3834 21012 3836
rect 21036 3834 21092 3836
rect 21116 3834 21172 3836
rect 21196 3834 21252 3836
rect 20956 3782 20982 3834
rect 20982 3782 21012 3834
rect 21036 3782 21046 3834
rect 21046 3782 21092 3834
rect 21116 3782 21162 3834
rect 21162 3782 21172 3834
rect 21196 3782 21226 3834
rect 21226 3782 21252 3834
rect 20956 3780 21012 3782
rect 21036 3780 21092 3782
rect 21116 3780 21172 3782
rect 21196 3780 21252 3782
rect 24398 20304 24454 20360
rect 24950 20168 25006 20224
rect 24214 19488 24270 19544
rect 25410 19896 25466 19952
rect 25226 19352 25282 19408
rect 25134 18808 25190 18864
rect 25042 15816 25098 15872
rect 24858 14592 24914 14648
rect 24766 13368 24822 13424
rect 24950 13912 25006 13968
rect 25318 15408 25374 15464
rect 25226 12960 25282 13016
rect 25134 12688 25190 12744
rect 25042 12144 25098 12200
rect 25410 14456 25466 14512
rect 25410 13368 25466 13424
rect 25318 10920 25374 10976
rect 24950 9968 25006 10024
rect 25594 19624 25650 19680
rect 25594 18264 25650 18320
rect 25502 11600 25558 11656
rect 25870 23024 25926 23080
rect 25778 21256 25834 21312
rect 25778 20476 25780 20496
rect 25780 20476 25832 20496
rect 25832 20476 25834 20496
rect 25778 20440 25834 20476
rect 25778 17040 25834 17096
rect 25956 21786 26012 21788
rect 26036 21786 26092 21788
rect 26116 21786 26172 21788
rect 26196 21786 26252 21788
rect 25956 21734 25982 21786
rect 25982 21734 26012 21786
rect 26036 21734 26046 21786
rect 26046 21734 26092 21786
rect 26116 21734 26162 21786
rect 26162 21734 26172 21786
rect 26196 21734 26226 21786
rect 26226 21734 26252 21786
rect 25956 21732 26012 21734
rect 26036 21732 26092 21734
rect 26116 21732 26172 21734
rect 26196 21732 26252 21734
rect 25956 20698 26012 20700
rect 26036 20698 26092 20700
rect 26116 20698 26172 20700
rect 26196 20698 26252 20700
rect 25956 20646 25982 20698
rect 25982 20646 26012 20698
rect 26036 20646 26046 20698
rect 26046 20646 26092 20698
rect 26116 20646 26162 20698
rect 26162 20646 26172 20698
rect 26196 20646 26226 20698
rect 26226 20646 26252 20698
rect 25956 20644 26012 20646
rect 26036 20644 26092 20646
rect 26116 20644 26172 20646
rect 26196 20644 26252 20646
rect 27710 20440 27766 20496
rect 26422 20304 26478 20360
rect 26698 20052 26754 20088
rect 26698 20032 26700 20052
rect 26700 20032 26752 20052
rect 26752 20032 26754 20052
rect 25956 19610 26012 19612
rect 26036 19610 26092 19612
rect 26116 19610 26172 19612
rect 26196 19610 26252 19612
rect 25956 19558 25982 19610
rect 25982 19558 26012 19610
rect 26036 19558 26046 19610
rect 26046 19558 26092 19610
rect 26116 19558 26162 19610
rect 26162 19558 26172 19610
rect 26196 19558 26226 19610
rect 26226 19558 26252 19610
rect 25956 19556 26012 19558
rect 26036 19556 26092 19558
rect 26116 19556 26172 19558
rect 26196 19556 26252 19558
rect 26882 19760 26938 19816
rect 26514 18672 26570 18728
rect 25956 18522 26012 18524
rect 26036 18522 26092 18524
rect 26116 18522 26172 18524
rect 26196 18522 26252 18524
rect 25956 18470 25982 18522
rect 25982 18470 26012 18522
rect 26036 18470 26046 18522
rect 26046 18470 26092 18522
rect 26116 18470 26162 18522
rect 26162 18470 26172 18522
rect 26196 18470 26226 18522
rect 26226 18470 26252 18522
rect 25956 18468 26012 18470
rect 26036 18468 26092 18470
rect 26116 18468 26172 18470
rect 26196 18468 26252 18470
rect 25956 17434 26012 17436
rect 26036 17434 26092 17436
rect 26116 17434 26172 17436
rect 26196 17434 26252 17436
rect 25956 17382 25982 17434
rect 25982 17382 26012 17434
rect 26036 17382 26046 17434
rect 26046 17382 26092 17434
rect 26116 17382 26162 17434
rect 26162 17382 26172 17434
rect 26196 17382 26226 17434
rect 26226 17382 26252 17434
rect 25956 17380 26012 17382
rect 26036 17380 26092 17382
rect 26116 17380 26172 17382
rect 26196 17380 26252 17382
rect 25956 16346 26012 16348
rect 26036 16346 26092 16348
rect 26116 16346 26172 16348
rect 26196 16346 26252 16348
rect 25956 16294 25982 16346
rect 25982 16294 26012 16346
rect 26036 16294 26046 16346
rect 26046 16294 26092 16346
rect 26116 16294 26162 16346
rect 26162 16294 26172 16346
rect 26196 16294 26226 16346
rect 26226 16294 26252 16346
rect 25956 16292 26012 16294
rect 26036 16292 26092 16294
rect 26116 16292 26172 16294
rect 26196 16292 26252 16294
rect 25870 16088 25926 16144
rect 25778 15272 25834 15328
rect 25686 11056 25742 11112
rect 25594 9016 25650 9072
rect 25956 15258 26012 15260
rect 26036 15258 26092 15260
rect 26116 15258 26172 15260
rect 26196 15258 26252 15260
rect 25956 15206 25982 15258
rect 25982 15206 26012 15258
rect 26036 15206 26046 15258
rect 26046 15206 26092 15258
rect 26116 15206 26162 15258
rect 26162 15206 26172 15258
rect 26196 15206 26226 15258
rect 26226 15206 26252 15258
rect 25956 15204 26012 15206
rect 26036 15204 26092 15206
rect 26116 15204 26172 15206
rect 26196 15204 26252 15206
rect 25956 14170 26012 14172
rect 26036 14170 26092 14172
rect 26116 14170 26172 14172
rect 26196 14170 26252 14172
rect 25956 14118 25982 14170
rect 25982 14118 26012 14170
rect 26036 14118 26046 14170
rect 26046 14118 26092 14170
rect 26116 14118 26162 14170
rect 26162 14118 26172 14170
rect 26196 14118 26226 14170
rect 26226 14118 26252 14170
rect 25956 14116 26012 14118
rect 26036 14116 26092 14118
rect 26116 14116 26172 14118
rect 26196 14116 26252 14118
rect 25870 13776 25926 13832
rect 25956 13082 26012 13084
rect 26036 13082 26092 13084
rect 26116 13082 26172 13084
rect 26196 13082 26252 13084
rect 25956 13030 25982 13082
rect 25982 13030 26012 13082
rect 26036 13030 26046 13082
rect 26046 13030 26092 13082
rect 26116 13030 26162 13082
rect 26162 13030 26172 13082
rect 26196 13030 26226 13082
rect 26226 13030 26252 13082
rect 25956 13028 26012 13030
rect 26036 13028 26092 13030
rect 26116 13028 26172 13030
rect 26196 13028 26252 13030
rect 25870 12280 25926 12336
rect 25778 8608 25834 8664
rect 25410 8336 25466 8392
rect 21362 8236 21364 8256
rect 21364 8236 21416 8256
rect 21416 8236 21418 8256
rect 21362 8200 21418 8236
rect 21914 8200 21970 8256
rect 24858 8200 24914 8256
rect 25956 11994 26012 11996
rect 26036 11994 26092 11996
rect 26116 11994 26172 11996
rect 26196 11994 26252 11996
rect 25956 11942 25982 11994
rect 25982 11942 26012 11994
rect 26036 11942 26046 11994
rect 26046 11942 26092 11994
rect 26116 11942 26162 11994
rect 26162 11942 26172 11994
rect 26196 11942 26226 11994
rect 26226 11942 26252 11994
rect 25956 11940 26012 11942
rect 26036 11940 26092 11942
rect 26116 11940 26172 11942
rect 26196 11940 26252 11942
rect 26422 11736 26478 11792
rect 26698 11600 26754 11656
rect 25956 10906 26012 10908
rect 26036 10906 26092 10908
rect 26116 10906 26172 10908
rect 26196 10906 26252 10908
rect 25956 10854 25982 10906
rect 25982 10854 26012 10906
rect 26036 10854 26046 10906
rect 26046 10854 26092 10906
rect 26116 10854 26162 10906
rect 26162 10854 26172 10906
rect 26196 10854 26226 10906
rect 26226 10854 26252 10906
rect 25956 10852 26012 10854
rect 26036 10852 26092 10854
rect 26116 10852 26172 10854
rect 26196 10852 26252 10854
rect 26606 11056 26662 11112
rect 26514 10648 26570 10704
rect 26422 10548 26424 10568
rect 26424 10548 26476 10568
rect 26476 10548 26478 10568
rect 26422 10512 26478 10548
rect 26606 10412 26608 10432
rect 26608 10412 26660 10432
rect 26660 10412 26662 10432
rect 26606 10376 26662 10412
rect 26790 10104 26846 10160
rect 26698 9832 26754 9888
rect 25956 9818 26012 9820
rect 26036 9818 26092 9820
rect 26116 9818 26172 9820
rect 26196 9818 26252 9820
rect 25956 9766 25982 9818
rect 25982 9766 26012 9818
rect 26036 9766 26046 9818
rect 26046 9766 26092 9818
rect 26116 9766 26162 9818
rect 26162 9766 26172 9818
rect 26196 9766 26226 9818
rect 26226 9766 26252 9818
rect 25956 9764 26012 9766
rect 26036 9764 26092 9766
rect 26116 9764 26172 9766
rect 26196 9764 26252 9766
rect 26606 9288 26662 9344
rect 26514 8880 26570 8936
rect 25956 8730 26012 8732
rect 26036 8730 26092 8732
rect 26116 8730 26172 8732
rect 26196 8730 26252 8732
rect 25956 8678 25982 8730
rect 25982 8678 26012 8730
rect 26036 8678 26046 8730
rect 26046 8678 26092 8730
rect 26116 8678 26162 8730
rect 26162 8678 26172 8730
rect 26196 8678 26226 8730
rect 26226 8678 26252 8730
rect 25956 8676 26012 8678
rect 26036 8676 26092 8678
rect 26116 8676 26172 8678
rect 26196 8676 26252 8678
rect 26698 8608 26754 8664
rect 26422 8472 26478 8528
rect 25870 7928 25926 7984
rect 25956 7642 26012 7644
rect 26036 7642 26092 7644
rect 26116 7642 26172 7644
rect 26196 7642 26252 7644
rect 25956 7590 25982 7642
rect 25982 7590 26012 7642
rect 26036 7590 26046 7642
rect 26046 7590 26092 7642
rect 26116 7590 26162 7642
rect 26162 7590 26172 7642
rect 26196 7590 26226 7642
rect 26226 7590 26252 7642
rect 25956 7588 26012 7590
rect 26036 7588 26092 7590
rect 26116 7588 26172 7590
rect 26196 7588 26252 7590
rect 26422 7384 26478 7440
rect 26698 7384 26754 7440
rect 26514 7248 26570 7304
rect 26606 6976 26662 7032
rect 26514 6860 26570 6896
rect 26514 6840 26516 6860
rect 26516 6840 26568 6860
rect 26568 6840 26570 6860
rect 25956 6554 26012 6556
rect 26036 6554 26092 6556
rect 26116 6554 26172 6556
rect 26196 6554 26252 6556
rect 25956 6502 25982 6554
rect 25982 6502 26012 6554
rect 26036 6502 26046 6554
rect 26046 6502 26092 6554
rect 26116 6502 26162 6554
rect 26162 6502 26172 6554
rect 26196 6502 26226 6554
rect 26226 6502 26252 6554
rect 25956 6500 26012 6502
rect 26036 6500 26092 6502
rect 26116 6500 26172 6502
rect 26196 6500 26252 6502
rect 26330 6296 26386 6352
rect 26606 6332 26608 6352
rect 26608 6332 26660 6352
rect 26660 6332 26662 6352
rect 26606 6296 26662 6332
rect 25318 5616 25374 5672
rect 25956 5466 26012 5468
rect 26036 5466 26092 5468
rect 26116 5466 26172 5468
rect 26196 5466 26252 5468
rect 25956 5414 25982 5466
rect 25982 5414 26012 5466
rect 26036 5414 26046 5466
rect 26046 5414 26092 5466
rect 26116 5414 26162 5466
rect 26162 5414 26172 5466
rect 26196 5414 26226 5466
rect 26226 5414 26252 5466
rect 25956 5412 26012 5414
rect 26036 5412 26092 5414
rect 26116 5412 26172 5414
rect 26196 5412 26252 5414
rect 21270 3576 21326 3632
rect 23202 3576 23258 3632
rect 22190 2896 22246 2952
rect 20956 2746 21012 2748
rect 21036 2746 21092 2748
rect 21116 2746 21172 2748
rect 21196 2746 21252 2748
rect 20956 2694 20982 2746
rect 20982 2694 21012 2746
rect 21036 2694 21046 2746
rect 21046 2694 21092 2746
rect 21116 2694 21162 2746
rect 21162 2694 21172 2746
rect 21196 2694 21226 2746
rect 21226 2694 21252 2746
rect 20956 2692 21012 2694
rect 21036 2692 21092 2694
rect 21116 2692 21172 2694
rect 21196 2692 21252 2694
rect 25318 3032 25374 3088
rect 25502 2896 25558 2952
rect 25956 4378 26012 4380
rect 26036 4378 26092 4380
rect 26116 4378 26172 4380
rect 26196 4378 26252 4380
rect 25956 4326 25982 4378
rect 25982 4326 26012 4378
rect 26036 4326 26046 4378
rect 26046 4326 26092 4378
rect 26116 4326 26162 4378
rect 26162 4326 26172 4378
rect 26196 4326 26226 4378
rect 26226 4326 26252 4378
rect 25956 4324 26012 4326
rect 26036 4324 26092 4326
rect 26116 4324 26172 4326
rect 26196 4324 26252 4326
rect 25956 3290 26012 3292
rect 26036 3290 26092 3292
rect 26116 3290 26172 3292
rect 26196 3290 26252 3292
rect 25956 3238 25982 3290
rect 25982 3238 26012 3290
rect 26036 3238 26046 3290
rect 26046 3238 26092 3290
rect 26116 3238 26162 3290
rect 26162 3238 26172 3290
rect 26196 3238 26226 3290
rect 26226 3238 26252 3290
rect 25956 3236 26012 3238
rect 26036 3236 26092 3238
rect 26116 3236 26172 3238
rect 26196 3236 26252 3238
rect 26514 6160 26570 6216
rect 26422 5752 26478 5808
rect 26698 5636 26754 5672
rect 26698 5616 26700 5636
rect 26700 5616 26752 5636
rect 26752 5616 26754 5636
rect 26422 5108 26424 5128
rect 26424 5108 26476 5128
rect 26476 5108 26478 5128
rect 26422 5072 26478 5108
rect 26606 5072 26662 5128
rect 29182 20032 29238 20088
rect 27526 9424 27582 9480
rect 27710 8336 27766 8392
rect 27250 6704 27306 6760
rect 28354 6704 28410 6760
rect 26882 5208 26938 5264
rect 26698 4428 26700 4448
rect 26700 4428 26752 4448
rect 26752 4428 26754 4448
rect 26698 4392 26754 4428
rect 26422 4020 26424 4040
rect 26424 4020 26476 4040
rect 26476 4020 26478 4040
rect 26422 3984 26478 4020
rect 26606 3884 26608 3904
rect 26608 3884 26660 3904
rect 26660 3884 26662 3904
rect 26606 3848 26662 3884
rect 26698 3340 26700 3360
rect 26700 3340 26752 3360
rect 26752 3340 26754 3360
rect 26698 3304 26754 3340
rect 25870 2760 25926 2816
rect 25778 2624 25834 2680
rect 24398 2508 24454 2544
rect 24398 2488 24400 2508
rect 24400 2488 24452 2508
rect 24452 2488 24454 2508
rect 25956 2202 26012 2204
rect 26036 2202 26092 2204
rect 26116 2202 26172 2204
rect 26196 2202 26252 2204
rect 25956 2150 25982 2202
rect 25982 2150 26012 2202
rect 26036 2150 26046 2202
rect 26046 2150 26092 2202
rect 26116 2150 26162 2202
rect 26162 2150 26172 2202
rect 26196 2150 26226 2202
rect 26226 2150 26252 2202
rect 25956 2148 26012 2150
rect 26036 2148 26092 2150
rect 26116 2148 26172 2150
rect 26196 2148 26252 2150
rect 24214 1944 24270 2000
rect 25226 1400 25282 1456
rect 2778 312 2834 368
rect 27342 2896 27398 2952
rect 27066 1400 27122 1456
rect 29366 2760 29422 2816
rect 26606 312 26662 368
<< metal3 >>
rect 0 23626 480 23656
rect 2957 23626 3023 23629
rect 0 23624 3023 23626
rect 0 23568 2962 23624
rect 3018 23568 3023 23624
rect 0 23566 3023 23568
rect 0 23536 480 23566
rect 2957 23563 3023 23566
rect 25681 23626 25747 23629
rect 29520 23626 30000 23656
rect 25681 23624 30000 23626
rect 25681 23568 25686 23624
rect 25742 23568 30000 23624
rect 25681 23566 30000 23568
rect 25681 23563 25747 23566
rect 29520 23536 30000 23566
rect 0 23082 480 23112
rect 3141 23082 3207 23085
rect 0 23080 3207 23082
rect 0 23024 3146 23080
rect 3202 23024 3207 23080
rect 0 23022 3207 23024
rect 0 22992 480 23022
rect 3141 23019 3207 23022
rect 25865 23082 25931 23085
rect 29520 23082 30000 23112
rect 25865 23080 30000 23082
rect 25865 23024 25870 23080
rect 25926 23024 30000 23080
rect 25865 23022 30000 23024
rect 25865 23019 25931 23022
rect 29520 22992 30000 23022
rect 0 22402 480 22432
rect 2865 22402 2931 22405
rect 0 22400 2931 22402
rect 0 22344 2870 22400
rect 2926 22344 2931 22400
rect 0 22342 2931 22344
rect 0 22312 480 22342
rect 2865 22339 2931 22342
rect 25497 22402 25563 22405
rect 29520 22402 30000 22432
rect 25497 22400 30000 22402
rect 25497 22344 25502 22400
rect 25558 22344 30000 22400
rect 25497 22342 30000 22344
rect 25497 22339 25563 22342
rect 29520 22312 30000 22342
rect 0 21858 480 21888
rect 3877 21858 3943 21861
rect 29520 21858 30000 21888
rect 0 21856 3943 21858
rect 0 21800 3882 21856
rect 3938 21800 3943 21856
rect 0 21798 3943 21800
rect 0 21768 480 21798
rect 3877 21795 3943 21798
rect 26374 21798 30000 21858
rect 5944 21792 6264 21793
rect 5944 21728 5952 21792
rect 6016 21728 6032 21792
rect 6096 21728 6112 21792
rect 6176 21728 6192 21792
rect 6256 21728 6264 21792
rect 5944 21727 6264 21728
rect 15944 21792 16264 21793
rect 15944 21728 15952 21792
rect 16016 21728 16032 21792
rect 16096 21728 16112 21792
rect 16176 21728 16192 21792
rect 16256 21728 16264 21792
rect 15944 21727 16264 21728
rect 25944 21792 26264 21793
rect 25944 21728 25952 21792
rect 26016 21728 26032 21792
rect 26096 21728 26112 21792
rect 26176 21728 26192 21792
rect 26256 21728 26264 21792
rect 25944 21727 26264 21728
rect 25405 21586 25471 21589
rect 26374 21586 26434 21798
rect 29520 21768 30000 21798
rect 25405 21584 26434 21586
rect 25405 21528 25410 21584
rect 25466 21528 26434 21584
rect 25405 21526 26434 21528
rect 25405 21523 25471 21526
rect 0 21314 480 21344
rect 3509 21314 3575 21317
rect 0 21312 3575 21314
rect 0 21256 3514 21312
rect 3570 21256 3575 21312
rect 0 21254 3575 21256
rect 0 21224 480 21254
rect 3509 21251 3575 21254
rect 25773 21314 25839 21317
rect 29520 21314 30000 21344
rect 25773 21312 30000 21314
rect 25773 21256 25778 21312
rect 25834 21256 30000 21312
rect 25773 21254 30000 21256
rect 25773 21251 25839 21254
rect 10944 21248 11264 21249
rect 10944 21184 10952 21248
rect 11016 21184 11032 21248
rect 11096 21184 11112 21248
rect 11176 21184 11192 21248
rect 11256 21184 11264 21248
rect 10944 21183 11264 21184
rect 20944 21248 21264 21249
rect 20944 21184 20952 21248
rect 21016 21184 21032 21248
rect 21096 21184 21112 21248
rect 21176 21184 21192 21248
rect 21256 21184 21264 21248
rect 29520 21224 30000 21254
rect 20944 21183 21264 21184
rect 5944 20704 6264 20705
rect 0 20634 480 20664
rect 5944 20640 5952 20704
rect 6016 20640 6032 20704
rect 6096 20640 6112 20704
rect 6176 20640 6192 20704
rect 6256 20640 6264 20704
rect 5944 20639 6264 20640
rect 15944 20704 16264 20705
rect 15944 20640 15952 20704
rect 16016 20640 16032 20704
rect 16096 20640 16112 20704
rect 16176 20640 16192 20704
rect 16256 20640 16264 20704
rect 15944 20639 16264 20640
rect 25944 20704 26264 20705
rect 25944 20640 25952 20704
rect 26016 20640 26032 20704
rect 26096 20640 26112 20704
rect 26176 20640 26192 20704
rect 26256 20640 26264 20704
rect 25944 20639 26264 20640
rect 3233 20634 3299 20637
rect 0 20632 3299 20634
rect 0 20576 3238 20632
rect 3294 20576 3299 20632
rect 0 20574 3299 20576
rect 0 20544 480 20574
rect 3233 20571 3299 20574
rect 18229 20634 18295 20637
rect 24669 20634 24735 20637
rect 29520 20634 30000 20664
rect 18229 20632 24735 20634
rect 18229 20576 18234 20632
rect 18290 20576 24674 20632
rect 24730 20576 24735 20632
rect 18229 20574 24735 20576
rect 18229 20571 18295 20574
rect 24669 20571 24735 20574
rect 27846 20574 30000 20634
rect 9673 20498 9739 20501
rect 16297 20498 16363 20501
rect 9673 20496 16363 20498
rect 9673 20440 9678 20496
rect 9734 20440 16302 20496
rect 16358 20440 16363 20496
rect 9673 20438 16363 20440
rect 9673 20435 9739 20438
rect 16297 20435 16363 20438
rect 16665 20498 16731 20501
rect 23197 20498 23263 20501
rect 16665 20496 23263 20498
rect 16665 20440 16670 20496
rect 16726 20440 23202 20496
rect 23258 20440 23263 20496
rect 16665 20438 23263 20440
rect 16665 20435 16731 20438
rect 23197 20435 23263 20438
rect 25773 20498 25839 20501
rect 27705 20498 27771 20501
rect 25773 20496 27771 20498
rect 25773 20440 25778 20496
rect 25834 20440 27710 20496
rect 27766 20440 27771 20496
rect 25773 20438 27771 20440
rect 25773 20435 25839 20438
rect 27705 20435 27771 20438
rect 7465 20362 7531 20365
rect 15377 20362 15443 20365
rect 7465 20360 11530 20362
rect 7465 20304 7470 20360
rect 7526 20304 11530 20360
rect 7465 20302 11530 20304
rect 7465 20299 7531 20302
rect 749 20226 815 20229
rect 7557 20226 7623 20229
rect 749 20224 7623 20226
rect 749 20168 754 20224
rect 810 20168 7562 20224
rect 7618 20168 7623 20224
rect 749 20166 7623 20168
rect 11470 20226 11530 20302
rect 12574 20360 15443 20362
rect 12574 20304 15382 20360
rect 15438 20304 15443 20360
rect 12574 20302 15443 20304
rect 12574 20226 12634 20302
rect 15377 20299 15443 20302
rect 15561 20362 15627 20365
rect 21725 20362 21791 20365
rect 15561 20360 21791 20362
rect 15561 20304 15566 20360
rect 15622 20304 21730 20360
rect 21786 20304 21791 20360
rect 15561 20302 21791 20304
rect 15561 20299 15627 20302
rect 21725 20299 21791 20302
rect 24393 20362 24459 20365
rect 26417 20362 26483 20365
rect 24393 20360 26483 20362
rect 24393 20304 24398 20360
rect 24454 20304 26422 20360
rect 26478 20304 26483 20360
rect 24393 20302 26483 20304
rect 24393 20299 24459 20302
rect 26417 20299 26483 20302
rect 11470 20166 12634 20226
rect 12709 20226 12775 20229
rect 19977 20226 20043 20229
rect 12709 20224 20043 20226
rect 12709 20168 12714 20224
rect 12770 20168 19982 20224
rect 20038 20168 20043 20224
rect 12709 20166 20043 20168
rect 749 20163 815 20166
rect 7557 20163 7623 20166
rect 12709 20163 12775 20166
rect 19977 20163 20043 20166
rect 24945 20226 25011 20229
rect 27846 20226 27906 20574
rect 29520 20544 30000 20574
rect 24945 20224 27906 20226
rect 24945 20168 24950 20224
rect 25006 20168 27906 20224
rect 24945 20166 27906 20168
rect 24945 20163 25011 20166
rect 10944 20160 11264 20161
rect 0 20090 480 20120
rect 10944 20096 10952 20160
rect 11016 20096 11032 20160
rect 11096 20096 11112 20160
rect 11176 20096 11192 20160
rect 11256 20096 11264 20160
rect 10944 20095 11264 20096
rect 20944 20160 21264 20161
rect 20944 20096 20952 20160
rect 21016 20096 21032 20160
rect 21096 20096 21112 20160
rect 21176 20096 21192 20160
rect 21256 20096 21264 20160
rect 20944 20095 21264 20096
rect 3601 20090 3667 20093
rect 0 20088 3667 20090
rect 0 20032 3606 20088
rect 3662 20032 3667 20088
rect 0 20030 3667 20032
rect 0 20000 480 20030
rect 3601 20027 3667 20030
rect 14181 20090 14247 20093
rect 20805 20090 20871 20093
rect 14181 20088 20871 20090
rect 14181 20032 14186 20088
rect 14242 20032 20810 20088
rect 20866 20032 20871 20088
rect 14181 20030 20871 20032
rect 14181 20027 14247 20030
rect 20805 20027 20871 20030
rect 26693 20090 26759 20093
rect 29177 20090 29243 20093
rect 29520 20090 30000 20120
rect 26693 20088 29243 20090
rect 26693 20032 26698 20088
rect 26754 20032 29182 20088
rect 29238 20032 29243 20088
rect 26693 20030 29243 20032
rect 26693 20027 26759 20030
rect 29177 20027 29243 20030
rect 29318 20030 30000 20090
rect 3693 19954 3759 19957
rect 16573 19954 16639 19957
rect 3693 19952 16639 19954
rect 3693 19896 3698 19952
rect 3754 19896 16578 19952
rect 16634 19896 16639 19952
rect 3693 19894 16639 19896
rect 3693 19891 3759 19894
rect 16573 19891 16639 19894
rect 25405 19954 25471 19957
rect 29318 19954 29378 20030
rect 29520 20000 30000 20030
rect 25405 19952 29378 19954
rect 25405 19896 25410 19952
rect 25466 19896 29378 19952
rect 25405 19894 29378 19896
rect 25405 19891 25471 19894
rect 2221 19818 2287 19821
rect 15469 19818 15535 19821
rect 2221 19816 15535 19818
rect 2221 19760 2226 19816
rect 2282 19760 15474 19816
rect 15530 19760 15535 19816
rect 2221 19758 15535 19760
rect 2221 19755 2287 19758
rect 15469 19755 15535 19758
rect 16297 19818 16363 19821
rect 26877 19818 26943 19821
rect 16297 19816 26943 19818
rect 16297 19760 16302 19816
rect 16358 19760 26882 19816
rect 26938 19760 26943 19816
rect 16297 19758 26943 19760
rect 16297 19755 16363 19758
rect 26877 19755 26943 19758
rect 7557 19682 7623 19685
rect 14273 19682 14339 19685
rect 7557 19680 14339 19682
rect 7557 19624 7562 19680
rect 7618 19624 14278 19680
rect 14334 19624 14339 19680
rect 7557 19622 14339 19624
rect 7557 19619 7623 19622
rect 14273 19619 14339 19622
rect 16573 19682 16639 19685
rect 19517 19682 19583 19685
rect 25589 19682 25655 19685
rect 16573 19680 25655 19682
rect 16573 19624 16578 19680
rect 16634 19624 19522 19680
rect 19578 19624 25594 19680
rect 25650 19624 25655 19680
rect 16573 19622 25655 19624
rect 16573 19619 16639 19622
rect 19517 19619 19583 19622
rect 25589 19619 25655 19622
rect 5944 19616 6264 19617
rect 5944 19552 5952 19616
rect 6016 19552 6032 19616
rect 6096 19552 6112 19616
rect 6176 19552 6192 19616
rect 6256 19552 6264 19616
rect 5944 19551 6264 19552
rect 15944 19616 16264 19617
rect 15944 19552 15952 19616
rect 16016 19552 16032 19616
rect 16096 19552 16112 19616
rect 16176 19552 16192 19616
rect 16256 19552 16264 19616
rect 15944 19551 16264 19552
rect 25944 19616 26264 19617
rect 25944 19552 25952 19616
rect 26016 19552 26032 19616
rect 26096 19552 26112 19616
rect 26176 19552 26192 19616
rect 26256 19552 26264 19616
rect 25944 19551 26264 19552
rect 18045 19546 18111 19549
rect 24209 19546 24275 19549
rect 16438 19544 24275 19546
rect 16438 19488 18050 19544
rect 18106 19488 24214 19544
rect 24270 19488 24275 19544
rect 16438 19486 24275 19488
rect 0 19410 480 19440
rect 3325 19410 3391 19413
rect 0 19408 3391 19410
rect 0 19352 3330 19408
rect 3386 19352 3391 19408
rect 0 19350 3391 19352
rect 0 19320 480 19350
rect 3325 19347 3391 19350
rect 5349 19410 5415 19413
rect 16438 19410 16498 19486
rect 18045 19483 18111 19486
rect 24209 19483 24275 19486
rect 5349 19408 16498 19410
rect 5349 19352 5354 19408
rect 5410 19352 16498 19408
rect 5349 19350 16498 19352
rect 25221 19410 25287 19413
rect 29520 19410 30000 19440
rect 25221 19408 30000 19410
rect 25221 19352 25226 19408
rect 25282 19352 30000 19408
rect 25221 19350 30000 19352
rect 5349 19347 5415 19350
rect 25221 19347 25287 19350
rect 29520 19320 30000 19350
rect 10944 19072 11264 19073
rect 10944 19008 10952 19072
rect 11016 19008 11032 19072
rect 11096 19008 11112 19072
rect 11176 19008 11192 19072
rect 11256 19008 11264 19072
rect 10944 19007 11264 19008
rect 20944 19072 21264 19073
rect 20944 19008 20952 19072
rect 21016 19008 21032 19072
rect 21096 19008 21112 19072
rect 21176 19008 21192 19072
rect 21256 19008 21264 19072
rect 20944 19007 21264 19008
rect 0 18866 480 18896
rect 3693 18866 3759 18869
rect 0 18864 3759 18866
rect 0 18808 3698 18864
rect 3754 18808 3759 18864
rect 0 18806 3759 18808
rect 0 18776 480 18806
rect 3693 18803 3759 18806
rect 25129 18866 25195 18869
rect 29520 18866 30000 18896
rect 25129 18864 30000 18866
rect 25129 18808 25134 18864
rect 25190 18808 30000 18864
rect 25129 18806 30000 18808
rect 25129 18803 25195 18806
rect 29520 18776 30000 18806
rect 8569 18730 8635 18733
rect 20713 18730 20779 18733
rect 26509 18730 26575 18733
rect 8569 18728 26575 18730
rect 8569 18672 8574 18728
rect 8630 18672 20718 18728
rect 20774 18672 26514 18728
rect 26570 18672 26575 18728
rect 8569 18670 26575 18672
rect 8569 18667 8635 18670
rect 20713 18667 20779 18670
rect 26509 18667 26575 18670
rect 5944 18528 6264 18529
rect 5944 18464 5952 18528
rect 6016 18464 6032 18528
rect 6096 18464 6112 18528
rect 6176 18464 6192 18528
rect 6256 18464 6264 18528
rect 5944 18463 6264 18464
rect 15944 18528 16264 18529
rect 15944 18464 15952 18528
rect 16016 18464 16032 18528
rect 16096 18464 16112 18528
rect 16176 18464 16192 18528
rect 16256 18464 16264 18528
rect 15944 18463 16264 18464
rect 25944 18528 26264 18529
rect 25944 18464 25952 18528
rect 26016 18464 26032 18528
rect 26096 18464 26112 18528
rect 26176 18464 26192 18528
rect 26256 18464 26264 18528
rect 25944 18463 26264 18464
rect 0 18322 480 18352
rect 5717 18322 5783 18325
rect 0 18320 5783 18322
rect 0 18264 5722 18320
rect 5778 18264 5783 18320
rect 0 18262 5783 18264
rect 0 18232 480 18262
rect 5717 18259 5783 18262
rect 25589 18322 25655 18325
rect 29520 18322 30000 18352
rect 25589 18320 30000 18322
rect 25589 18264 25594 18320
rect 25650 18264 30000 18320
rect 25589 18262 30000 18264
rect 25589 18259 25655 18262
rect 29520 18232 30000 18262
rect 10944 17984 11264 17985
rect 10944 17920 10952 17984
rect 11016 17920 11032 17984
rect 11096 17920 11112 17984
rect 11176 17920 11192 17984
rect 11256 17920 11264 17984
rect 10944 17919 11264 17920
rect 20944 17984 21264 17985
rect 20944 17920 20952 17984
rect 21016 17920 21032 17984
rect 21096 17920 21112 17984
rect 21176 17920 21192 17984
rect 21256 17920 21264 17984
rect 20944 17919 21264 17920
rect 0 17642 480 17672
rect 3785 17642 3851 17645
rect 29520 17642 30000 17672
rect 0 17640 3851 17642
rect 0 17584 3790 17640
rect 3846 17584 3851 17640
rect 0 17582 3851 17584
rect 0 17552 480 17582
rect 3785 17579 3851 17582
rect 29318 17582 30000 17642
rect 5944 17440 6264 17441
rect 5944 17376 5952 17440
rect 6016 17376 6032 17440
rect 6096 17376 6112 17440
rect 6176 17376 6192 17440
rect 6256 17376 6264 17440
rect 5944 17375 6264 17376
rect 15944 17440 16264 17441
rect 15944 17376 15952 17440
rect 16016 17376 16032 17440
rect 16096 17376 16112 17440
rect 16176 17376 16192 17440
rect 16256 17376 16264 17440
rect 15944 17375 16264 17376
rect 25944 17440 26264 17441
rect 25944 17376 25952 17440
rect 26016 17376 26032 17440
rect 26096 17376 26112 17440
rect 26176 17376 26192 17440
rect 26256 17376 26264 17440
rect 25944 17375 26264 17376
rect 29318 17234 29378 17582
rect 29520 17552 30000 17582
rect 25638 17174 29378 17234
rect 0 17098 480 17128
rect 3509 17098 3575 17101
rect 0 17096 3575 17098
rect 0 17040 3514 17096
rect 3570 17040 3575 17096
rect 0 17038 3575 17040
rect 0 17008 480 17038
rect 3509 17035 3575 17038
rect 11697 17098 11763 17101
rect 25638 17098 25698 17174
rect 11697 17096 25698 17098
rect 11697 17040 11702 17096
rect 11758 17040 25698 17096
rect 11697 17038 25698 17040
rect 25773 17098 25839 17101
rect 29520 17098 30000 17128
rect 25773 17096 30000 17098
rect 25773 17040 25778 17096
rect 25834 17040 30000 17096
rect 25773 17038 30000 17040
rect 11697 17035 11763 17038
rect 25773 17035 25839 17038
rect 29520 17008 30000 17038
rect 10944 16896 11264 16897
rect 10944 16832 10952 16896
rect 11016 16832 11032 16896
rect 11096 16832 11112 16896
rect 11176 16832 11192 16896
rect 11256 16832 11264 16896
rect 10944 16831 11264 16832
rect 20944 16896 21264 16897
rect 20944 16832 20952 16896
rect 21016 16832 21032 16896
rect 21096 16832 21112 16896
rect 21176 16832 21192 16896
rect 21256 16832 21264 16896
rect 20944 16831 21264 16832
rect 0 16418 480 16448
rect 3417 16418 3483 16421
rect 29520 16418 30000 16448
rect 0 16416 3483 16418
rect 0 16360 3422 16416
rect 3478 16360 3483 16416
rect 0 16358 3483 16360
rect 0 16328 480 16358
rect 3417 16355 3483 16358
rect 26374 16358 30000 16418
rect 5944 16352 6264 16353
rect 5944 16288 5952 16352
rect 6016 16288 6032 16352
rect 6096 16288 6112 16352
rect 6176 16288 6192 16352
rect 6256 16288 6264 16352
rect 5944 16287 6264 16288
rect 15944 16352 16264 16353
rect 15944 16288 15952 16352
rect 16016 16288 16032 16352
rect 16096 16288 16112 16352
rect 16176 16288 16192 16352
rect 16256 16288 16264 16352
rect 15944 16287 16264 16288
rect 25944 16352 26264 16353
rect 25944 16288 25952 16352
rect 26016 16288 26032 16352
rect 26096 16288 26112 16352
rect 26176 16288 26192 16352
rect 26256 16288 26264 16352
rect 25944 16287 26264 16288
rect 25865 16146 25931 16149
rect 26374 16146 26434 16358
rect 29520 16328 30000 16358
rect 25865 16144 26434 16146
rect 25865 16088 25870 16144
rect 25926 16088 26434 16144
rect 25865 16086 26434 16088
rect 25865 16083 25931 16086
rect 0 15874 480 15904
rect 9949 15874 10015 15877
rect 0 15872 10015 15874
rect 0 15816 9954 15872
rect 10010 15816 10015 15872
rect 0 15814 10015 15816
rect 0 15784 480 15814
rect 9949 15811 10015 15814
rect 25037 15874 25103 15877
rect 29520 15874 30000 15904
rect 25037 15872 30000 15874
rect 25037 15816 25042 15872
rect 25098 15816 30000 15872
rect 25037 15814 30000 15816
rect 25037 15811 25103 15814
rect 10944 15808 11264 15809
rect 10944 15744 10952 15808
rect 11016 15744 11032 15808
rect 11096 15744 11112 15808
rect 11176 15744 11192 15808
rect 11256 15744 11264 15808
rect 10944 15743 11264 15744
rect 20944 15808 21264 15809
rect 20944 15744 20952 15808
rect 21016 15744 21032 15808
rect 21096 15744 21112 15808
rect 21176 15744 21192 15808
rect 21256 15744 21264 15808
rect 29520 15784 30000 15814
rect 20944 15743 21264 15744
rect 25313 15466 25379 15469
rect 25313 15464 26434 15466
rect 25313 15408 25318 15464
rect 25374 15408 26434 15464
rect 25313 15406 26434 15408
rect 25313 15403 25379 15406
rect 0 15330 480 15360
rect 2773 15330 2839 15333
rect 0 15328 2839 15330
rect 0 15272 2778 15328
rect 2834 15272 2839 15328
rect 0 15270 2839 15272
rect 0 15240 480 15270
rect 2773 15267 2839 15270
rect 17493 15330 17559 15333
rect 25773 15330 25839 15333
rect 17493 15328 25839 15330
rect 17493 15272 17498 15328
rect 17554 15272 25778 15328
rect 25834 15272 25839 15328
rect 17493 15270 25839 15272
rect 26374 15330 26434 15406
rect 29520 15330 30000 15360
rect 26374 15270 30000 15330
rect 17493 15267 17559 15270
rect 25773 15267 25839 15270
rect 5944 15264 6264 15265
rect 5944 15200 5952 15264
rect 6016 15200 6032 15264
rect 6096 15200 6112 15264
rect 6176 15200 6192 15264
rect 6256 15200 6264 15264
rect 5944 15199 6264 15200
rect 15944 15264 16264 15265
rect 15944 15200 15952 15264
rect 16016 15200 16032 15264
rect 16096 15200 16112 15264
rect 16176 15200 16192 15264
rect 16256 15200 16264 15264
rect 15944 15199 16264 15200
rect 25944 15264 26264 15265
rect 25944 15200 25952 15264
rect 26016 15200 26032 15264
rect 26096 15200 26112 15264
rect 26176 15200 26192 15264
rect 26256 15200 26264 15264
rect 29520 15240 30000 15270
rect 25944 15199 26264 15200
rect 10944 14720 11264 14721
rect 0 14650 480 14680
rect 10944 14656 10952 14720
rect 11016 14656 11032 14720
rect 11096 14656 11112 14720
rect 11176 14656 11192 14720
rect 11256 14656 11264 14720
rect 10944 14655 11264 14656
rect 20944 14720 21264 14721
rect 20944 14656 20952 14720
rect 21016 14656 21032 14720
rect 21096 14656 21112 14720
rect 21176 14656 21192 14720
rect 21256 14656 21264 14720
rect 20944 14655 21264 14656
rect 2957 14650 3023 14653
rect 0 14648 3023 14650
rect 0 14592 2962 14648
rect 3018 14592 3023 14648
rect 0 14590 3023 14592
rect 0 14560 480 14590
rect 2957 14587 3023 14590
rect 24853 14650 24919 14653
rect 29520 14650 30000 14680
rect 24853 14648 30000 14650
rect 24853 14592 24858 14648
rect 24914 14592 30000 14648
rect 24853 14590 30000 14592
rect 24853 14587 24919 14590
rect 29520 14560 30000 14590
rect 16297 14514 16363 14517
rect 25405 14514 25471 14517
rect 16297 14512 25471 14514
rect 16297 14456 16302 14512
rect 16358 14456 25410 14512
rect 25466 14456 25471 14512
rect 16297 14454 25471 14456
rect 16297 14451 16363 14454
rect 25405 14451 25471 14454
rect 5944 14176 6264 14177
rect 0 14106 480 14136
rect 5944 14112 5952 14176
rect 6016 14112 6032 14176
rect 6096 14112 6112 14176
rect 6176 14112 6192 14176
rect 6256 14112 6264 14176
rect 5944 14111 6264 14112
rect 15944 14176 16264 14177
rect 15944 14112 15952 14176
rect 16016 14112 16032 14176
rect 16096 14112 16112 14176
rect 16176 14112 16192 14176
rect 16256 14112 16264 14176
rect 15944 14111 16264 14112
rect 25944 14176 26264 14177
rect 25944 14112 25952 14176
rect 26016 14112 26032 14176
rect 26096 14112 26112 14176
rect 26176 14112 26192 14176
rect 26256 14112 26264 14176
rect 25944 14111 26264 14112
rect 3877 14106 3943 14109
rect 29520 14106 30000 14136
rect 0 14104 3943 14106
rect 0 14048 3882 14104
rect 3938 14048 3943 14104
rect 0 14046 3943 14048
rect 0 14016 480 14046
rect 3877 14043 3943 14046
rect 26374 14046 30000 14106
rect 24945 13970 25011 13973
rect 26374 13970 26434 14046
rect 29520 14016 30000 14046
rect 24945 13968 26434 13970
rect 24945 13912 24950 13968
rect 25006 13912 26434 13968
rect 24945 13910 26434 13912
rect 24945 13907 25011 13910
rect 18321 13834 18387 13837
rect 25865 13834 25931 13837
rect 18321 13832 25931 13834
rect 18321 13776 18326 13832
rect 18382 13776 25870 13832
rect 25926 13776 25931 13832
rect 18321 13774 25931 13776
rect 18321 13771 18387 13774
rect 25865 13771 25931 13774
rect 10944 13632 11264 13633
rect 10944 13568 10952 13632
rect 11016 13568 11032 13632
rect 11096 13568 11112 13632
rect 11176 13568 11192 13632
rect 11256 13568 11264 13632
rect 10944 13567 11264 13568
rect 20944 13632 21264 13633
rect 20944 13568 20952 13632
rect 21016 13568 21032 13632
rect 21096 13568 21112 13632
rect 21176 13568 21192 13632
rect 21256 13568 21264 13632
rect 20944 13567 21264 13568
rect 0 13426 480 13456
rect 3049 13426 3115 13429
rect 0 13424 3115 13426
rect 0 13368 3054 13424
rect 3110 13368 3115 13424
rect 0 13366 3115 13368
rect 0 13336 480 13366
rect 3049 13363 3115 13366
rect 10133 13426 10199 13429
rect 24761 13426 24827 13429
rect 10133 13424 24827 13426
rect 10133 13368 10138 13424
rect 10194 13368 24766 13424
rect 24822 13368 24827 13424
rect 10133 13366 24827 13368
rect 10133 13363 10199 13366
rect 24761 13363 24827 13366
rect 25405 13426 25471 13429
rect 29520 13426 30000 13456
rect 25405 13424 30000 13426
rect 25405 13368 25410 13424
rect 25466 13368 30000 13424
rect 25405 13366 30000 13368
rect 25405 13363 25471 13366
rect 29520 13336 30000 13366
rect 9305 13290 9371 13293
rect 9305 13288 17234 13290
rect 9305 13232 9310 13288
rect 9366 13232 17234 13288
rect 9305 13230 17234 13232
rect 9305 13227 9371 13230
rect 5944 13088 6264 13089
rect 5944 13024 5952 13088
rect 6016 13024 6032 13088
rect 6096 13024 6112 13088
rect 6176 13024 6192 13088
rect 6256 13024 6264 13088
rect 5944 13023 6264 13024
rect 15944 13088 16264 13089
rect 15944 13024 15952 13088
rect 16016 13024 16032 13088
rect 16096 13024 16112 13088
rect 16176 13024 16192 13088
rect 16256 13024 16264 13088
rect 15944 13023 16264 13024
rect 8569 13018 8635 13021
rect 13813 13018 13879 13021
rect 3742 12958 5826 13018
rect 0 12882 480 12912
rect 1393 12882 1459 12885
rect 3742 12882 3802 12958
rect 0 12822 1226 12882
rect 0 12792 480 12822
rect 1166 12746 1226 12822
rect 1393 12880 3802 12882
rect 1393 12824 1398 12880
rect 1454 12824 3802 12880
rect 1393 12822 3802 12824
rect 3969 12882 4035 12885
rect 5766 12882 5826 12958
rect 8569 13016 13879 13018
rect 8569 12960 8574 13016
rect 8630 12960 13818 13016
rect 13874 12960 13879 13016
rect 8569 12958 13879 12960
rect 17174 13018 17234 13230
rect 25944 13088 26264 13089
rect 25944 13024 25952 13088
rect 26016 13024 26032 13088
rect 26096 13024 26112 13088
rect 26176 13024 26192 13088
rect 26256 13024 26264 13088
rect 25944 13023 26264 13024
rect 25221 13018 25287 13021
rect 17174 13016 25287 13018
rect 17174 12960 25226 13016
rect 25282 12960 25287 13016
rect 17174 12958 25287 12960
rect 8569 12955 8635 12958
rect 13813 12955 13879 12958
rect 25221 12955 25287 12958
rect 10041 12882 10107 12885
rect 3969 12880 4354 12882
rect 3969 12824 3974 12880
rect 4030 12824 4354 12880
rect 3969 12822 4354 12824
rect 5766 12880 10107 12882
rect 5766 12824 10046 12880
rect 10102 12824 10107 12880
rect 5766 12822 10107 12824
rect 1393 12819 1459 12822
rect 3969 12819 4035 12822
rect 4061 12746 4127 12749
rect 1166 12744 4127 12746
rect 1166 12688 4066 12744
rect 4122 12688 4127 12744
rect 1166 12686 4127 12688
rect 4294 12746 4354 12822
rect 10041 12819 10107 12822
rect 19241 12882 19307 12885
rect 29520 12882 30000 12912
rect 19241 12880 30000 12882
rect 19241 12824 19246 12880
rect 19302 12824 30000 12880
rect 19241 12822 30000 12824
rect 19241 12819 19307 12822
rect 29520 12792 30000 12822
rect 25129 12746 25195 12749
rect 4294 12744 25195 12746
rect 4294 12688 25134 12744
rect 25190 12688 25195 12744
rect 4294 12686 25195 12688
rect 4061 12683 4127 12686
rect 25129 12683 25195 12686
rect 10944 12544 11264 12545
rect 10944 12480 10952 12544
rect 11016 12480 11032 12544
rect 11096 12480 11112 12544
rect 11176 12480 11192 12544
rect 11256 12480 11264 12544
rect 10944 12479 11264 12480
rect 20944 12544 21264 12545
rect 20944 12480 20952 12544
rect 21016 12480 21032 12544
rect 21096 12480 21112 12544
rect 21176 12480 21192 12544
rect 21256 12480 21264 12544
rect 20944 12479 21264 12480
rect 3325 12472 3391 12477
rect 3325 12416 3330 12472
rect 3386 12416 3391 12472
rect 3325 12411 3391 12416
rect 3785 12474 3851 12477
rect 4061 12474 4127 12477
rect 20161 12474 20227 12477
rect 3785 12472 4127 12474
rect 3785 12416 3790 12472
rect 3846 12416 4066 12472
rect 4122 12416 4127 12472
rect 3785 12414 4127 12416
rect 3785 12411 3851 12414
rect 4061 12411 4127 12414
rect 20118 12472 20227 12474
rect 20118 12416 20166 12472
rect 20222 12416 20227 12472
rect 20118 12411 20227 12416
rect 0 12338 480 12368
rect 3328 12338 3388 12411
rect 9857 12338 9923 12341
rect 0 12278 2514 12338
rect 3328 12336 9923 12338
rect 3328 12280 9862 12336
rect 9918 12280 9923 12336
rect 3328 12278 9923 12280
rect 20118 12338 20178 12411
rect 20253 12338 20319 12341
rect 20118 12336 20319 12338
rect 20118 12280 20258 12336
rect 20314 12280 20319 12336
rect 20118 12278 20319 12280
rect 0 12248 480 12278
rect 0 11658 480 11688
rect 1577 11658 1643 11661
rect 0 11656 1643 11658
rect 0 11600 1582 11656
rect 1638 11600 1643 11656
rect 0 11598 1643 11600
rect 0 11568 480 11598
rect 1577 11595 1643 11598
rect 0 11114 480 11144
rect 1393 11114 1459 11117
rect 0 11112 1459 11114
rect 0 11056 1398 11112
rect 1454 11056 1459 11112
rect 0 11054 1459 11056
rect 2454 11114 2514 12278
rect 9857 12275 9923 12278
rect 20253 12275 20319 12278
rect 25865 12338 25931 12341
rect 29520 12338 30000 12368
rect 25865 12336 30000 12338
rect 25865 12280 25870 12336
rect 25926 12280 30000 12336
rect 25865 12278 30000 12280
rect 25865 12275 25931 12278
rect 29520 12248 30000 12278
rect 4337 12202 4403 12205
rect 10225 12202 10291 12205
rect 4337 12200 10291 12202
rect 4337 12144 4342 12200
rect 4398 12144 10230 12200
rect 10286 12144 10291 12200
rect 4337 12142 10291 12144
rect 4337 12139 4403 12142
rect 10225 12139 10291 12142
rect 12157 12202 12223 12205
rect 25037 12202 25103 12205
rect 12157 12200 25103 12202
rect 12157 12144 12162 12200
rect 12218 12144 25042 12200
rect 25098 12144 25103 12200
rect 12157 12142 25103 12144
rect 12157 12139 12223 12142
rect 25037 12139 25103 12142
rect 5944 12000 6264 12001
rect 5944 11936 5952 12000
rect 6016 11936 6032 12000
rect 6096 11936 6112 12000
rect 6176 11936 6192 12000
rect 6256 11936 6264 12000
rect 5944 11935 6264 11936
rect 15944 12000 16264 12001
rect 15944 11936 15952 12000
rect 16016 11936 16032 12000
rect 16096 11936 16112 12000
rect 16176 11936 16192 12000
rect 16256 11936 16264 12000
rect 15944 11935 16264 11936
rect 25944 12000 26264 12001
rect 25944 11936 25952 12000
rect 26016 11936 26032 12000
rect 26096 11936 26112 12000
rect 26176 11936 26192 12000
rect 26256 11936 26264 12000
rect 25944 11935 26264 11936
rect 2773 11794 2839 11797
rect 3233 11794 3299 11797
rect 9397 11794 9463 11797
rect 26417 11794 26483 11797
rect 2773 11792 5826 11794
rect 2773 11736 2778 11792
rect 2834 11736 3238 11792
rect 3294 11736 5826 11792
rect 2773 11734 5826 11736
rect 2773 11731 2839 11734
rect 3233 11731 3299 11734
rect 2681 11658 2747 11661
rect 5533 11658 5599 11661
rect 2681 11656 5599 11658
rect 2681 11600 2686 11656
rect 2742 11600 5538 11656
rect 5594 11600 5599 11656
rect 2681 11598 5599 11600
rect 5766 11658 5826 11734
rect 9397 11792 26483 11794
rect 9397 11736 9402 11792
rect 9458 11736 26422 11792
rect 26478 11736 26483 11792
rect 9397 11734 26483 11736
rect 9397 11731 9463 11734
rect 26417 11731 26483 11734
rect 25497 11658 25563 11661
rect 5766 11656 25563 11658
rect 5766 11600 25502 11656
rect 25558 11600 25563 11656
rect 5766 11598 25563 11600
rect 2681 11595 2747 11598
rect 5533 11595 5599 11598
rect 25497 11595 25563 11598
rect 26693 11658 26759 11661
rect 29520 11658 30000 11688
rect 26693 11656 30000 11658
rect 26693 11600 26698 11656
rect 26754 11600 30000 11656
rect 26693 11598 30000 11600
rect 26693 11595 26759 11598
rect 29520 11568 30000 11598
rect 10944 11456 11264 11457
rect 10944 11392 10952 11456
rect 11016 11392 11032 11456
rect 11096 11392 11112 11456
rect 11176 11392 11192 11456
rect 11256 11392 11264 11456
rect 10944 11391 11264 11392
rect 20944 11456 21264 11457
rect 20944 11392 20952 11456
rect 21016 11392 21032 11456
rect 21096 11392 21112 11456
rect 21176 11392 21192 11456
rect 21256 11392 21264 11456
rect 20944 11391 21264 11392
rect 3141 11114 3207 11117
rect 2454 11112 3207 11114
rect 2454 11056 3146 11112
rect 3202 11056 3207 11112
rect 2454 11054 3207 11056
rect 0 11024 480 11054
rect 1393 11051 1459 11054
rect 3141 11051 3207 11054
rect 16205 11114 16271 11117
rect 25681 11114 25747 11117
rect 16205 11112 25747 11114
rect 16205 11056 16210 11112
rect 16266 11056 25686 11112
rect 25742 11056 25747 11112
rect 16205 11054 25747 11056
rect 16205 11051 16271 11054
rect 25681 11051 25747 11054
rect 26601 11114 26667 11117
rect 29520 11114 30000 11144
rect 26601 11112 30000 11114
rect 26601 11056 26606 11112
rect 26662 11056 30000 11112
rect 26601 11054 30000 11056
rect 26601 11051 26667 11054
rect 29520 11024 30000 11054
rect 17125 10978 17191 10981
rect 25313 10978 25379 10981
rect 17125 10976 25379 10978
rect 17125 10920 17130 10976
rect 17186 10920 25318 10976
rect 25374 10920 25379 10976
rect 17125 10918 25379 10920
rect 17125 10915 17191 10918
rect 25313 10915 25379 10918
rect 5944 10912 6264 10913
rect 5944 10848 5952 10912
rect 6016 10848 6032 10912
rect 6096 10848 6112 10912
rect 6176 10848 6192 10912
rect 6256 10848 6264 10912
rect 5944 10847 6264 10848
rect 15944 10912 16264 10913
rect 15944 10848 15952 10912
rect 16016 10848 16032 10912
rect 16096 10848 16112 10912
rect 16176 10848 16192 10912
rect 16256 10848 16264 10912
rect 15944 10847 16264 10848
rect 25944 10912 26264 10913
rect 25944 10848 25952 10912
rect 26016 10848 26032 10912
rect 26096 10848 26112 10912
rect 26176 10848 26192 10912
rect 26256 10848 26264 10912
rect 25944 10847 26264 10848
rect 17309 10842 17375 10845
rect 18689 10842 18755 10845
rect 17309 10840 18755 10842
rect 17309 10784 17314 10840
rect 17370 10784 18694 10840
rect 18750 10784 18755 10840
rect 17309 10782 18755 10784
rect 17309 10779 17375 10782
rect 18689 10779 18755 10782
rect 9489 10706 9555 10709
rect 12341 10706 12407 10709
rect 9489 10704 12407 10706
rect 9489 10648 9494 10704
rect 9550 10648 12346 10704
rect 12402 10648 12407 10704
rect 9489 10646 12407 10648
rect 9489 10643 9555 10646
rect 12341 10643 12407 10646
rect 15653 10706 15719 10709
rect 26509 10706 26575 10709
rect 15653 10704 26575 10706
rect 15653 10648 15658 10704
rect 15714 10648 26514 10704
rect 26570 10648 26575 10704
rect 15653 10646 26575 10648
rect 15653 10643 15719 10646
rect 26509 10643 26575 10646
rect 9581 10570 9647 10573
rect 26417 10570 26483 10573
rect 9581 10568 26483 10570
rect 9581 10512 9586 10568
rect 9642 10512 26422 10568
rect 26478 10512 26483 10568
rect 9581 10510 26483 10512
rect 9581 10507 9647 10510
rect 26417 10507 26483 10510
rect 0 10434 480 10464
rect 1577 10434 1643 10437
rect 0 10432 1643 10434
rect 0 10376 1582 10432
rect 1638 10376 1643 10432
rect 0 10374 1643 10376
rect 0 10344 480 10374
rect 1577 10371 1643 10374
rect 3141 10434 3207 10437
rect 6453 10434 6519 10437
rect 10501 10434 10567 10437
rect 3141 10432 10567 10434
rect 3141 10376 3146 10432
rect 3202 10376 6458 10432
rect 6514 10376 10506 10432
rect 10562 10376 10567 10432
rect 3141 10374 10567 10376
rect 3141 10371 3207 10374
rect 6453 10371 6519 10374
rect 10501 10371 10567 10374
rect 26601 10434 26667 10437
rect 29520 10434 30000 10464
rect 26601 10432 30000 10434
rect 26601 10376 26606 10432
rect 26662 10376 30000 10432
rect 26601 10374 30000 10376
rect 26601 10371 26667 10374
rect 10944 10368 11264 10369
rect 10944 10304 10952 10368
rect 11016 10304 11032 10368
rect 11096 10304 11112 10368
rect 11176 10304 11192 10368
rect 11256 10304 11264 10368
rect 10944 10303 11264 10304
rect 20944 10368 21264 10369
rect 20944 10304 20952 10368
rect 21016 10304 21032 10368
rect 21096 10304 21112 10368
rect 21176 10304 21192 10368
rect 21256 10304 21264 10368
rect 29520 10344 30000 10374
rect 20944 10303 21264 10304
rect 3417 10298 3483 10301
rect 12157 10298 12223 10301
rect 17125 10298 17191 10301
rect 3417 10296 6930 10298
rect 3417 10240 3422 10296
rect 3478 10240 6930 10296
rect 3417 10238 6930 10240
rect 3417 10235 3483 10238
rect 4521 10162 4587 10165
rect 6870 10162 6930 10238
rect 12157 10296 17191 10298
rect 12157 10240 12162 10296
rect 12218 10240 17130 10296
rect 17186 10240 17191 10296
rect 12157 10238 17191 10240
rect 12157 10235 12223 10238
rect 17125 10235 17191 10238
rect 17401 10162 17467 10165
rect 18321 10162 18387 10165
rect 26785 10162 26851 10165
rect 4521 10160 6746 10162
rect 4521 10104 4526 10160
rect 4582 10104 6746 10160
rect 4521 10102 6746 10104
rect 6870 10160 26851 10162
rect 6870 10104 17406 10160
rect 17462 10104 18326 10160
rect 18382 10104 26790 10160
rect 26846 10104 26851 10160
rect 6870 10102 26851 10104
rect 4521 10099 4587 10102
rect 2037 10026 2103 10029
rect 2865 10026 2931 10029
rect 2037 10024 2931 10026
rect 2037 9968 2042 10024
rect 2098 9968 2870 10024
rect 2926 9968 2931 10024
rect 2037 9966 2931 9968
rect 6686 10026 6746 10102
rect 17401 10099 17467 10102
rect 18321 10099 18387 10102
rect 26785 10099 26851 10102
rect 13261 10026 13327 10029
rect 16573 10026 16639 10029
rect 6686 10024 16639 10026
rect 6686 9968 13266 10024
rect 13322 9968 16578 10024
rect 16634 9968 16639 10024
rect 6686 9966 16639 9968
rect 2037 9963 2103 9966
rect 2865 9963 2931 9966
rect 13261 9963 13327 9966
rect 16573 9963 16639 9966
rect 18965 10026 19031 10029
rect 24945 10026 25011 10029
rect 18965 10024 25011 10026
rect 18965 9968 18970 10024
rect 19026 9968 24950 10024
rect 25006 9968 25011 10024
rect 18965 9966 25011 9968
rect 18965 9963 19031 9966
rect 24945 9963 25011 9966
rect 0 9890 480 9920
rect 1485 9890 1551 9893
rect 0 9888 1551 9890
rect 0 9832 1490 9888
rect 1546 9832 1551 9888
rect 0 9830 1551 9832
rect 0 9800 480 9830
rect 1485 9827 1551 9830
rect 3601 9890 3667 9893
rect 5533 9890 5599 9893
rect 3601 9888 5599 9890
rect 3601 9832 3606 9888
rect 3662 9832 5538 9888
rect 5594 9832 5599 9888
rect 3601 9830 5599 9832
rect 3601 9827 3667 9830
rect 5533 9827 5599 9830
rect 9581 9890 9647 9893
rect 12249 9890 12315 9893
rect 9581 9888 12315 9890
rect 9581 9832 9586 9888
rect 9642 9832 12254 9888
rect 12310 9832 12315 9888
rect 9581 9830 12315 9832
rect 9581 9827 9647 9830
rect 12249 9827 12315 9830
rect 26693 9890 26759 9893
rect 29520 9890 30000 9920
rect 26693 9888 30000 9890
rect 26693 9832 26698 9888
rect 26754 9832 30000 9888
rect 26693 9830 30000 9832
rect 26693 9827 26759 9830
rect 5944 9824 6264 9825
rect 5944 9760 5952 9824
rect 6016 9760 6032 9824
rect 6096 9760 6112 9824
rect 6176 9760 6192 9824
rect 6256 9760 6264 9824
rect 5944 9759 6264 9760
rect 15944 9824 16264 9825
rect 15944 9760 15952 9824
rect 16016 9760 16032 9824
rect 16096 9760 16112 9824
rect 16176 9760 16192 9824
rect 16256 9760 16264 9824
rect 15944 9759 16264 9760
rect 25944 9824 26264 9825
rect 25944 9760 25952 9824
rect 26016 9760 26032 9824
rect 26096 9760 26112 9824
rect 26176 9760 26192 9824
rect 26256 9760 26264 9824
rect 29520 9800 30000 9830
rect 25944 9759 26264 9760
rect 1669 9754 1735 9757
rect 3693 9754 3759 9757
rect 1669 9752 3759 9754
rect 1669 9696 1674 9752
rect 1730 9696 3698 9752
rect 3754 9696 3759 9752
rect 1669 9694 3759 9696
rect 1669 9691 1735 9694
rect 3693 9691 3759 9694
rect 3877 9754 3943 9757
rect 12157 9754 12223 9757
rect 3877 9752 5826 9754
rect 3877 9696 3882 9752
rect 3938 9696 5826 9752
rect 3877 9694 5826 9696
rect 3877 9691 3943 9694
rect 2589 9618 2655 9621
rect 5766 9618 5826 9694
rect 6502 9752 12223 9754
rect 6502 9696 12162 9752
rect 12218 9696 12223 9752
rect 6502 9694 12223 9696
rect 6502 9618 6562 9694
rect 12157 9691 12223 9694
rect 2589 9616 3434 9618
rect 2589 9560 2594 9616
rect 2650 9560 3434 9616
rect 2589 9558 3434 9560
rect 5766 9558 6562 9618
rect 7741 9618 7807 9621
rect 10869 9618 10935 9621
rect 7741 9616 10935 9618
rect 7741 9560 7746 9616
rect 7802 9560 10874 9616
rect 10930 9560 10935 9616
rect 7741 9558 10935 9560
rect 2589 9555 2655 9558
rect 0 9346 480 9376
rect 1393 9346 1459 9349
rect 0 9344 1459 9346
rect 0 9288 1398 9344
rect 1454 9288 1459 9344
rect 0 9286 1459 9288
rect 3374 9346 3434 9558
rect 7741 9555 7807 9558
rect 10869 9555 10935 9558
rect 3509 9482 3575 9485
rect 17769 9482 17835 9485
rect 27521 9482 27587 9485
rect 3509 9480 27587 9482
rect 3509 9424 3514 9480
rect 3570 9424 17774 9480
rect 17830 9424 27526 9480
rect 27582 9424 27587 9480
rect 3509 9422 27587 9424
rect 3509 9419 3575 9422
rect 17769 9419 17835 9422
rect 27521 9419 27587 9422
rect 10041 9346 10107 9349
rect 3374 9344 10107 9346
rect 3374 9288 10046 9344
rect 10102 9288 10107 9344
rect 3374 9286 10107 9288
rect 0 9256 480 9286
rect 1393 9283 1459 9286
rect 10041 9283 10107 9286
rect 11329 9346 11395 9349
rect 19977 9346 20043 9349
rect 11329 9344 20043 9346
rect 11329 9288 11334 9344
rect 11390 9288 19982 9344
rect 20038 9288 20043 9344
rect 11329 9286 20043 9288
rect 11329 9283 11395 9286
rect 19977 9283 20043 9286
rect 26601 9346 26667 9349
rect 29520 9346 30000 9376
rect 26601 9344 30000 9346
rect 26601 9288 26606 9344
rect 26662 9288 30000 9344
rect 26601 9286 30000 9288
rect 26601 9283 26667 9286
rect 10944 9280 11264 9281
rect 10944 9216 10952 9280
rect 11016 9216 11032 9280
rect 11096 9216 11112 9280
rect 11176 9216 11192 9280
rect 11256 9216 11264 9280
rect 10944 9215 11264 9216
rect 20944 9280 21264 9281
rect 20944 9216 20952 9280
rect 21016 9216 21032 9280
rect 21096 9216 21112 9280
rect 21176 9216 21192 9280
rect 21256 9216 21264 9280
rect 29520 9256 30000 9286
rect 20944 9215 21264 9216
rect 14917 9210 14983 9213
rect 16665 9210 16731 9213
rect 14917 9208 16731 9210
rect 14917 9152 14922 9208
rect 14978 9152 16670 9208
rect 16726 9152 16731 9208
rect 14917 9150 16731 9152
rect 14917 9147 14983 9150
rect 16665 9147 16731 9150
rect 7557 9074 7623 9077
rect 25589 9074 25655 9077
rect 7557 9072 25655 9074
rect 7557 9016 7562 9072
rect 7618 9016 25594 9072
rect 25650 9016 25655 9072
rect 7557 9014 25655 9016
rect 7557 9011 7623 9014
rect 25589 9011 25655 9014
rect 2037 8938 2103 8941
rect 11513 8938 11579 8941
rect 26509 8940 26575 8941
rect 26509 8938 26556 8940
rect 2037 8936 11579 8938
rect 2037 8880 2042 8936
rect 2098 8880 11518 8936
rect 11574 8880 11579 8936
rect 2037 8878 11579 8880
rect 26464 8936 26556 8938
rect 26464 8880 26514 8936
rect 26464 8878 26556 8880
rect 2037 8875 2103 8878
rect 11513 8875 11579 8878
rect 26509 8876 26556 8878
rect 26620 8876 26626 8940
rect 26509 8875 26575 8876
rect 5944 8736 6264 8737
rect 0 8666 480 8696
rect 5944 8672 5952 8736
rect 6016 8672 6032 8736
rect 6096 8672 6112 8736
rect 6176 8672 6192 8736
rect 6256 8672 6264 8736
rect 5944 8671 6264 8672
rect 15944 8736 16264 8737
rect 15944 8672 15952 8736
rect 16016 8672 16032 8736
rect 16096 8672 16112 8736
rect 16176 8672 16192 8736
rect 16256 8672 16264 8736
rect 15944 8671 16264 8672
rect 25944 8736 26264 8737
rect 25944 8672 25952 8736
rect 26016 8672 26032 8736
rect 26096 8672 26112 8736
rect 26176 8672 26192 8736
rect 26256 8672 26264 8736
rect 25944 8671 26264 8672
rect 1577 8666 1643 8669
rect 15469 8666 15535 8669
rect 0 8664 1643 8666
rect 0 8608 1582 8664
rect 1638 8608 1643 8664
rect 0 8606 1643 8608
rect 0 8576 480 8606
rect 1577 8603 1643 8606
rect 6502 8664 15535 8666
rect 6502 8608 15474 8664
rect 15530 8608 15535 8664
rect 6502 8606 15535 8608
rect 3141 8530 3207 8533
rect 6502 8530 6562 8606
rect 15469 8603 15535 8606
rect 16757 8666 16823 8669
rect 25773 8666 25839 8669
rect 16757 8664 25839 8666
rect 16757 8608 16762 8664
rect 16818 8608 25778 8664
rect 25834 8608 25839 8664
rect 16757 8606 25839 8608
rect 16757 8603 16823 8606
rect 25773 8603 25839 8606
rect 26693 8666 26759 8669
rect 29520 8666 30000 8696
rect 26693 8664 30000 8666
rect 26693 8608 26698 8664
rect 26754 8608 30000 8664
rect 26693 8606 30000 8608
rect 26693 8603 26759 8606
rect 29520 8576 30000 8606
rect 7189 8532 7255 8533
rect 7189 8530 7236 8532
rect 3141 8528 6562 8530
rect 3141 8472 3146 8528
rect 3202 8472 6562 8528
rect 3141 8470 6562 8472
rect 7144 8528 7236 8530
rect 7144 8472 7194 8528
rect 7144 8470 7236 8472
rect 3141 8467 3207 8470
rect 7189 8468 7236 8470
rect 7300 8468 7306 8532
rect 10777 8530 10843 8533
rect 26417 8530 26483 8533
rect 10777 8528 26483 8530
rect 10777 8472 10782 8528
rect 10838 8472 26422 8528
rect 26478 8472 26483 8528
rect 10777 8470 26483 8472
rect 7189 8467 7255 8468
rect 10777 8467 10843 8470
rect 26417 8467 26483 8470
rect 2405 8394 2471 8397
rect 7649 8394 7715 8397
rect 2405 8392 7715 8394
rect 2405 8336 2410 8392
rect 2466 8336 7654 8392
rect 7710 8336 7715 8392
rect 2405 8334 7715 8336
rect 2405 8331 2471 8334
rect 7649 8331 7715 8334
rect 19977 8394 20043 8397
rect 25405 8394 25471 8397
rect 19977 8392 25471 8394
rect 19977 8336 19982 8392
rect 20038 8336 25410 8392
rect 25466 8336 25471 8392
rect 19977 8334 25471 8336
rect 19977 8331 20043 8334
rect 25405 8331 25471 8334
rect 27705 8394 27771 8397
rect 27705 8392 28642 8394
rect 27705 8336 27710 8392
rect 27766 8336 28642 8392
rect 27705 8334 28642 8336
rect 27705 8331 27771 8334
rect 2037 8258 2103 8261
rect 9029 8258 9095 8261
rect 20805 8258 20871 8261
rect 2037 8256 9095 8258
rect 2037 8200 2042 8256
rect 2098 8200 9034 8256
rect 9090 8200 9095 8256
rect 2037 8198 9095 8200
rect 2037 8195 2103 8198
rect 9029 8195 9095 8198
rect 11470 8256 20871 8258
rect 11470 8200 20810 8256
rect 20866 8200 20871 8256
rect 11470 8198 20871 8200
rect 10944 8192 11264 8193
rect 0 8122 480 8152
rect 10944 8128 10952 8192
rect 11016 8128 11032 8192
rect 11096 8128 11112 8192
rect 11176 8128 11192 8192
rect 11256 8128 11264 8192
rect 10944 8127 11264 8128
rect 2681 8122 2747 8125
rect 0 8120 2747 8122
rect 0 8064 2686 8120
rect 2742 8064 2747 8120
rect 0 8062 2747 8064
rect 0 8032 480 8062
rect 2681 8059 2747 8062
rect 3785 8122 3851 8125
rect 6361 8122 6427 8125
rect 3785 8120 6427 8122
rect 3785 8064 3790 8120
rect 3846 8064 6366 8120
rect 6422 8064 6427 8120
rect 3785 8062 6427 8064
rect 3785 8059 3851 8062
rect 6361 8059 6427 8062
rect 6269 7986 6335 7989
rect 11470 7986 11530 8198
rect 20805 8195 20871 8198
rect 21357 8258 21423 8261
rect 21909 8258 21975 8261
rect 24853 8258 24919 8261
rect 21357 8256 24919 8258
rect 21357 8200 21362 8256
rect 21418 8200 21914 8256
rect 21970 8200 24858 8256
rect 24914 8200 24919 8256
rect 21357 8198 24919 8200
rect 21357 8195 21423 8198
rect 21909 8195 21975 8198
rect 24853 8195 24919 8198
rect 20944 8192 21264 8193
rect 20944 8128 20952 8192
rect 21016 8128 21032 8192
rect 21096 8128 21112 8192
rect 21176 8128 21192 8192
rect 21256 8128 21264 8192
rect 20944 8127 21264 8128
rect 12249 8122 12315 8125
rect 14733 8122 14799 8125
rect 12249 8120 14799 8122
rect 12249 8064 12254 8120
rect 12310 8064 14738 8120
rect 14794 8064 14799 8120
rect 12249 8062 14799 8064
rect 28582 8122 28642 8334
rect 29520 8122 30000 8152
rect 28582 8062 30000 8122
rect 12249 8059 12315 8062
rect 14733 8059 14799 8062
rect 29520 8032 30000 8062
rect 6269 7984 11530 7986
rect 6269 7928 6274 7984
rect 6330 7928 11530 7984
rect 6269 7926 11530 7928
rect 11605 7986 11671 7989
rect 11789 7986 11855 7989
rect 19885 7986 19951 7989
rect 25865 7986 25931 7989
rect 11605 7984 25931 7986
rect 11605 7928 11610 7984
rect 11666 7928 11794 7984
rect 11850 7928 19890 7984
rect 19946 7928 25870 7984
rect 25926 7928 25931 7984
rect 11605 7926 25931 7928
rect 6269 7923 6335 7926
rect 11605 7923 11671 7926
rect 11789 7923 11855 7926
rect 19885 7923 19951 7926
rect 25865 7923 25931 7926
rect 3417 7850 3483 7853
rect 16941 7850 17007 7853
rect 3417 7848 17007 7850
rect 3417 7792 3422 7848
rect 3478 7792 16946 7848
rect 17002 7792 17007 7848
rect 3417 7790 17007 7792
rect 3417 7787 3483 7790
rect 16941 7787 17007 7790
rect 6361 7714 6427 7717
rect 11237 7714 11303 7717
rect 6361 7712 11303 7714
rect 6361 7656 6366 7712
rect 6422 7656 11242 7712
rect 11298 7656 11303 7712
rect 6361 7654 11303 7656
rect 6361 7651 6427 7654
rect 11237 7651 11303 7654
rect 5944 7648 6264 7649
rect 5944 7584 5952 7648
rect 6016 7584 6032 7648
rect 6096 7584 6112 7648
rect 6176 7584 6192 7648
rect 6256 7584 6264 7648
rect 5944 7583 6264 7584
rect 15944 7648 16264 7649
rect 15944 7584 15952 7648
rect 16016 7584 16032 7648
rect 16096 7584 16112 7648
rect 16176 7584 16192 7648
rect 16256 7584 16264 7648
rect 15944 7583 16264 7584
rect 25944 7648 26264 7649
rect 25944 7584 25952 7648
rect 26016 7584 26032 7648
rect 26096 7584 26112 7648
rect 26176 7584 26192 7648
rect 26256 7584 26264 7648
rect 25944 7583 26264 7584
rect 13353 7578 13419 7581
rect 6502 7576 13419 7578
rect 6502 7520 13358 7576
rect 13414 7520 13419 7576
rect 6502 7518 13419 7520
rect 0 7442 480 7472
rect 1577 7442 1643 7445
rect 0 7440 1643 7442
rect 0 7384 1582 7440
rect 1638 7384 1643 7440
rect 0 7382 1643 7384
rect 0 7352 480 7382
rect 1577 7379 1643 7382
rect 4981 7442 5047 7445
rect 6502 7442 6562 7518
rect 13353 7515 13419 7518
rect 4981 7440 6562 7442
rect 4981 7384 4986 7440
rect 5042 7384 6562 7440
rect 4981 7382 6562 7384
rect 9213 7442 9279 7445
rect 11053 7442 11119 7445
rect 9213 7440 11119 7442
rect 9213 7384 9218 7440
rect 9274 7384 11058 7440
rect 11114 7384 11119 7440
rect 9213 7382 11119 7384
rect 4981 7379 5047 7382
rect 9213 7379 9279 7382
rect 11053 7379 11119 7382
rect 11237 7442 11303 7445
rect 26417 7442 26483 7445
rect 11237 7440 26483 7442
rect 11237 7384 11242 7440
rect 11298 7384 26422 7440
rect 26478 7384 26483 7440
rect 11237 7382 26483 7384
rect 11237 7379 11303 7382
rect 26417 7379 26483 7382
rect 26693 7442 26759 7445
rect 29520 7442 30000 7472
rect 26693 7440 30000 7442
rect 26693 7384 26698 7440
rect 26754 7384 30000 7440
rect 26693 7382 30000 7384
rect 26693 7379 26759 7382
rect 29520 7352 30000 7382
rect 2405 7306 2471 7309
rect 15469 7306 15535 7309
rect 2405 7304 15535 7306
rect 2405 7248 2410 7304
rect 2466 7248 15474 7304
rect 15530 7248 15535 7304
rect 2405 7246 15535 7248
rect 2405 7243 2471 7246
rect 15469 7243 15535 7246
rect 16941 7306 17007 7309
rect 26509 7306 26575 7309
rect 16941 7304 26575 7306
rect 16941 7248 16946 7304
rect 17002 7248 26514 7304
rect 26570 7248 26575 7304
rect 16941 7246 26575 7248
rect 16941 7243 17007 7246
rect 26509 7243 26575 7246
rect 10944 7104 11264 7105
rect 10944 7040 10952 7104
rect 11016 7040 11032 7104
rect 11096 7040 11112 7104
rect 11176 7040 11192 7104
rect 11256 7040 11264 7104
rect 10944 7039 11264 7040
rect 20944 7104 21264 7105
rect 20944 7040 20952 7104
rect 21016 7040 21032 7104
rect 21096 7040 21112 7104
rect 21176 7040 21192 7104
rect 21256 7040 21264 7104
rect 20944 7039 21264 7040
rect 6361 7034 6427 7037
rect 10777 7034 10843 7037
rect 6361 7032 10843 7034
rect 6361 6976 6366 7032
rect 6422 6976 10782 7032
rect 10838 6976 10843 7032
rect 6361 6974 10843 6976
rect 6361 6971 6427 6974
rect 10777 6971 10843 6974
rect 13353 7034 13419 7037
rect 19057 7034 19123 7037
rect 13353 7032 19123 7034
rect 13353 6976 13358 7032
rect 13414 6976 19062 7032
rect 19118 6976 19123 7032
rect 13353 6974 19123 6976
rect 13353 6971 13419 6974
rect 19057 6971 19123 6974
rect 26601 7034 26667 7037
rect 26601 7032 26802 7034
rect 26601 6976 26606 7032
rect 26662 6976 26802 7032
rect 26601 6974 26802 6976
rect 26601 6971 26667 6974
rect 0 6898 480 6928
rect 1577 6898 1643 6901
rect 0 6896 1643 6898
rect 0 6840 1582 6896
rect 1638 6840 1643 6896
rect 0 6838 1643 6840
rect 0 6808 480 6838
rect 1577 6835 1643 6838
rect 2037 6898 2103 6901
rect 6545 6898 6611 6901
rect 2037 6896 6611 6898
rect 2037 6840 2042 6896
rect 2098 6840 6550 6896
rect 6606 6840 6611 6896
rect 2037 6838 6611 6840
rect 2037 6835 2103 6838
rect 6545 6835 6611 6838
rect 9857 6898 9923 6901
rect 26509 6898 26575 6901
rect 9857 6896 26575 6898
rect 9857 6840 9862 6896
rect 9918 6840 26514 6896
rect 26570 6840 26575 6896
rect 9857 6838 26575 6840
rect 26742 6898 26802 6974
rect 29520 6898 30000 6928
rect 26742 6838 30000 6898
rect 9857 6835 9923 6838
rect 26509 6835 26575 6838
rect 29520 6808 30000 6838
rect 3049 6762 3115 6765
rect 19609 6762 19675 6765
rect 3049 6760 19675 6762
rect 3049 6704 3054 6760
rect 3110 6704 19614 6760
rect 19670 6704 19675 6760
rect 3049 6702 19675 6704
rect 3049 6699 3115 6702
rect 19609 6699 19675 6702
rect 27245 6762 27311 6765
rect 28349 6762 28415 6765
rect 27245 6760 28415 6762
rect 27245 6704 27250 6760
rect 27306 6704 28354 6760
rect 28410 6704 28415 6760
rect 27245 6702 28415 6704
rect 27245 6699 27311 6702
rect 28349 6699 28415 6702
rect 3325 6626 3391 6629
rect 5625 6626 5691 6629
rect 3325 6624 5691 6626
rect 3325 6568 3330 6624
rect 3386 6568 5630 6624
rect 5686 6568 5691 6624
rect 3325 6566 5691 6568
rect 3325 6563 3391 6566
rect 5625 6563 5691 6566
rect 5944 6560 6264 6561
rect 5944 6496 5952 6560
rect 6016 6496 6032 6560
rect 6096 6496 6112 6560
rect 6176 6496 6192 6560
rect 6256 6496 6264 6560
rect 5944 6495 6264 6496
rect 15944 6560 16264 6561
rect 15944 6496 15952 6560
rect 16016 6496 16032 6560
rect 16096 6496 16112 6560
rect 16176 6496 16192 6560
rect 16256 6496 16264 6560
rect 15944 6495 16264 6496
rect 25944 6560 26264 6561
rect 25944 6496 25952 6560
rect 26016 6496 26032 6560
rect 26096 6496 26112 6560
rect 26176 6496 26192 6560
rect 26256 6496 26264 6560
rect 25944 6495 26264 6496
rect 12341 6490 12407 6493
rect 6502 6488 12407 6490
rect 6502 6432 12346 6488
rect 12402 6432 12407 6488
rect 6502 6430 12407 6432
rect 0 6354 480 6384
rect 1577 6354 1643 6357
rect 0 6352 1643 6354
rect 0 6296 1582 6352
rect 1638 6296 1643 6352
rect 0 6294 1643 6296
rect 0 6264 480 6294
rect 1577 6291 1643 6294
rect 4613 6354 4679 6357
rect 6502 6354 6562 6430
rect 12341 6427 12407 6430
rect 4613 6352 6562 6354
rect 4613 6296 4618 6352
rect 4674 6296 6562 6352
rect 4613 6294 6562 6296
rect 6821 6354 6887 6357
rect 11421 6354 11487 6357
rect 6821 6352 11487 6354
rect 6821 6296 6826 6352
rect 6882 6296 11426 6352
rect 11482 6296 11487 6352
rect 6821 6294 11487 6296
rect 4613 6291 4679 6294
rect 6821 6291 6887 6294
rect 11421 6291 11487 6294
rect 11881 6354 11947 6357
rect 19793 6354 19859 6357
rect 26325 6354 26391 6357
rect 11881 6352 26391 6354
rect 11881 6296 11886 6352
rect 11942 6296 19798 6352
rect 19854 6296 26330 6352
rect 26386 6296 26391 6352
rect 11881 6294 26391 6296
rect 11881 6291 11947 6294
rect 19793 6291 19859 6294
rect 26325 6291 26391 6294
rect 26601 6354 26667 6357
rect 29520 6354 30000 6384
rect 26601 6352 30000 6354
rect 26601 6296 26606 6352
rect 26662 6296 30000 6352
rect 26601 6294 30000 6296
rect 26601 6291 26667 6294
rect 29520 6264 30000 6294
rect 11053 6218 11119 6221
rect 26509 6218 26575 6221
rect 11053 6216 26575 6218
rect 11053 6160 11058 6216
rect 11114 6160 26514 6216
rect 26570 6160 26575 6216
rect 11053 6158 26575 6160
rect 11053 6155 11119 6158
rect 26509 6155 26575 6158
rect 5073 6082 5139 6085
rect 7005 6082 7071 6085
rect 5073 6080 7071 6082
rect 5073 6024 5078 6080
rect 5134 6024 7010 6080
rect 7066 6024 7071 6080
rect 5073 6022 7071 6024
rect 5073 6019 5139 6022
rect 7005 6019 7071 6022
rect 11421 6082 11487 6085
rect 20805 6082 20871 6085
rect 11421 6080 20871 6082
rect 11421 6024 11426 6080
rect 11482 6024 20810 6080
rect 20866 6024 20871 6080
rect 11421 6022 20871 6024
rect 11421 6019 11487 6022
rect 20805 6019 20871 6022
rect 10944 6016 11264 6017
rect 10944 5952 10952 6016
rect 11016 5952 11032 6016
rect 11096 5952 11112 6016
rect 11176 5952 11192 6016
rect 11256 5952 11264 6016
rect 10944 5951 11264 5952
rect 20944 6016 21264 6017
rect 20944 5952 20952 6016
rect 21016 5952 21032 6016
rect 21096 5952 21112 6016
rect 21176 5952 21192 6016
rect 21256 5952 21264 6016
rect 20944 5951 21264 5952
rect 2405 5946 2471 5949
rect 10685 5946 10751 5949
rect 2405 5944 10751 5946
rect 2405 5888 2410 5944
rect 2466 5888 10690 5944
rect 10746 5888 10751 5944
rect 2405 5886 10751 5888
rect 2405 5883 2471 5886
rect 10685 5883 10751 5886
rect 12893 5946 12959 5949
rect 19149 5946 19215 5949
rect 12893 5944 19215 5946
rect 12893 5888 12898 5944
rect 12954 5888 19154 5944
rect 19210 5888 19215 5944
rect 12893 5886 19215 5888
rect 12893 5883 12959 5886
rect 19149 5883 19215 5886
rect 5809 5810 5875 5813
rect 26417 5810 26483 5813
rect 5809 5808 26483 5810
rect 5809 5752 5814 5808
rect 5870 5752 26422 5808
rect 26478 5752 26483 5808
rect 5809 5750 26483 5752
rect 5809 5747 5875 5750
rect 26417 5747 26483 5750
rect 0 5674 480 5704
rect 1577 5674 1643 5677
rect 0 5672 1643 5674
rect 0 5616 1582 5672
rect 1638 5616 1643 5672
rect 0 5614 1643 5616
rect 0 5584 480 5614
rect 1577 5611 1643 5614
rect 20805 5674 20871 5677
rect 25313 5674 25379 5677
rect 20805 5672 25379 5674
rect 20805 5616 20810 5672
rect 20866 5616 25318 5672
rect 25374 5616 25379 5672
rect 20805 5614 25379 5616
rect 20805 5611 20871 5614
rect 25313 5611 25379 5614
rect 26693 5674 26759 5677
rect 29520 5674 30000 5704
rect 26693 5672 30000 5674
rect 26693 5616 26698 5672
rect 26754 5616 30000 5672
rect 26693 5614 30000 5616
rect 26693 5611 26759 5614
rect 29520 5584 30000 5614
rect 5944 5472 6264 5473
rect 5944 5408 5952 5472
rect 6016 5408 6032 5472
rect 6096 5408 6112 5472
rect 6176 5408 6192 5472
rect 6256 5408 6264 5472
rect 5944 5407 6264 5408
rect 15944 5472 16264 5473
rect 15944 5408 15952 5472
rect 16016 5408 16032 5472
rect 16096 5408 16112 5472
rect 16176 5408 16192 5472
rect 16256 5408 16264 5472
rect 15944 5407 16264 5408
rect 25944 5472 26264 5473
rect 25944 5408 25952 5472
rect 26016 5408 26032 5472
rect 26096 5408 26112 5472
rect 26176 5408 26192 5472
rect 26256 5408 26264 5472
rect 25944 5407 26264 5408
rect 6637 5402 6703 5405
rect 9765 5402 9831 5405
rect 6637 5400 15762 5402
rect 6637 5344 6642 5400
rect 6698 5344 9770 5400
rect 9826 5344 15762 5400
rect 6637 5342 15762 5344
rect 6637 5339 6703 5342
rect 9765 5339 9831 5342
rect 3141 5266 3207 5269
rect 15469 5266 15535 5269
rect 3141 5264 15535 5266
rect 3141 5208 3146 5264
rect 3202 5208 15474 5264
rect 15530 5208 15535 5264
rect 3141 5206 15535 5208
rect 15702 5266 15762 5342
rect 19977 5266 20043 5269
rect 26877 5266 26943 5269
rect 15702 5264 26943 5266
rect 15702 5208 19982 5264
rect 20038 5208 26882 5264
rect 26938 5208 26943 5264
rect 15702 5206 26943 5208
rect 3141 5203 3207 5206
rect 15469 5203 15535 5206
rect 19977 5203 20043 5206
rect 26877 5203 26943 5206
rect 0 5130 480 5160
rect 2681 5130 2747 5133
rect 0 5128 2747 5130
rect 0 5072 2686 5128
rect 2742 5072 2747 5128
rect 0 5070 2747 5072
rect 0 5040 480 5070
rect 2681 5067 2747 5070
rect 4061 5130 4127 5133
rect 15377 5130 15443 5133
rect 4061 5128 15443 5130
rect 4061 5072 4066 5128
rect 4122 5072 15382 5128
rect 15438 5072 15443 5128
rect 4061 5070 15443 5072
rect 4061 5067 4127 5070
rect 15377 5067 15443 5070
rect 19609 5130 19675 5133
rect 26417 5130 26483 5133
rect 19609 5128 26483 5130
rect 19609 5072 19614 5128
rect 19670 5072 26422 5128
rect 26478 5072 26483 5128
rect 19609 5070 26483 5072
rect 19609 5067 19675 5070
rect 26417 5067 26483 5070
rect 26601 5130 26667 5133
rect 29520 5130 30000 5160
rect 26601 5128 30000 5130
rect 26601 5072 26606 5128
rect 26662 5072 30000 5128
rect 26601 5070 30000 5072
rect 26601 5067 26667 5070
rect 29520 5040 30000 5070
rect 10944 4928 11264 4929
rect 10944 4864 10952 4928
rect 11016 4864 11032 4928
rect 11096 4864 11112 4928
rect 11176 4864 11192 4928
rect 11256 4864 11264 4928
rect 10944 4863 11264 4864
rect 20944 4928 21264 4929
rect 20944 4864 20952 4928
rect 21016 4864 21032 4928
rect 21096 4864 21112 4928
rect 21176 4864 21192 4928
rect 21256 4864 21264 4928
rect 20944 4863 21264 4864
rect 2037 4858 2103 4861
rect 6361 4858 6427 4861
rect 2037 4856 6427 4858
rect 2037 4800 2042 4856
rect 2098 4800 6366 4856
rect 6422 4800 6427 4856
rect 2037 4798 6427 4800
rect 2037 4795 2103 4798
rect 6361 4795 6427 4798
rect 15929 4858 15995 4861
rect 18321 4858 18387 4861
rect 15929 4856 18387 4858
rect 15929 4800 15934 4856
rect 15990 4800 18326 4856
rect 18382 4800 18387 4856
rect 15929 4798 18387 4800
rect 15929 4795 15995 4798
rect 18321 4795 18387 4798
rect 0 4450 480 4480
rect 1577 4450 1643 4453
rect 0 4448 1643 4450
rect 0 4392 1582 4448
rect 1638 4392 1643 4448
rect 0 4390 1643 4392
rect 0 4360 480 4390
rect 1577 4387 1643 4390
rect 26693 4450 26759 4453
rect 29520 4450 30000 4480
rect 26693 4448 30000 4450
rect 26693 4392 26698 4448
rect 26754 4392 30000 4448
rect 26693 4390 30000 4392
rect 26693 4387 26759 4390
rect 5944 4384 6264 4385
rect 5944 4320 5952 4384
rect 6016 4320 6032 4384
rect 6096 4320 6112 4384
rect 6176 4320 6192 4384
rect 6256 4320 6264 4384
rect 5944 4319 6264 4320
rect 15944 4384 16264 4385
rect 15944 4320 15952 4384
rect 16016 4320 16032 4384
rect 16096 4320 16112 4384
rect 16176 4320 16192 4384
rect 16256 4320 16264 4384
rect 15944 4319 16264 4320
rect 25944 4384 26264 4385
rect 25944 4320 25952 4384
rect 26016 4320 26032 4384
rect 26096 4320 26112 4384
rect 26176 4320 26192 4384
rect 26256 4320 26264 4384
rect 29520 4360 30000 4390
rect 25944 4319 26264 4320
rect 2405 4178 2471 4181
rect 18597 4178 18663 4181
rect 2405 4176 18663 4178
rect 2405 4120 2410 4176
rect 2466 4120 18602 4176
rect 18658 4120 18663 4176
rect 2405 4118 18663 4120
rect 2405 4115 2471 4118
rect 18597 4115 18663 4118
rect 4613 4042 4679 4045
rect 9397 4042 9463 4045
rect 4613 4040 9463 4042
rect 4613 3984 4618 4040
rect 4674 3984 9402 4040
rect 9458 3984 9463 4040
rect 4613 3982 9463 3984
rect 4613 3979 4679 3982
rect 9397 3979 9463 3982
rect 10409 4042 10475 4045
rect 26417 4042 26483 4045
rect 10409 4040 26483 4042
rect 10409 3984 10414 4040
rect 10470 3984 26422 4040
rect 26478 3984 26483 4040
rect 10409 3982 26483 3984
rect 10409 3979 10475 3982
rect 26417 3979 26483 3982
rect 0 3906 480 3936
rect 1577 3906 1643 3909
rect 0 3904 1643 3906
rect 0 3848 1582 3904
rect 1638 3848 1643 3904
rect 0 3846 1643 3848
rect 0 3816 480 3846
rect 1577 3843 1643 3846
rect 3141 3906 3207 3909
rect 7189 3906 7255 3909
rect 3141 3904 7255 3906
rect 3141 3848 3146 3904
rect 3202 3848 7194 3904
rect 7250 3848 7255 3904
rect 3141 3846 7255 3848
rect 3141 3843 3207 3846
rect 7189 3843 7255 3846
rect 26601 3906 26667 3909
rect 29520 3906 30000 3936
rect 26601 3904 30000 3906
rect 26601 3848 26606 3904
rect 26662 3848 30000 3904
rect 26601 3846 30000 3848
rect 26601 3843 26667 3846
rect 10944 3840 11264 3841
rect 10944 3776 10952 3840
rect 11016 3776 11032 3840
rect 11096 3776 11112 3840
rect 11176 3776 11192 3840
rect 11256 3776 11264 3840
rect 10944 3775 11264 3776
rect 20944 3840 21264 3841
rect 20944 3776 20952 3840
rect 21016 3776 21032 3840
rect 21096 3776 21112 3840
rect 21176 3776 21192 3840
rect 21256 3776 21264 3840
rect 29520 3816 30000 3846
rect 20944 3775 21264 3776
rect 8109 3634 8175 3637
rect 12065 3634 12131 3637
rect 8109 3632 12131 3634
rect 8109 3576 8114 3632
rect 8170 3576 12070 3632
rect 12126 3576 12131 3632
rect 21265 3634 21331 3637
rect 23197 3634 23263 3637
rect 21265 3632 23263 3634
rect 18137 3600 18203 3603
rect 8109 3574 12131 3576
rect 8109 3571 8175 3574
rect 12065 3571 12131 3574
rect 17910 3598 18203 3600
rect 17910 3542 18142 3598
rect 18198 3542 18203 3598
rect 21265 3576 21270 3632
rect 21326 3576 23202 3632
rect 23258 3576 23263 3632
rect 21265 3574 23263 3576
rect 21265 3571 21331 3574
rect 23197 3571 23263 3574
rect 17910 3540 18203 3542
rect 2037 3498 2103 3501
rect 6269 3498 6335 3501
rect 2037 3496 6335 3498
rect 2037 3440 2042 3496
rect 2098 3440 6274 3496
rect 6330 3440 6335 3496
rect 2037 3438 6335 3440
rect 2037 3435 2103 3438
rect 6269 3435 6335 3438
rect 11881 3498 11947 3501
rect 17910 3498 17970 3540
rect 18137 3537 18203 3540
rect 11881 3496 17970 3498
rect 11881 3440 11886 3496
rect 11942 3440 17970 3496
rect 11881 3438 17970 3440
rect 11881 3435 11947 3438
rect 0 3362 480 3392
rect 1577 3362 1643 3365
rect 0 3360 1643 3362
rect 0 3304 1582 3360
rect 1638 3304 1643 3360
rect 0 3302 1643 3304
rect 0 3272 480 3302
rect 1577 3299 1643 3302
rect 26693 3362 26759 3365
rect 29520 3362 30000 3392
rect 26693 3360 30000 3362
rect 26693 3304 26698 3360
rect 26754 3304 30000 3360
rect 26693 3302 30000 3304
rect 26693 3299 26759 3302
rect 5944 3296 6264 3297
rect 5944 3232 5952 3296
rect 6016 3232 6032 3296
rect 6096 3232 6112 3296
rect 6176 3232 6192 3296
rect 6256 3232 6264 3296
rect 5944 3231 6264 3232
rect 15944 3296 16264 3297
rect 15944 3232 15952 3296
rect 16016 3232 16032 3296
rect 16096 3232 16112 3296
rect 16176 3232 16192 3296
rect 16256 3232 16264 3296
rect 15944 3231 16264 3232
rect 25944 3296 26264 3297
rect 25944 3232 25952 3296
rect 26016 3232 26032 3296
rect 26096 3232 26112 3296
rect 26176 3232 26192 3296
rect 26256 3232 26264 3296
rect 29520 3272 30000 3302
rect 25944 3231 26264 3232
rect 11881 3226 11947 3229
rect 13813 3226 13879 3229
rect 11881 3224 13879 3226
rect 11881 3168 11886 3224
rect 11942 3168 13818 3224
rect 13874 3168 13879 3224
rect 11881 3166 13879 3168
rect 11881 3163 11947 3166
rect 13813 3163 13879 3166
rect 4153 3090 4219 3093
rect 14365 3090 14431 3093
rect 4153 3088 14431 3090
rect 4153 3032 4158 3088
rect 4214 3032 14370 3088
rect 14426 3032 14431 3088
rect 4153 3030 14431 3032
rect 4153 3027 4219 3030
rect 14365 3027 14431 3030
rect 20529 3090 20595 3093
rect 25313 3090 25379 3093
rect 20529 3088 25379 3090
rect 20529 3032 20534 3088
rect 20590 3032 25318 3088
rect 25374 3032 25379 3088
rect 20529 3030 25379 3032
rect 20529 3027 20595 3030
rect 25313 3027 25379 3030
rect 8293 2954 8359 2957
rect 13169 2954 13235 2957
rect 8293 2952 13235 2954
rect 8293 2896 8298 2952
rect 8354 2896 13174 2952
rect 13230 2896 13235 2952
rect 8293 2894 13235 2896
rect 8293 2891 8359 2894
rect 13169 2891 13235 2894
rect 20253 2954 20319 2957
rect 22185 2954 22251 2957
rect 20253 2952 22251 2954
rect 20253 2896 20258 2952
rect 20314 2896 22190 2952
rect 22246 2896 22251 2952
rect 20253 2894 22251 2896
rect 20253 2891 20319 2894
rect 22185 2891 22251 2894
rect 25497 2954 25563 2957
rect 27337 2954 27403 2957
rect 25497 2952 27403 2954
rect 25497 2896 25502 2952
rect 25558 2896 27342 2952
rect 27398 2896 27403 2952
rect 25497 2894 27403 2896
rect 25497 2891 25563 2894
rect 27337 2891 27403 2894
rect 565 2818 631 2821
rect 2957 2818 3023 2821
rect 565 2816 3023 2818
rect 565 2760 570 2816
rect 626 2760 2962 2816
rect 3018 2760 3023 2816
rect 565 2758 3023 2760
rect 565 2755 631 2758
rect 2957 2755 3023 2758
rect 13353 2818 13419 2821
rect 14917 2818 14983 2821
rect 13353 2816 14983 2818
rect 13353 2760 13358 2816
rect 13414 2760 14922 2816
rect 14978 2760 14983 2816
rect 13353 2758 14983 2760
rect 13353 2755 13419 2758
rect 14917 2755 14983 2758
rect 25865 2818 25931 2821
rect 29361 2818 29427 2821
rect 25865 2816 29427 2818
rect 25865 2760 25870 2816
rect 25926 2760 29366 2816
rect 29422 2760 29427 2816
rect 25865 2758 29427 2760
rect 25865 2755 25931 2758
rect 29361 2755 29427 2758
rect 10944 2752 11264 2753
rect 0 2682 480 2712
rect 10944 2688 10952 2752
rect 11016 2688 11032 2752
rect 11096 2688 11112 2752
rect 11176 2688 11192 2752
rect 11256 2688 11264 2752
rect 10944 2687 11264 2688
rect 20944 2752 21264 2753
rect 20944 2688 20952 2752
rect 21016 2688 21032 2752
rect 21096 2688 21112 2752
rect 21176 2688 21192 2752
rect 21256 2688 21264 2752
rect 20944 2687 21264 2688
rect 1577 2682 1643 2685
rect 0 2680 1643 2682
rect 0 2624 1582 2680
rect 1638 2624 1643 2680
rect 0 2622 1643 2624
rect 0 2592 480 2622
rect 1577 2619 1643 2622
rect 4889 2682 4955 2685
rect 8017 2682 8083 2685
rect 4889 2680 8083 2682
rect 4889 2624 4894 2680
rect 4950 2624 8022 2680
rect 8078 2624 8083 2680
rect 4889 2622 8083 2624
rect 4889 2619 4955 2622
rect 8017 2619 8083 2622
rect 25773 2682 25839 2685
rect 29520 2682 30000 2712
rect 25773 2680 30000 2682
rect 25773 2624 25778 2680
rect 25834 2624 30000 2680
rect 25773 2622 30000 2624
rect 25773 2619 25839 2622
rect 29520 2592 30000 2622
rect 18229 2546 18295 2549
rect 24393 2546 24459 2549
rect 18229 2544 24459 2546
rect 18229 2488 18234 2544
rect 18290 2488 24398 2544
rect 24454 2488 24459 2544
rect 18229 2486 24459 2488
rect 18229 2483 18295 2486
rect 24393 2483 24459 2486
rect 19241 2410 19307 2413
rect 19241 2408 27906 2410
rect 19241 2352 19246 2408
rect 19302 2352 27906 2408
rect 19241 2350 27906 2352
rect 19241 2347 19307 2350
rect 5944 2208 6264 2209
rect 0 2138 480 2168
rect 5944 2144 5952 2208
rect 6016 2144 6032 2208
rect 6096 2144 6112 2208
rect 6176 2144 6192 2208
rect 6256 2144 6264 2208
rect 5944 2143 6264 2144
rect 15944 2208 16264 2209
rect 15944 2144 15952 2208
rect 16016 2144 16032 2208
rect 16096 2144 16112 2208
rect 16176 2144 16192 2208
rect 16256 2144 16264 2208
rect 15944 2143 16264 2144
rect 25944 2208 26264 2209
rect 25944 2144 25952 2208
rect 26016 2144 26032 2208
rect 26096 2144 26112 2208
rect 26176 2144 26192 2208
rect 26256 2144 26264 2208
rect 25944 2143 26264 2144
rect 2681 2138 2747 2141
rect 0 2136 2747 2138
rect 0 2080 2686 2136
rect 2742 2080 2747 2136
rect 0 2078 2747 2080
rect 27846 2138 27906 2350
rect 29520 2138 30000 2168
rect 27846 2078 30000 2138
rect 0 2048 480 2078
rect 2681 2075 2747 2078
rect 29520 2048 30000 2078
rect 15653 2002 15719 2005
rect 24209 2002 24275 2005
rect 15653 2000 24275 2002
rect 15653 1944 15658 2000
rect 15714 1944 24214 2000
rect 24270 1944 24275 2000
rect 15653 1942 24275 1944
rect 15653 1939 15719 1942
rect 24209 1939 24275 1942
rect 0 1458 480 1488
rect 2865 1458 2931 1461
rect 0 1456 2931 1458
rect 0 1400 2870 1456
rect 2926 1400 2931 1456
rect 0 1398 2931 1400
rect 0 1368 480 1398
rect 2865 1395 2931 1398
rect 17861 1458 17927 1461
rect 25221 1458 25287 1461
rect 17861 1456 25287 1458
rect 17861 1400 17866 1456
rect 17922 1400 25226 1456
rect 25282 1400 25287 1456
rect 17861 1398 25287 1400
rect 17861 1395 17927 1398
rect 25221 1395 25287 1398
rect 27061 1458 27127 1461
rect 29520 1458 30000 1488
rect 27061 1456 30000 1458
rect 27061 1400 27066 1456
rect 27122 1400 30000 1456
rect 27061 1398 30000 1400
rect 27061 1395 27127 1398
rect 29520 1368 30000 1398
rect 0 914 480 944
rect 4061 914 4127 917
rect 0 912 4127 914
rect 0 856 4066 912
rect 4122 856 4127 912
rect 0 854 4127 856
rect 0 824 480 854
rect 4061 851 4127 854
rect 19149 914 19215 917
rect 29520 914 30000 944
rect 19149 912 30000 914
rect 19149 856 19154 912
rect 19210 856 30000 912
rect 19149 854 30000 856
rect 19149 851 19215 854
rect 29520 824 30000 854
rect 0 370 480 400
rect 2773 370 2839 373
rect 0 368 2839 370
rect 0 312 2778 368
rect 2834 312 2839 368
rect 0 310 2839 312
rect 0 280 480 310
rect 2773 307 2839 310
rect 26601 370 26667 373
rect 29520 370 30000 400
rect 26601 368 30000 370
rect 26601 312 26606 368
rect 26662 312 30000 368
rect 26601 310 30000 312
rect 26601 307 26667 310
rect 29520 280 30000 310
<< via3 >>
rect 5952 21788 6016 21792
rect 5952 21732 5956 21788
rect 5956 21732 6012 21788
rect 6012 21732 6016 21788
rect 5952 21728 6016 21732
rect 6032 21788 6096 21792
rect 6032 21732 6036 21788
rect 6036 21732 6092 21788
rect 6092 21732 6096 21788
rect 6032 21728 6096 21732
rect 6112 21788 6176 21792
rect 6112 21732 6116 21788
rect 6116 21732 6172 21788
rect 6172 21732 6176 21788
rect 6112 21728 6176 21732
rect 6192 21788 6256 21792
rect 6192 21732 6196 21788
rect 6196 21732 6252 21788
rect 6252 21732 6256 21788
rect 6192 21728 6256 21732
rect 15952 21788 16016 21792
rect 15952 21732 15956 21788
rect 15956 21732 16012 21788
rect 16012 21732 16016 21788
rect 15952 21728 16016 21732
rect 16032 21788 16096 21792
rect 16032 21732 16036 21788
rect 16036 21732 16092 21788
rect 16092 21732 16096 21788
rect 16032 21728 16096 21732
rect 16112 21788 16176 21792
rect 16112 21732 16116 21788
rect 16116 21732 16172 21788
rect 16172 21732 16176 21788
rect 16112 21728 16176 21732
rect 16192 21788 16256 21792
rect 16192 21732 16196 21788
rect 16196 21732 16252 21788
rect 16252 21732 16256 21788
rect 16192 21728 16256 21732
rect 25952 21788 26016 21792
rect 25952 21732 25956 21788
rect 25956 21732 26012 21788
rect 26012 21732 26016 21788
rect 25952 21728 26016 21732
rect 26032 21788 26096 21792
rect 26032 21732 26036 21788
rect 26036 21732 26092 21788
rect 26092 21732 26096 21788
rect 26032 21728 26096 21732
rect 26112 21788 26176 21792
rect 26112 21732 26116 21788
rect 26116 21732 26172 21788
rect 26172 21732 26176 21788
rect 26112 21728 26176 21732
rect 26192 21788 26256 21792
rect 26192 21732 26196 21788
rect 26196 21732 26252 21788
rect 26252 21732 26256 21788
rect 26192 21728 26256 21732
rect 10952 21244 11016 21248
rect 10952 21188 10956 21244
rect 10956 21188 11012 21244
rect 11012 21188 11016 21244
rect 10952 21184 11016 21188
rect 11032 21244 11096 21248
rect 11032 21188 11036 21244
rect 11036 21188 11092 21244
rect 11092 21188 11096 21244
rect 11032 21184 11096 21188
rect 11112 21244 11176 21248
rect 11112 21188 11116 21244
rect 11116 21188 11172 21244
rect 11172 21188 11176 21244
rect 11112 21184 11176 21188
rect 11192 21244 11256 21248
rect 11192 21188 11196 21244
rect 11196 21188 11252 21244
rect 11252 21188 11256 21244
rect 11192 21184 11256 21188
rect 20952 21244 21016 21248
rect 20952 21188 20956 21244
rect 20956 21188 21012 21244
rect 21012 21188 21016 21244
rect 20952 21184 21016 21188
rect 21032 21244 21096 21248
rect 21032 21188 21036 21244
rect 21036 21188 21092 21244
rect 21092 21188 21096 21244
rect 21032 21184 21096 21188
rect 21112 21244 21176 21248
rect 21112 21188 21116 21244
rect 21116 21188 21172 21244
rect 21172 21188 21176 21244
rect 21112 21184 21176 21188
rect 21192 21244 21256 21248
rect 21192 21188 21196 21244
rect 21196 21188 21252 21244
rect 21252 21188 21256 21244
rect 21192 21184 21256 21188
rect 5952 20700 6016 20704
rect 5952 20644 5956 20700
rect 5956 20644 6012 20700
rect 6012 20644 6016 20700
rect 5952 20640 6016 20644
rect 6032 20700 6096 20704
rect 6032 20644 6036 20700
rect 6036 20644 6092 20700
rect 6092 20644 6096 20700
rect 6032 20640 6096 20644
rect 6112 20700 6176 20704
rect 6112 20644 6116 20700
rect 6116 20644 6172 20700
rect 6172 20644 6176 20700
rect 6112 20640 6176 20644
rect 6192 20700 6256 20704
rect 6192 20644 6196 20700
rect 6196 20644 6252 20700
rect 6252 20644 6256 20700
rect 6192 20640 6256 20644
rect 15952 20700 16016 20704
rect 15952 20644 15956 20700
rect 15956 20644 16012 20700
rect 16012 20644 16016 20700
rect 15952 20640 16016 20644
rect 16032 20700 16096 20704
rect 16032 20644 16036 20700
rect 16036 20644 16092 20700
rect 16092 20644 16096 20700
rect 16032 20640 16096 20644
rect 16112 20700 16176 20704
rect 16112 20644 16116 20700
rect 16116 20644 16172 20700
rect 16172 20644 16176 20700
rect 16112 20640 16176 20644
rect 16192 20700 16256 20704
rect 16192 20644 16196 20700
rect 16196 20644 16252 20700
rect 16252 20644 16256 20700
rect 16192 20640 16256 20644
rect 25952 20700 26016 20704
rect 25952 20644 25956 20700
rect 25956 20644 26012 20700
rect 26012 20644 26016 20700
rect 25952 20640 26016 20644
rect 26032 20700 26096 20704
rect 26032 20644 26036 20700
rect 26036 20644 26092 20700
rect 26092 20644 26096 20700
rect 26032 20640 26096 20644
rect 26112 20700 26176 20704
rect 26112 20644 26116 20700
rect 26116 20644 26172 20700
rect 26172 20644 26176 20700
rect 26112 20640 26176 20644
rect 26192 20700 26256 20704
rect 26192 20644 26196 20700
rect 26196 20644 26252 20700
rect 26252 20644 26256 20700
rect 26192 20640 26256 20644
rect 10952 20156 11016 20160
rect 10952 20100 10956 20156
rect 10956 20100 11012 20156
rect 11012 20100 11016 20156
rect 10952 20096 11016 20100
rect 11032 20156 11096 20160
rect 11032 20100 11036 20156
rect 11036 20100 11092 20156
rect 11092 20100 11096 20156
rect 11032 20096 11096 20100
rect 11112 20156 11176 20160
rect 11112 20100 11116 20156
rect 11116 20100 11172 20156
rect 11172 20100 11176 20156
rect 11112 20096 11176 20100
rect 11192 20156 11256 20160
rect 11192 20100 11196 20156
rect 11196 20100 11252 20156
rect 11252 20100 11256 20156
rect 11192 20096 11256 20100
rect 20952 20156 21016 20160
rect 20952 20100 20956 20156
rect 20956 20100 21012 20156
rect 21012 20100 21016 20156
rect 20952 20096 21016 20100
rect 21032 20156 21096 20160
rect 21032 20100 21036 20156
rect 21036 20100 21092 20156
rect 21092 20100 21096 20156
rect 21032 20096 21096 20100
rect 21112 20156 21176 20160
rect 21112 20100 21116 20156
rect 21116 20100 21172 20156
rect 21172 20100 21176 20156
rect 21112 20096 21176 20100
rect 21192 20156 21256 20160
rect 21192 20100 21196 20156
rect 21196 20100 21252 20156
rect 21252 20100 21256 20156
rect 21192 20096 21256 20100
rect 5952 19612 6016 19616
rect 5952 19556 5956 19612
rect 5956 19556 6012 19612
rect 6012 19556 6016 19612
rect 5952 19552 6016 19556
rect 6032 19612 6096 19616
rect 6032 19556 6036 19612
rect 6036 19556 6092 19612
rect 6092 19556 6096 19612
rect 6032 19552 6096 19556
rect 6112 19612 6176 19616
rect 6112 19556 6116 19612
rect 6116 19556 6172 19612
rect 6172 19556 6176 19612
rect 6112 19552 6176 19556
rect 6192 19612 6256 19616
rect 6192 19556 6196 19612
rect 6196 19556 6252 19612
rect 6252 19556 6256 19612
rect 6192 19552 6256 19556
rect 15952 19612 16016 19616
rect 15952 19556 15956 19612
rect 15956 19556 16012 19612
rect 16012 19556 16016 19612
rect 15952 19552 16016 19556
rect 16032 19612 16096 19616
rect 16032 19556 16036 19612
rect 16036 19556 16092 19612
rect 16092 19556 16096 19612
rect 16032 19552 16096 19556
rect 16112 19612 16176 19616
rect 16112 19556 16116 19612
rect 16116 19556 16172 19612
rect 16172 19556 16176 19612
rect 16112 19552 16176 19556
rect 16192 19612 16256 19616
rect 16192 19556 16196 19612
rect 16196 19556 16252 19612
rect 16252 19556 16256 19612
rect 16192 19552 16256 19556
rect 25952 19612 26016 19616
rect 25952 19556 25956 19612
rect 25956 19556 26012 19612
rect 26012 19556 26016 19612
rect 25952 19552 26016 19556
rect 26032 19612 26096 19616
rect 26032 19556 26036 19612
rect 26036 19556 26092 19612
rect 26092 19556 26096 19612
rect 26032 19552 26096 19556
rect 26112 19612 26176 19616
rect 26112 19556 26116 19612
rect 26116 19556 26172 19612
rect 26172 19556 26176 19612
rect 26112 19552 26176 19556
rect 26192 19612 26256 19616
rect 26192 19556 26196 19612
rect 26196 19556 26252 19612
rect 26252 19556 26256 19612
rect 26192 19552 26256 19556
rect 10952 19068 11016 19072
rect 10952 19012 10956 19068
rect 10956 19012 11012 19068
rect 11012 19012 11016 19068
rect 10952 19008 11016 19012
rect 11032 19068 11096 19072
rect 11032 19012 11036 19068
rect 11036 19012 11092 19068
rect 11092 19012 11096 19068
rect 11032 19008 11096 19012
rect 11112 19068 11176 19072
rect 11112 19012 11116 19068
rect 11116 19012 11172 19068
rect 11172 19012 11176 19068
rect 11112 19008 11176 19012
rect 11192 19068 11256 19072
rect 11192 19012 11196 19068
rect 11196 19012 11252 19068
rect 11252 19012 11256 19068
rect 11192 19008 11256 19012
rect 20952 19068 21016 19072
rect 20952 19012 20956 19068
rect 20956 19012 21012 19068
rect 21012 19012 21016 19068
rect 20952 19008 21016 19012
rect 21032 19068 21096 19072
rect 21032 19012 21036 19068
rect 21036 19012 21092 19068
rect 21092 19012 21096 19068
rect 21032 19008 21096 19012
rect 21112 19068 21176 19072
rect 21112 19012 21116 19068
rect 21116 19012 21172 19068
rect 21172 19012 21176 19068
rect 21112 19008 21176 19012
rect 21192 19068 21256 19072
rect 21192 19012 21196 19068
rect 21196 19012 21252 19068
rect 21252 19012 21256 19068
rect 21192 19008 21256 19012
rect 5952 18524 6016 18528
rect 5952 18468 5956 18524
rect 5956 18468 6012 18524
rect 6012 18468 6016 18524
rect 5952 18464 6016 18468
rect 6032 18524 6096 18528
rect 6032 18468 6036 18524
rect 6036 18468 6092 18524
rect 6092 18468 6096 18524
rect 6032 18464 6096 18468
rect 6112 18524 6176 18528
rect 6112 18468 6116 18524
rect 6116 18468 6172 18524
rect 6172 18468 6176 18524
rect 6112 18464 6176 18468
rect 6192 18524 6256 18528
rect 6192 18468 6196 18524
rect 6196 18468 6252 18524
rect 6252 18468 6256 18524
rect 6192 18464 6256 18468
rect 15952 18524 16016 18528
rect 15952 18468 15956 18524
rect 15956 18468 16012 18524
rect 16012 18468 16016 18524
rect 15952 18464 16016 18468
rect 16032 18524 16096 18528
rect 16032 18468 16036 18524
rect 16036 18468 16092 18524
rect 16092 18468 16096 18524
rect 16032 18464 16096 18468
rect 16112 18524 16176 18528
rect 16112 18468 16116 18524
rect 16116 18468 16172 18524
rect 16172 18468 16176 18524
rect 16112 18464 16176 18468
rect 16192 18524 16256 18528
rect 16192 18468 16196 18524
rect 16196 18468 16252 18524
rect 16252 18468 16256 18524
rect 16192 18464 16256 18468
rect 25952 18524 26016 18528
rect 25952 18468 25956 18524
rect 25956 18468 26012 18524
rect 26012 18468 26016 18524
rect 25952 18464 26016 18468
rect 26032 18524 26096 18528
rect 26032 18468 26036 18524
rect 26036 18468 26092 18524
rect 26092 18468 26096 18524
rect 26032 18464 26096 18468
rect 26112 18524 26176 18528
rect 26112 18468 26116 18524
rect 26116 18468 26172 18524
rect 26172 18468 26176 18524
rect 26112 18464 26176 18468
rect 26192 18524 26256 18528
rect 26192 18468 26196 18524
rect 26196 18468 26252 18524
rect 26252 18468 26256 18524
rect 26192 18464 26256 18468
rect 10952 17980 11016 17984
rect 10952 17924 10956 17980
rect 10956 17924 11012 17980
rect 11012 17924 11016 17980
rect 10952 17920 11016 17924
rect 11032 17980 11096 17984
rect 11032 17924 11036 17980
rect 11036 17924 11092 17980
rect 11092 17924 11096 17980
rect 11032 17920 11096 17924
rect 11112 17980 11176 17984
rect 11112 17924 11116 17980
rect 11116 17924 11172 17980
rect 11172 17924 11176 17980
rect 11112 17920 11176 17924
rect 11192 17980 11256 17984
rect 11192 17924 11196 17980
rect 11196 17924 11252 17980
rect 11252 17924 11256 17980
rect 11192 17920 11256 17924
rect 20952 17980 21016 17984
rect 20952 17924 20956 17980
rect 20956 17924 21012 17980
rect 21012 17924 21016 17980
rect 20952 17920 21016 17924
rect 21032 17980 21096 17984
rect 21032 17924 21036 17980
rect 21036 17924 21092 17980
rect 21092 17924 21096 17980
rect 21032 17920 21096 17924
rect 21112 17980 21176 17984
rect 21112 17924 21116 17980
rect 21116 17924 21172 17980
rect 21172 17924 21176 17980
rect 21112 17920 21176 17924
rect 21192 17980 21256 17984
rect 21192 17924 21196 17980
rect 21196 17924 21252 17980
rect 21252 17924 21256 17980
rect 21192 17920 21256 17924
rect 5952 17436 6016 17440
rect 5952 17380 5956 17436
rect 5956 17380 6012 17436
rect 6012 17380 6016 17436
rect 5952 17376 6016 17380
rect 6032 17436 6096 17440
rect 6032 17380 6036 17436
rect 6036 17380 6092 17436
rect 6092 17380 6096 17436
rect 6032 17376 6096 17380
rect 6112 17436 6176 17440
rect 6112 17380 6116 17436
rect 6116 17380 6172 17436
rect 6172 17380 6176 17436
rect 6112 17376 6176 17380
rect 6192 17436 6256 17440
rect 6192 17380 6196 17436
rect 6196 17380 6252 17436
rect 6252 17380 6256 17436
rect 6192 17376 6256 17380
rect 15952 17436 16016 17440
rect 15952 17380 15956 17436
rect 15956 17380 16012 17436
rect 16012 17380 16016 17436
rect 15952 17376 16016 17380
rect 16032 17436 16096 17440
rect 16032 17380 16036 17436
rect 16036 17380 16092 17436
rect 16092 17380 16096 17436
rect 16032 17376 16096 17380
rect 16112 17436 16176 17440
rect 16112 17380 16116 17436
rect 16116 17380 16172 17436
rect 16172 17380 16176 17436
rect 16112 17376 16176 17380
rect 16192 17436 16256 17440
rect 16192 17380 16196 17436
rect 16196 17380 16252 17436
rect 16252 17380 16256 17436
rect 16192 17376 16256 17380
rect 25952 17436 26016 17440
rect 25952 17380 25956 17436
rect 25956 17380 26012 17436
rect 26012 17380 26016 17436
rect 25952 17376 26016 17380
rect 26032 17436 26096 17440
rect 26032 17380 26036 17436
rect 26036 17380 26092 17436
rect 26092 17380 26096 17436
rect 26032 17376 26096 17380
rect 26112 17436 26176 17440
rect 26112 17380 26116 17436
rect 26116 17380 26172 17436
rect 26172 17380 26176 17436
rect 26112 17376 26176 17380
rect 26192 17436 26256 17440
rect 26192 17380 26196 17436
rect 26196 17380 26252 17436
rect 26252 17380 26256 17436
rect 26192 17376 26256 17380
rect 10952 16892 11016 16896
rect 10952 16836 10956 16892
rect 10956 16836 11012 16892
rect 11012 16836 11016 16892
rect 10952 16832 11016 16836
rect 11032 16892 11096 16896
rect 11032 16836 11036 16892
rect 11036 16836 11092 16892
rect 11092 16836 11096 16892
rect 11032 16832 11096 16836
rect 11112 16892 11176 16896
rect 11112 16836 11116 16892
rect 11116 16836 11172 16892
rect 11172 16836 11176 16892
rect 11112 16832 11176 16836
rect 11192 16892 11256 16896
rect 11192 16836 11196 16892
rect 11196 16836 11252 16892
rect 11252 16836 11256 16892
rect 11192 16832 11256 16836
rect 20952 16892 21016 16896
rect 20952 16836 20956 16892
rect 20956 16836 21012 16892
rect 21012 16836 21016 16892
rect 20952 16832 21016 16836
rect 21032 16892 21096 16896
rect 21032 16836 21036 16892
rect 21036 16836 21092 16892
rect 21092 16836 21096 16892
rect 21032 16832 21096 16836
rect 21112 16892 21176 16896
rect 21112 16836 21116 16892
rect 21116 16836 21172 16892
rect 21172 16836 21176 16892
rect 21112 16832 21176 16836
rect 21192 16892 21256 16896
rect 21192 16836 21196 16892
rect 21196 16836 21252 16892
rect 21252 16836 21256 16892
rect 21192 16832 21256 16836
rect 5952 16348 6016 16352
rect 5952 16292 5956 16348
rect 5956 16292 6012 16348
rect 6012 16292 6016 16348
rect 5952 16288 6016 16292
rect 6032 16348 6096 16352
rect 6032 16292 6036 16348
rect 6036 16292 6092 16348
rect 6092 16292 6096 16348
rect 6032 16288 6096 16292
rect 6112 16348 6176 16352
rect 6112 16292 6116 16348
rect 6116 16292 6172 16348
rect 6172 16292 6176 16348
rect 6112 16288 6176 16292
rect 6192 16348 6256 16352
rect 6192 16292 6196 16348
rect 6196 16292 6252 16348
rect 6252 16292 6256 16348
rect 6192 16288 6256 16292
rect 15952 16348 16016 16352
rect 15952 16292 15956 16348
rect 15956 16292 16012 16348
rect 16012 16292 16016 16348
rect 15952 16288 16016 16292
rect 16032 16348 16096 16352
rect 16032 16292 16036 16348
rect 16036 16292 16092 16348
rect 16092 16292 16096 16348
rect 16032 16288 16096 16292
rect 16112 16348 16176 16352
rect 16112 16292 16116 16348
rect 16116 16292 16172 16348
rect 16172 16292 16176 16348
rect 16112 16288 16176 16292
rect 16192 16348 16256 16352
rect 16192 16292 16196 16348
rect 16196 16292 16252 16348
rect 16252 16292 16256 16348
rect 16192 16288 16256 16292
rect 25952 16348 26016 16352
rect 25952 16292 25956 16348
rect 25956 16292 26012 16348
rect 26012 16292 26016 16348
rect 25952 16288 26016 16292
rect 26032 16348 26096 16352
rect 26032 16292 26036 16348
rect 26036 16292 26092 16348
rect 26092 16292 26096 16348
rect 26032 16288 26096 16292
rect 26112 16348 26176 16352
rect 26112 16292 26116 16348
rect 26116 16292 26172 16348
rect 26172 16292 26176 16348
rect 26112 16288 26176 16292
rect 26192 16348 26256 16352
rect 26192 16292 26196 16348
rect 26196 16292 26252 16348
rect 26252 16292 26256 16348
rect 26192 16288 26256 16292
rect 10952 15804 11016 15808
rect 10952 15748 10956 15804
rect 10956 15748 11012 15804
rect 11012 15748 11016 15804
rect 10952 15744 11016 15748
rect 11032 15804 11096 15808
rect 11032 15748 11036 15804
rect 11036 15748 11092 15804
rect 11092 15748 11096 15804
rect 11032 15744 11096 15748
rect 11112 15804 11176 15808
rect 11112 15748 11116 15804
rect 11116 15748 11172 15804
rect 11172 15748 11176 15804
rect 11112 15744 11176 15748
rect 11192 15804 11256 15808
rect 11192 15748 11196 15804
rect 11196 15748 11252 15804
rect 11252 15748 11256 15804
rect 11192 15744 11256 15748
rect 20952 15804 21016 15808
rect 20952 15748 20956 15804
rect 20956 15748 21012 15804
rect 21012 15748 21016 15804
rect 20952 15744 21016 15748
rect 21032 15804 21096 15808
rect 21032 15748 21036 15804
rect 21036 15748 21092 15804
rect 21092 15748 21096 15804
rect 21032 15744 21096 15748
rect 21112 15804 21176 15808
rect 21112 15748 21116 15804
rect 21116 15748 21172 15804
rect 21172 15748 21176 15804
rect 21112 15744 21176 15748
rect 21192 15804 21256 15808
rect 21192 15748 21196 15804
rect 21196 15748 21252 15804
rect 21252 15748 21256 15804
rect 21192 15744 21256 15748
rect 5952 15260 6016 15264
rect 5952 15204 5956 15260
rect 5956 15204 6012 15260
rect 6012 15204 6016 15260
rect 5952 15200 6016 15204
rect 6032 15260 6096 15264
rect 6032 15204 6036 15260
rect 6036 15204 6092 15260
rect 6092 15204 6096 15260
rect 6032 15200 6096 15204
rect 6112 15260 6176 15264
rect 6112 15204 6116 15260
rect 6116 15204 6172 15260
rect 6172 15204 6176 15260
rect 6112 15200 6176 15204
rect 6192 15260 6256 15264
rect 6192 15204 6196 15260
rect 6196 15204 6252 15260
rect 6252 15204 6256 15260
rect 6192 15200 6256 15204
rect 15952 15260 16016 15264
rect 15952 15204 15956 15260
rect 15956 15204 16012 15260
rect 16012 15204 16016 15260
rect 15952 15200 16016 15204
rect 16032 15260 16096 15264
rect 16032 15204 16036 15260
rect 16036 15204 16092 15260
rect 16092 15204 16096 15260
rect 16032 15200 16096 15204
rect 16112 15260 16176 15264
rect 16112 15204 16116 15260
rect 16116 15204 16172 15260
rect 16172 15204 16176 15260
rect 16112 15200 16176 15204
rect 16192 15260 16256 15264
rect 16192 15204 16196 15260
rect 16196 15204 16252 15260
rect 16252 15204 16256 15260
rect 16192 15200 16256 15204
rect 25952 15260 26016 15264
rect 25952 15204 25956 15260
rect 25956 15204 26012 15260
rect 26012 15204 26016 15260
rect 25952 15200 26016 15204
rect 26032 15260 26096 15264
rect 26032 15204 26036 15260
rect 26036 15204 26092 15260
rect 26092 15204 26096 15260
rect 26032 15200 26096 15204
rect 26112 15260 26176 15264
rect 26112 15204 26116 15260
rect 26116 15204 26172 15260
rect 26172 15204 26176 15260
rect 26112 15200 26176 15204
rect 26192 15260 26256 15264
rect 26192 15204 26196 15260
rect 26196 15204 26252 15260
rect 26252 15204 26256 15260
rect 26192 15200 26256 15204
rect 10952 14716 11016 14720
rect 10952 14660 10956 14716
rect 10956 14660 11012 14716
rect 11012 14660 11016 14716
rect 10952 14656 11016 14660
rect 11032 14716 11096 14720
rect 11032 14660 11036 14716
rect 11036 14660 11092 14716
rect 11092 14660 11096 14716
rect 11032 14656 11096 14660
rect 11112 14716 11176 14720
rect 11112 14660 11116 14716
rect 11116 14660 11172 14716
rect 11172 14660 11176 14716
rect 11112 14656 11176 14660
rect 11192 14716 11256 14720
rect 11192 14660 11196 14716
rect 11196 14660 11252 14716
rect 11252 14660 11256 14716
rect 11192 14656 11256 14660
rect 20952 14716 21016 14720
rect 20952 14660 20956 14716
rect 20956 14660 21012 14716
rect 21012 14660 21016 14716
rect 20952 14656 21016 14660
rect 21032 14716 21096 14720
rect 21032 14660 21036 14716
rect 21036 14660 21092 14716
rect 21092 14660 21096 14716
rect 21032 14656 21096 14660
rect 21112 14716 21176 14720
rect 21112 14660 21116 14716
rect 21116 14660 21172 14716
rect 21172 14660 21176 14716
rect 21112 14656 21176 14660
rect 21192 14716 21256 14720
rect 21192 14660 21196 14716
rect 21196 14660 21252 14716
rect 21252 14660 21256 14716
rect 21192 14656 21256 14660
rect 5952 14172 6016 14176
rect 5952 14116 5956 14172
rect 5956 14116 6012 14172
rect 6012 14116 6016 14172
rect 5952 14112 6016 14116
rect 6032 14172 6096 14176
rect 6032 14116 6036 14172
rect 6036 14116 6092 14172
rect 6092 14116 6096 14172
rect 6032 14112 6096 14116
rect 6112 14172 6176 14176
rect 6112 14116 6116 14172
rect 6116 14116 6172 14172
rect 6172 14116 6176 14172
rect 6112 14112 6176 14116
rect 6192 14172 6256 14176
rect 6192 14116 6196 14172
rect 6196 14116 6252 14172
rect 6252 14116 6256 14172
rect 6192 14112 6256 14116
rect 15952 14172 16016 14176
rect 15952 14116 15956 14172
rect 15956 14116 16012 14172
rect 16012 14116 16016 14172
rect 15952 14112 16016 14116
rect 16032 14172 16096 14176
rect 16032 14116 16036 14172
rect 16036 14116 16092 14172
rect 16092 14116 16096 14172
rect 16032 14112 16096 14116
rect 16112 14172 16176 14176
rect 16112 14116 16116 14172
rect 16116 14116 16172 14172
rect 16172 14116 16176 14172
rect 16112 14112 16176 14116
rect 16192 14172 16256 14176
rect 16192 14116 16196 14172
rect 16196 14116 16252 14172
rect 16252 14116 16256 14172
rect 16192 14112 16256 14116
rect 25952 14172 26016 14176
rect 25952 14116 25956 14172
rect 25956 14116 26012 14172
rect 26012 14116 26016 14172
rect 25952 14112 26016 14116
rect 26032 14172 26096 14176
rect 26032 14116 26036 14172
rect 26036 14116 26092 14172
rect 26092 14116 26096 14172
rect 26032 14112 26096 14116
rect 26112 14172 26176 14176
rect 26112 14116 26116 14172
rect 26116 14116 26172 14172
rect 26172 14116 26176 14172
rect 26112 14112 26176 14116
rect 26192 14172 26256 14176
rect 26192 14116 26196 14172
rect 26196 14116 26252 14172
rect 26252 14116 26256 14172
rect 26192 14112 26256 14116
rect 10952 13628 11016 13632
rect 10952 13572 10956 13628
rect 10956 13572 11012 13628
rect 11012 13572 11016 13628
rect 10952 13568 11016 13572
rect 11032 13628 11096 13632
rect 11032 13572 11036 13628
rect 11036 13572 11092 13628
rect 11092 13572 11096 13628
rect 11032 13568 11096 13572
rect 11112 13628 11176 13632
rect 11112 13572 11116 13628
rect 11116 13572 11172 13628
rect 11172 13572 11176 13628
rect 11112 13568 11176 13572
rect 11192 13628 11256 13632
rect 11192 13572 11196 13628
rect 11196 13572 11252 13628
rect 11252 13572 11256 13628
rect 11192 13568 11256 13572
rect 20952 13628 21016 13632
rect 20952 13572 20956 13628
rect 20956 13572 21012 13628
rect 21012 13572 21016 13628
rect 20952 13568 21016 13572
rect 21032 13628 21096 13632
rect 21032 13572 21036 13628
rect 21036 13572 21092 13628
rect 21092 13572 21096 13628
rect 21032 13568 21096 13572
rect 21112 13628 21176 13632
rect 21112 13572 21116 13628
rect 21116 13572 21172 13628
rect 21172 13572 21176 13628
rect 21112 13568 21176 13572
rect 21192 13628 21256 13632
rect 21192 13572 21196 13628
rect 21196 13572 21252 13628
rect 21252 13572 21256 13628
rect 21192 13568 21256 13572
rect 5952 13084 6016 13088
rect 5952 13028 5956 13084
rect 5956 13028 6012 13084
rect 6012 13028 6016 13084
rect 5952 13024 6016 13028
rect 6032 13084 6096 13088
rect 6032 13028 6036 13084
rect 6036 13028 6092 13084
rect 6092 13028 6096 13084
rect 6032 13024 6096 13028
rect 6112 13084 6176 13088
rect 6112 13028 6116 13084
rect 6116 13028 6172 13084
rect 6172 13028 6176 13084
rect 6112 13024 6176 13028
rect 6192 13084 6256 13088
rect 6192 13028 6196 13084
rect 6196 13028 6252 13084
rect 6252 13028 6256 13084
rect 6192 13024 6256 13028
rect 15952 13084 16016 13088
rect 15952 13028 15956 13084
rect 15956 13028 16012 13084
rect 16012 13028 16016 13084
rect 15952 13024 16016 13028
rect 16032 13084 16096 13088
rect 16032 13028 16036 13084
rect 16036 13028 16092 13084
rect 16092 13028 16096 13084
rect 16032 13024 16096 13028
rect 16112 13084 16176 13088
rect 16112 13028 16116 13084
rect 16116 13028 16172 13084
rect 16172 13028 16176 13084
rect 16112 13024 16176 13028
rect 16192 13084 16256 13088
rect 16192 13028 16196 13084
rect 16196 13028 16252 13084
rect 16252 13028 16256 13084
rect 16192 13024 16256 13028
rect 25952 13084 26016 13088
rect 25952 13028 25956 13084
rect 25956 13028 26012 13084
rect 26012 13028 26016 13084
rect 25952 13024 26016 13028
rect 26032 13084 26096 13088
rect 26032 13028 26036 13084
rect 26036 13028 26092 13084
rect 26092 13028 26096 13084
rect 26032 13024 26096 13028
rect 26112 13084 26176 13088
rect 26112 13028 26116 13084
rect 26116 13028 26172 13084
rect 26172 13028 26176 13084
rect 26112 13024 26176 13028
rect 26192 13084 26256 13088
rect 26192 13028 26196 13084
rect 26196 13028 26252 13084
rect 26252 13028 26256 13084
rect 26192 13024 26256 13028
rect 10952 12540 11016 12544
rect 10952 12484 10956 12540
rect 10956 12484 11012 12540
rect 11012 12484 11016 12540
rect 10952 12480 11016 12484
rect 11032 12540 11096 12544
rect 11032 12484 11036 12540
rect 11036 12484 11092 12540
rect 11092 12484 11096 12540
rect 11032 12480 11096 12484
rect 11112 12540 11176 12544
rect 11112 12484 11116 12540
rect 11116 12484 11172 12540
rect 11172 12484 11176 12540
rect 11112 12480 11176 12484
rect 11192 12540 11256 12544
rect 11192 12484 11196 12540
rect 11196 12484 11252 12540
rect 11252 12484 11256 12540
rect 11192 12480 11256 12484
rect 20952 12540 21016 12544
rect 20952 12484 20956 12540
rect 20956 12484 21012 12540
rect 21012 12484 21016 12540
rect 20952 12480 21016 12484
rect 21032 12540 21096 12544
rect 21032 12484 21036 12540
rect 21036 12484 21092 12540
rect 21092 12484 21096 12540
rect 21032 12480 21096 12484
rect 21112 12540 21176 12544
rect 21112 12484 21116 12540
rect 21116 12484 21172 12540
rect 21172 12484 21176 12540
rect 21112 12480 21176 12484
rect 21192 12540 21256 12544
rect 21192 12484 21196 12540
rect 21196 12484 21252 12540
rect 21252 12484 21256 12540
rect 21192 12480 21256 12484
rect 5952 11996 6016 12000
rect 5952 11940 5956 11996
rect 5956 11940 6012 11996
rect 6012 11940 6016 11996
rect 5952 11936 6016 11940
rect 6032 11996 6096 12000
rect 6032 11940 6036 11996
rect 6036 11940 6092 11996
rect 6092 11940 6096 11996
rect 6032 11936 6096 11940
rect 6112 11996 6176 12000
rect 6112 11940 6116 11996
rect 6116 11940 6172 11996
rect 6172 11940 6176 11996
rect 6112 11936 6176 11940
rect 6192 11996 6256 12000
rect 6192 11940 6196 11996
rect 6196 11940 6252 11996
rect 6252 11940 6256 11996
rect 6192 11936 6256 11940
rect 15952 11996 16016 12000
rect 15952 11940 15956 11996
rect 15956 11940 16012 11996
rect 16012 11940 16016 11996
rect 15952 11936 16016 11940
rect 16032 11996 16096 12000
rect 16032 11940 16036 11996
rect 16036 11940 16092 11996
rect 16092 11940 16096 11996
rect 16032 11936 16096 11940
rect 16112 11996 16176 12000
rect 16112 11940 16116 11996
rect 16116 11940 16172 11996
rect 16172 11940 16176 11996
rect 16112 11936 16176 11940
rect 16192 11996 16256 12000
rect 16192 11940 16196 11996
rect 16196 11940 16252 11996
rect 16252 11940 16256 11996
rect 16192 11936 16256 11940
rect 25952 11996 26016 12000
rect 25952 11940 25956 11996
rect 25956 11940 26012 11996
rect 26012 11940 26016 11996
rect 25952 11936 26016 11940
rect 26032 11996 26096 12000
rect 26032 11940 26036 11996
rect 26036 11940 26092 11996
rect 26092 11940 26096 11996
rect 26032 11936 26096 11940
rect 26112 11996 26176 12000
rect 26112 11940 26116 11996
rect 26116 11940 26172 11996
rect 26172 11940 26176 11996
rect 26112 11936 26176 11940
rect 26192 11996 26256 12000
rect 26192 11940 26196 11996
rect 26196 11940 26252 11996
rect 26252 11940 26256 11996
rect 26192 11936 26256 11940
rect 10952 11452 11016 11456
rect 10952 11396 10956 11452
rect 10956 11396 11012 11452
rect 11012 11396 11016 11452
rect 10952 11392 11016 11396
rect 11032 11452 11096 11456
rect 11032 11396 11036 11452
rect 11036 11396 11092 11452
rect 11092 11396 11096 11452
rect 11032 11392 11096 11396
rect 11112 11452 11176 11456
rect 11112 11396 11116 11452
rect 11116 11396 11172 11452
rect 11172 11396 11176 11452
rect 11112 11392 11176 11396
rect 11192 11452 11256 11456
rect 11192 11396 11196 11452
rect 11196 11396 11252 11452
rect 11252 11396 11256 11452
rect 11192 11392 11256 11396
rect 20952 11452 21016 11456
rect 20952 11396 20956 11452
rect 20956 11396 21012 11452
rect 21012 11396 21016 11452
rect 20952 11392 21016 11396
rect 21032 11452 21096 11456
rect 21032 11396 21036 11452
rect 21036 11396 21092 11452
rect 21092 11396 21096 11452
rect 21032 11392 21096 11396
rect 21112 11452 21176 11456
rect 21112 11396 21116 11452
rect 21116 11396 21172 11452
rect 21172 11396 21176 11452
rect 21112 11392 21176 11396
rect 21192 11452 21256 11456
rect 21192 11396 21196 11452
rect 21196 11396 21252 11452
rect 21252 11396 21256 11452
rect 21192 11392 21256 11396
rect 5952 10908 6016 10912
rect 5952 10852 5956 10908
rect 5956 10852 6012 10908
rect 6012 10852 6016 10908
rect 5952 10848 6016 10852
rect 6032 10908 6096 10912
rect 6032 10852 6036 10908
rect 6036 10852 6092 10908
rect 6092 10852 6096 10908
rect 6032 10848 6096 10852
rect 6112 10908 6176 10912
rect 6112 10852 6116 10908
rect 6116 10852 6172 10908
rect 6172 10852 6176 10908
rect 6112 10848 6176 10852
rect 6192 10908 6256 10912
rect 6192 10852 6196 10908
rect 6196 10852 6252 10908
rect 6252 10852 6256 10908
rect 6192 10848 6256 10852
rect 15952 10908 16016 10912
rect 15952 10852 15956 10908
rect 15956 10852 16012 10908
rect 16012 10852 16016 10908
rect 15952 10848 16016 10852
rect 16032 10908 16096 10912
rect 16032 10852 16036 10908
rect 16036 10852 16092 10908
rect 16092 10852 16096 10908
rect 16032 10848 16096 10852
rect 16112 10908 16176 10912
rect 16112 10852 16116 10908
rect 16116 10852 16172 10908
rect 16172 10852 16176 10908
rect 16112 10848 16176 10852
rect 16192 10908 16256 10912
rect 16192 10852 16196 10908
rect 16196 10852 16252 10908
rect 16252 10852 16256 10908
rect 16192 10848 16256 10852
rect 25952 10908 26016 10912
rect 25952 10852 25956 10908
rect 25956 10852 26012 10908
rect 26012 10852 26016 10908
rect 25952 10848 26016 10852
rect 26032 10908 26096 10912
rect 26032 10852 26036 10908
rect 26036 10852 26092 10908
rect 26092 10852 26096 10908
rect 26032 10848 26096 10852
rect 26112 10908 26176 10912
rect 26112 10852 26116 10908
rect 26116 10852 26172 10908
rect 26172 10852 26176 10908
rect 26112 10848 26176 10852
rect 26192 10908 26256 10912
rect 26192 10852 26196 10908
rect 26196 10852 26252 10908
rect 26252 10852 26256 10908
rect 26192 10848 26256 10852
rect 10952 10364 11016 10368
rect 10952 10308 10956 10364
rect 10956 10308 11012 10364
rect 11012 10308 11016 10364
rect 10952 10304 11016 10308
rect 11032 10364 11096 10368
rect 11032 10308 11036 10364
rect 11036 10308 11092 10364
rect 11092 10308 11096 10364
rect 11032 10304 11096 10308
rect 11112 10364 11176 10368
rect 11112 10308 11116 10364
rect 11116 10308 11172 10364
rect 11172 10308 11176 10364
rect 11112 10304 11176 10308
rect 11192 10364 11256 10368
rect 11192 10308 11196 10364
rect 11196 10308 11252 10364
rect 11252 10308 11256 10364
rect 11192 10304 11256 10308
rect 20952 10364 21016 10368
rect 20952 10308 20956 10364
rect 20956 10308 21012 10364
rect 21012 10308 21016 10364
rect 20952 10304 21016 10308
rect 21032 10364 21096 10368
rect 21032 10308 21036 10364
rect 21036 10308 21092 10364
rect 21092 10308 21096 10364
rect 21032 10304 21096 10308
rect 21112 10364 21176 10368
rect 21112 10308 21116 10364
rect 21116 10308 21172 10364
rect 21172 10308 21176 10364
rect 21112 10304 21176 10308
rect 21192 10364 21256 10368
rect 21192 10308 21196 10364
rect 21196 10308 21252 10364
rect 21252 10308 21256 10364
rect 21192 10304 21256 10308
rect 5952 9820 6016 9824
rect 5952 9764 5956 9820
rect 5956 9764 6012 9820
rect 6012 9764 6016 9820
rect 5952 9760 6016 9764
rect 6032 9820 6096 9824
rect 6032 9764 6036 9820
rect 6036 9764 6092 9820
rect 6092 9764 6096 9820
rect 6032 9760 6096 9764
rect 6112 9820 6176 9824
rect 6112 9764 6116 9820
rect 6116 9764 6172 9820
rect 6172 9764 6176 9820
rect 6112 9760 6176 9764
rect 6192 9820 6256 9824
rect 6192 9764 6196 9820
rect 6196 9764 6252 9820
rect 6252 9764 6256 9820
rect 6192 9760 6256 9764
rect 15952 9820 16016 9824
rect 15952 9764 15956 9820
rect 15956 9764 16012 9820
rect 16012 9764 16016 9820
rect 15952 9760 16016 9764
rect 16032 9820 16096 9824
rect 16032 9764 16036 9820
rect 16036 9764 16092 9820
rect 16092 9764 16096 9820
rect 16032 9760 16096 9764
rect 16112 9820 16176 9824
rect 16112 9764 16116 9820
rect 16116 9764 16172 9820
rect 16172 9764 16176 9820
rect 16112 9760 16176 9764
rect 16192 9820 16256 9824
rect 16192 9764 16196 9820
rect 16196 9764 16252 9820
rect 16252 9764 16256 9820
rect 16192 9760 16256 9764
rect 25952 9820 26016 9824
rect 25952 9764 25956 9820
rect 25956 9764 26012 9820
rect 26012 9764 26016 9820
rect 25952 9760 26016 9764
rect 26032 9820 26096 9824
rect 26032 9764 26036 9820
rect 26036 9764 26092 9820
rect 26092 9764 26096 9820
rect 26032 9760 26096 9764
rect 26112 9820 26176 9824
rect 26112 9764 26116 9820
rect 26116 9764 26172 9820
rect 26172 9764 26176 9820
rect 26112 9760 26176 9764
rect 26192 9820 26256 9824
rect 26192 9764 26196 9820
rect 26196 9764 26252 9820
rect 26252 9764 26256 9820
rect 26192 9760 26256 9764
rect 10952 9276 11016 9280
rect 10952 9220 10956 9276
rect 10956 9220 11012 9276
rect 11012 9220 11016 9276
rect 10952 9216 11016 9220
rect 11032 9276 11096 9280
rect 11032 9220 11036 9276
rect 11036 9220 11092 9276
rect 11092 9220 11096 9276
rect 11032 9216 11096 9220
rect 11112 9276 11176 9280
rect 11112 9220 11116 9276
rect 11116 9220 11172 9276
rect 11172 9220 11176 9276
rect 11112 9216 11176 9220
rect 11192 9276 11256 9280
rect 11192 9220 11196 9276
rect 11196 9220 11252 9276
rect 11252 9220 11256 9276
rect 11192 9216 11256 9220
rect 20952 9276 21016 9280
rect 20952 9220 20956 9276
rect 20956 9220 21012 9276
rect 21012 9220 21016 9276
rect 20952 9216 21016 9220
rect 21032 9276 21096 9280
rect 21032 9220 21036 9276
rect 21036 9220 21092 9276
rect 21092 9220 21096 9276
rect 21032 9216 21096 9220
rect 21112 9276 21176 9280
rect 21112 9220 21116 9276
rect 21116 9220 21172 9276
rect 21172 9220 21176 9276
rect 21112 9216 21176 9220
rect 21192 9276 21256 9280
rect 21192 9220 21196 9276
rect 21196 9220 21252 9276
rect 21252 9220 21256 9276
rect 21192 9216 21256 9220
rect 26556 8936 26620 8940
rect 26556 8880 26570 8936
rect 26570 8880 26620 8936
rect 26556 8876 26620 8880
rect 5952 8732 6016 8736
rect 5952 8676 5956 8732
rect 5956 8676 6012 8732
rect 6012 8676 6016 8732
rect 5952 8672 6016 8676
rect 6032 8732 6096 8736
rect 6032 8676 6036 8732
rect 6036 8676 6092 8732
rect 6092 8676 6096 8732
rect 6032 8672 6096 8676
rect 6112 8732 6176 8736
rect 6112 8676 6116 8732
rect 6116 8676 6172 8732
rect 6172 8676 6176 8732
rect 6112 8672 6176 8676
rect 6192 8732 6256 8736
rect 6192 8676 6196 8732
rect 6196 8676 6252 8732
rect 6252 8676 6256 8732
rect 6192 8672 6256 8676
rect 15952 8732 16016 8736
rect 15952 8676 15956 8732
rect 15956 8676 16012 8732
rect 16012 8676 16016 8732
rect 15952 8672 16016 8676
rect 16032 8732 16096 8736
rect 16032 8676 16036 8732
rect 16036 8676 16092 8732
rect 16092 8676 16096 8732
rect 16032 8672 16096 8676
rect 16112 8732 16176 8736
rect 16112 8676 16116 8732
rect 16116 8676 16172 8732
rect 16172 8676 16176 8732
rect 16112 8672 16176 8676
rect 16192 8732 16256 8736
rect 16192 8676 16196 8732
rect 16196 8676 16252 8732
rect 16252 8676 16256 8732
rect 16192 8672 16256 8676
rect 25952 8732 26016 8736
rect 25952 8676 25956 8732
rect 25956 8676 26012 8732
rect 26012 8676 26016 8732
rect 25952 8672 26016 8676
rect 26032 8732 26096 8736
rect 26032 8676 26036 8732
rect 26036 8676 26092 8732
rect 26092 8676 26096 8732
rect 26032 8672 26096 8676
rect 26112 8732 26176 8736
rect 26112 8676 26116 8732
rect 26116 8676 26172 8732
rect 26172 8676 26176 8732
rect 26112 8672 26176 8676
rect 26192 8732 26256 8736
rect 26192 8676 26196 8732
rect 26196 8676 26252 8732
rect 26252 8676 26256 8732
rect 26192 8672 26256 8676
rect 7236 8528 7300 8532
rect 7236 8472 7250 8528
rect 7250 8472 7300 8528
rect 7236 8468 7300 8472
rect 10952 8188 11016 8192
rect 10952 8132 10956 8188
rect 10956 8132 11012 8188
rect 11012 8132 11016 8188
rect 10952 8128 11016 8132
rect 11032 8188 11096 8192
rect 11032 8132 11036 8188
rect 11036 8132 11092 8188
rect 11092 8132 11096 8188
rect 11032 8128 11096 8132
rect 11112 8188 11176 8192
rect 11112 8132 11116 8188
rect 11116 8132 11172 8188
rect 11172 8132 11176 8188
rect 11112 8128 11176 8132
rect 11192 8188 11256 8192
rect 11192 8132 11196 8188
rect 11196 8132 11252 8188
rect 11252 8132 11256 8188
rect 11192 8128 11256 8132
rect 20952 8188 21016 8192
rect 20952 8132 20956 8188
rect 20956 8132 21012 8188
rect 21012 8132 21016 8188
rect 20952 8128 21016 8132
rect 21032 8188 21096 8192
rect 21032 8132 21036 8188
rect 21036 8132 21092 8188
rect 21092 8132 21096 8188
rect 21032 8128 21096 8132
rect 21112 8188 21176 8192
rect 21112 8132 21116 8188
rect 21116 8132 21172 8188
rect 21172 8132 21176 8188
rect 21112 8128 21176 8132
rect 21192 8188 21256 8192
rect 21192 8132 21196 8188
rect 21196 8132 21252 8188
rect 21252 8132 21256 8188
rect 21192 8128 21256 8132
rect 5952 7644 6016 7648
rect 5952 7588 5956 7644
rect 5956 7588 6012 7644
rect 6012 7588 6016 7644
rect 5952 7584 6016 7588
rect 6032 7644 6096 7648
rect 6032 7588 6036 7644
rect 6036 7588 6092 7644
rect 6092 7588 6096 7644
rect 6032 7584 6096 7588
rect 6112 7644 6176 7648
rect 6112 7588 6116 7644
rect 6116 7588 6172 7644
rect 6172 7588 6176 7644
rect 6112 7584 6176 7588
rect 6192 7644 6256 7648
rect 6192 7588 6196 7644
rect 6196 7588 6252 7644
rect 6252 7588 6256 7644
rect 6192 7584 6256 7588
rect 15952 7644 16016 7648
rect 15952 7588 15956 7644
rect 15956 7588 16012 7644
rect 16012 7588 16016 7644
rect 15952 7584 16016 7588
rect 16032 7644 16096 7648
rect 16032 7588 16036 7644
rect 16036 7588 16092 7644
rect 16092 7588 16096 7644
rect 16032 7584 16096 7588
rect 16112 7644 16176 7648
rect 16112 7588 16116 7644
rect 16116 7588 16172 7644
rect 16172 7588 16176 7644
rect 16112 7584 16176 7588
rect 16192 7644 16256 7648
rect 16192 7588 16196 7644
rect 16196 7588 16252 7644
rect 16252 7588 16256 7644
rect 16192 7584 16256 7588
rect 25952 7644 26016 7648
rect 25952 7588 25956 7644
rect 25956 7588 26012 7644
rect 26012 7588 26016 7644
rect 25952 7584 26016 7588
rect 26032 7644 26096 7648
rect 26032 7588 26036 7644
rect 26036 7588 26092 7644
rect 26092 7588 26096 7644
rect 26032 7584 26096 7588
rect 26112 7644 26176 7648
rect 26112 7588 26116 7644
rect 26116 7588 26172 7644
rect 26172 7588 26176 7644
rect 26112 7584 26176 7588
rect 26192 7644 26256 7648
rect 26192 7588 26196 7644
rect 26196 7588 26252 7644
rect 26252 7588 26256 7644
rect 26192 7584 26256 7588
rect 10952 7100 11016 7104
rect 10952 7044 10956 7100
rect 10956 7044 11012 7100
rect 11012 7044 11016 7100
rect 10952 7040 11016 7044
rect 11032 7100 11096 7104
rect 11032 7044 11036 7100
rect 11036 7044 11092 7100
rect 11092 7044 11096 7100
rect 11032 7040 11096 7044
rect 11112 7100 11176 7104
rect 11112 7044 11116 7100
rect 11116 7044 11172 7100
rect 11172 7044 11176 7100
rect 11112 7040 11176 7044
rect 11192 7100 11256 7104
rect 11192 7044 11196 7100
rect 11196 7044 11252 7100
rect 11252 7044 11256 7100
rect 11192 7040 11256 7044
rect 20952 7100 21016 7104
rect 20952 7044 20956 7100
rect 20956 7044 21012 7100
rect 21012 7044 21016 7100
rect 20952 7040 21016 7044
rect 21032 7100 21096 7104
rect 21032 7044 21036 7100
rect 21036 7044 21092 7100
rect 21092 7044 21096 7100
rect 21032 7040 21096 7044
rect 21112 7100 21176 7104
rect 21112 7044 21116 7100
rect 21116 7044 21172 7100
rect 21172 7044 21176 7100
rect 21112 7040 21176 7044
rect 21192 7100 21256 7104
rect 21192 7044 21196 7100
rect 21196 7044 21252 7100
rect 21252 7044 21256 7100
rect 21192 7040 21256 7044
rect 5952 6556 6016 6560
rect 5952 6500 5956 6556
rect 5956 6500 6012 6556
rect 6012 6500 6016 6556
rect 5952 6496 6016 6500
rect 6032 6556 6096 6560
rect 6032 6500 6036 6556
rect 6036 6500 6092 6556
rect 6092 6500 6096 6556
rect 6032 6496 6096 6500
rect 6112 6556 6176 6560
rect 6112 6500 6116 6556
rect 6116 6500 6172 6556
rect 6172 6500 6176 6556
rect 6112 6496 6176 6500
rect 6192 6556 6256 6560
rect 6192 6500 6196 6556
rect 6196 6500 6252 6556
rect 6252 6500 6256 6556
rect 6192 6496 6256 6500
rect 15952 6556 16016 6560
rect 15952 6500 15956 6556
rect 15956 6500 16012 6556
rect 16012 6500 16016 6556
rect 15952 6496 16016 6500
rect 16032 6556 16096 6560
rect 16032 6500 16036 6556
rect 16036 6500 16092 6556
rect 16092 6500 16096 6556
rect 16032 6496 16096 6500
rect 16112 6556 16176 6560
rect 16112 6500 16116 6556
rect 16116 6500 16172 6556
rect 16172 6500 16176 6556
rect 16112 6496 16176 6500
rect 16192 6556 16256 6560
rect 16192 6500 16196 6556
rect 16196 6500 16252 6556
rect 16252 6500 16256 6556
rect 16192 6496 16256 6500
rect 25952 6556 26016 6560
rect 25952 6500 25956 6556
rect 25956 6500 26012 6556
rect 26012 6500 26016 6556
rect 25952 6496 26016 6500
rect 26032 6556 26096 6560
rect 26032 6500 26036 6556
rect 26036 6500 26092 6556
rect 26092 6500 26096 6556
rect 26032 6496 26096 6500
rect 26112 6556 26176 6560
rect 26112 6500 26116 6556
rect 26116 6500 26172 6556
rect 26172 6500 26176 6556
rect 26112 6496 26176 6500
rect 26192 6556 26256 6560
rect 26192 6500 26196 6556
rect 26196 6500 26252 6556
rect 26252 6500 26256 6556
rect 26192 6496 26256 6500
rect 10952 6012 11016 6016
rect 10952 5956 10956 6012
rect 10956 5956 11012 6012
rect 11012 5956 11016 6012
rect 10952 5952 11016 5956
rect 11032 6012 11096 6016
rect 11032 5956 11036 6012
rect 11036 5956 11092 6012
rect 11092 5956 11096 6012
rect 11032 5952 11096 5956
rect 11112 6012 11176 6016
rect 11112 5956 11116 6012
rect 11116 5956 11172 6012
rect 11172 5956 11176 6012
rect 11112 5952 11176 5956
rect 11192 6012 11256 6016
rect 11192 5956 11196 6012
rect 11196 5956 11252 6012
rect 11252 5956 11256 6012
rect 11192 5952 11256 5956
rect 20952 6012 21016 6016
rect 20952 5956 20956 6012
rect 20956 5956 21012 6012
rect 21012 5956 21016 6012
rect 20952 5952 21016 5956
rect 21032 6012 21096 6016
rect 21032 5956 21036 6012
rect 21036 5956 21092 6012
rect 21092 5956 21096 6012
rect 21032 5952 21096 5956
rect 21112 6012 21176 6016
rect 21112 5956 21116 6012
rect 21116 5956 21172 6012
rect 21172 5956 21176 6012
rect 21112 5952 21176 5956
rect 21192 6012 21256 6016
rect 21192 5956 21196 6012
rect 21196 5956 21252 6012
rect 21252 5956 21256 6012
rect 21192 5952 21256 5956
rect 5952 5468 6016 5472
rect 5952 5412 5956 5468
rect 5956 5412 6012 5468
rect 6012 5412 6016 5468
rect 5952 5408 6016 5412
rect 6032 5468 6096 5472
rect 6032 5412 6036 5468
rect 6036 5412 6092 5468
rect 6092 5412 6096 5468
rect 6032 5408 6096 5412
rect 6112 5468 6176 5472
rect 6112 5412 6116 5468
rect 6116 5412 6172 5468
rect 6172 5412 6176 5468
rect 6112 5408 6176 5412
rect 6192 5468 6256 5472
rect 6192 5412 6196 5468
rect 6196 5412 6252 5468
rect 6252 5412 6256 5468
rect 6192 5408 6256 5412
rect 15952 5468 16016 5472
rect 15952 5412 15956 5468
rect 15956 5412 16012 5468
rect 16012 5412 16016 5468
rect 15952 5408 16016 5412
rect 16032 5468 16096 5472
rect 16032 5412 16036 5468
rect 16036 5412 16092 5468
rect 16092 5412 16096 5468
rect 16032 5408 16096 5412
rect 16112 5468 16176 5472
rect 16112 5412 16116 5468
rect 16116 5412 16172 5468
rect 16172 5412 16176 5468
rect 16112 5408 16176 5412
rect 16192 5468 16256 5472
rect 16192 5412 16196 5468
rect 16196 5412 16252 5468
rect 16252 5412 16256 5468
rect 16192 5408 16256 5412
rect 25952 5468 26016 5472
rect 25952 5412 25956 5468
rect 25956 5412 26012 5468
rect 26012 5412 26016 5468
rect 25952 5408 26016 5412
rect 26032 5468 26096 5472
rect 26032 5412 26036 5468
rect 26036 5412 26092 5468
rect 26092 5412 26096 5468
rect 26032 5408 26096 5412
rect 26112 5468 26176 5472
rect 26112 5412 26116 5468
rect 26116 5412 26172 5468
rect 26172 5412 26176 5468
rect 26112 5408 26176 5412
rect 26192 5468 26256 5472
rect 26192 5412 26196 5468
rect 26196 5412 26252 5468
rect 26252 5412 26256 5468
rect 26192 5408 26256 5412
rect 10952 4924 11016 4928
rect 10952 4868 10956 4924
rect 10956 4868 11012 4924
rect 11012 4868 11016 4924
rect 10952 4864 11016 4868
rect 11032 4924 11096 4928
rect 11032 4868 11036 4924
rect 11036 4868 11092 4924
rect 11092 4868 11096 4924
rect 11032 4864 11096 4868
rect 11112 4924 11176 4928
rect 11112 4868 11116 4924
rect 11116 4868 11172 4924
rect 11172 4868 11176 4924
rect 11112 4864 11176 4868
rect 11192 4924 11256 4928
rect 11192 4868 11196 4924
rect 11196 4868 11252 4924
rect 11252 4868 11256 4924
rect 11192 4864 11256 4868
rect 20952 4924 21016 4928
rect 20952 4868 20956 4924
rect 20956 4868 21012 4924
rect 21012 4868 21016 4924
rect 20952 4864 21016 4868
rect 21032 4924 21096 4928
rect 21032 4868 21036 4924
rect 21036 4868 21092 4924
rect 21092 4868 21096 4924
rect 21032 4864 21096 4868
rect 21112 4924 21176 4928
rect 21112 4868 21116 4924
rect 21116 4868 21172 4924
rect 21172 4868 21176 4924
rect 21112 4864 21176 4868
rect 21192 4924 21256 4928
rect 21192 4868 21196 4924
rect 21196 4868 21252 4924
rect 21252 4868 21256 4924
rect 21192 4864 21256 4868
rect 5952 4380 6016 4384
rect 5952 4324 5956 4380
rect 5956 4324 6012 4380
rect 6012 4324 6016 4380
rect 5952 4320 6016 4324
rect 6032 4380 6096 4384
rect 6032 4324 6036 4380
rect 6036 4324 6092 4380
rect 6092 4324 6096 4380
rect 6032 4320 6096 4324
rect 6112 4380 6176 4384
rect 6112 4324 6116 4380
rect 6116 4324 6172 4380
rect 6172 4324 6176 4380
rect 6112 4320 6176 4324
rect 6192 4380 6256 4384
rect 6192 4324 6196 4380
rect 6196 4324 6252 4380
rect 6252 4324 6256 4380
rect 6192 4320 6256 4324
rect 15952 4380 16016 4384
rect 15952 4324 15956 4380
rect 15956 4324 16012 4380
rect 16012 4324 16016 4380
rect 15952 4320 16016 4324
rect 16032 4380 16096 4384
rect 16032 4324 16036 4380
rect 16036 4324 16092 4380
rect 16092 4324 16096 4380
rect 16032 4320 16096 4324
rect 16112 4380 16176 4384
rect 16112 4324 16116 4380
rect 16116 4324 16172 4380
rect 16172 4324 16176 4380
rect 16112 4320 16176 4324
rect 16192 4380 16256 4384
rect 16192 4324 16196 4380
rect 16196 4324 16252 4380
rect 16252 4324 16256 4380
rect 16192 4320 16256 4324
rect 25952 4380 26016 4384
rect 25952 4324 25956 4380
rect 25956 4324 26012 4380
rect 26012 4324 26016 4380
rect 25952 4320 26016 4324
rect 26032 4380 26096 4384
rect 26032 4324 26036 4380
rect 26036 4324 26092 4380
rect 26092 4324 26096 4380
rect 26032 4320 26096 4324
rect 26112 4380 26176 4384
rect 26112 4324 26116 4380
rect 26116 4324 26172 4380
rect 26172 4324 26176 4380
rect 26112 4320 26176 4324
rect 26192 4380 26256 4384
rect 26192 4324 26196 4380
rect 26196 4324 26252 4380
rect 26252 4324 26256 4380
rect 26192 4320 26256 4324
rect 10952 3836 11016 3840
rect 10952 3780 10956 3836
rect 10956 3780 11012 3836
rect 11012 3780 11016 3836
rect 10952 3776 11016 3780
rect 11032 3836 11096 3840
rect 11032 3780 11036 3836
rect 11036 3780 11092 3836
rect 11092 3780 11096 3836
rect 11032 3776 11096 3780
rect 11112 3836 11176 3840
rect 11112 3780 11116 3836
rect 11116 3780 11172 3836
rect 11172 3780 11176 3836
rect 11112 3776 11176 3780
rect 11192 3836 11256 3840
rect 11192 3780 11196 3836
rect 11196 3780 11252 3836
rect 11252 3780 11256 3836
rect 11192 3776 11256 3780
rect 20952 3836 21016 3840
rect 20952 3780 20956 3836
rect 20956 3780 21012 3836
rect 21012 3780 21016 3836
rect 20952 3776 21016 3780
rect 21032 3836 21096 3840
rect 21032 3780 21036 3836
rect 21036 3780 21092 3836
rect 21092 3780 21096 3836
rect 21032 3776 21096 3780
rect 21112 3836 21176 3840
rect 21112 3780 21116 3836
rect 21116 3780 21172 3836
rect 21172 3780 21176 3836
rect 21112 3776 21176 3780
rect 21192 3836 21256 3840
rect 21192 3780 21196 3836
rect 21196 3780 21252 3836
rect 21252 3780 21256 3836
rect 21192 3776 21256 3780
rect 5952 3292 6016 3296
rect 5952 3236 5956 3292
rect 5956 3236 6012 3292
rect 6012 3236 6016 3292
rect 5952 3232 6016 3236
rect 6032 3292 6096 3296
rect 6032 3236 6036 3292
rect 6036 3236 6092 3292
rect 6092 3236 6096 3292
rect 6032 3232 6096 3236
rect 6112 3292 6176 3296
rect 6112 3236 6116 3292
rect 6116 3236 6172 3292
rect 6172 3236 6176 3292
rect 6112 3232 6176 3236
rect 6192 3292 6256 3296
rect 6192 3236 6196 3292
rect 6196 3236 6252 3292
rect 6252 3236 6256 3292
rect 6192 3232 6256 3236
rect 15952 3292 16016 3296
rect 15952 3236 15956 3292
rect 15956 3236 16012 3292
rect 16012 3236 16016 3292
rect 15952 3232 16016 3236
rect 16032 3292 16096 3296
rect 16032 3236 16036 3292
rect 16036 3236 16092 3292
rect 16092 3236 16096 3292
rect 16032 3232 16096 3236
rect 16112 3292 16176 3296
rect 16112 3236 16116 3292
rect 16116 3236 16172 3292
rect 16172 3236 16176 3292
rect 16112 3232 16176 3236
rect 16192 3292 16256 3296
rect 16192 3236 16196 3292
rect 16196 3236 16252 3292
rect 16252 3236 16256 3292
rect 16192 3232 16256 3236
rect 25952 3292 26016 3296
rect 25952 3236 25956 3292
rect 25956 3236 26012 3292
rect 26012 3236 26016 3292
rect 25952 3232 26016 3236
rect 26032 3292 26096 3296
rect 26032 3236 26036 3292
rect 26036 3236 26092 3292
rect 26092 3236 26096 3292
rect 26032 3232 26096 3236
rect 26112 3292 26176 3296
rect 26112 3236 26116 3292
rect 26116 3236 26172 3292
rect 26172 3236 26176 3292
rect 26112 3232 26176 3236
rect 26192 3292 26256 3296
rect 26192 3236 26196 3292
rect 26196 3236 26252 3292
rect 26252 3236 26256 3292
rect 26192 3232 26256 3236
rect 10952 2748 11016 2752
rect 10952 2692 10956 2748
rect 10956 2692 11012 2748
rect 11012 2692 11016 2748
rect 10952 2688 11016 2692
rect 11032 2748 11096 2752
rect 11032 2692 11036 2748
rect 11036 2692 11092 2748
rect 11092 2692 11096 2748
rect 11032 2688 11096 2692
rect 11112 2748 11176 2752
rect 11112 2692 11116 2748
rect 11116 2692 11172 2748
rect 11172 2692 11176 2748
rect 11112 2688 11176 2692
rect 11192 2748 11256 2752
rect 11192 2692 11196 2748
rect 11196 2692 11252 2748
rect 11252 2692 11256 2748
rect 11192 2688 11256 2692
rect 20952 2748 21016 2752
rect 20952 2692 20956 2748
rect 20956 2692 21012 2748
rect 21012 2692 21016 2748
rect 20952 2688 21016 2692
rect 21032 2748 21096 2752
rect 21032 2692 21036 2748
rect 21036 2692 21092 2748
rect 21092 2692 21096 2748
rect 21032 2688 21096 2692
rect 21112 2748 21176 2752
rect 21112 2692 21116 2748
rect 21116 2692 21172 2748
rect 21172 2692 21176 2748
rect 21112 2688 21176 2692
rect 21192 2748 21256 2752
rect 21192 2692 21196 2748
rect 21196 2692 21252 2748
rect 21252 2692 21256 2748
rect 21192 2688 21256 2692
rect 5952 2204 6016 2208
rect 5952 2148 5956 2204
rect 5956 2148 6012 2204
rect 6012 2148 6016 2204
rect 5952 2144 6016 2148
rect 6032 2204 6096 2208
rect 6032 2148 6036 2204
rect 6036 2148 6092 2204
rect 6092 2148 6096 2204
rect 6032 2144 6096 2148
rect 6112 2204 6176 2208
rect 6112 2148 6116 2204
rect 6116 2148 6172 2204
rect 6172 2148 6176 2204
rect 6112 2144 6176 2148
rect 6192 2204 6256 2208
rect 6192 2148 6196 2204
rect 6196 2148 6252 2204
rect 6252 2148 6256 2204
rect 6192 2144 6256 2148
rect 15952 2204 16016 2208
rect 15952 2148 15956 2204
rect 15956 2148 16012 2204
rect 16012 2148 16016 2204
rect 15952 2144 16016 2148
rect 16032 2204 16096 2208
rect 16032 2148 16036 2204
rect 16036 2148 16092 2204
rect 16092 2148 16096 2204
rect 16032 2144 16096 2148
rect 16112 2204 16176 2208
rect 16112 2148 16116 2204
rect 16116 2148 16172 2204
rect 16172 2148 16176 2204
rect 16112 2144 16176 2148
rect 16192 2204 16256 2208
rect 16192 2148 16196 2204
rect 16196 2148 16252 2204
rect 16252 2148 16256 2204
rect 16192 2144 16256 2148
rect 25952 2204 26016 2208
rect 25952 2148 25956 2204
rect 25956 2148 26012 2204
rect 26012 2148 26016 2204
rect 25952 2144 26016 2148
rect 26032 2204 26096 2208
rect 26032 2148 26036 2204
rect 26036 2148 26092 2204
rect 26092 2148 26096 2204
rect 26032 2144 26096 2148
rect 26112 2204 26176 2208
rect 26112 2148 26116 2204
rect 26116 2148 26172 2204
rect 26172 2148 26176 2204
rect 26112 2144 26176 2148
rect 26192 2204 26256 2208
rect 26192 2148 26196 2204
rect 26196 2148 26252 2204
rect 26252 2148 26256 2204
rect 26192 2144 26256 2148
<< metal4 >>
rect 5944 21792 6264 21808
rect 5944 21728 5952 21792
rect 6016 21728 6032 21792
rect 6096 21728 6112 21792
rect 6176 21728 6192 21792
rect 6256 21728 6264 21792
rect 5944 20704 6264 21728
rect 5944 20640 5952 20704
rect 6016 20640 6032 20704
rect 6096 20640 6112 20704
rect 6176 20640 6192 20704
rect 6256 20640 6264 20704
rect 5944 19616 6264 20640
rect 5944 19552 5952 19616
rect 6016 19552 6032 19616
rect 6096 19552 6112 19616
rect 6176 19552 6192 19616
rect 6256 19552 6264 19616
rect 5944 18528 6264 19552
rect 5944 18464 5952 18528
rect 6016 18464 6032 18528
rect 6096 18464 6112 18528
rect 6176 18464 6192 18528
rect 6256 18464 6264 18528
rect 5944 17440 6264 18464
rect 5944 17376 5952 17440
rect 6016 17376 6032 17440
rect 6096 17376 6112 17440
rect 6176 17376 6192 17440
rect 6256 17376 6264 17440
rect 5944 16352 6264 17376
rect 5944 16288 5952 16352
rect 6016 16288 6032 16352
rect 6096 16288 6112 16352
rect 6176 16288 6192 16352
rect 6256 16288 6264 16352
rect 5944 15264 6264 16288
rect 5944 15200 5952 15264
rect 6016 15200 6032 15264
rect 6096 15200 6112 15264
rect 6176 15200 6192 15264
rect 6256 15200 6264 15264
rect 5944 14176 6264 15200
rect 5944 14112 5952 14176
rect 6016 14112 6032 14176
rect 6096 14112 6112 14176
rect 6176 14112 6192 14176
rect 6256 14112 6264 14176
rect 5944 13088 6264 14112
rect 5944 13024 5952 13088
rect 6016 13024 6032 13088
rect 6096 13024 6112 13088
rect 6176 13024 6192 13088
rect 6256 13024 6264 13088
rect 5944 12000 6264 13024
rect 5944 11936 5952 12000
rect 6016 11936 6032 12000
rect 6096 11936 6112 12000
rect 6176 11936 6192 12000
rect 6256 11936 6264 12000
rect 5944 10912 6264 11936
rect 5944 10848 5952 10912
rect 6016 10848 6032 10912
rect 6096 10848 6112 10912
rect 6176 10848 6192 10912
rect 6256 10848 6264 10912
rect 5944 9824 6264 10848
rect 5944 9760 5952 9824
rect 6016 9760 6032 9824
rect 6096 9760 6112 9824
rect 6176 9760 6192 9824
rect 6256 9760 6264 9824
rect 5944 8736 6264 9760
rect 5944 8672 5952 8736
rect 6016 8672 6032 8736
rect 6096 8672 6112 8736
rect 6176 8672 6192 8736
rect 6256 8672 6264 8736
rect 5944 7648 6264 8672
rect 10944 21248 11264 21808
rect 10944 21184 10952 21248
rect 11016 21184 11032 21248
rect 11096 21184 11112 21248
rect 11176 21184 11192 21248
rect 11256 21184 11264 21248
rect 10944 20160 11264 21184
rect 10944 20096 10952 20160
rect 11016 20096 11032 20160
rect 11096 20096 11112 20160
rect 11176 20096 11192 20160
rect 11256 20096 11264 20160
rect 10944 19072 11264 20096
rect 10944 19008 10952 19072
rect 11016 19008 11032 19072
rect 11096 19008 11112 19072
rect 11176 19008 11192 19072
rect 11256 19008 11264 19072
rect 10944 17984 11264 19008
rect 10944 17920 10952 17984
rect 11016 17920 11032 17984
rect 11096 17920 11112 17984
rect 11176 17920 11192 17984
rect 11256 17920 11264 17984
rect 10944 16896 11264 17920
rect 10944 16832 10952 16896
rect 11016 16832 11032 16896
rect 11096 16832 11112 16896
rect 11176 16832 11192 16896
rect 11256 16832 11264 16896
rect 10944 15808 11264 16832
rect 10944 15744 10952 15808
rect 11016 15744 11032 15808
rect 11096 15744 11112 15808
rect 11176 15744 11192 15808
rect 11256 15744 11264 15808
rect 10944 14720 11264 15744
rect 10944 14656 10952 14720
rect 11016 14656 11032 14720
rect 11096 14656 11112 14720
rect 11176 14656 11192 14720
rect 11256 14656 11264 14720
rect 10944 13632 11264 14656
rect 10944 13568 10952 13632
rect 11016 13568 11032 13632
rect 11096 13568 11112 13632
rect 11176 13568 11192 13632
rect 11256 13568 11264 13632
rect 10944 12544 11264 13568
rect 10944 12480 10952 12544
rect 11016 12480 11032 12544
rect 11096 12480 11112 12544
rect 11176 12480 11192 12544
rect 11256 12480 11264 12544
rect 10944 11456 11264 12480
rect 10944 11392 10952 11456
rect 11016 11392 11032 11456
rect 11096 11392 11112 11456
rect 11176 11392 11192 11456
rect 11256 11392 11264 11456
rect 10944 10368 11264 11392
rect 10944 10304 10952 10368
rect 11016 10304 11032 10368
rect 11096 10304 11112 10368
rect 11176 10304 11192 10368
rect 11256 10304 11264 10368
rect 10944 9280 11264 10304
rect 10944 9216 10952 9280
rect 11016 9216 11032 9280
rect 11096 9216 11112 9280
rect 11176 9216 11192 9280
rect 11256 9216 11264 9280
rect 5944 7584 5952 7648
rect 6016 7584 6032 7648
rect 6096 7584 6112 7648
rect 6176 7584 6192 7648
rect 6256 7584 6264 7648
rect 5944 6560 6264 7584
rect 5944 6496 5952 6560
rect 6016 6496 6032 6560
rect 6096 6496 6112 6560
rect 6176 6496 6192 6560
rect 6256 6496 6264 6560
rect 5944 5472 6264 6496
rect 5944 5408 5952 5472
rect 6016 5408 6032 5472
rect 6096 5408 6112 5472
rect 6176 5408 6192 5472
rect 6256 5408 6264 5472
rect 5944 4384 6264 5408
rect 5944 4320 5952 4384
rect 6016 4320 6032 4384
rect 6096 4320 6112 4384
rect 6176 4320 6192 4384
rect 6256 4320 6264 4384
rect 5944 3296 6264 4320
rect 5944 3232 5952 3296
rect 6016 3232 6032 3296
rect 6096 3232 6112 3296
rect 6176 3232 6192 3296
rect 6256 3232 6264 3296
rect 5944 2208 6264 3232
rect 5944 2144 5952 2208
rect 6016 2144 6032 2208
rect 6096 2144 6112 2208
rect 6176 2144 6192 2208
rect 6256 2144 6264 2208
rect 5944 2128 6264 2144
rect 10944 8192 11264 9216
rect 10944 8128 10952 8192
rect 11016 8128 11032 8192
rect 11096 8128 11112 8192
rect 11176 8128 11192 8192
rect 11256 8128 11264 8192
rect 10944 7104 11264 8128
rect 10944 7040 10952 7104
rect 11016 7040 11032 7104
rect 11096 7040 11112 7104
rect 11176 7040 11192 7104
rect 11256 7040 11264 7104
rect 10944 6016 11264 7040
rect 10944 5952 10952 6016
rect 11016 5952 11032 6016
rect 11096 5952 11112 6016
rect 11176 5952 11192 6016
rect 11256 5952 11264 6016
rect 10944 4928 11264 5952
rect 10944 4864 10952 4928
rect 11016 4864 11032 4928
rect 11096 4864 11112 4928
rect 11176 4864 11192 4928
rect 11256 4864 11264 4928
rect 10944 3840 11264 4864
rect 10944 3776 10952 3840
rect 11016 3776 11032 3840
rect 11096 3776 11112 3840
rect 11176 3776 11192 3840
rect 11256 3776 11264 3840
rect 10944 2752 11264 3776
rect 10944 2688 10952 2752
rect 11016 2688 11032 2752
rect 11096 2688 11112 2752
rect 11176 2688 11192 2752
rect 11256 2688 11264 2752
rect 10944 2128 11264 2688
rect 15944 21792 16264 21808
rect 15944 21728 15952 21792
rect 16016 21728 16032 21792
rect 16096 21728 16112 21792
rect 16176 21728 16192 21792
rect 16256 21728 16264 21792
rect 15944 20704 16264 21728
rect 15944 20640 15952 20704
rect 16016 20640 16032 20704
rect 16096 20640 16112 20704
rect 16176 20640 16192 20704
rect 16256 20640 16264 20704
rect 15944 19616 16264 20640
rect 15944 19552 15952 19616
rect 16016 19552 16032 19616
rect 16096 19552 16112 19616
rect 16176 19552 16192 19616
rect 16256 19552 16264 19616
rect 15944 18528 16264 19552
rect 15944 18464 15952 18528
rect 16016 18464 16032 18528
rect 16096 18464 16112 18528
rect 16176 18464 16192 18528
rect 16256 18464 16264 18528
rect 15944 17440 16264 18464
rect 15944 17376 15952 17440
rect 16016 17376 16032 17440
rect 16096 17376 16112 17440
rect 16176 17376 16192 17440
rect 16256 17376 16264 17440
rect 15944 16352 16264 17376
rect 15944 16288 15952 16352
rect 16016 16288 16032 16352
rect 16096 16288 16112 16352
rect 16176 16288 16192 16352
rect 16256 16288 16264 16352
rect 15944 15264 16264 16288
rect 15944 15200 15952 15264
rect 16016 15200 16032 15264
rect 16096 15200 16112 15264
rect 16176 15200 16192 15264
rect 16256 15200 16264 15264
rect 15944 14176 16264 15200
rect 15944 14112 15952 14176
rect 16016 14112 16032 14176
rect 16096 14112 16112 14176
rect 16176 14112 16192 14176
rect 16256 14112 16264 14176
rect 15944 13088 16264 14112
rect 15944 13024 15952 13088
rect 16016 13024 16032 13088
rect 16096 13024 16112 13088
rect 16176 13024 16192 13088
rect 16256 13024 16264 13088
rect 15944 12000 16264 13024
rect 15944 11936 15952 12000
rect 16016 11936 16032 12000
rect 16096 11936 16112 12000
rect 16176 11936 16192 12000
rect 16256 11936 16264 12000
rect 15944 10912 16264 11936
rect 15944 10848 15952 10912
rect 16016 10848 16032 10912
rect 16096 10848 16112 10912
rect 16176 10848 16192 10912
rect 16256 10848 16264 10912
rect 15944 9824 16264 10848
rect 15944 9760 15952 9824
rect 16016 9760 16032 9824
rect 16096 9760 16112 9824
rect 16176 9760 16192 9824
rect 16256 9760 16264 9824
rect 15944 8736 16264 9760
rect 15944 8672 15952 8736
rect 16016 8672 16032 8736
rect 16096 8672 16112 8736
rect 16176 8672 16192 8736
rect 16256 8672 16264 8736
rect 15944 7648 16264 8672
rect 15944 7584 15952 7648
rect 16016 7584 16032 7648
rect 16096 7584 16112 7648
rect 16176 7584 16192 7648
rect 16256 7584 16264 7648
rect 15944 6560 16264 7584
rect 15944 6496 15952 6560
rect 16016 6496 16032 6560
rect 16096 6496 16112 6560
rect 16176 6496 16192 6560
rect 16256 6496 16264 6560
rect 15944 5472 16264 6496
rect 15944 5408 15952 5472
rect 16016 5408 16032 5472
rect 16096 5408 16112 5472
rect 16176 5408 16192 5472
rect 16256 5408 16264 5472
rect 15944 4384 16264 5408
rect 15944 4320 15952 4384
rect 16016 4320 16032 4384
rect 16096 4320 16112 4384
rect 16176 4320 16192 4384
rect 16256 4320 16264 4384
rect 15944 3296 16264 4320
rect 15944 3232 15952 3296
rect 16016 3232 16032 3296
rect 16096 3232 16112 3296
rect 16176 3232 16192 3296
rect 16256 3232 16264 3296
rect 15944 2208 16264 3232
rect 15944 2144 15952 2208
rect 16016 2144 16032 2208
rect 16096 2144 16112 2208
rect 16176 2144 16192 2208
rect 16256 2144 16264 2208
rect 15944 2128 16264 2144
rect 20944 21248 21264 21808
rect 20944 21184 20952 21248
rect 21016 21184 21032 21248
rect 21096 21184 21112 21248
rect 21176 21184 21192 21248
rect 21256 21184 21264 21248
rect 20944 20160 21264 21184
rect 20944 20096 20952 20160
rect 21016 20096 21032 20160
rect 21096 20096 21112 20160
rect 21176 20096 21192 20160
rect 21256 20096 21264 20160
rect 20944 19072 21264 20096
rect 20944 19008 20952 19072
rect 21016 19008 21032 19072
rect 21096 19008 21112 19072
rect 21176 19008 21192 19072
rect 21256 19008 21264 19072
rect 20944 17984 21264 19008
rect 20944 17920 20952 17984
rect 21016 17920 21032 17984
rect 21096 17920 21112 17984
rect 21176 17920 21192 17984
rect 21256 17920 21264 17984
rect 20944 16896 21264 17920
rect 20944 16832 20952 16896
rect 21016 16832 21032 16896
rect 21096 16832 21112 16896
rect 21176 16832 21192 16896
rect 21256 16832 21264 16896
rect 20944 15808 21264 16832
rect 20944 15744 20952 15808
rect 21016 15744 21032 15808
rect 21096 15744 21112 15808
rect 21176 15744 21192 15808
rect 21256 15744 21264 15808
rect 20944 14720 21264 15744
rect 20944 14656 20952 14720
rect 21016 14656 21032 14720
rect 21096 14656 21112 14720
rect 21176 14656 21192 14720
rect 21256 14656 21264 14720
rect 20944 13632 21264 14656
rect 20944 13568 20952 13632
rect 21016 13568 21032 13632
rect 21096 13568 21112 13632
rect 21176 13568 21192 13632
rect 21256 13568 21264 13632
rect 20944 12544 21264 13568
rect 20944 12480 20952 12544
rect 21016 12480 21032 12544
rect 21096 12480 21112 12544
rect 21176 12480 21192 12544
rect 21256 12480 21264 12544
rect 20944 11456 21264 12480
rect 20944 11392 20952 11456
rect 21016 11392 21032 11456
rect 21096 11392 21112 11456
rect 21176 11392 21192 11456
rect 21256 11392 21264 11456
rect 20944 10368 21264 11392
rect 20944 10304 20952 10368
rect 21016 10304 21032 10368
rect 21096 10304 21112 10368
rect 21176 10304 21192 10368
rect 21256 10304 21264 10368
rect 20944 9280 21264 10304
rect 20944 9216 20952 9280
rect 21016 9216 21032 9280
rect 21096 9216 21112 9280
rect 21176 9216 21192 9280
rect 21256 9216 21264 9280
rect 20944 8192 21264 9216
rect 20944 8128 20952 8192
rect 21016 8128 21032 8192
rect 21096 8128 21112 8192
rect 21176 8128 21192 8192
rect 21256 8128 21264 8192
rect 20944 7104 21264 8128
rect 20944 7040 20952 7104
rect 21016 7040 21032 7104
rect 21096 7040 21112 7104
rect 21176 7040 21192 7104
rect 21256 7040 21264 7104
rect 20944 6016 21264 7040
rect 20944 5952 20952 6016
rect 21016 5952 21032 6016
rect 21096 5952 21112 6016
rect 21176 5952 21192 6016
rect 21256 5952 21264 6016
rect 20944 4928 21264 5952
rect 20944 4864 20952 4928
rect 21016 4864 21032 4928
rect 21096 4864 21112 4928
rect 21176 4864 21192 4928
rect 21256 4864 21264 4928
rect 20944 3840 21264 4864
rect 20944 3776 20952 3840
rect 21016 3776 21032 3840
rect 21096 3776 21112 3840
rect 21176 3776 21192 3840
rect 21256 3776 21264 3840
rect 20944 2752 21264 3776
rect 20944 2688 20952 2752
rect 21016 2688 21032 2752
rect 21096 2688 21112 2752
rect 21176 2688 21192 2752
rect 21256 2688 21264 2752
rect 20944 2128 21264 2688
rect 25944 21792 26264 21808
rect 25944 21728 25952 21792
rect 26016 21728 26032 21792
rect 26096 21728 26112 21792
rect 26176 21728 26192 21792
rect 26256 21728 26264 21792
rect 25944 20704 26264 21728
rect 25944 20640 25952 20704
rect 26016 20640 26032 20704
rect 26096 20640 26112 20704
rect 26176 20640 26192 20704
rect 26256 20640 26264 20704
rect 25944 19616 26264 20640
rect 25944 19552 25952 19616
rect 26016 19552 26032 19616
rect 26096 19552 26112 19616
rect 26176 19552 26192 19616
rect 26256 19552 26264 19616
rect 25944 18528 26264 19552
rect 25944 18464 25952 18528
rect 26016 18464 26032 18528
rect 26096 18464 26112 18528
rect 26176 18464 26192 18528
rect 26256 18464 26264 18528
rect 25944 17440 26264 18464
rect 25944 17376 25952 17440
rect 26016 17376 26032 17440
rect 26096 17376 26112 17440
rect 26176 17376 26192 17440
rect 26256 17376 26264 17440
rect 25944 16352 26264 17376
rect 25944 16288 25952 16352
rect 26016 16288 26032 16352
rect 26096 16288 26112 16352
rect 26176 16288 26192 16352
rect 26256 16288 26264 16352
rect 25944 15264 26264 16288
rect 25944 15200 25952 15264
rect 26016 15200 26032 15264
rect 26096 15200 26112 15264
rect 26176 15200 26192 15264
rect 26256 15200 26264 15264
rect 25944 14176 26264 15200
rect 25944 14112 25952 14176
rect 26016 14112 26032 14176
rect 26096 14112 26112 14176
rect 26176 14112 26192 14176
rect 26256 14112 26264 14176
rect 25944 13088 26264 14112
rect 25944 13024 25952 13088
rect 26016 13024 26032 13088
rect 26096 13024 26112 13088
rect 26176 13024 26192 13088
rect 26256 13024 26264 13088
rect 25944 12000 26264 13024
rect 25944 11936 25952 12000
rect 26016 11936 26032 12000
rect 26096 11936 26112 12000
rect 26176 11936 26192 12000
rect 26256 11936 26264 12000
rect 25944 10912 26264 11936
rect 25944 10848 25952 10912
rect 26016 10848 26032 10912
rect 26096 10848 26112 10912
rect 26176 10848 26192 10912
rect 26256 10848 26264 10912
rect 25944 9824 26264 10848
rect 25944 9760 25952 9824
rect 26016 9760 26032 9824
rect 26096 9760 26112 9824
rect 26176 9760 26192 9824
rect 26256 9760 26264 9824
rect 25944 8736 26264 9760
rect 26555 8940 26621 8941
rect 26555 8876 26556 8940
rect 26620 8876 26621 8940
rect 26555 8875 26621 8876
rect 25944 8672 25952 8736
rect 26016 8672 26032 8736
rect 26096 8672 26112 8736
rect 26176 8672 26192 8736
rect 26256 8672 26264 8736
rect 25944 7648 26264 8672
rect 26558 8618 26618 8875
rect 25944 7584 25952 7648
rect 26016 7584 26032 7648
rect 26096 7584 26112 7648
rect 26176 7584 26192 7648
rect 26256 7584 26264 7648
rect 25944 6560 26264 7584
rect 25944 6496 25952 6560
rect 26016 6496 26032 6560
rect 26096 6496 26112 6560
rect 26176 6496 26192 6560
rect 26256 6496 26264 6560
rect 25944 5472 26264 6496
rect 25944 5408 25952 5472
rect 26016 5408 26032 5472
rect 26096 5408 26112 5472
rect 26176 5408 26192 5472
rect 26256 5408 26264 5472
rect 25944 4384 26264 5408
rect 25944 4320 25952 4384
rect 26016 4320 26032 4384
rect 26096 4320 26112 4384
rect 26176 4320 26192 4384
rect 26256 4320 26264 4384
rect 25944 3296 26264 4320
rect 25944 3232 25952 3296
rect 26016 3232 26032 3296
rect 26096 3232 26112 3296
rect 26176 3232 26192 3296
rect 26256 3232 26264 3296
rect 25944 2208 26264 3232
rect 25944 2144 25952 2208
rect 26016 2144 26032 2208
rect 26096 2144 26112 2208
rect 26176 2144 26192 2208
rect 26256 2144 26264 2208
rect 25944 2128 26264 2144
<< via4 >>
rect 7150 8532 7386 8618
rect 7150 8468 7236 8532
rect 7236 8468 7300 8532
rect 7300 8468 7386 8532
rect 7150 8382 7386 8468
rect 26470 8382 26706 8618
<< metal5 >>
rect 7108 8618 26748 8660
rect 7108 8382 7150 8618
rect 7386 8382 26470 8618
rect 26706 8382 26748 8618
rect 7108 8340 26748 8382
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _15_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_11 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2116 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_7 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1748 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13
timestamp 1604681595
transform 1 0 2300 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9
timestamp 1604681595
transform 1 0 1932 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0__A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2116 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__15__A
timestamp 1604681595
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_17 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2668 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__16__A
timestamp 1604681595
transform 1 0 2484 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2668 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_23 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3220 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27
timestamp 1604681595
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23
timestamp 1604681595
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 3312 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_34
timestamp 1604681595
transform 1 0 4232 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_30
timestamp 1604681595
transform 1 0 3864 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 4048 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38
timestamp 1604681595
transform 1 0 4600 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 4784 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__18__A
timestamp 1604681595
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _18_
timestamp 1604681595
transform 1 0 4600 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_52 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5888 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_48
timestamp 1604681595
transform 1 0 5520 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_42
timestamp 1604681595
transform 1 0 4968 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 5704 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 5336 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_62
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_60
timestamp 1604681595
transform 1 0 6624 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58
timestamp 1604681595
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1604681595
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_mode_io__5.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_mode_io__5.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_42 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4968 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_mode_io__0.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 7268 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  ltile_mode_io__5.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_mode_io__0.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 7084 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_82
timestamp 1604681595
transform 1 0 8648 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_90
timestamp 1604681595
transform 1 0 9384 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_86
timestamp 1604681595
transform 1 0 9016 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89
timestamp 1604681595
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86
timestamp 1604681595
transform 1 0 9016 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_mode_io__2.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9568 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_mode_io__1.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1604681595
transform 1 0 9200 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_mode_io__1.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_102
timestamp 1604681595
transform 1 0 10488 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_94
timestamp 1604681595
transform 1 0 9752 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1604681595
transform 1 0 10672 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_mode_io__2.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9936 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1604681595
transform 1 0 10120 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_mode_io__1.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_1_114
timestamp 1604681595
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_106
timestamp 1604681595
transform 1 0 10856 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113
timestamp 1604681595
transform 1 0 11500 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1604681595
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1604681595
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_mode_io__4.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117
timestamp 1604681595
transform 1 0 11868 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_118
timestamp 1604681595
transform 1 0 11960 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_mode_io__4.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120
timestamp 1604681595
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_123
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_mode_io__3.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12604 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_mode_io__4.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1604681595
transform 1 0 13156 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1604681595
transform 1 0 14260 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1604681595
transform 1 0 13708 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_mode_io__3.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 12972 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_144
timestamp 1604681595
transform 1 0 14352 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_127
timestamp 1604681595
transform 1 0 12788 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_135
timestamp 1604681595
transform 1 0 13524 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_139
timestamp 1604681595
transform 1 0 13892 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_147
timestamp 1604681595
transform 1 0 14628 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_152
timestamp 1604681595
transform 1 0 15088 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1604681595
transform 1 0 14812 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_164
timestamp 1604681595
transform 1 0 16192 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_160
timestamp 1604681595
transform 1 0 15824 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1604681595
transform 1 0 16008 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_163
timestamp 1604681595
transform 1 0 16100 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_151
timestamp 1604681595
transform 1 0 14996 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1604681595
transform 1 0 16744 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1604681595
transform 1 0 17296 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_174
timestamp 1604681595
transform 1 0 17112 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_178
timestamp 1604681595
transform 1 0 17480 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_187
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_175
timestamp 1604681595
transform 1 0 17204 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_184
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1604681595
transform 1 0 19044 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1604681595
transform 1 0 19044 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1604681595
transform 1 0 19596 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1604681595
transform 1 0 19596 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_199
timestamp 1604681595
transform 1 0 19412 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_203
timestamp 1604681595
transform 1 0 19780 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_192
timestamp 1604681595
transform 1 0 18768 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_199
timestamp 1604681595
transform 1 0 19412 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_203
timestamp 1604681595
transform 1 0 19780 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1604681595
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_218
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_215
timestamp 1604681595
transform 1 0 20884 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_227
timestamp 1604681595
transform 1 0 21988 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1604681595
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1604681595
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_230
timestamp 1604681595
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_242
timestamp 1604681595
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_249
timestamp 1604681595
transform 1 0 24012 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_239
timestamp 1604681595
transform 1 0 23092 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_243
timestamp 1604681595
transform 1 0 23460 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_245
timestamp 1604681595
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1604681595
transform 1 0 25300 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1604681595
transform 1 0 24380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1604681595
transform 1 0 25668 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1604681595
transform 1 0 25852 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1604681595
transform 1 0 24932 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_257
timestamp 1604681595
transform 1 0 24748 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_261
timestamp 1604681595
transform 1 0 25116 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_257
timestamp 1604681595
transform 1 0 24748 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_267
timestamp 1604681595
transform 1 0 25668 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_279
timestamp 1604681595
transform 1 0 26772 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_271
timestamp 1604681595
transform 1 0 26036 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_271
timestamp 1604681595
transform 1 0 26036 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1604681595
transform 1 0 26956 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1604681595
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1604681595
transform 1 0 26404 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1604681595
transform 1 0 26864 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_283
timestamp 1604681595
transform 1 0 27140 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_288
timestamp 1604681595
transform 1 0 27600 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_284
timestamp 1604681595
transform 1 0 27232 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A
timestamp 1604681595
transform 1 0 27324 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1604681595
transform 1 0 27416 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_287
timestamp 1604681595
transform 1 0 27508 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 28888 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 28888 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_296
timestamp 1604681595
transform 1 0 28336 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _14_
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _16_
timestamp 1604681595
transform 1 0 2484 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__14__A
timestamp 1604681595
transform 1 0 1932 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_7
timestamp 1604681595
transform 1 0 1748 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_11
timestamp 1604681595
transform 1 0 2116 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_19
timestamp 1604681595
transform 1 0 2852 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 5336 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_2_44
timestamp 1604681595
transform 1 0 5152 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1604681595
transform 1 0 8188 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_mode_io__0.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 7268 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_65
timestamp 1604681595
transform 1 0 7084 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_69
timestamp 1604681595
transform 1 0 7452 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_81
timestamp 1604681595
transform 1 0 8556 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  ltile_mode_io__2.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9936 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_89
timestamp 1604681595
transform 1 0 9292 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_93
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  ltile_mode_io__3.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12420 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_2_115
timestamp 1604681595
transform 1 0 11684 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_142
timestamp 1604681595
transform 1 0 14168 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_150
timestamp 1604681595
transform 1 0 14904 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1604681595
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1604681595
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1604681595
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1604681595
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_215
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_227
timestamp 1604681595
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_239
timestamp 1604681595
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_251
timestamp 1604681595
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_263
timestamp 1604681595
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1604681595
transform 1 0 26496 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_280
timestamp 1604681595
transform 1 0 26864 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 28888 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_292
timestamp 1604681595
transform 1 0 27968 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_298
timestamp 1604681595
transform 1 0 28520 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _13_
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _17_
timestamp 1604681595
transform 1 0 2484 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__13__A
timestamp 1604681595
transform 1 0 1932 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__12__A
timestamp 1604681595
transform 1 0 2300 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_7
timestamp 1604681595
transform 1 0 1748 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_11
timestamp 1604681595
transform 1 0 2116 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_19
timestamp 1604681595
transform 1 0 2852 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4692 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__17__A
timestamp 1604681595
transform 1 0 3036 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 4048 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 4508 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_23
timestamp 1604681595
transform 1 0 3220 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_31
timestamp 1604681595
transform 1 0 3956 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_34
timestamp 1604681595
transform 1 0 4232 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 5612 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_45
timestamp 1604681595
transform 1 0 5244 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_51
timestamp 1604681595
transform 1 0 5796 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_55
timestamp 1604681595
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1604681595
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1604681595
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1604681595
transform 1 0 9752 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1604681595
transform 1 0 10304 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 10672 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_86
timestamp 1604681595
transform 1 0 9016 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_98
timestamp 1604681595
transform 1 0 10120 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_102
timestamp 1604681595
transform 1 0 10488 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 11040 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_106
timestamp 1604681595
transform 1 0 10856 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1604681595
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1604681595
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 16100 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1604681595
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_159
timestamp 1604681595
transform 1 0 15732 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_165
timestamp 1604681595
transform 1 0 16284 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 16468 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_169
timestamp 1604681595
transform 1 0 16652 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_181
timestamp 1604681595
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1604681595
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1604681595
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_220
timestamp 1604681595
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_232
timestamp 1604681595
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_245
timestamp 1604681595
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1604681595
transform 1 0 25300 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_257
timestamp 1604681595
transform 1 0 24748 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_265
timestamp 1604681595
transform 1 0 25484 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1604681595
transform 1 0 26404 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__33__A
timestamp 1604681595
transform 1 0 26956 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__32__A
timestamp 1604681595
transform 1 0 27324 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_273
timestamp 1604681595
transform 1 0 26220 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_279
timestamp 1604681595
transform 1 0 26772 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_283
timestamp 1604681595
transform 1 0 27140 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_287
timestamp 1604681595
transform 1 0 27508 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 28888 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _12_
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_7
timestamp 1604681595
transform 1 0 1748 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_19
timestamp 1604681595
transform 1 0 2852 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_38
timestamp 1604681595
transform 1 0 4600 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5980 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_4_50
timestamp 1604681595
transform 1 0 5704 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_62
timestamp 1604681595
transform 1 0 6808 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6992 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7360 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_66
timestamp 1604681595
transform 1 0 7176 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_70
timestamp 1604681595
transform 1 0 7544 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_82
timestamp 1604681595
transform 1 0 8648 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 10672 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_93
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_101
timestamp 1604681595
transform 1 0 10396 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_123
timestamp 1604681595
transform 1 0 12420 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_135
timestamp 1604681595
transform 1 0 13524 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_143
timestamp 1604681595
transform 1 0 14260 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_154
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_152
timestamp 1604681595
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_148
timestamp 1604681595
transform 1 0 14720 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14536 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 15456 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_162
timestamp 1604681595
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_158
timestamp 1604681595
transform 1 0 15640 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 15824 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 16100 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 18308 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_182
timestamp 1604681595
transform 1 0 17848 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_186
timestamp 1604681595
transform 1 0 18216 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 18676 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_189
timestamp 1604681595
transform 1 0 18492 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_193
timestamp 1604681595
transform 1 0 18860 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_205
timestamp 1604681595
transform 1 0 19964 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_213
timestamp 1604681595
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_215
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_227
timestamp 1604681595
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_239
timestamp 1604681595
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1604681595
transform 1 0 25300 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_251
timestamp 1604681595
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_267
timestamp 1604681595
transform 1 0 25668 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1604681595
transform 1 0 26496 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_280
timestamp 1604681595
transform 1 0 26864 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 28888 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_292
timestamp 1604681595
transform 1 0 27968 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_298
timestamp 1604681595
transform 1 0 28520 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _19_
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1604681595
transform 1 0 2484 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__19__A
timestamp 1604681595
transform 1 0 1932 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1604681595
transform 1 0 2300 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_7
timestamp 1604681595
transform 1 0 1748 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_11
timestamp 1604681595
transform 1 0 2116 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_19
timestamp 1604681595
transform 1 0 2852 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__78__A
timestamp 1604681595
transform 1 0 3036 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_23
timestamp 1604681595
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_35
timestamp 1604681595
transform 1 0 4324 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_49
timestamp 1604681595
transform 1 0 5612 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_45
timestamp 1604681595
transform 1 0 5244 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 5060 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 5796 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 5428 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1604681595
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_53
timestamp 1604681595
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 8556 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 8372 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_71
timestamp 1604681595
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_75
timestamp 1604681595
transform 1 0 8004 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1604681595
transform 1 0 9384 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 9200 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_84
timestamp 1604681595
transform 1 0 8832 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_99
timestamp 1604681595
transform 1 0 10212 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11224 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_107
timestamp 1604681595
transform 1 0 10948 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_112
timestamp 1604681595
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_116
timestamp 1604681595
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1604681595
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_123
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 12788 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 13156 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 14352 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 13524 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_129
timestamp 1604681595
transform 1 0 12972 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_133
timestamp 1604681595
transform 1 0 13340 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_137
timestamp 1604681595
transform 1 0 13708 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_143
timestamp 1604681595
transform 1 0 14260 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 14536 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_5_165
timestamp 1604681595
transform 1 0 16284 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18308 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 16468 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1604681595
transform 1 0 16652 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_184
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 19320 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 19688 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 20056 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_196
timestamp 1604681595
transform 1 0 19136 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_200
timestamp 1604681595
transform 1 0 19504 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_204
timestamp 1604681595
transform 1 0 19872 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1604681595
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_220
timestamp 1604681595
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_232
timestamp 1604681595
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_245
timestamp 1604681595
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_257
timestamp 1604681595
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_269
timestamp 1604681595
transform 1 0 25852 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _31_
timestamp 1604681595
transform 1 0 26404 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__31__A
timestamp 1604681595
transform 1 0 26956 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__30__A
timestamp 1604681595
transform 1 0 27324 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_279
timestamp 1604681595
transform 1 0 26772 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_283
timestamp 1604681595
transform 1 0 27140 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_287
timestamp 1604681595
transform 1 0 27508 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 28888 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_7
timestamp 1604681595
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1604681595
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_11
timestamp 1604681595
transform 1 0 2116 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1604681595
transform 1 0 2300 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1604681595
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_19
timestamp 1604681595
transform 1 0 2852 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_7
timestamp 1604681595
transform 1 0 1748 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_30
timestamp 1604681595
transform 1 0 3864 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_27
timestamp 1604681595
transform 1 0 3588 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 3680 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 4232 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_32
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_34
timestamp 1604681595
transform 1 0 4232 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 4600 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_36
timestamp 1604681595
transform 1 0 4416 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_40
timestamp 1604681595
transform 1 0 4784 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4600 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_7_51
timestamp 1604681595
transform 1 0 5796 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_47
timestamp 1604681595
transform 1 0 5428 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_44
timestamp 1604681595
transform 1 0 5152 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 4968 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 5428 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_7_58
timestamp 1604681595
transform 1 0 6440 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1604681595
transform 1 0 6072 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_60
timestamp 1604681595
transform 1 0 6624 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_56
timestamp 1604681595
transform 1 0 6256 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 6440 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 6256 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 5888 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_62
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 7544 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6992 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 7360 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_73
timestamp 1604681595
transform 1 0 7820 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_93
timestamp 1604681595
transform 1 0 9660 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_89
timestamp 1604681595
transform 1 0 9292 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_93
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_89
timestamp 1604681595
transform 1 0 9292 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_85
timestamp 1604681595
transform 1 0 8924 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_100
timestamp 1604681595
transform 1 0 10304 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_96
timestamp 1604681595
transform 1 0 9936 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_101
timestamp 1604681595
transform 1 0 10396 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 10212 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 9752 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 10120 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10488 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10672 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10672 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_7_113
timestamp 1604681595
transform 1 0 11500 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_106
timestamp 1604681595
transform 1 0 10856 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 11040 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 11224 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_123
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_118
timestamp 1604681595
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_123
timestamp 1604681595
transform 1 0 12420 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_119
timestamp 1604681595
transform 1 0 12052 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 12236 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12604 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12788 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12788 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 14352 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_136
timestamp 1604681595
transform 1 0 13616 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_136
timestamp 1604681595
transform 1 0 13616 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_147
timestamp 1604681595
transform 1 0 14628 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_154
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_152
timestamp 1604681595
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_148
timestamp 1604681595
transform 1 0 14720 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 14812 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1604681595
transform 1 0 15364 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_7_163
timestamp 1604681595
transform 1 0 16100 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_151
timestamp 1604681595
transform 1 0 14996 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_164
timestamp 1604681595
transform 1 0 16192 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_176
timestamp 1604681595
transform 1 0 17296 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_172
timestamp 1604681595
transform 1 0 16928 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_169
timestamp 1604681595
transform 1 0 16652 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 16744 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 17112 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_184
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_180
timestamp 1604681595
transform 1 0 17664 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 18216 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_176
timestamp 1604681595
transform 1 0 17296 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_197
timestamp 1604681595
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_196
timestamp 1604681595
transform 1 0 19136 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_190
timestamp 1604681595
transform 1 0 18584 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 18400 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 19228 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18400 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_201
timestamp 1604681595
transform 1 0 19596 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_206
timestamp 1604681595
transform 1 0 20056 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19780 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19964 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 21528 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 21344 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 21528 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_215
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_221
timestamp 1604681595
transform 1 0 21436 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_224
timestamp 1604681595
transform 1 0 21712 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_214
timestamp 1604681595
transform 1 0 20792 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_236
timestamp 1604681595
transform 1 0 22816 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_248
timestamp 1604681595
transform 1 0 23920 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_231
timestamp 1604681595
transform 1 0 22356 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_243
timestamp 1604681595
transform 1 0 23460 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_245
timestamp 1604681595
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_260
timestamp 1604681595
transform 1 0 25024 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_257
timestamp 1604681595
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_269
timestamp 1604681595
transform 1 0 25852 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_279
timestamp 1604681595
transform 1 0 26772 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_272
timestamp 1604681595
transform 1 0 26128 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__29__A
timestamp 1604681595
transform 1 0 26956 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _30_
timestamp 1604681595
transform 1 0 26496 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _29_
timestamp 1604681595
transform 1 0 26404 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_283
timestamp 1604681595
transform 1 0 27140 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__27__A
timestamp 1604681595
transform 1 0 27324 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_287
timestamp 1604681595
transform 1 0 27508 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_280
timestamp 1604681595
transform 1 0 26864 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 28888 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 28888 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_292
timestamp 1604681595
transform 1 0 27968 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_298
timestamp 1604681595
transform 1 0 28520 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_7
timestamp 1604681595
transform 1 0 1748 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_19
timestamp 1604681595
transform 1 0 2852 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 3312 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_23
timestamp 1604681595
transform 1 0 3220 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_26
timestamp 1604681595
transform 1 0 3496 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_30
timestamp 1604681595
transform 1 0 3864 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_41
timestamp 1604681595
transform 1 0 4876 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 5888 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_8_49
timestamp 1604681595
transform 1 0 5612 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_61
timestamp 1604681595
transform 1 0 6716 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 6900 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 7544 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_65
timestamp 1604681595
transform 1 0 7084 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_69
timestamp 1604681595
transform 1 0 7452 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_72
timestamp 1604681595
transform 1 0 7728 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10212 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 9844 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_84
timestamp 1604681595
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_88
timestamp 1604681595
transform 1 0 9200 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_93
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_97
timestamp 1604681595
transform 1 0 10028 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_2_
timestamp 1604681595
transform 1 0 11776 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 11224 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 11592 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_108
timestamp 1604681595
transform 1 0 11040 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_112
timestamp 1604681595
transform 1 0 11408 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_125
timestamp 1604681595
transform 1 0 12604 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12788 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13156 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_129
timestamp 1604681595
transform 1 0 12972 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_133
timestamp 1604681595
transform 1 0 13340 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_145
timestamp 1604681595
transform 1 0 14444 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 16284 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 15824 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_154
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_8_162
timestamp 1604681595
transform 1 0 16008 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 17112 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_8_167
timestamp 1604681595
transform 1 0 16468 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_173
timestamp 1604681595
transform 1 0 17020 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19964 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_193
timestamp 1604681595
transform 1 0 18860 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_207
timestamp 1604681595
transform 1 0 20148 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 21528 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1604681595
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_215
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_221
timestamp 1604681595
transform 1 0 21436 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_224
timestamp 1604681595
transform 1 0 21712 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_236
timestamp 1604681595
transform 1 0 22816 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_248
timestamp 1604681595
transform 1 0 23920 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_260
timestamp 1604681595
transform 1 0 25024 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _27_
timestamp 1604681595
transform 1 0 26496 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_272
timestamp 1604681595
transform 1 0 26128 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_280
timestamp 1604681595
transform 1 0 26864 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 28888 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_292
timestamp 1604681595
transform 1 0 27968 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_298
timestamp 1604681595
transform 1 0 28520 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1604681595
transform 1 0 1932 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1604681595
transform 1 0 2300 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_7
timestamp 1604681595
transform 1 0 1748 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_11
timestamp 1604681595
transform 1 0 2116 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_15
timestamp 1604681595
transform 1 0 2484 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 3312 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 3128 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_21
timestamp 1604681595
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_43
timestamp 1604681595
transform 1 0 5060 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1604681595
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_71
timestamp 1604681595
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_75
timestamp 1604681595
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_79
timestamp 1604681595
transform 1 0 8372 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_83
timestamp 1604681595
transform 1 0 8740 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 10396 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1604681595
transform 1 0 9568 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1604681595
transform 1 0 9016 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 8832 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_89
timestamp 1604681595
transform 1 0 9292 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1604681595
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_123
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 13340 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 13156 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1604681595
transform 1 0 15824 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 15640 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_152
timestamp 1604681595
transform 1 0 15088 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_156
timestamp 1604681595
transform 1 0 15456 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 16836 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1604681595
transform 1 0 16652 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_173
timestamp 1604681595
transform 1 0 17020 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_181
timestamp 1604681595
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 19964 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 19780 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_196
timestamp 1604681595
transform 1 0 19136 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_201
timestamp 1604681595
transform 1 0 19596 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_214
timestamp 1604681595
transform 1 0 20792 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_226
timestamp 1604681595
transform 1 0 21896 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_238
timestamp 1604681595
transform 1 0 23000 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_245
timestamp 1604681595
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_257
timestamp 1604681595
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_269
timestamp 1604681595
transform 1 0 25852 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _28_
timestamp 1604681595
transform 1 0 26404 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__28__A
timestamp 1604681595
transform 1 0 26956 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__25__A
timestamp 1604681595
transform 1 0 27324 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_279
timestamp 1604681595
transform 1 0 26772 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_283
timestamp 1604681595
transform 1 0 27140 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_287
timestamp 1604681595
transform 1 0 27508 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 28888 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_7
timestamp 1604681595
transform 1 0 1748 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_19
timestamp 1604681595
transform 1 0 2852 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1604681595
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1604681595
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_56
timestamp 1604681595
transform 1 0 6256 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_62
timestamp 1604681595
transform 1 0 6808 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 7084 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 6900 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 10396 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 9844 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_84
timestamp 1604681595
transform 1 0 8832 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_97
timestamp 1604681595
transform 1 0 10028 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_103
timestamp 1604681595
transform 1 0 10580 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 11224 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 10764 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_107
timestamp 1604681595
transform 1 0 10948 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 13340 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_130
timestamp 1604681595
transform 1 0 13064 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_135
timestamp 1604681595
transform 1 0 13524 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1604681595
transform 1 0 16284 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 15824 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_147
timestamp 1604681595
transform 1 0 14628 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_10_154
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_10_162
timestamp 1604681595
transform 1 0 16008 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _10_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 17848 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 18308 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_174
timestamp 1604681595
transform 1 0 17112 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_185
timestamp 1604681595
transform 1 0 18124 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 19964 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 19136 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1604681595
transform 1 0 18492 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1604681595
transform 1 0 19044 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_198
timestamp 1604681595
transform 1 0 19320 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_204
timestamp 1604681595
transform 1 0 19872 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_207
timestamp 1604681595
transform 1 0 20148 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_213
timestamp 1604681595
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_215
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_227
timestamp 1604681595
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_239
timestamp 1604681595
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_251
timestamp 1604681595
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_263
timestamp 1604681595
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _25_
timestamp 1604681595
transform 1 0 26496 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_280
timestamp 1604681595
transform 1 0 26864 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 28888 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_292
timestamp 1604681595
transform 1 0 27968 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_298
timestamp 1604681595
transform 1 0 28520 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1604681595
transform 1 0 2484 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1604681595
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1604681595
transform 1 0 2300 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_7
timestamp 1604681595
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_11
timestamp 1604681595
transform 1 0 2116 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_19
timestamp 1604681595
transform 1 0 2852 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 3772 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1604681595
transform 1 0 3036 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 3588 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_23
timestamp 1604681595
transform 1 0 3220 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_48
timestamp 1604681595
transform 1 0 5520 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_54
timestamp 1604681595
transform 1 0 6072 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1604681595
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_62
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _06_
timestamp 1604681595
transform 1 0 8740 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 7176 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 6992 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 8556 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_75
timestamp 1604681595
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_79
timestamp 1604681595
transform 1 0 8372 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 10212 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_86
timestamp 1604681595
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_98
timestamp 1604681595
transform 1 0 10120 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_101
timestamp 1604681595
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _11_
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1604681595
transform 1 0 10764 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_114
timestamp 1604681595
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_118
timestamp 1604681595
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1604681595
transform 1 0 13524 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 13984 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_126
timestamp 1604681595
transform 1 0 12696 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_134
timestamp 1604681595
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_138
timestamp 1604681595
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_142
timestamp 1604681595
transform 1 0 14168 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1604681595
transform 1 0 16284 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 16100 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 15732 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 15272 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 14904 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_152
timestamp 1604681595
transform 1 0 15088 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_156
timestamp 1604681595
transform 1 0 15456 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_161
timestamp 1604681595
transform 1 0 15916 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 18308 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 17296 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_174
timestamp 1604681595
transform 1 0 17112 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_178
timestamp 1604681595
transform 1 0 17480 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_182
timestamp 1604681595
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_184
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 19136 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 18952 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_189
timestamp 1604681595
transform 1 0 18492 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_193
timestamp 1604681595
transform 1 0 18860 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_215
timestamp 1604681595
transform 1 0 20884 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_227
timestamp 1604681595
transform 1 0 21988 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_239
timestamp 1604681595
transform 1 0 23092 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_243
timestamp 1604681595
transform 1 0 23460 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_245
timestamp 1604681595
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_257
timestamp 1604681595
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_269
timestamp 1604681595
transform 1 0 25852 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _24_
timestamp 1604681595
transform 1 0 26404 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _26_
timestamp 1604681595
transform 1 0 27508 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__24__A
timestamp 1604681595
transform 1 0 26956 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__23__A
timestamp 1604681595
transform 1 0 27324 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_279
timestamp 1604681595
transform 1 0 26772 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_283
timestamp 1604681595
transform 1 0 27140 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_291
timestamp 1604681595
transform 1 0 27876 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 28888 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__26__A
timestamp 1604681595
transform 1 0 28060 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_295
timestamp 1604681595
transform 1 0 28244 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 2392 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2944 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_7
timestamp 1604681595
transform 1 0 1748 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_13
timestamp 1604681595
transform 1 0 2300 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_16
timestamp 1604681595
transform 1 0 2576 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4508 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3312 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_22
timestamp 1604681595
transform 1 0 3128 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_26
timestamp 1604681595
transform 1 0 3496 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_30
timestamp 1604681595
transform 1 0 3864 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_32
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_36
timestamp 1604681595
transform 1 0 4416 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_39
timestamp 1604681595
transform 1 0 4692 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_51
timestamp 1604681595
transform 1 0 5796 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 7084 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_63
timestamp 1604681595
transform 1 0 6900 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_74
timestamp 1604681595
transform 1 0 7912 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_86
timestamp 1604681595
transform 1 0 9016 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_93
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1604681595
transform 1 0 11040 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 10764 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_107
timestamp 1604681595
transform 1 0 10948 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_117
timestamp 1604681595
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 14352 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_129
timestamp 1604681595
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_141
timestamp 1604681595
transform 1 0 14076 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_146
timestamp 1604681595
transform 1 0 14536 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_152
timestamp 1604681595
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 18308 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 17848 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_173
timestamp 1604681595
transform 1 0 17020 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_181
timestamp 1604681595
transform 1 0 17756 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_184
timestamp 1604681595
transform 1 0 18032 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_206
timestamp 1604681595
transform 1 0 20056 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_215
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_227
timestamp 1604681595
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_239
timestamp 1604681595
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_251
timestamp 1604681595
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_263
timestamp 1604681595
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _23_
timestamp 1604681595
transform 1 0 26496 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_280
timestamp 1604681595
transform 1 0 26864 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 28888 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_292
timestamp 1604681595
transform 1 0 27968 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_298
timestamp 1604681595
transform 1 0 28520 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_7
timestamp 1604681595
transform 1 0 1748 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_7
timestamp 1604681595
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 1840 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1604681595
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_10
timestamp 1604681595
transform 1 0 2024 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_16
timestamp 1604681595
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_11
timestamp 1604681595
transform 1 0 2116 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 2760 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_2_
timestamp 1604681595
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2944 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1604681595
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_23
timestamp 1604681595
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_29
timestamp 1604681595
transform 1 0 3772 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_36
timestamp 1604681595
transform 1 0 4416 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_32
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_33
timestamp 1604681595
transform 1 0 4140 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3956 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 4232 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4324 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4508 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 5152 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 5520 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 5888 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_46
timestamp 1604681595
transform 1 0 5336 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_50
timestamp 1604681595
transform 1 0 5704 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_54
timestamp 1604681595
transform 1 0 6072 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_60
timestamp 1604681595
transform 1 0 6624 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_62
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 7544 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 8188 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_73
timestamp 1604681595
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_77
timestamp 1604681595
transform 1 0 8188 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_63
timestamp 1604681595
transform 1 0 6900 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_75
timestamp 1604681595
transform 1 0 8004 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_79
timestamp 1604681595
transform 1 0 8372 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_93
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1604681595
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_99
timestamp 1604681595
transform 1 0 10212 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_104
timestamp 1604681595
transform 1 0 10672 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_101
timestamp 1604681595
transform 1 0 10396 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 10304 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 10488 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10488 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_13_89
timestamp 1604681595
transform 1 0 9292 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 10856 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 11224 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_108
timestamp 1604681595
transform 1 0 11040 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_112
timestamp 1604681595
transform 1 0 11408 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1604681595
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_111
timestamp 1604681595
transform 1 0 11316 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_123
timestamp 1604681595
transform 1 0 12420 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1604681595
transform 1 0 14352 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 14168 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 14352 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 13892 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_135
timestamp 1604681595
transform 1 0 13524 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_141
timestamp 1604681595
transform 1 0 14076 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_135
timestamp 1604681595
transform 1 0 13524 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_141
timestamp 1604681595
transform 1 0 14076 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_154
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_149
timestamp 1604681595
transform 1 0 14812 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_153
timestamp 1604681595
transform 1 0 15180 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 15364 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 14536 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_162
timestamp 1604681595
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_158
timestamp 1604681595
transform 1 0 15640 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_165
timestamp 1604681595
transform 1 0 16284 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_161
timestamp 1604681595
transform 1 0 15916 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_157
timestamp 1604681595
transform 1 0 15548 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 15732 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 16100 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 15456 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16100 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_14_176
timestamp 1604681595
transform 1 0 17296 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_172
timestamp 1604681595
transform 1 0 16928 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_175
timestamp 1604681595
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_169
timestamp 1604681595
transform 1 0 16652 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 16468 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17112 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 17020 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_179
timestamp 1604681595
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1604681595
transform 1 0 17848 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 18860 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 19412 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_193
timestamp 1604681595
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_197
timestamp 1604681595
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_201
timestamp 1604681595
transform 1 0 19596 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_191
timestamp 1604681595
transform 1 0 18676 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_195
timestamp 1604681595
transform 1 0 19044 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_207
timestamp 1604681595
transform 1 0 20148 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_213
timestamp 1604681595
transform 1 0 20700 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1604681595
transform 1 0 21804 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1604681595
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_215
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_227
timestamp 1604681595
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_237
timestamp 1604681595
transform 1 0 22908 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_243
timestamp 1604681595
transform 1 0 23460 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_245
timestamp 1604681595
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_239
timestamp 1604681595
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_257
timestamp 1604681595
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_269
timestamp 1604681595
transform 1 0 25852 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_251
timestamp 1604681595
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_263
timestamp 1604681595
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1604681595
transform 1 0 26956 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_276
timestamp 1604681595
transform 1 0 26496 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_288
timestamp 1604681595
transform 1 0 27600 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 28888 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 28888 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_293
timestamp 1604681595
transform 1 0 28060 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_14_296
timestamp 1604681595
transform 1 0 28336 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 2484 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 2300 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1604681595
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_7
timestamp 1604681595
transform 1 0 1748 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_11
timestamp 1604681595
transform 1 0 2116 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 4048 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 3496 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_24
timestamp 1604681595
transform 1 0 3312 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_28
timestamp 1604681595
transform 1 0 3680 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_41
timestamp 1604681595
transform 1 0 4876 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_53
timestamp 1604681595
transform 1 0 5980 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_62
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 8188 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6992 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 7360 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_66
timestamp 1604681595
transform 1 0 7176 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_70
timestamp 1604681595
transform 1 0 7544 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_74
timestamp 1604681595
transform 1 0 7912 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10672 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10488 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_96
timestamp 1604681595
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_100
timestamp 1604681595
transform 1 0 10304 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 11684 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 12052 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1604681595
transform 1 0 11500 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_117
timestamp 1604681595
transform 1 0 11868 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1604681595
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_123
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 13892 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 13708 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_135
timestamp 1604681595
transform 1 0 13524 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_158
timestamp 1604681595
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_162
timestamp 1604681595
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_175
timestamp 1604681595
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_179
timestamp 1604681595
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19780 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_193
timestamp 1604681595
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_197
timestamp 1604681595
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_201
timestamp 1604681595
transform 1 0 19596 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_205
timestamp 1604681595
transform 1 0 19964 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_217
timestamp 1604681595
transform 1 0 21068 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_229
timestamp 1604681595
transform 1 0 22172 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_241
timestamp 1604681595
transform 1 0 23276 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_245
timestamp 1604681595
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_257
timestamp 1604681595
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_269
timestamp 1604681595
transform 1 0 25852 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _22_
timestamp 1604681595
transform 1 0 26404 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__22__A
timestamp 1604681595
transform 1 0 26956 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__20__A
timestamp 1604681595
transform 1 0 27324 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_279
timestamp 1604681595
transform 1 0 26772 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_283
timestamp 1604681595
transform 1 0 27140 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_287
timestamp 1604681595
transform 1 0 27508 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 28888 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2208 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_8
timestamp 1604681595
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_21
timestamp 1604681595
transform 1 0 3036 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_25
timestamp 1604681595
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1604681595
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 6624 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1604681595
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_56
timestamp 1604681595
transform 1 0 6256 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 8556 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_79
timestamp 1604681595
transform 1 0 8372 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_83
timestamp 1604681595
transform 1 0 8740 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_2_
timestamp 1604681595
transform 1 0 10396 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10028 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 8924 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_87
timestamp 1604681595
transform 1 0 9108 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_93
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_99
timestamp 1604681595
transform 1 0 10212 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11408 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_110
timestamp 1604681595
transform 1 0 11224 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_114
timestamp 1604681595
transform 1 0 11592 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 14168 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_126
timestamp 1604681595
transform 1 0 12696 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_138
timestamp 1604681595
transform 1 0 13800 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_144
timestamp 1604681595
transform 1 0 14352 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16376 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_152
timestamp 1604681595
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_163
timestamp 1604681595
transform 1 0 16100 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18032 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16744 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_168
timestamp 1604681595
transform 1 0 16560 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_172
timestamp 1604681595
transform 1 0 16928 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_193
timestamp 1604681595
transform 1 0 18860 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_205
timestamp 1604681595
transform 1 0 19964 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_213
timestamp 1604681595
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_215
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_227
timestamp 1604681595
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_239
timestamp 1604681595
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_251
timestamp 1604681595
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_263
timestamp 1604681595
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _20_
timestamp 1604681595
transform 1 0 26496 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_280
timestamp 1604681595
transform 1 0 26864 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 28888 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_292
timestamp 1604681595
transform 1 0 27968 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_298
timestamp 1604681595
transform 1 0 28520 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1604681595
transform 1 0 2116 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_7
timestamp 1604681595
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_20
timestamp 1604681595
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1604681595
transform 1 0 3680 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 3128 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 3496 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 4692 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_24
timestamp 1604681595
transform 1 0 3312 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_37
timestamp 1604681595
transform 1 0 4508 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_41
timestamp 1604681595
transform 1 0 4876 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 5428 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 5796 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_49
timestamp 1604681595
transform 1 0 5612 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_53
timestamp 1604681595
transform 1 0 5980 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_62
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 8464 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 7268 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_66
timestamp 1604681595
transform 1 0 7176 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_69
timestamp 1604681595
transform 1 0 7452 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_73
timestamp 1604681595
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_77
timestamp 1604681595
transform 1 0 8188 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10028 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 9476 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_89
timestamp 1604681595
transform 1 0 9292 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_93
timestamp 1604681595
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11040 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11408 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_106
timestamp 1604681595
transform 1 0 10856 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1604681595
transform 1 0 11224 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_114
timestamp 1604681595
transform 1 0 11592 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1604681595
transform 1 0 14168 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 13984 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_135
timestamp 1604681595
transform 1 0 13524 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_139
timestamp 1604681595
transform 1 0 13892 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1604681595
transform 1 0 15732 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 15548 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 15180 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_151
timestamp 1604681595
transform 1 0 14996 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_155
timestamp 1604681595
transform 1 0 15364 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 17296 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 17664 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_168
timestamp 1604681595
transform 1 0 16560 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_178
timestamp 1604681595
transform 1 0 17480 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_182
timestamp 1604681595
transform 1 0 17848 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1604681595
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_208
timestamp 1604681595
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_220
timestamp 1604681595
transform 1 0 21344 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_232
timestamp 1604681595
transform 1 0 22448 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_245
timestamp 1604681595
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_257
timestamp 1604681595
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_269
timestamp 1604681595
transform 1 0 25852 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _21_
timestamp 1604681595
transform 1 0 26404 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__21__A
timestamp 1604681595
transform 1 0 26956 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_279
timestamp 1604681595
transform 1 0 26772 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_283
timestamp 1604681595
transform 1 0 27140 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 28888 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_295
timestamp 1604681595
transform 1 0 28244 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1604681595
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1604681595
transform 1 0 1564 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 2116 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_7
timestamp 1604681595
transform 1 0 1748 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_13
timestamp 1604681595
transform 1 0 2300 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 4232 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_23
timestamp 1604681595
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1604681595
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_32
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_36
timestamp 1604681595
transform 1 0 4416 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 5428 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_18_44
timestamp 1604681595
transform 1 0 5152 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 7820 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_66
timestamp 1604681595
transform 1 0 7176 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_72
timestamp 1604681595
transform 1 0 7728 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9936 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_84
timestamp 1604681595
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_88
timestamp 1604681595
transform 1 0 9200 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_93
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 10948 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 11316 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_105
timestamp 1604681595
transform 1 0 10764 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_109
timestamp 1604681595
transform 1 0 11132 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_113
timestamp 1604681595
transform 1 0 11500 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_121
timestamp 1604681595
transform 1 0 12236 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_125
timestamp 1604681595
transform 1 0 12604 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 14168 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_137
timestamp 1604681595
transform 1 0 13708 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_141
timestamp 1604681595
transform 1 0 14076 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_144
timestamp 1604681595
transform 1 0 14352 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _09_
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 15732 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_152
timestamp 1604681595
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_157
timestamp 1604681595
transform 1 0 15548 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_161
timestamp 1604681595
transform 1 0 15916 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 17296 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_18_173
timestamp 1604681595
transform 1 0 17020 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_195
timestamp 1604681595
transform 1 0 19044 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_207
timestamp 1604681595
transform 1 0 20148 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_213
timestamp 1604681595
transform 1 0 20700 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_215
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_227
timestamp 1604681595
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_239
timestamp 1604681595
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_251
timestamp 1604681595
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_263
timestamp 1604681595
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_276
timestamp 1604681595
transform 1 0 26496 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_288
timestamp 1604681595
transform 1 0 27600 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 28888 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_296
timestamp 1604681595
transform 1 0 28336 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_7
timestamp 1604681595
transform 1 0 1748 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 1932 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_18
timestamp 1604681595
transform 1 0 2760 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_11
timestamp 1604681595
transform 1 0 2116 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 2944 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 2300 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1604681595
transform 1 0 2484 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _07_
timestamp 1604681595
transform 1 0 2484 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 4232 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 4048 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_24
timestamp 1604681595
transform 1 0 3312 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_22
timestamp 1604681595
transform 1 0 3128 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_30
timestamp 1604681595
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_53
timestamp 1604681595
transform 1 0 5980 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1604681595
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1604681595
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _08_
timestamp 1604681595
transform 1 0 8556 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_74
timestamp 1604681595
transform 1 0 7912 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_82
timestamp 1604681595
transform 1 0 8648 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1604681595
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_80
timestamp 1604681595
transform 1 0 8464 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_88
timestamp 1604681595
transform 1 0 9200 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_84
timestamp 1604681595
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 8832 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1604681595
transform 1 0 9016 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_102
timestamp 1604681595
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_99
timestamp 1604681595
transform 1 0 10212 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_95
timestamp 1604681595
transform 1 0 9844 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 10028 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1604681595
transform 1 0 10580 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_110
timestamp 1604681595
transform 1 0 11224 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_106
timestamp 1604681595
transform 1 0 10856 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_112
timestamp 1604681595
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 11040 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_116
timestamp 1604681595
transform 1 0 11776 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 11316 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_19_142
timestamp 1604681595
transform 1 0 14168 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_130
timestamp 1604681595
transform 1 0 13064 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_142
timestamp 1604681595
transform 1 0 14168 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 15272 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 15088 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14720 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_150
timestamp 1604681595
transform 1 0 14904 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_150
timestamp 1604681595
transform 1 0 14904 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_166
timestamp 1604681595
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_173
timestamp 1604681595
transform 1 0 17020 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_181
timestamp 1604681595
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_178
timestamp 1604681595
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1604681595
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1604681595
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_190
timestamp 1604681595
transform 1 0 18584 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_202
timestamp 1604681595
transform 1 0 19688 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_220
timestamp 1604681595
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_215
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_227
timestamp 1604681595
transform 1 0 21988 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_232
timestamp 1604681595
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_245
timestamp 1604681595
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_239
timestamp 1604681595
transform 1 0 23092 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_257
timestamp 1604681595
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_269
timestamp 1604681595
transform 1 0 25852 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_251
timestamp 1604681595
transform 1 0 24196 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_263
timestamp 1604681595
transform 1 0 25300 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1604681595
transform 1 0 26956 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_276
timestamp 1604681595
transform 1 0 26496 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_288
timestamp 1604681595
transform 1 0 27600 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 28888 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 28888 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_293
timestamp 1604681595
transform 1 0 28060 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_20_296
timestamp 1604681595
transform 1 0 28336 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1604681595
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1604681595
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1604681595
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1604681595
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1604681595
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_74
timestamp 1604681595
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_86
timestamp 1604681595
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_98
timestamp 1604681595
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_110
timestamp 1604681595
transform 1 0 11224 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_135
timestamp 1604681595
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_147
timestamp 1604681595
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_159
timestamp 1604681595
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_171
timestamp 1604681595
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1604681595
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1604681595
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_220
timestamp 1604681595
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_232
timestamp 1604681595
transform 1 0 22448 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_245
timestamp 1604681595
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_257
timestamp 1604681595
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_269
timestamp 1604681595
transform 1 0 25852 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1604681595
transform 1 0 26956 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 28888 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_293
timestamp 1604681595
transform 1 0 28060 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1604681595
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1604681595
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1604681595
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1604681595
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_68
timestamp 1604681595
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_80
timestamp 1604681595
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_93
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_105
timestamp 1604681595
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_117
timestamp 1604681595
transform 1 0 11868 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_129
timestamp 1604681595
transform 1 0 12972 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1604681595
transform 1 0 14076 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_154
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_166
timestamp 1604681595
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_178
timestamp 1604681595
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_190
timestamp 1604681595
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_202
timestamp 1604681595
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_215
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_227
timestamp 1604681595
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_239
timestamp 1604681595
transform 1 0 23092 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_251
timestamp 1604681595
transform 1 0 24196 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_263
timestamp 1604681595
transform 1 0 25300 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_276
timestamp 1604681595
transform 1 0 26496 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_288
timestamp 1604681595
transform 1 0 27600 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 28888 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_296
timestamp 1604681595
transform 1 0 28336 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1604681595
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1604681595
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1604681595
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1604681595
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_74
timestamp 1604681595
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_86
timestamp 1604681595
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_98
timestamp 1604681595
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_110
timestamp 1604681595
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1604681595
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_147
timestamp 1604681595
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_159
timestamp 1604681595
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_171
timestamp 1604681595
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1604681595
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1604681595
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_220
timestamp 1604681595
transform 1 0 21344 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_232
timestamp 1604681595
transform 1 0 22448 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_245
timestamp 1604681595
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_257
timestamp 1604681595
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_269
timestamp 1604681595
transform 1 0 25852 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1604681595
transform 1 0 26956 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 28888 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_293
timestamp 1604681595
transform 1 0 28060 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1604681595
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1604681595
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1604681595
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1604681595
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1604681595
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_80
timestamp 1604681595
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1604681595
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_117
timestamp 1604681595
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_129
timestamp 1604681595
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1604681595
transform 1 0 14076 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1604681595
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1604681595
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1604681595
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_202
timestamp 1604681595
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_215
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_227
timestamp 1604681595
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_239
timestamp 1604681595
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_251
timestamp 1604681595
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_263
timestamp 1604681595
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_276
timestamp 1604681595
transform 1 0 26496 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_288
timestamp 1604681595
transform 1 0 27600 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 28888 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_296
timestamp 1604681595
transform 1 0 28336 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1604681595
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1604681595
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1604681595
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1604681595
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1604681595
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1604681595
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1604681595
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_98
timestamp 1604681595
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1604681595
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_135
timestamp 1604681595
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_147
timestamp 1604681595
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_159
timestamp 1604681595
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_171
timestamp 1604681595
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1604681595
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1604681595
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_220
timestamp 1604681595
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_232
timestamp 1604681595
transform 1 0 22448 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_245
timestamp 1604681595
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_257
timestamp 1604681595
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_269
timestamp 1604681595
transform 1 0 25852 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1604681595
transform 1 0 26956 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 28888 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_293
timestamp 1604681595
transform 1 0 28060 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1604681595
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1604681595
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1604681595
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1604681595
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1604681595
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1604681595
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1604681595
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1604681595
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1604681595
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1604681595
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1604681595
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_74
timestamp 1604681595
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_86
timestamp 1604681595
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_98
timestamp 1604681595
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1604681595
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_117
timestamp 1604681595
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_110
timestamp 1604681595
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_129
timestamp 1604681595
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1604681595
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_135
timestamp 1604681595
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1604681595
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_147
timestamp 1604681595
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_159
timestamp 1604681595
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1604681595
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_171
timestamp 1604681595
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_190
timestamp 1604681595
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_202
timestamp 1604681595
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1604681595
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1604681595
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_215
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_227
timestamp 1604681595
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_220
timestamp 1604681595
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_239
timestamp 1604681595
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_232
timestamp 1604681595
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_245
timestamp 1604681595
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_251
timestamp 1604681595
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_263
timestamp 1604681595
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_257
timestamp 1604681595
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_269
timestamp 1604681595
transform 1 0 25852 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_276
timestamp 1604681595
transform 1 0 26496 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_288
timestamp 1604681595
transform 1 0 27600 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1604681595
transform 1 0 26956 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 28888 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 28888 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_296
timestamp 1604681595
transform 1 0 28336 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_293
timestamp 1604681595
transform 1 0 28060 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1604681595
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1604681595
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1604681595
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1604681595
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1604681595
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_80
timestamp 1604681595
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_93
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_105
timestamp 1604681595
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_117
timestamp 1604681595
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_129
timestamp 1604681595
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1604681595
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1604681595
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1604681595
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1604681595
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_202
timestamp 1604681595
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_215
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_227
timestamp 1604681595
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_239
timestamp 1604681595
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_251
timestamp 1604681595
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_263
timestamp 1604681595
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_276
timestamp 1604681595
transform 1 0 26496 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_288
timestamp 1604681595
transform 1 0 27600 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 28888 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_296
timestamp 1604681595
transform 1 0 28336 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1604681595
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1604681595
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1604681595
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1604681595
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1604681595
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_74
timestamp 1604681595
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_86
timestamp 1604681595
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_98
timestamp 1604681595
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_110
timestamp 1604681595
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_135
timestamp 1604681595
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_147
timestamp 1604681595
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_159
timestamp 1604681595
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_171
timestamp 1604681595
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1604681595
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1604681595
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_220
timestamp 1604681595
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_232
timestamp 1604681595
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_245
timestamp 1604681595
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_257
timestamp 1604681595
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_269
timestamp 1604681595
transform 1 0 25852 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1604681595
transform 1 0 26956 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 28888 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_293
timestamp 1604681595
transform 1 0 28060 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1604681595
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1604681595
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1604681595
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1604681595
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1604681595
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_80
timestamp 1604681595
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_105
timestamp 1604681595
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_117
timestamp 1604681595
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_129
timestamp 1604681595
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1604681595
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_166
timestamp 1604681595
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_178
timestamp 1604681595
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_190
timestamp 1604681595
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_202
timestamp 1604681595
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_215
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_227
timestamp 1604681595
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_239
timestamp 1604681595
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_251
timestamp 1604681595
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_263
timestamp 1604681595
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_276
timestamp 1604681595
transform 1 0 26496 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_288
timestamp 1604681595
transform 1 0 27600 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 28888 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_296
timestamp 1604681595
transform 1 0 28336 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1604681595
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1604681595
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1604681595
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1604681595
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1604681595
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_86
timestamp 1604681595
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_98
timestamp 1604681595
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_110
timestamp 1604681595
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_135
timestamp 1604681595
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1604681595
transform 1 0 15272 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1604681595
transform 1 0 16376 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_147
timestamp 1604681595
transform 1 0 14628 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_153
timestamp 1604681595
transform 1 0 15180 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_156
timestamp 1604681595
transform 1 0 15456 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_164
timestamp 1604681595
transform 1 0 16192 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_168
timestamp 1604681595
transform 1 0 16560 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_180
timestamp 1604681595
transform 1 0 17664 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1604681595
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1604681595
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_220
timestamp 1604681595
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_232
timestamp 1604681595
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_245
timestamp 1604681595
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_257
timestamp 1604681595
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_269
timestamp 1604681595
transform 1 0 25852 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1604681595
transform 1 0 26496 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_275
timestamp 1604681595
transform 1 0 26404 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_278
timestamp 1604681595
transform 1 0 26680 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_290
timestamp 1604681595
transform 1 0 27784 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 28888 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_298
timestamp 1604681595
transform 1 0 28520 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1604681595
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1604681595
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1604681595
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1604681595
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_68
timestamp 1604681595
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_80
timestamp 1604681595
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_105
timestamp 1604681595
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_117
timestamp 1604681595
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_129
timestamp 1604681595
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1604681595
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1604681595
transform 1 0 16376 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_158
timestamp 1604681595
transform 1 0 15640 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_170
timestamp 1604681595
transform 1 0 16744 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_182
timestamp 1604681595
transform 1 0 17848 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_194
timestamp 1604681595
transform 1 0 18952 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_206
timestamp 1604681595
transform 1 0 20056 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_215
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_227
timestamp 1604681595
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_239
timestamp 1604681595
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_251
timestamp 1604681595
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_263
timestamp 1604681595
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1604681595
transform 1 0 26496 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_280
timestamp 1604681595
transform 1 0 26864 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 28888 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_292
timestamp 1604681595
transform 1 0 27968 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_298
timestamp 1604681595
transform 1 0 28520 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1604681595
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1604681595
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1604681595
transform 1 0 4692 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1604681595
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1604681595
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1604681595
transform 1 0 5244 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_43
timestamp 1604681595
transform 1 0 5060 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_47
timestamp 1604681595
transform 1 0 5428 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1604681595
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1604681595
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1604681595
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1604681595
transform 1 0 7912 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1604681595
transform 1 0 7360 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1604681595
transform 1 0 8464 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_66
timestamp 1604681595
transform 1 0 7176 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_70
timestamp 1604681595
transform 1 0 7544 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_78
timestamp 1604681595
transform 1 0 8280 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_82
timestamp 1604681595
transform 1 0 8648 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_68
timestamp 1604681595
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_80
timestamp 1604681595
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1604681595
transform 1 0 9936 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_94
timestamp 1604681595
transform 1 0 9752 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_100
timestamp 1604681595
transform 1 0 10304 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_112
timestamp 1604681595
transform 1 0 11408 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_120
timestamp 1604681595
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_123
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_105
timestamp 1604681595
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_117
timestamp 1604681595
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1604681595
transform 1 0 14076 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_135
timestamp 1604681595
transform 1 0 13524 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_145
timestamp 1604681595
transform 1 0 14444 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_129
timestamp 1604681595
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1604681595
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1604681595
transform 1 0 15364 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1604681595
transform 1 0 14628 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1604681595
transform 1 0 15916 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_149
timestamp 1604681595
transform 1 0 14812 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_159
timestamp 1604681595
transform 1 0 15732 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_163
timestamp 1604681595
transform 1 0 16100 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_154
timestamp 1604681595
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_166
timestamp 1604681595
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1604681595
transform 1 0 16468 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1604681595
transform 1 0 18032 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1604681595
transform 1 0 17020 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_171
timestamp 1604681595
transform 1 0 16836 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_175
timestamp 1604681595
transform 1 0 17204 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_178
timestamp 1604681595
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1604681595
transform 1 0 19964 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1604681595
transform 1 0 18584 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_188
timestamp 1604681595
transform 1 0 18400 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_192
timestamp 1604681595
transform 1 0 18768 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_204
timestamp 1604681595
transform 1 0 19872 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_190
timestamp 1604681595
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_202
timestamp 1604681595
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_213
timestamp 1604681595
transform 1 0 20700 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_209
timestamp 1604681595
transform 1 0 20332 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1604681595
transform 1 0 20516 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1604681595
transform 1 0 21068 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_221
timestamp 1604681595
transform 1 0 21436 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1604681595
transform 1 0 21620 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_227
timestamp 1604681595
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_215
timestamp 1604681595
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_225
timestamp 1604681595
transform 1 0 21804 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_237
timestamp 1604681595
transform 1 0 22908 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_243
timestamp 1604681595
transform 1 0 23460 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_245
timestamp 1604681595
transform 1 0 23644 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_239
timestamp 1604681595
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1604681595
transform 1 0 24196 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1604681595
transform 1 0 25576 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1604681595
transform 1 0 24748 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_255
timestamp 1604681595
transform 1 0 24564 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_259
timestamp 1604681595
transform 1 0 24932 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_265
timestamp 1604681595
transform 1 0 25484 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_270
timestamp 1604681595
transform 1 0 25944 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_251
timestamp 1604681595
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_263
timestamp 1604681595
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1604681595
transform 1 0 26680 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1604681595
transform 1 0 27232 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1604681595
transform 1 0 26128 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_274
timestamp 1604681595
transform 1 0 26312 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_282
timestamp 1604681595
transform 1 0 27048 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_286
timestamp 1604681595
transform 1 0 27416 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_276
timestamp 1604681595
transform 1 0 26496 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_288
timestamp 1604681595
transform 1 0 27600 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 28888 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 28888 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_298
timestamp 1604681595
transform 1 0 28520 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_296
timestamp 1604681595
transform 1 0 28336 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1604681595
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 3956 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_27
timestamp 1604681595
transform 1 0 3588 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_32
timestamp 1604681595
transform 1 0 4048 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_44
timestamp 1604681595
transform 1 0 5152 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_56
timestamp 1604681595
transform 1 0 6256 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_63
timestamp 1604681595
transform 1 0 6900 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_75
timestamp 1604681595
transform 1 0 8004 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 9660 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_87
timestamp 1604681595
transform 1 0 9108 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_94
timestamp 1604681595
transform 1 0 9752 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 12512 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_106
timestamp 1604681595
transform 1 0 10856 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_118
timestamp 1604681595
transform 1 0 11960 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1604681595
transform 1 0 12604 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1604681595
transform 1 0 13708 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 15364 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_149
timestamp 1604681595
transform 1 0 14812 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_156
timestamp 1604681595
transform 1 0 15456 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 18216 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_168
timestamp 1604681595
transform 1 0 16560 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_180
timestamp 1604681595
transform 1 0 17664 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_187
timestamp 1604681595
transform 1 0 18308 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_199
timestamp 1604681595
transform 1 0 19412 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 21068 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_211
timestamp 1604681595
transform 1 0 20516 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_218
timestamp 1604681595
transform 1 0 21160 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 23920 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_230
timestamp 1604681595
transform 1 0 22264 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_242
timestamp 1604681595
transform 1 0 23368 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_249
timestamp 1604681595
transform 1 0 24012 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_261
timestamp 1604681595
transform 1 0 25116 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 26772 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1604681595
transform 1 0 26220 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_280
timestamp 1604681595
transform 1 0 26864 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 28888 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_292
timestamp 1604681595
transform 1 0 27968 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_298
timestamp 1604681595
transform 1 0 28520 0 1 21216
box -38 -48 130 592
<< labels >>
rlabel metal2 s 28354 0 28410 480 6 SC_IN_BOT
port 0 nsew default input
rlabel metal2 s 9678 23520 9734 24000 6 SC_IN_TOP
port 1 nsew default input
rlabel metal2 s 29366 0 29422 480 6 SC_OUT_BOT
port 2 nsew default tristate
rlabel metal2 s 11242 23520 11298 24000 6 SC_OUT_TOP
port 3 nsew default tristate
rlabel metal2 s 478 0 534 480 6 bottom_grid_pin_0_
port 4 nsew default tristate
rlabel metal2 s 5630 0 5686 480 6 bottom_grid_pin_10_
port 5 nsew default tristate
rlabel metal2 s 1490 0 1546 480 6 bottom_grid_pin_2_
port 6 nsew default tristate
rlabel metal2 s 2502 0 2558 480 6 bottom_grid_pin_4_
port 7 nsew default tristate
rlabel metal2 s 3514 0 3570 480 6 bottom_grid_pin_6_
port 8 nsew default tristate
rlabel metal2 s 4526 0 4582 480 6 bottom_grid_pin_8_
port 9 nsew default tristate
rlabel metal2 s 6642 0 6698 480 6 ccff_head
port 10 nsew default input
rlabel metal2 s 7654 0 7710 480 6 ccff_tail
port 11 nsew default tristate
rlabel metal3 s 0 12248 480 12368 6 chanx_left_in[0]
port 12 nsew default input
rlabel metal3 s 0 18232 480 18352 6 chanx_left_in[10]
port 13 nsew default input
rlabel metal3 s 0 18776 480 18896 6 chanx_left_in[11]
port 14 nsew default input
rlabel metal3 s 0 19320 480 19440 6 chanx_left_in[12]
port 15 nsew default input
rlabel metal3 s 0 20000 480 20120 6 chanx_left_in[13]
port 16 nsew default input
rlabel metal3 s 0 20544 480 20664 6 chanx_left_in[14]
port 17 nsew default input
rlabel metal3 s 0 21224 480 21344 6 chanx_left_in[15]
port 18 nsew default input
rlabel metal3 s 0 21768 480 21888 6 chanx_left_in[16]
port 19 nsew default input
rlabel metal3 s 0 22312 480 22432 6 chanx_left_in[17]
port 20 nsew default input
rlabel metal3 s 0 22992 480 23112 6 chanx_left_in[18]
port 21 nsew default input
rlabel metal3 s 0 23536 480 23656 6 chanx_left_in[19]
port 22 nsew default input
rlabel metal3 s 0 12792 480 12912 6 chanx_left_in[1]
port 23 nsew default input
rlabel metal3 s 0 13336 480 13456 6 chanx_left_in[2]
port 24 nsew default input
rlabel metal3 s 0 14016 480 14136 6 chanx_left_in[3]
port 25 nsew default input
rlabel metal3 s 0 14560 480 14680 6 chanx_left_in[4]
port 26 nsew default input
rlabel metal3 s 0 15240 480 15360 6 chanx_left_in[5]
port 27 nsew default input
rlabel metal3 s 0 15784 480 15904 6 chanx_left_in[6]
port 28 nsew default input
rlabel metal3 s 0 16328 480 16448 6 chanx_left_in[7]
port 29 nsew default input
rlabel metal3 s 0 17008 480 17128 6 chanx_left_in[8]
port 30 nsew default input
rlabel metal3 s 0 17552 480 17672 6 chanx_left_in[9]
port 31 nsew default input
rlabel metal3 s 0 280 480 400 6 chanx_left_out[0]
port 32 nsew default tristate
rlabel metal3 s 0 6264 480 6384 6 chanx_left_out[10]
port 33 nsew default tristate
rlabel metal3 s 0 6808 480 6928 6 chanx_left_out[11]
port 34 nsew default tristate
rlabel metal3 s 0 7352 480 7472 6 chanx_left_out[12]
port 35 nsew default tristate
rlabel metal3 s 0 8032 480 8152 6 chanx_left_out[13]
port 36 nsew default tristate
rlabel metal3 s 0 8576 480 8696 6 chanx_left_out[14]
port 37 nsew default tristate
rlabel metal3 s 0 9256 480 9376 6 chanx_left_out[15]
port 38 nsew default tristate
rlabel metal3 s 0 9800 480 9920 6 chanx_left_out[16]
port 39 nsew default tristate
rlabel metal3 s 0 10344 480 10464 6 chanx_left_out[17]
port 40 nsew default tristate
rlabel metal3 s 0 11024 480 11144 6 chanx_left_out[18]
port 41 nsew default tristate
rlabel metal3 s 0 11568 480 11688 6 chanx_left_out[19]
port 42 nsew default tristate
rlabel metal3 s 0 824 480 944 6 chanx_left_out[1]
port 43 nsew default tristate
rlabel metal3 s 0 1368 480 1488 6 chanx_left_out[2]
port 44 nsew default tristate
rlabel metal3 s 0 2048 480 2168 6 chanx_left_out[3]
port 45 nsew default tristate
rlabel metal3 s 0 2592 480 2712 6 chanx_left_out[4]
port 46 nsew default tristate
rlabel metal3 s 0 3272 480 3392 6 chanx_left_out[5]
port 47 nsew default tristate
rlabel metal3 s 0 3816 480 3936 6 chanx_left_out[6]
port 48 nsew default tristate
rlabel metal3 s 0 4360 480 4480 6 chanx_left_out[7]
port 49 nsew default tristate
rlabel metal3 s 0 5040 480 5160 6 chanx_left_out[8]
port 50 nsew default tristate
rlabel metal3 s 0 5584 480 5704 6 chanx_left_out[9]
port 51 nsew default tristate
rlabel metal3 s 29520 12248 30000 12368 6 chanx_right_in[0]
port 52 nsew default input
rlabel metal3 s 29520 18232 30000 18352 6 chanx_right_in[10]
port 53 nsew default input
rlabel metal3 s 29520 18776 30000 18896 6 chanx_right_in[11]
port 54 nsew default input
rlabel metal3 s 29520 19320 30000 19440 6 chanx_right_in[12]
port 55 nsew default input
rlabel metal3 s 29520 20000 30000 20120 6 chanx_right_in[13]
port 56 nsew default input
rlabel metal3 s 29520 20544 30000 20664 6 chanx_right_in[14]
port 57 nsew default input
rlabel metal3 s 29520 21224 30000 21344 6 chanx_right_in[15]
port 58 nsew default input
rlabel metal3 s 29520 21768 30000 21888 6 chanx_right_in[16]
port 59 nsew default input
rlabel metal3 s 29520 22312 30000 22432 6 chanx_right_in[17]
port 60 nsew default input
rlabel metal3 s 29520 22992 30000 23112 6 chanx_right_in[18]
port 61 nsew default input
rlabel metal3 s 29520 23536 30000 23656 6 chanx_right_in[19]
port 62 nsew default input
rlabel metal3 s 29520 12792 30000 12912 6 chanx_right_in[1]
port 63 nsew default input
rlabel metal3 s 29520 13336 30000 13456 6 chanx_right_in[2]
port 64 nsew default input
rlabel metal3 s 29520 14016 30000 14136 6 chanx_right_in[3]
port 65 nsew default input
rlabel metal3 s 29520 14560 30000 14680 6 chanx_right_in[4]
port 66 nsew default input
rlabel metal3 s 29520 15240 30000 15360 6 chanx_right_in[5]
port 67 nsew default input
rlabel metal3 s 29520 15784 30000 15904 6 chanx_right_in[6]
port 68 nsew default input
rlabel metal3 s 29520 16328 30000 16448 6 chanx_right_in[7]
port 69 nsew default input
rlabel metal3 s 29520 17008 30000 17128 6 chanx_right_in[8]
port 70 nsew default input
rlabel metal3 s 29520 17552 30000 17672 6 chanx_right_in[9]
port 71 nsew default input
rlabel metal3 s 29520 280 30000 400 6 chanx_right_out[0]
port 72 nsew default tristate
rlabel metal3 s 29520 6264 30000 6384 6 chanx_right_out[10]
port 73 nsew default tristate
rlabel metal3 s 29520 6808 30000 6928 6 chanx_right_out[11]
port 74 nsew default tristate
rlabel metal3 s 29520 7352 30000 7472 6 chanx_right_out[12]
port 75 nsew default tristate
rlabel metal3 s 29520 8032 30000 8152 6 chanx_right_out[13]
port 76 nsew default tristate
rlabel metal3 s 29520 8576 30000 8696 6 chanx_right_out[14]
port 77 nsew default tristate
rlabel metal3 s 29520 9256 30000 9376 6 chanx_right_out[15]
port 78 nsew default tristate
rlabel metal3 s 29520 9800 30000 9920 6 chanx_right_out[16]
port 79 nsew default tristate
rlabel metal3 s 29520 10344 30000 10464 6 chanx_right_out[17]
port 80 nsew default tristate
rlabel metal3 s 29520 11024 30000 11144 6 chanx_right_out[18]
port 81 nsew default tristate
rlabel metal3 s 29520 11568 30000 11688 6 chanx_right_out[19]
port 82 nsew default tristate
rlabel metal3 s 29520 824 30000 944 6 chanx_right_out[1]
port 83 nsew default tristate
rlabel metal3 s 29520 1368 30000 1488 6 chanx_right_out[2]
port 84 nsew default tristate
rlabel metal3 s 29520 2048 30000 2168 6 chanx_right_out[3]
port 85 nsew default tristate
rlabel metal3 s 29520 2592 30000 2712 6 chanx_right_out[4]
port 86 nsew default tristate
rlabel metal3 s 29520 3272 30000 3392 6 chanx_right_out[5]
port 87 nsew default tristate
rlabel metal3 s 29520 3816 30000 3936 6 chanx_right_out[6]
port 88 nsew default tristate
rlabel metal3 s 29520 4360 30000 4480 6 chanx_right_out[7]
port 89 nsew default tristate
rlabel metal3 s 29520 5040 30000 5160 6 chanx_right_out[8]
port 90 nsew default tristate
rlabel metal3 s 29520 5584 30000 5704 6 chanx_right_out[9]
port 91 nsew default tristate
rlabel metal2 s 9770 0 9826 480 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[0]
port 92 nsew default tristate
rlabel metal2 s 10782 0 10838 480 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[1]
port 93 nsew default tristate
rlabel metal2 s 11794 0 11850 480 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[2]
port 94 nsew default tristate
rlabel metal2 s 12806 0 12862 480 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[3]
port 95 nsew default tristate
rlabel metal2 s 13910 0 13966 480 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[4]
port 96 nsew default tristate
rlabel metal2 s 14922 0 14978 480 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[5]
port 97 nsew default tristate
rlabel metal2 s 15934 0 15990 480 6 gfpga_pad_EMBEDDED_IO_SOC_IN[0]
port 98 nsew default input
rlabel metal2 s 16946 0 17002 480 6 gfpga_pad_EMBEDDED_IO_SOC_IN[1]
port 99 nsew default input
rlabel metal2 s 18050 0 18106 480 6 gfpga_pad_EMBEDDED_IO_SOC_IN[2]
port 100 nsew default input
rlabel metal2 s 19062 0 19118 480 6 gfpga_pad_EMBEDDED_IO_SOC_IN[3]
port 101 nsew default input
rlabel metal2 s 20074 0 20130 480 6 gfpga_pad_EMBEDDED_IO_SOC_IN[4]
port 102 nsew default input
rlabel metal2 s 21086 0 21142 480 6 gfpga_pad_EMBEDDED_IO_SOC_IN[5]
port 103 nsew default input
rlabel metal2 s 22190 0 22246 480 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[0]
port 104 nsew default tristate
rlabel metal2 s 23202 0 23258 480 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[1]
port 105 nsew default tristate
rlabel metal2 s 24214 0 24270 480 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[2]
port 106 nsew default tristate
rlabel metal2 s 25226 0 25282 480 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[3]
port 107 nsew default tristate
rlabel metal2 s 26330 0 26386 480 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[4]
port 108 nsew default tristate
rlabel metal2 s 27342 0 27398 480 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[5]
port 109 nsew default tristate
rlabel metal2 s 8666 0 8722 480 6 prog_clk
port 110 nsew default input
rlabel metal2 s 12714 23520 12770 24000 6 top_width_0_height_0__pin_0_
port 111 nsew default input
rlabel metal2 s 20166 23520 20222 24000 6 top_width_0_height_0__pin_10_
port 112 nsew default input
rlabel metal2 s 29182 23520 29238 24000 6 top_width_0_height_0__pin_11_lower
port 113 nsew default tristate
rlabel metal2 s 8206 23520 8262 24000 6 top_width_0_height_0__pin_11_upper
port 114 nsew default tristate
rlabel metal2 s 21730 23520 21786 24000 6 top_width_0_height_0__pin_1_lower
port 115 nsew default tristate
rlabel metal2 s 754 23520 810 24000 6 top_width_0_height_0__pin_1_upper
port 116 nsew default tristate
rlabel metal2 s 14186 23520 14242 24000 6 top_width_0_height_0__pin_2_
port 117 nsew default input
rlabel metal2 s 23202 23520 23258 24000 6 top_width_0_height_0__pin_3_lower
port 118 nsew default tristate
rlabel metal2 s 2226 23520 2282 24000 6 top_width_0_height_0__pin_3_upper
port 119 nsew default tristate
rlabel metal2 s 15750 23520 15806 24000 6 top_width_0_height_0__pin_4_
port 120 nsew default input
rlabel metal2 s 24674 23520 24730 24000 6 top_width_0_height_0__pin_5_lower
port 121 nsew default tristate
rlabel metal2 s 3698 23520 3754 24000 6 top_width_0_height_0__pin_5_upper
port 122 nsew default tristate
rlabel metal2 s 17222 23520 17278 24000 6 top_width_0_height_0__pin_6_
port 123 nsew default input
rlabel metal2 s 26238 23520 26294 24000 6 top_width_0_height_0__pin_7_lower
port 124 nsew default tristate
rlabel metal2 s 5170 23520 5226 24000 6 top_width_0_height_0__pin_7_upper
port 125 nsew default tristate
rlabel metal2 s 18694 23520 18750 24000 6 top_width_0_height_0__pin_8_
port 126 nsew default input
rlabel metal2 s 27710 23520 27766 24000 6 top_width_0_height_0__pin_9_lower
port 127 nsew default tristate
rlabel metal2 s 6734 23520 6790 24000 6 top_width_0_height_0__pin_9_upper
port 128 nsew default tristate
rlabel metal4 s 5944 2128 6264 21808 6 VPWR
port 129 nsew default input
rlabel metal4 s 10944 2128 11264 21808 6 VGND
port 130 nsew default input
<< properties >>
string FIXED_BBOX 0 0 30000 24000
<< end >>
