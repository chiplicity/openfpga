magic
tech sky130A
magscale 1 2
timestamp 1608156581
<< obsli1 >>
rect 1104 2159 21620 20145
<< obsm1 >>
rect 198 1300 22158 21140
<< metal2 >>
rect 202 22000 258 22800
rect 570 22000 626 22800
rect 1030 22000 1086 22800
rect 1398 22000 1454 22800
rect 1858 22000 1914 22800
rect 2226 22000 2282 22800
rect 2686 22000 2742 22800
rect 3146 22000 3202 22800
rect 3514 22000 3570 22800
rect 3974 22000 4030 22800
rect 4342 22000 4398 22800
rect 4802 22000 4858 22800
rect 5262 22000 5318 22800
rect 5630 22000 5686 22800
rect 6090 22000 6146 22800
rect 6458 22000 6514 22800
rect 6918 22000 6974 22800
rect 7378 22000 7434 22800
rect 7746 22000 7802 22800
rect 8206 22000 8262 22800
rect 8574 22000 8630 22800
rect 9034 22000 9090 22800
rect 9494 22000 9550 22800
rect 9862 22000 9918 22800
rect 10322 22000 10378 22800
rect 10690 22000 10746 22800
rect 11150 22000 11206 22800
rect 11610 22000 11666 22800
rect 11978 22000 12034 22800
rect 12438 22000 12494 22800
rect 12806 22000 12862 22800
rect 13266 22000 13322 22800
rect 13634 22000 13690 22800
rect 14094 22000 14150 22800
rect 14554 22000 14610 22800
rect 14922 22000 14978 22800
rect 15382 22000 15438 22800
rect 15750 22000 15806 22800
rect 16210 22000 16266 22800
rect 16670 22000 16726 22800
rect 17038 22000 17094 22800
rect 17498 22000 17554 22800
rect 17866 22000 17922 22800
rect 18326 22000 18382 22800
rect 18786 22000 18842 22800
rect 19154 22000 19210 22800
rect 19614 22000 19670 22800
rect 19982 22000 20038 22800
rect 20442 22000 20498 22800
rect 20902 22000 20958 22800
rect 21270 22000 21326 22800
rect 21730 22000 21786 22800
rect 22098 22000 22154 22800
rect 22558 22000 22614 22800
rect 2226 0 2282 800
rect 6734 0 6790 800
rect 11334 0 11390 800
rect 15842 0 15898 800
rect 20442 0 20498 800
<< obsm2 >>
rect 314 21944 514 22545
rect 682 21944 974 22545
rect 1142 21944 1342 22545
rect 1510 21944 1802 22545
rect 1970 21944 2170 22545
rect 2338 21944 2630 22545
rect 2798 21944 3090 22545
rect 3258 21944 3458 22545
rect 3626 21944 3918 22545
rect 4086 21944 4286 22545
rect 4454 21944 4746 22545
rect 4914 21944 5206 22545
rect 5374 21944 5574 22545
rect 5742 21944 6034 22545
rect 6202 21944 6402 22545
rect 6570 21944 6862 22545
rect 7030 21944 7322 22545
rect 7490 21944 7690 22545
rect 7858 21944 8150 22545
rect 8318 21944 8518 22545
rect 8686 21944 8978 22545
rect 9146 21944 9438 22545
rect 9606 21944 9806 22545
rect 9974 21944 10266 22545
rect 10434 21944 10634 22545
rect 10802 21944 11094 22545
rect 11262 21944 11554 22545
rect 11722 21944 11922 22545
rect 12090 21944 12382 22545
rect 12550 21944 12750 22545
rect 12918 21944 13210 22545
rect 13378 21944 13578 22545
rect 13746 21944 14038 22545
rect 14206 21944 14498 22545
rect 14666 21944 14866 22545
rect 15034 21944 15326 22545
rect 15494 21944 15694 22545
rect 15862 21944 16154 22545
rect 16322 21944 16614 22545
rect 16782 21944 16982 22545
rect 17150 21944 17442 22545
rect 17610 21944 17810 22545
rect 17978 21944 18270 22545
rect 18438 21944 18730 22545
rect 18898 21944 19098 22545
rect 19266 21944 19558 22545
rect 19726 21944 19926 22545
rect 20094 21944 20386 22545
rect 20554 21944 20846 22545
rect 21014 21944 21214 22545
rect 21382 21944 21674 22545
rect 21842 21944 22042 22545
rect 22210 21944 22502 22545
rect 204 856 22600 21944
rect 204 167 2170 856
rect 2338 167 6678 856
rect 6846 167 11278 856
rect 11446 167 15786 856
rect 15954 167 20386 856
rect 20554 167 22600 856
<< metal3 >>
rect 0 22448 800 22568
rect 22000 22448 22800 22568
rect 0 22040 800 22160
rect 22000 22040 22800 22160
rect 0 21496 800 21616
rect 22000 21496 22800 21616
rect 0 21088 800 21208
rect 22000 21088 22800 21208
rect 0 20544 800 20664
rect 22000 20544 22800 20664
rect 0 20136 800 20256
rect 22000 20136 22800 20256
rect 0 19728 800 19848
rect 22000 19728 22800 19848
rect 0 19184 800 19304
rect 22000 19184 22800 19304
rect 0 18776 800 18896
rect 22000 18776 22800 18896
rect 0 18232 800 18352
rect 22000 18232 22800 18352
rect 0 17824 800 17944
rect 22000 17824 22800 17944
rect 0 17280 800 17400
rect 22000 17280 22800 17400
rect 0 16872 800 16992
rect 22000 16872 22800 16992
rect 0 16464 800 16584
rect 22000 16464 22800 16584
rect 0 15920 800 16040
rect 22000 15920 22800 16040
rect 0 15512 800 15632
rect 22000 15512 22800 15632
rect 0 14968 800 15088
rect 22000 14968 22800 15088
rect 0 14560 800 14680
rect 22000 14560 22800 14680
rect 0 14016 800 14136
rect 22000 14016 22800 14136
rect 0 13608 800 13728
rect 22000 13608 22800 13728
rect 0 13200 800 13320
rect 22000 13200 22800 13320
rect 0 12656 800 12776
rect 22000 12656 22800 12776
rect 0 12248 800 12368
rect 22000 12248 22800 12368
rect 0 11704 800 11824
rect 22000 11704 22800 11824
rect 0 11296 800 11416
rect 22000 11296 22800 11416
rect 0 10752 800 10872
rect 22000 10752 22800 10872
rect 0 10344 800 10464
rect 22000 10344 22800 10464
rect 0 9936 800 10056
rect 22000 9936 22800 10056
rect 0 9392 800 9512
rect 22000 9392 22800 9512
rect 0 8984 800 9104
rect 22000 8984 22800 9104
rect 0 8440 800 8560
rect 22000 8440 22800 8560
rect 0 8032 800 8152
rect 22000 8032 22800 8152
rect 0 7488 800 7608
rect 22000 7488 22800 7608
rect 0 7080 800 7200
rect 22000 7080 22800 7200
rect 0 6672 800 6792
rect 22000 6672 22800 6792
rect 0 6128 800 6248
rect 22000 6128 22800 6248
rect 0 5720 800 5840
rect 22000 5720 22800 5840
rect 0 5176 800 5296
rect 22000 5176 22800 5296
rect 0 4768 800 4888
rect 22000 4768 22800 4888
rect 0 4224 800 4344
rect 22000 4224 22800 4344
rect 0 3816 800 3936
rect 22000 3816 22800 3936
rect 0 3408 800 3528
rect 22000 3408 22800 3528
rect 0 2864 800 2984
rect 22000 2864 22800 2984
rect 0 2456 800 2576
rect 22000 2456 22800 2576
rect 0 1912 800 2032
rect 22000 1912 22800 2032
rect 0 1504 800 1624
rect 22000 1504 22800 1624
rect 0 960 800 1080
rect 22000 960 22800 1080
rect 0 552 800 672
rect 22000 552 22800 672
rect 0 144 800 264
rect 22000 144 22800 264
<< obsm3 >>
rect 880 22368 21920 22541
rect 798 22240 22000 22368
rect 880 21960 21920 22240
rect 798 21696 22000 21960
rect 880 21416 21920 21696
rect 798 21288 22000 21416
rect 880 21008 21920 21288
rect 798 20744 22000 21008
rect 880 20464 21920 20744
rect 798 20336 22000 20464
rect 880 20056 21920 20336
rect 798 19928 22000 20056
rect 880 19648 21920 19928
rect 798 19384 22000 19648
rect 880 19104 21920 19384
rect 798 18976 22000 19104
rect 880 18696 21920 18976
rect 798 18432 22000 18696
rect 880 18152 21920 18432
rect 798 18024 22000 18152
rect 880 17744 21920 18024
rect 798 17480 22000 17744
rect 880 17200 21920 17480
rect 798 17072 22000 17200
rect 880 16792 21920 17072
rect 798 16664 22000 16792
rect 880 16384 21920 16664
rect 798 16120 22000 16384
rect 880 15840 21920 16120
rect 798 15712 22000 15840
rect 880 15432 21920 15712
rect 798 15168 22000 15432
rect 880 14888 21920 15168
rect 798 14760 22000 14888
rect 880 14480 21920 14760
rect 798 14216 22000 14480
rect 880 13936 21920 14216
rect 798 13808 22000 13936
rect 880 13528 21920 13808
rect 798 13400 22000 13528
rect 880 13120 21920 13400
rect 798 12856 22000 13120
rect 880 12576 21920 12856
rect 798 12448 22000 12576
rect 880 12168 21920 12448
rect 798 11904 22000 12168
rect 880 11624 21920 11904
rect 798 11496 22000 11624
rect 880 11216 21920 11496
rect 798 10952 22000 11216
rect 880 10672 21920 10952
rect 798 10544 22000 10672
rect 880 10264 21920 10544
rect 798 10136 22000 10264
rect 880 9856 21920 10136
rect 798 9592 22000 9856
rect 880 9312 21920 9592
rect 798 9184 22000 9312
rect 880 8904 21920 9184
rect 798 8640 22000 8904
rect 880 8360 21920 8640
rect 798 8232 22000 8360
rect 880 7952 21920 8232
rect 798 7688 22000 7952
rect 880 7408 21920 7688
rect 798 7280 22000 7408
rect 880 7000 21920 7280
rect 798 6872 22000 7000
rect 880 6592 21920 6872
rect 798 6328 22000 6592
rect 880 6048 21920 6328
rect 798 5920 22000 6048
rect 880 5640 21920 5920
rect 798 5376 22000 5640
rect 880 5096 21920 5376
rect 798 4968 22000 5096
rect 880 4688 21920 4968
rect 798 4424 22000 4688
rect 880 4144 21920 4424
rect 798 4016 22000 4144
rect 880 3736 21920 4016
rect 798 3608 22000 3736
rect 880 3328 21920 3608
rect 798 3064 22000 3328
rect 880 2784 21920 3064
rect 798 2656 22000 2784
rect 880 2376 21920 2656
rect 798 2112 22000 2376
rect 880 1832 21920 2112
rect 798 1704 22000 1832
rect 880 1424 21920 1704
rect 798 1160 22000 1424
rect 880 880 21920 1160
rect 798 752 22000 880
rect 880 472 21920 752
rect 798 344 22000 472
rect 880 171 21920 344
<< metal4 >>
rect 4376 2128 4696 20176
rect 7808 2128 8128 20176
<< obsm4 >>
rect 11099 2128 19261 20176
<< labels >>
rlabel metal2 s 202 22000 258 22800 6 SC_IN_TOP
port 1 nsew default input
rlabel metal2 s 22558 22000 22614 22800 6 SC_OUT_TOP
port 2 nsew default output
rlabel metal2 s 4342 22000 4398 22800 6 Test_en_N_out
port 3 nsew default output
rlabel metal2 s 20442 0 20498 800 6 Test_en_S_in
port 4 nsew default input
rlabel metal2 s 2226 0 2282 800 6 ccff_head
port 5 nsew default input
rlabel metal2 s 6734 0 6790 800 6 ccff_tail
port 6 nsew default output
rlabel metal3 s 0 4224 800 4344 6 chanx_left_in[0]
port 7 nsew default input
rlabel metal3 s 0 8984 800 9104 6 chanx_left_in[10]
port 8 nsew default input
rlabel metal3 s 0 9392 800 9512 6 chanx_left_in[11]
port 9 nsew default input
rlabel metal3 s 0 9936 800 10056 6 chanx_left_in[12]
port 10 nsew default input
rlabel metal3 s 0 10344 800 10464 6 chanx_left_in[13]
port 11 nsew default input
rlabel metal3 s 0 10752 800 10872 6 chanx_left_in[14]
port 12 nsew default input
rlabel metal3 s 0 11296 800 11416 6 chanx_left_in[15]
port 13 nsew default input
rlabel metal3 s 0 11704 800 11824 6 chanx_left_in[16]
port 14 nsew default input
rlabel metal3 s 0 12248 800 12368 6 chanx_left_in[17]
port 15 nsew default input
rlabel metal3 s 0 12656 800 12776 6 chanx_left_in[18]
port 16 nsew default input
rlabel metal3 s 0 13200 800 13320 6 chanx_left_in[19]
port 17 nsew default input
rlabel metal3 s 0 4768 800 4888 6 chanx_left_in[1]
port 18 nsew default input
rlabel metal3 s 0 5176 800 5296 6 chanx_left_in[2]
port 19 nsew default input
rlabel metal3 s 0 5720 800 5840 6 chanx_left_in[3]
port 20 nsew default input
rlabel metal3 s 0 6128 800 6248 6 chanx_left_in[4]
port 21 nsew default input
rlabel metal3 s 0 6672 800 6792 6 chanx_left_in[5]
port 22 nsew default input
rlabel metal3 s 0 7080 800 7200 6 chanx_left_in[6]
port 23 nsew default input
rlabel metal3 s 0 7488 800 7608 6 chanx_left_in[7]
port 24 nsew default input
rlabel metal3 s 0 8032 800 8152 6 chanx_left_in[8]
port 25 nsew default input
rlabel metal3 s 0 8440 800 8560 6 chanx_left_in[9]
port 26 nsew default input
rlabel metal3 s 0 13608 800 13728 6 chanx_left_out[0]
port 27 nsew default output
rlabel metal3 s 0 18232 800 18352 6 chanx_left_out[10]
port 28 nsew default output
rlabel metal3 s 0 18776 800 18896 6 chanx_left_out[11]
port 29 nsew default output
rlabel metal3 s 0 19184 800 19304 6 chanx_left_out[12]
port 30 nsew default output
rlabel metal3 s 0 19728 800 19848 6 chanx_left_out[13]
port 31 nsew default output
rlabel metal3 s 0 20136 800 20256 6 chanx_left_out[14]
port 32 nsew default output
rlabel metal3 s 0 20544 800 20664 6 chanx_left_out[15]
port 33 nsew default output
rlabel metal3 s 0 21088 800 21208 6 chanx_left_out[16]
port 34 nsew default output
rlabel metal3 s 0 21496 800 21616 6 chanx_left_out[17]
port 35 nsew default output
rlabel metal3 s 0 22040 800 22160 6 chanx_left_out[18]
port 36 nsew default output
rlabel metal3 s 0 22448 800 22568 6 chanx_left_out[19]
port 37 nsew default output
rlabel metal3 s 0 14016 800 14136 6 chanx_left_out[1]
port 38 nsew default output
rlabel metal3 s 0 14560 800 14680 6 chanx_left_out[2]
port 39 nsew default output
rlabel metal3 s 0 14968 800 15088 6 chanx_left_out[3]
port 40 nsew default output
rlabel metal3 s 0 15512 800 15632 6 chanx_left_out[4]
port 41 nsew default output
rlabel metal3 s 0 15920 800 16040 6 chanx_left_out[5]
port 42 nsew default output
rlabel metal3 s 0 16464 800 16584 6 chanx_left_out[6]
port 43 nsew default output
rlabel metal3 s 0 16872 800 16992 6 chanx_left_out[7]
port 44 nsew default output
rlabel metal3 s 0 17280 800 17400 6 chanx_left_out[8]
port 45 nsew default output
rlabel metal3 s 0 17824 800 17944 6 chanx_left_out[9]
port 46 nsew default output
rlabel metal3 s 22000 4224 22800 4344 6 chanx_right_in[0]
port 47 nsew default input
rlabel metal3 s 22000 8984 22800 9104 6 chanx_right_in[10]
port 48 nsew default input
rlabel metal3 s 22000 9392 22800 9512 6 chanx_right_in[11]
port 49 nsew default input
rlabel metal3 s 22000 9936 22800 10056 6 chanx_right_in[12]
port 50 nsew default input
rlabel metal3 s 22000 10344 22800 10464 6 chanx_right_in[13]
port 51 nsew default input
rlabel metal3 s 22000 10752 22800 10872 6 chanx_right_in[14]
port 52 nsew default input
rlabel metal3 s 22000 11296 22800 11416 6 chanx_right_in[15]
port 53 nsew default input
rlabel metal3 s 22000 11704 22800 11824 6 chanx_right_in[16]
port 54 nsew default input
rlabel metal3 s 22000 12248 22800 12368 6 chanx_right_in[17]
port 55 nsew default input
rlabel metal3 s 22000 12656 22800 12776 6 chanx_right_in[18]
port 56 nsew default input
rlabel metal3 s 22000 13200 22800 13320 6 chanx_right_in[19]
port 57 nsew default input
rlabel metal3 s 22000 4768 22800 4888 6 chanx_right_in[1]
port 58 nsew default input
rlabel metal3 s 22000 5176 22800 5296 6 chanx_right_in[2]
port 59 nsew default input
rlabel metal3 s 22000 5720 22800 5840 6 chanx_right_in[3]
port 60 nsew default input
rlabel metal3 s 22000 6128 22800 6248 6 chanx_right_in[4]
port 61 nsew default input
rlabel metal3 s 22000 6672 22800 6792 6 chanx_right_in[5]
port 62 nsew default input
rlabel metal3 s 22000 7080 22800 7200 6 chanx_right_in[6]
port 63 nsew default input
rlabel metal3 s 22000 7488 22800 7608 6 chanx_right_in[7]
port 64 nsew default input
rlabel metal3 s 22000 8032 22800 8152 6 chanx_right_in[8]
port 65 nsew default input
rlabel metal3 s 22000 8440 22800 8560 6 chanx_right_in[9]
port 66 nsew default input
rlabel metal3 s 22000 13608 22800 13728 6 chanx_right_out[0]
port 67 nsew default output
rlabel metal3 s 22000 18232 22800 18352 6 chanx_right_out[10]
port 68 nsew default output
rlabel metal3 s 22000 18776 22800 18896 6 chanx_right_out[11]
port 69 nsew default output
rlabel metal3 s 22000 19184 22800 19304 6 chanx_right_out[12]
port 70 nsew default output
rlabel metal3 s 22000 19728 22800 19848 6 chanx_right_out[13]
port 71 nsew default output
rlabel metal3 s 22000 20136 22800 20256 6 chanx_right_out[14]
port 72 nsew default output
rlabel metal3 s 22000 20544 22800 20664 6 chanx_right_out[15]
port 73 nsew default output
rlabel metal3 s 22000 21088 22800 21208 6 chanx_right_out[16]
port 74 nsew default output
rlabel metal3 s 22000 21496 22800 21616 6 chanx_right_out[17]
port 75 nsew default output
rlabel metal3 s 22000 22040 22800 22160 6 chanx_right_out[18]
port 76 nsew default output
rlabel metal3 s 22000 22448 22800 22568 6 chanx_right_out[19]
port 77 nsew default output
rlabel metal3 s 22000 14016 22800 14136 6 chanx_right_out[1]
port 78 nsew default output
rlabel metal3 s 22000 14560 22800 14680 6 chanx_right_out[2]
port 79 nsew default output
rlabel metal3 s 22000 14968 22800 15088 6 chanx_right_out[3]
port 80 nsew default output
rlabel metal3 s 22000 15512 22800 15632 6 chanx_right_out[4]
port 81 nsew default output
rlabel metal3 s 22000 15920 22800 16040 6 chanx_right_out[5]
port 82 nsew default output
rlabel metal3 s 22000 16464 22800 16584 6 chanx_right_out[6]
port 83 nsew default output
rlabel metal3 s 22000 16872 22800 16992 6 chanx_right_out[7]
port 84 nsew default output
rlabel metal3 s 22000 17280 22800 17400 6 chanx_right_out[8]
port 85 nsew default output
rlabel metal3 s 22000 17824 22800 17944 6 chanx_right_out[9]
port 86 nsew default output
rlabel metal2 s 5630 22000 5686 22800 6 chany_top_in[0]
port 87 nsew default input
rlabel metal2 s 9862 22000 9918 22800 6 chany_top_in[10]
port 88 nsew default input
rlabel metal2 s 10322 22000 10378 22800 6 chany_top_in[11]
port 89 nsew default input
rlabel metal2 s 10690 22000 10746 22800 6 chany_top_in[12]
port 90 nsew default input
rlabel metal2 s 11150 22000 11206 22800 6 chany_top_in[13]
port 91 nsew default input
rlabel metal2 s 11610 22000 11666 22800 6 chany_top_in[14]
port 92 nsew default input
rlabel metal2 s 11978 22000 12034 22800 6 chany_top_in[15]
port 93 nsew default input
rlabel metal2 s 12438 22000 12494 22800 6 chany_top_in[16]
port 94 nsew default input
rlabel metal2 s 12806 22000 12862 22800 6 chany_top_in[17]
port 95 nsew default input
rlabel metal2 s 13266 22000 13322 22800 6 chany_top_in[18]
port 96 nsew default input
rlabel metal2 s 13634 22000 13690 22800 6 chany_top_in[19]
port 97 nsew default input
rlabel metal2 s 6090 22000 6146 22800 6 chany_top_in[1]
port 98 nsew default input
rlabel metal2 s 6458 22000 6514 22800 6 chany_top_in[2]
port 99 nsew default input
rlabel metal2 s 6918 22000 6974 22800 6 chany_top_in[3]
port 100 nsew default input
rlabel metal2 s 7378 22000 7434 22800 6 chany_top_in[4]
port 101 nsew default input
rlabel metal2 s 7746 22000 7802 22800 6 chany_top_in[5]
port 102 nsew default input
rlabel metal2 s 8206 22000 8262 22800 6 chany_top_in[6]
port 103 nsew default input
rlabel metal2 s 8574 22000 8630 22800 6 chany_top_in[7]
port 104 nsew default input
rlabel metal2 s 9034 22000 9090 22800 6 chany_top_in[8]
port 105 nsew default input
rlabel metal2 s 9494 22000 9550 22800 6 chany_top_in[9]
port 106 nsew default input
rlabel metal2 s 14094 22000 14150 22800 6 chany_top_out[0]
port 107 nsew default output
rlabel metal2 s 18326 22000 18382 22800 6 chany_top_out[10]
port 108 nsew default output
rlabel metal2 s 18786 22000 18842 22800 6 chany_top_out[11]
port 109 nsew default output
rlabel metal2 s 19154 22000 19210 22800 6 chany_top_out[12]
port 110 nsew default output
rlabel metal2 s 19614 22000 19670 22800 6 chany_top_out[13]
port 111 nsew default output
rlabel metal2 s 19982 22000 20038 22800 6 chany_top_out[14]
port 112 nsew default output
rlabel metal2 s 20442 22000 20498 22800 6 chany_top_out[15]
port 113 nsew default output
rlabel metal2 s 20902 22000 20958 22800 6 chany_top_out[16]
port 114 nsew default output
rlabel metal2 s 21270 22000 21326 22800 6 chany_top_out[17]
port 115 nsew default output
rlabel metal2 s 21730 22000 21786 22800 6 chany_top_out[18]
port 116 nsew default output
rlabel metal2 s 22098 22000 22154 22800 6 chany_top_out[19]
port 117 nsew default output
rlabel metal2 s 14554 22000 14610 22800 6 chany_top_out[1]
port 118 nsew default output
rlabel metal2 s 14922 22000 14978 22800 6 chany_top_out[2]
port 119 nsew default output
rlabel metal2 s 15382 22000 15438 22800 6 chany_top_out[3]
port 120 nsew default output
rlabel metal2 s 15750 22000 15806 22800 6 chany_top_out[4]
port 121 nsew default output
rlabel metal2 s 16210 22000 16266 22800 6 chany_top_out[5]
port 122 nsew default output
rlabel metal2 s 16670 22000 16726 22800 6 chany_top_out[6]
port 123 nsew default output
rlabel metal2 s 17038 22000 17094 22800 6 chany_top_out[7]
port 124 nsew default output
rlabel metal2 s 17498 22000 17554 22800 6 chany_top_out[8]
port 125 nsew default output
rlabel metal2 s 17866 22000 17922 22800 6 chany_top_out[9]
port 126 nsew default output
rlabel metal2 s 4802 22000 4858 22800 6 clk_3_N_out
port 127 nsew default output
rlabel metal2 s 15842 0 15898 800 6 clk_3_S_in
port 128 nsew default input
rlabel metal3 s 0 2456 800 2576 6 left_bottom_grid_pin_11_
port 129 nsew default input
rlabel metal3 s 0 2864 800 2984 6 left_bottom_grid_pin_13_
port 130 nsew default input
rlabel metal3 s 0 3408 800 3528 6 left_bottom_grid_pin_15_
port 131 nsew default input
rlabel metal3 s 0 3816 800 3936 6 left_bottom_grid_pin_17_
port 132 nsew default input
rlabel metal3 s 0 144 800 264 6 left_bottom_grid_pin_1_
port 133 nsew default input
rlabel metal3 s 0 552 800 672 6 left_bottom_grid_pin_3_
port 134 nsew default input
rlabel metal3 s 0 960 800 1080 6 left_bottom_grid_pin_5_
port 135 nsew default input
rlabel metal3 s 0 1504 800 1624 6 left_bottom_grid_pin_7_
port 136 nsew default input
rlabel metal3 s 0 1912 800 2032 6 left_bottom_grid_pin_9_
port 137 nsew default input
rlabel metal2 s 3974 22000 4030 22800 6 prog_clk_0_N_in
port 138 nsew default input
rlabel metal2 s 5262 22000 5318 22800 6 prog_clk_3_N_out
port 139 nsew default output
rlabel metal2 s 11334 0 11390 800 6 prog_clk_3_S_in
port 140 nsew default input
rlabel metal3 s 22000 2456 22800 2576 6 right_bottom_grid_pin_11_
port 141 nsew default input
rlabel metal3 s 22000 2864 22800 2984 6 right_bottom_grid_pin_13_
port 142 nsew default input
rlabel metal3 s 22000 3408 22800 3528 6 right_bottom_grid_pin_15_
port 143 nsew default input
rlabel metal3 s 22000 3816 22800 3936 6 right_bottom_grid_pin_17_
port 144 nsew default input
rlabel metal3 s 22000 144 22800 264 6 right_bottom_grid_pin_1_
port 145 nsew default input
rlabel metal3 s 22000 552 22800 672 6 right_bottom_grid_pin_3_
port 146 nsew default input
rlabel metal3 s 22000 960 22800 1080 6 right_bottom_grid_pin_5_
port 147 nsew default input
rlabel metal3 s 22000 1504 22800 1624 6 right_bottom_grid_pin_7_
port 148 nsew default input
rlabel metal3 s 22000 1912 22800 2032 6 right_bottom_grid_pin_9_
port 149 nsew default input
rlabel metal2 s 570 22000 626 22800 6 top_left_grid_pin_42_
port 150 nsew default input
rlabel metal2 s 1030 22000 1086 22800 6 top_left_grid_pin_43_
port 151 nsew default input
rlabel metal2 s 1398 22000 1454 22800 6 top_left_grid_pin_44_
port 152 nsew default input
rlabel metal2 s 1858 22000 1914 22800 6 top_left_grid_pin_45_
port 153 nsew default input
rlabel metal2 s 2226 22000 2282 22800 6 top_left_grid_pin_46_
port 154 nsew default input
rlabel metal2 s 2686 22000 2742 22800 6 top_left_grid_pin_47_
port 155 nsew default input
rlabel metal2 s 3146 22000 3202 22800 6 top_left_grid_pin_48_
port 156 nsew default input
rlabel metal2 s 3514 22000 3570 22800 6 top_left_grid_pin_49_
port 157 nsew default input
rlabel metal4 s 4376 2128 4696 20176 6 VPWR
port 158 nsew power input
rlabel metal4 s 7808 2128 8128 20176 6 VGND
port 159 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 22800 22800
string LEFview TRUE
<< end >>
