* NGSPICE file created from sb_1__1_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand2_4 abstract view
.subckt scs8hd_nand2_4 A B Y vgnd vpwr
.ends

.subckt sb_1__1_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] bottom_left_grid_pin_13_ bottom_right_grid_pin_11_ chanx_left_in[0] chanx_left_in[1]
+ chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6]
+ chanx_left_in[7] chanx_left_in[8] chanx_left_out[0] chanx_left_out[1] chanx_left_out[2]
+ chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7]
+ chanx_left_out[8] chanx_right_in[0] chanx_right_in[1] chanx_right_in[2] chanx_right_in[3]
+ chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7] chanx_right_in[8]
+ chanx_right_out[0] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4]
+ chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chany_bottom_in[0]
+ chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5]
+ chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_out[0] chany_bottom_out[1]
+ chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5]
+ chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8] chany_top_in[0] chany_top_in[1]
+ chany_top_in[2] chany_top_in[3] chany_top_in[4] chany_top_in[5] chany_top_in[6]
+ chany_top_in[7] chany_top_in[8] chany_top_out[0] chany_top_out[1] chany_top_out[2]
+ chany_top_out[3] chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7]
+ chany_top_out[8] data_in enable left_bottom_grid_pin_12_ left_top_grid_pin_10_ right_bottom_grid_pin_12_
+ right_top_grid_pin_10_ top_left_grid_pin_13_ top_right_grid_pin_11_ vpwr vgnd
XFILLER_39_233 vgnd vpwr scs8hd_decap_4
XFILLER_39_222 vgnd vpwr scs8hd_decap_4
XFILLER_22_133 vgnd vpwr scs8hd_fill_1
XFILLER_7_7 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[4] mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_100 vpwr vgnd scs8hd_fill_2
XFILLER_9_137 vpwr vgnd scs8hd_fill_2
XFILLER_13_144 vpwr vgnd scs8hd_fill_2
XFILLER_13_199 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__113__B _045_/Y vgnd vpwr scs8hd_diode_2
XFILLER_36_236 vgnd vpwr scs8hd_decap_12
XFILLER_36_203 vgnd vpwr scs8hd_decap_8
XFILLER_3_89 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_11_ mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_left_track_1.LATCH_6_.latch data_in mem_left_track_1.LATCH_6_.latch/Q _116_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_158 vgnd vpwr scs8hd_fill_1
XFILLER_12_10 vpwr vgnd scs8hd_fill_2
XFILLER_12_32 vgnd vpwr scs8hd_decap_3
XFILLER_12_65 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB _138_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_258 vgnd vpwr scs8hd_decap_12
XANTENNA__108__B _104_/X vgnd vpwr scs8hd_diode_2
XANTENNA__124__A _124_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_173 vpwr vgnd scs8hd_fill_2
XFILLER_5_151 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_184 vgnd vpwr scs8hd_decap_4
XFILLER_24_228 vgnd vpwr scs8hd_decap_4
XFILLER_24_206 vgnd vpwr scs8hd_decap_6
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _161_/HI mem_bottom_track_17.LATCH_2_.latch/Q
+ mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_track_1.LATCH_4_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
X_200_ chany_bottom_in[6] chany_top_out[7] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_right_track_16.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_131_ _094_/A _129_/B _131_/Y vgnd vpwr scs8hd_nor2_4
X_062_ _064_/A _092_/A _062_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_53 vpwr vgnd scs8hd_fill_2
XFILLER_2_154 vpwr vgnd scs8hd_fill_2
XFILLER_0_79 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__119__A _059_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_11 vpwr vgnd scs8hd_fill_2
XFILLER_9_44 vpwr vgnd scs8hd_fill_2
XFILLER_9_99 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _194_/A vgnd vpwr scs8hd_inv_1
Xmem_bottom_track_17.LATCH_2_.latch data_in mem_bottom_track_17.LATCH_2_.latch/Q _150_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_209 vgnd vpwr scs8hd_decap_3
XFILLER_20_253 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_34_41 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB _062_/Y vgnd vpwr scs8hd_diode_2
X_114_ address[4] _139_/B _139_/C _114_/D _121_/B vgnd vpwr scs8hd_or4_4
XFILLER_7_257 vgnd vpwr scs8hd_decap_12
X_045_ address[6] _045_/Y vgnd vpwr scs8hd_inv_8
Xmux_left_track_9.INVTX1_3_.scs8hd_inv_1 chanx_right_in[1] mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__121__B _121_/B vgnd vpwr scs8hd_diode_2
XFILLER_38_106 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_track_16.LATCH_4_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_9.INVTX1_6_.scs8hd_inv_1 chanx_left_in[2] mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_0.LATCH_5_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_2_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_37_161 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.INVTX1_7_.scs8hd_inv_1 chanx_left_in[7] mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__116__B _121_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__132__A _046_/Y vgnd vpwr scs8hd_diode_2
XFILLER_13_3 vgnd vpwr scs8hd_fill_1
XFILLER_19_150 vpwr vgnd scs8hd_fill_2
Xmem_right_track_8.LATCH_1_.latch data_in mem_right_track_8.LATCH_1_.latch/Q _093_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__042__A address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_208 vpwr vgnd scs8hd_fill_2
XFILLER_25_164 vpwr vgnd scs8hd_fill_2
XFILLER_17_109 vpwr vgnd scs8hd_fill_2
XFILLER_40_145 vgnd vpwr scs8hd_decap_8
XFILLER_31_53 vgnd vpwr scs8hd_decap_4
XFILLER_25_197 vpwr vgnd scs8hd_fill_2
XFILLER_0_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.LATCH_4_.latch_SLEEPB _127_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__127__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_186 vpwr vgnd scs8hd_fill_2
XFILLER_16_197 vgnd vpwr scs8hd_decap_4
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_212 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_39_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _161_/HI vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_145 vgnd vpwr scs8hd_decap_8
XFILLER_9_116 vpwr vgnd scs8hd_fill_2
XFILLER_13_123 vgnd vpwr scs8hd_decap_4
XFILLER_42_63 vgnd vpwr scs8hd_decap_12
XFILLER_3_35 vgnd vpwr scs8hd_decap_3
Xmux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_8_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_6_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_36_248 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.INVTX1_3_.scs8hd_inv_1 chanx_right_in[7] mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_204 vpwr vgnd scs8hd_fill_2
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_248 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_12_88 vpwr vgnd scs8hd_fill_2
XFILLER_37_96 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_204 vpwr vgnd scs8hd_fill_2
XFILLER_26_270 vgnd vpwr scs8hd_decap_4
XANTENNA__124__B _129_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_3_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__140__A _126_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_8.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[0] mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_32_273 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__050__A address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.LATCH_6_.latch data_in mem_top_track_8.LATCH_6_.latch/Q _069_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_0.LATCH_6_.latch data_in mem_right_track_0.LATCH_6_.latch/Q _078_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_130_ _064_/B _129_/B _130_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 _171_/HI mem_top_track_8.LATCH_7_.latch/Q
+ mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_15_218 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_061_ address[2] _059_/B address[0] _092_/A vgnd vpwr scs8hd_or3_4
XANTENNA_mem_right_track_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_2_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__119__B _121_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_2_.latch/Q mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_23 vpwr vgnd scs8hd_fill_2
XANTENNA__135__A _059_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_6_.latch_SLEEPB _097_/Y vgnd vpwr scs8hd_diode_2
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
XANTENNA__045__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_18_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_32 vgnd vpwr scs8hd_fill_1
XFILLER_34_75 vgnd vpwr scs8hd_decap_6
X_113_ address[5] _045_/Y _114_/D vgnd vpwr scs8hd_or2_4
X_044_ address[0] _063_/C vgnd vpwr scs8hd_inv_8
XANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB _122_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[6] mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_37_195 vgnd vpwr scs8hd_decap_6
XFILLER_37_140 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1_A bottom_right_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_8_.scs8hd_inv_1 chanx_left_in[8] mux_top_track_8.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_4_239 vgnd vpwr scs8hd_decap_12
XFILLER_20_77 vpwr vgnd scs8hd_fill_2
XFILLER_20_88 vpwr vgnd scs8hd_fill_2
XFILLER_29_75 vpwr vgnd scs8hd_fill_2
XFILLER_29_20 vpwr vgnd scs8hd_fill_2
XFILLER_28_173 vpwr vgnd scs8hd_fill_2
XANTENNA__132__B address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB _145_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_173 vpwr vgnd scs8hd_fill_2
XFILLER_19_195 vgnd vpwr scs8hd_fill_1
XFILLER_34_198 vgnd vpwr scs8hd_decap_8
XFILLER_34_165 vgnd vpwr scs8hd_decap_3
XFILLER_34_143 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_121 vgnd vpwr scs8hd_fill_1
XFILLER_31_21 vpwr vgnd scs8hd_fill_2
XFILLER_15_88 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_3_.latch/Q mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_275 vpwr vgnd scs8hd_fill_2
XFILLER_16_121 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__127__B _129_/B vgnd vpwr scs8hd_diode_2
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_17.INVTX1_1_.scs8hd_inv_1 chany_top_in[5] mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__A _092_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_102 vpwr vgnd scs8hd_fill_2
XANTENNA__053__A _053_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_10 vpwr vgnd scs8hd_fill_2
XFILLER_26_87 vgnd vpwr scs8hd_decap_3
XFILLER_26_43 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_113 vpwr vgnd scs8hd_fill_2
XFILLER_13_157 vpwr vgnd scs8hd_fill_2
XFILLER_13_179 vpwr vgnd scs8hd_fill_2
XFILLER_42_75 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _190_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__138__A _094_/A vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.LATCH_7_.latch data_in mem_left_track_9.LATCH_7_.latch/Q _124_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_27_227 vpwr vgnd scs8hd_fill_2
XANTENNA__048__A enable vgnd vpwr scs8hd_diode_2
XFILLER_10_127 vpwr vgnd scs8hd_fill_2
XFILLER_12_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_75 vgnd vpwr scs8hd_decap_4
XFILLER_37_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__140__B _143_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_241 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.INVTX1_7_.scs8hd_inv_1 chanx_left_in[0] mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__050__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_23_252 vgnd vpwr scs8hd_decap_3
XFILLER_23_33 vpwr vgnd scs8hd_fill_2
X_060_ _064_/A _059_/X _060_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_99 vpwr vgnd scs8hd_fill_2
XFILLER_3_3 vgnd vpwr scs8hd_decap_12
XFILLER_0_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_37 vpwr vgnd scs8hd_fill_2
X_189_ _189_/A chanx_right_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_9_57 vpwr vgnd scs8hd_fill_2
XANTENNA__135__B _134_/B vgnd vpwr scs8hd_diode_2
XFILLER_36_3 vgnd vpwr scs8hd_decap_8
XANTENNA__151__A _064_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_2_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA__061__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_34_54 vpwr vgnd scs8hd_fill_2
XFILLER_34_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_55 vpwr vgnd scs8hd_fill_2
XFILLER_18_88 vpwr vgnd scs8hd_fill_2
X_043_ address[1] _059_/B vgnd vpwr scs8hd_inv_8
XFILLER_11_222 vpwr vgnd scs8hd_fill_2
XFILLER_11_233 vpwr vgnd scs8hd_fill_2
X_112_ _094_/A _104_/X _112_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__146__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_6_270 vgnd vpwr scs8hd_decap_4
XFILLER_37_174 vpwr vgnd scs8hd_fill_2
XANTENNA__056__A _064_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_8_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_6_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_23 vpwr vgnd scs8hd_fill_2
XFILLER_20_45 vpwr vgnd scs8hd_fill_2
XFILLER_6_36 vgnd vpwr scs8hd_fill_1
XFILLER_6_69 vgnd vpwr scs8hd_decap_6
XFILLER_20_6 vpwr vgnd scs8hd_fill_2
XANTENNA__132__C _139_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_177 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_158 vpwr vgnd scs8hd_fill_2
XFILLER_25_177 vgnd vpwr scs8hd_decap_4
XFILLER_25_111 vgnd vpwr scs8hd_decap_8
XFILLER_15_12 vpwr vgnd scs8hd_fill_2
XFILLER_31_99 vgnd vpwr scs8hd_decap_4
XFILLER_31_77 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A _160_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_144 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_8.LATCH_5_.latch_SLEEPB _089_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_31_147 vpwr vgnd scs8hd_fill_2
XFILLER_31_114 vpwr vgnd scs8hd_fill_2
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__B _143_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_114 vgnd vpwr scs8hd_fill_1
XANTENNA__053__B _059_/B vgnd vpwr scs8hd_diode_2
XFILLER_42_87 vgnd vpwr scs8hd_decap_6
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_3_48 vgnd vpwr scs8hd_fill_1
XFILLER_3_15 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.INVTX1_4_.scs8hd_inv_1 chanx_right_in[8] mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__138__B _134_/B vgnd vpwr scs8hd_diode_2
XANTENNA__154__A _126_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_180 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__064__A _064_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_46 vpwr vgnd scs8hd_fill_2
XFILLER_37_32 vpwr vgnd scs8hd_fill_2
XFILLER_41_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_228 vgnd vpwr scs8hd_decap_4
XFILLER_5_121 vgnd vpwr scs8hd_fill_1
Xmem_top_track_0.LATCH_0_.latch data_in mem_top_track_0.LATCH_0_.latch/Q _066_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_198 vgnd vpwr scs8hd_decap_12
XFILLER_5_132 vpwr vgnd scs8hd_fill_2
XANTENNA__149__A _059_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_32_253 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_track_17.LATCH_3_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_right_track_8.LATCH_7_.latch data_in mem_right_track_8.LATCH_7_.latch/Q _087_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_91 vgnd vpwr scs8hd_fill_1
XANTENNA__059__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_23_242 vpwr vgnd scs8hd_fill_2
XFILLER_23_78 vgnd vpwr scs8hd_decap_3
XFILLER_23_12 vpwr vgnd scs8hd_fill_2
XFILLER_2_102 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_17.LATCH_3_.latch data_in mem_left_track_17.LATCH_3_.latch/Q _156_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_69 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
X_188_ chanx_left_in[0] chanx_right_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_29_3 vpwr vgnd scs8hd_fill_2
XANTENNA__151__B _152_/B vgnd vpwr scs8hd_diode_2
XANTENNA__061__B _059_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_3_.latch/Q mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_23 vpwr vgnd scs8hd_fill_2
XFILLER_34_88 vpwr vgnd scs8hd_fill_2
XFILLER_18_78 vpwr vgnd scs8hd_fill_2
X_042_ address[2] _053_/A vgnd vpwr scs8hd_inv_8
XANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB _083_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
X_111_ _064_/B _104_/X _111_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_245 vpwr vgnd scs8hd_fill_2
XANTENNA__146__B address[3] vgnd vpwr scs8hd_diode_2
XFILLER_37_120 vpwr vgnd scs8hd_fill_2
XFILLER_29_109 vgnd vpwr scs8hd_fill_1
XFILLER_1_81 vpwr vgnd scs8hd_fill_2
XANTENNA__056__B _126_/A vgnd vpwr scs8hd_diode_2
XANTENNA__072__A _059_/X vgnd vpwr scs8hd_diode_2
XFILLER_29_44 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_88 vpwr vgnd scs8hd_fill_2
XFILLER_29_55 vgnd vpwr scs8hd_decap_4
XFILLER_28_186 vgnd vpwr scs8hd_decap_6
XFILLER_28_131 vpwr vgnd scs8hd_fill_2
XFILLER_6_15 vgnd vpwr scs8hd_decap_3
XFILLER_6_48 vgnd vpwr scs8hd_decap_8
XANTENNA__132__D _051_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__157__A _092_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_2_.latch data_in mem_bottom_track_1.LATCH_2_.latch/Q _101_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_25_123 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_3_.latch_SLEEPB _072_/Y vgnd vpwr scs8hd_diode_2
XFILLER_25_145 vpwr vgnd scs8hd_fill_2
XFILLER_15_35 vpwr vgnd scs8hd_fill_2
XFILLER_15_57 vpwr vgnd scs8hd_fill_2
XANTENNA__067__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_31_34 vpwr vgnd scs8hd_fill_2
XFILLER_0_200 vpwr vgnd scs8hd_fill_2
XFILLER_16_167 vpwr vgnd scs8hd_fill_2
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_259 vpwr vgnd scs8hd_fill_2
XFILLER_39_237 vgnd vpwr scs8hd_fill_1
XFILLER_39_204 vgnd vpwr scs8hd_decap_8
XFILLER_11_3 vpwr vgnd scs8hd_fill_2
XFILLER_22_126 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__053__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_30_192 vgnd vpwr scs8hd_fill_1
Xmem_left_track_1.LATCH_1_.latch data_in mem_left_track_1.LATCH_1_.latch/Q _121_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_78 vgnd vpwr scs8hd_decap_3
XFILLER_26_67 vpwr vgnd scs8hd_fill_2
XFILLER_26_23 vpwr vgnd scs8hd_fill_2
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XFILLER_3_27 vgnd vpwr scs8hd_decap_8
XANTENNA__154__B _153_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_163 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__064__B _064_/B vgnd vpwr scs8hd_diode_2
Xmem_right_track_16.LATCH_2_.latch data_in mem_right_track_16.LATCH_2_.latch/Q _143_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__080__A _118_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_12_69 vpwr vgnd scs8hd_fill_2
XFILLER_37_11 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_16.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_41_232 vgnd vpwr scs8hd_decap_12
XFILLER_37_99 vgnd vpwr scs8hd_fill_1
XFILLER_5_155 vpwr vgnd scs8hd_fill_2
XFILLER_5_177 vgnd vpwr scs8hd_decap_6
XANTENNA__149__B _152_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XFILLER_32_265 vgnd vpwr scs8hd_decap_8
XFILLER_32_210 vgnd vpwr scs8hd_decap_4
XFILLER_4_81 vpwr vgnd scs8hd_fill_2
XANTENNA__059__B _059_/B vgnd vpwr scs8hd_diode_2
XFILLER_23_210 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__075__A _094_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_158 vgnd vpwr scs8hd_decap_12
XFILLER_2_114 vgnd vpwr scs8hd_decap_12
XFILLER_9_15 vpwr vgnd scs8hd_fill_2
XFILLER_9_48 vpwr vgnd scs8hd_fill_2
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
X_187_ chanx_left_in[1] chanx_right_out[2] vgnd vpwr scs8hd_buf_2
Xmux_left_track_9.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_9.INVTX1_3_.scs8hd_inv_1 chanx_right_in[3] mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_224 vpwr vgnd scs8hd_fill_2
XANTENNA__061__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_34_23 vgnd vpwr scs8hd_decap_4
X_110_ _092_/A _104_/X _110_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_217 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__146__C _139_/C vgnd vpwr scs8hd_diode_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[6] mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_37_187 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__072__B _067_/X vgnd vpwr scs8hd_diode_2
XFILLER_28_154 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.LATCH_7_.latch_SLEEPB _105_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_220 vgnd vpwr scs8hd_decap_12
XFILLER_10_91 vgnd vpwr scs8hd_fill_1
XFILLER_13_7 vpwr vgnd scs8hd_fill_2
XFILLER_19_110 vpwr vgnd scs8hd_fill_2
XFILLER_19_132 vgnd vpwr scs8hd_decap_3
XFILLER_19_154 vpwr vgnd scs8hd_fill_2
XFILLER_34_157 vpwr vgnd scs8hd_fill_2
XFILLER_34_102 vgnd vpwr scs8hd_decap_8
XANTENNA__157__B _153_/X vgnd vpwr scs8hd_diode_2
XFILLER_19_187 vpwr vgnd scs8hd_fill_2
XANTENNA__173__A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB _130_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_105 vpwr vgnd scs8hd_fill_2
XANTENNA__083__A _064_/B vgnd vpwr scs8hd_diode_2
XANTENNA__067__B _139_/B vgnd vpwr scs8hd_diode_2
XFILLER_24_190 vgnd vpwr scs8hd_fill_1
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_7_92 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_13_ mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_127 vgnd vpwr scs8hd_fill_1
XANTENNA__078__A _116_/A vgnd vpwr scs8hd_diode_2
XFILLER_42_56 vgnd vpwr scs8hd_decap_6
XFILLER_21_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_90 vpwr vgnd scs8hd_fill_2
XFILLER_27_208 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__080__B _081_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_37_45 vpwr vgnd scs8hd_fill_2
XFILLER_18_208 vgnd vpwr scs8hd_decap_4
XFILLER_26_274 vgnd vpwr scs8hd_fill_1
XFILLER_26_241 vgnd vpwr scs8hd_decap_8
Xmem_right_track_0.LATCH_1_.latch data_in mem_right_track_0.LATCH_1_.latch/Q _083_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_top_track_8.LATCH_1_.latch data_in mem_top_track_8.LATCH_1_.latch/Q _074_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_263 vgnd vpwr scs8hd_decap_12
XANTENNA__181__A _181_/A vgnd vpwr scs8hd_diode_2
XANTENNA__059__C _063_/C vgnd vpwr scs8hd_diode_2
XANTENNA__075__B _067_/X vgnd vpwr scs8hd_diode_2
XANTENNA__091__A _059_/X vgnd vpwr scs8hd_diode_2
XFILLER_2_126 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_3_.latch_SLEEPB _100_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_27 vpwr vgnd scs8hd_fill_2
X_186_ chanx_left_in[2] chanx_right_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_1_181 vpwr vgnd scs8hd_fill_2
XFILLER_1_192 vgnd vpwr scs8hd_fill_1
XANTENNA__176__A _176_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.INVTX1_3_.scs8hd_inv_1 chanx_right_in[0] mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_bottom_track_1.INVTX1_6_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_36 vpwr vgnd scs8hd_fill_2
XFILLER_34_46 vpwr vgnd scs8hd_fill_2
XANTENNA__086__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_1_3 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[5] mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_169_ _169_/HI _169_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__146__D _114_/D vgnd vpwr scs8hd_diode_2
XFILLER_37_144 vpwr vgnd scs8hd_fill_2
XFILLER_1_72 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_24 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_28 vgnd vpwr scs8hd_fill_1
Xmux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_2_.latch/Q mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_232 vgnd vpwr scs8hd_decap_12
XFILLER_19_177 vgnd vpwr scs8hd_decap_6
XFILLER_42_180 vgnd vpwr scs8hd_decap_6
XFILLER_34_125 vgnd vpwr scs8hd_decap_3
Xmem_top_track_0.LATCH_6_.latch data_in mem_top_track_0.LATCH_6_.latch/Q _054_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmem_bottom_track_9.LATCH_3_.latch data_in mem_bottom_track_9.LATCH_3_.latch/Q _109_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__067__C _139_/C vgnd vpwr scs8hd_diode_2
XFILLER_33_180 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__083__B _081_/B vgnd vpwr scs8hd_diode_2
XFILLER_0_224 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_125 vpwr vgnd scs8hd_fill_2
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_track_0.LATCH_4_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_106 vpwr vgnd scs8hd_fill_2
XPHY_0 vgnd vpwr scs8hd_decap_3
XFILLER_30_150 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__184__A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.LATCH_2_.latch data_in mem_left_track_9.LATCH_2_.latch/Q _129_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_7_71 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_3_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__078__B _081_/B vgnd vpwr scs8hd_diode_2
XANTENNA__094__A _094_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_47 vpwr vgnd scs8hd_fill_2
XFILLER_13_117 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_0.LATCH_7_.latch_SLEEPB _052_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_150 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.INVTX1_8_.scs8hd_inv_1 left_bottom_grid_pin_12_ mux_left_track_9.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_121 vpwr vgnd scs8hd_fill_2
XFILLER_12_150 vgnd vpwr scs8hd_decap_3
XFILLER_8_198 vpwr vgnd scs8hd_fill_2
XANTENNA__179__A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_12_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.LATCH_4_.latch_SLEEPB _148_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_57 vpwr vgnd scs8hd_fill_2
XANTENNA__089__A _126_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[1] mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_top_track_16.LATCH_3_.latch data_in mem_top_track_16.LATCH_3_.latch/Q _135_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_41_245 vgnd vpwr scs8hd_decap_12
XFILLER_5_168 vgnd vpwr scs8hd_decap_3
XFILLER_5_113 vgnd vpwr scs8hd_decap_6
XFILLER_17_231 vgnd vpwr scs8hd_fill_1
XFILLER_17_242 vpwr vgnd scs8hd_fill_2
XFILLER_17_275 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_190 vgnd vpwr scs8hd_decap_12
XFILLER_23_234 vpwr vgnd scs8hd_fill_2
XFILLER_23_223 vpwr vgnd scs8hd_fill_2
XFILLER_23_201 vpwr vgnd scs8hd_fill_2
XFILLER_23_37 vpwr vgnd scs8hd_fill_2
XANTENNA__091__B _094_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
X_185_ _185_/A chanx_right_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_13_81 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA__192__A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_20_259 vgnd vpwr scs8hd_decap_12
XANTENNA__086__B address[3] vgnd vpwr scs8hd_diode_2
XFILLER_18_59 vpwr vgnd scs8hd_fill_2
XFILLER_34_58 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_8_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_11_226 vpwr vgnd scs8hd_fill_2
XFILLER_11_237 vpwr vgnd scs8hd_fill_2
Xmem_left_track_1.LATCH_7_.latch data_in mem_left_track_1.LATCH_7_.latch/Q _115_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_track_0.INVTX1_8_.scs8hd_inv_1 chanx_left_in[4] mux_top_track_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_168_ _168_/HI _168_/LO vgnd vpwr scs8hd_conb_1
XFILLER_24_80 vgnd vpwr scs8hd_fill_1
XFILLER_6_274 vgnd vpwr scs8hd_fill_1
XFILLER_27_3 vpwr vgnd scs8hd_fill_2
X_099_ _118_/A _095_/X _099_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_37_178 vpwr vgnd scs8hd_fill_2
XFILLER_37_123 vgnd vpwr scs8hd_decap_4
XFILLER_1_51 vgnd vpwr scs8hd_decap_8
XFILLER_1_62 vgnd vpwr scs8hd_decap_3
XANTENNA__187__A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_8_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_6_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_27 vpwr vgnd scs8hd_fill_2
XANTENNA__097__A _116_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_93 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_8.LATCH_2_.latch_SLEEPB _092_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_16 vpwr vgnd scs8hd_fill_2
XANTENNA__067__D _051_/D vgnd vpwr scs8hd_diode_2
XFILLER_31_59 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_17.LATCH_3_.latch data_in mem_bottom_track_17.LATCH_3_.latch/Q _149_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_31_118 vpwr vgnd scs8hd_fill_2
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_229 vpwr vgnd scs8hd_fill_2
XFILLER_39_218 vpwr vgnd scs8hd_fill_2
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_30_184 vgnd vpwr scs8hd_decap_8
XFILLER_38_251 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.INVTX1_1_.scs8hd_inv_1 chany_top_in[6] mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__094__B _094_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_5_.latch_SLEEPB _117_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_173 vpwr vgnd scs8hd_fill_2
XFILLER_32_80 vgnd vpwr scs8hd_decap_3
XFILLER_8_133 vgnd vpwr scs8hd_fill_1
XFILLER_8_188 vgnd vpwr scs8hd_fill_1
XFILLER_12_184 vpwr vgnd scs8hd_fill_2
XFILLER_35_232 vpwr vgnd scs8hd_fill_2
XANTENNA__195__A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA__089__B _094_/B vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_track_1.LATCH_5_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmem_right_track_8.LATCH_2_.latch data_in mem_right_track_8.LATCH_2_.latch/Q _092_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
XFILLER_26_210 vpwr vgnd scs8hd_fill_2
XFILLER_41_257 vgnd vpwr scs8hd_decap_12
XFILLER_5_136 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_5_.latch_SLEEPB _140_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_210 vpwr vgnd scs8hd_fill_2
XFILLER_32_224 vpwr vgnd scs8hd_fill_2
XFILLER_4_62 vgnd vpwr scs8hd_decap_4
XFILLER_23_257 vgnd vpwr scs8hd_decap_12
XFILLER_23_16 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_2_.latch/Q mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_139 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[8] mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[5] mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_202 vpwr vgnd scs8hd_fill_2
XFILLER_14_224 vpwr vgnd scs8hd_fill_2
XFILLER_14_235 vgnd vpwr scs8hd_decap_12
X_184_ chanx_left_in[4] chanx_right_out[5] vgnd vpwr scs8hd_buf_2
Xmux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_track_16.LATCH_5_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_60 vgnd vpwr scs8hd_fill_1
XFILLER_29_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_8_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_6_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_right_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_3_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_9.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_27 vpwr vgnd scs8hd_fill_2
XANTENNA__086__C _139_/C vgnd vpwr scs8hd_diode_2
XFILLER_11_205 vpwr vgnd scs8hd_fill_2
XFILLER_11_249 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_167_ _167_/HI _167_/LO vgnd vpwr scs8hd_conb_1
X_098_ _126_/A _095_/X _098_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_260 vgnd vpwr scs8hd_decap_12
XFILLER_37_113 vgnd vpwr scs8hd_fill_1
XFILLER_37_157 vpwr vgnd scs8hd_fill_2
XFILLER_1_85 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_102 vpwr vgnd scs8hd_fill_2
XANTENNA__097__B _095_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.LATCH_3_.latch_SLEEPB _156_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB _075_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_72 vgnd vpwr scs8hd_fill_1
XFILLER_10_83 vpwr vgnd scs8hd_fill_2
Xmem_right_track_0.LATCH_7_.latch data_in mem_right_track_0.LATCH_7_.latch/Q _077_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.LATCH_7_.latch data_in mem_top_track_8.LATCH_7_.latch/Q _068_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_19_70 vpwr vgnd scs8hd_fill_2
XFILLER_19_92 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__198__A _198_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_119 vpwr vgnd scs8hd_fill_2
XFILLER_33_160 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_127 vgnd vpwr scs8hd_decap_3
XFILLER_15_39 vgnd vpwr scs8hd_decap_3
XFILLER_18_190 vgnd vpwr scs8hd_fill_1
XFILLER_31_38 vgnd vpwr scs8hd_decap_4
XFILLER_0_259 vpwr vgnd scs8hd_fill_2
XFILLER_0_204 vgnd vpwr scs8hd_decap_12
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _170_/HI mem_top_track_16.LATCH_2_.latch/Q
+ mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 _165_/HI mem_left_track_9.LATCH_7_.latch/Q
+ mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_21_71 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_2_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_38_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_26_27 vpwr vgnd scs8hd_fill_2
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XFILLER_21_141 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_263 vgnd vpwr scs8hd_decap_12
XFILLER_29_252 vpwr vgnd scs8hd_fill_2
XFILLER_29_230 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _164_/HI mem_left_track_17.LATCH_2_.latch/Q
+ mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_16_82 vpwr vgnd scs8hd_fill_2
XFILLER_16_93 vpwr vgnd scs8hd_fill_2
XFILLER_8_145 vgnd vpwr scs8hd_decap_6
XFILLER_12_163 vgnd vpwr scs8hd_decap_3
XFILLER_35_211 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_3_.latch/Q mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_92 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.tap_buf4_0_.scs8hd_inv_1 mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _180_/A vgnd vpwr scs8hd_inv_1
XFILLER_4_85 vgnd vpwr scs8hd_decap_6
XFILLER_4_41 vpwr vgnd scs8hd_fill_2
XFILLER_23_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_19 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_9.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_247 vgnd vpwr scs8hd_decap_12
X_183_ chanx_left_in[5] chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_13_72 vgnd vpwr scs8hd_decap_3
XFILLER_1_184 vgnd vpwr scs8hd_decap_8
XFILLER_38_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_206 vgnd vpwr scs8hd_decap_6
XFILLER_20_228 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__086__D _139_/D vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_track_17.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
X_097_ _116_/A _095_/X _097_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_272 vgnd vpwr scs8hd_decap_3
X_166_ _166_/HI _166_/LO vgnd vpwr scs8hd_conb_1
XFILLER_34_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.LATCH_4_.latch_SLEEPB _108_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.INVTX1_8_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_28_169 vpwr vgnd scs8hd_fill_2
XFILLER_28_158 vpwr vgnd scs8hd_fill_2
XFILLER_28_114 vpwr vgnd scs8hd_fill_2
XFILLER_36_191 vgnd vpwr scs8hd_decap_4
XFILLER_3_257 vgnd vpwr scs8hd_decap_12
XFILLER_10_51 vgnd vpwr scs8hd_decap_3
XFILLER_19_114 vpwr vgnd scs8hd_fill_2
XFILLER_35_81 vpwr vgnd scs8hd_fill_2
XFILLER_34_139 vpwr vgnd scs8hd_fill_2
XFILLER_19_169 vpwr vgnd scs8hd_fill_2
X_149_ _059_/X _152_/B _149_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_40_109 vgnd vpwr scs8hd_decap_8
XFILLER_33_172 vpwr vgnd scs8hd_fill_2
XFILLER_31_17 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_29 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_249 vgnd vpwr scs8hd_decap_6
XFILLER_0_216 vgnd vpwr scs8hd_fill_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_106 vgnd vpwr scs8hd_decap_12
XFILLER_24_183 vgnd vpwr scs8hd_decap_4
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_21_83 vgnd vpwr scs8hd_decap_3
XFILLER_21_50 vpwr vgnd scs8hd_fill_2
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_15_150 vpwr vgnd scs8hd_fill_2
XFILLER_7_52 vgnd vpwr scs8hd_decap_6
XFILLER_7_96 vgnd vpwr scs8hd_decap_4
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XFILLER_21_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_6_.latch_SLEEPB _078_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_275 vpwr vgnd scs8hd_fill_2
XFILLER_16_50 vpwr vgnd scs8hd_fill_2
XFILLER_16_61 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_197 vpwr vgnd scs8hd_fill_2
XFILLER_35_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_49 vpwr vgnd scs8hd_fill_2
XFILLER_5_105 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_234 vgnd vpwr scs8hd_decap_8
XFILLER_17_245 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB _103_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_248 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_270 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_1.INVTX1_3_.scs8hd_inv_1 chanx_right_in[5] mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_259 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_182_ chanx_left_in[6] chanx_right_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_13_62 vgnd vpwr scs8hd_fill_1
XFILLER_38_81 vpwr vgnd scs8hd_fill_2
XFILLER_1_130 vpwr vgnd scs8hd_fill_2
XFILLER_1_141 vpwr vgnd scs8hd_fill_2
XFILLER_1_196 vpwr vgnd scs8hd_fill_2
XANTENNA__100__A _059_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_241 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_2_.scs8hd_inv_1 chanx_right_in[6] mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 _160_/HI mem_bottom_track_1.LATCH_7_.latch/Q
+ mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_165_ _165_/HI _165_/LO vgnd vpwr scs8hd_conb_1
XFILLER_24_72 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB _136_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_93 vgnd vpwr scs8hd_decap_8
X_096_ _124_/A _095_/X _096_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_76 vgnd vpwr scs8hd_fill_1
Xmem_top_track_0.LATCH_1_.latch data_in mem_top_track_0.LATCH_1_.latch/Q _064_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_28 vgnd vpwr scs8hd_fill_1
XFILLER_28_148 vgnd vpwr scs8hd_decap_3
XFILLER_3_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_19_83 vpwr vgnd scs8hd_fill_2
XFILLER_19_137 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_148_ _118_/A _152_/B _148_/Y vgnd vpwr scs8hd_nor2_4
X_079_ _126_/A _081_/B _079_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_107 vpwr vgnd scs8hd_fill_2
XFILLER_33_184 vgnd vpwr scs8hd_decap_3
XFILLER_33_151 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_17.LATCH_4_.latch data_in mem_left_track_17.LATCH_4_.latch/Q _155_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_0_228 vgnd vpwr scs8hd_decap_12
XFILLER_24_151 vpwr vgnd scs8hd_fill_2
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_8.INVTX1_2_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_95 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB _058_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[0] mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_30_154 vpwr vgnd scs8hd_fill_2
XFILLER_30_121 vpwr vgnd scs8hd_fill_2
XPHY_4 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_9.INVTX1_8_.scs8hd_inv_1 chanx_left_in[8] mux_bottom_track_9.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_195 vpwr vgnd scs8hd_fill_2
XFILLER_7_31 vpwr vgnd scs8hd_fill_2
XFILLER_7_75 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_left_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_21_165 vpwr vgnd scs8hd_fill_2
XFILLER_8_125 vpwr vgnd scs8hd_fill_2
XFILLER_32_72 vpwr vgnd scs8hd_fill_2
XFILLER_32_50 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB _151_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_1_.scs8hd_inv_1 chany_top_in[6] mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__103__A _094_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_35_257 vgnd vpwr scs8hd_decap_12
XFILLER_35_224 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_track_17.LATCH_4_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_37_28 vpwr vgnd scs8hd_fill_2
XFILLER_26_224 vpwr vgnd scs8hd_fill_2
XFILLER_26_202 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_3_.latch data_in mem_bottom_track_1.LATCH_3_.latch/Q _100_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_40_271 vgnd vpwr scs8hd_decap_4
XFILLER_4_32 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_bottom_track_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_6_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_260 vgnd vpwr scs8hd_decap_12
XFILLER_23_238 vpwr vgnd scs8hd_fill_2
XFILLER_23_227 vpwr vgnd scs8hd_fill_2
XFILLER_23_205 vgnd vpwr scs8hd_decap_3
X_181_ _181_/A chanx_right_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_13_30 vpwr vgnd scs8hd_fill_2
XFILLER_1_120 vpwr vgnd scs8hd_fill_2
XFILLER_13_96 vpwr vgnd scs8hd_fill_2
XFILLER_38_93 vpwr vgnd scs8hd_fill_2
XFILLER_38_60 vgnd vpwr scs8hd_fill_1
Xmem_left_track_1.LATCH_2_.latch data_in mem_left_track_1.LATCH_2_.latch/Q _120_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__100__B _095_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[4] mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_34_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__201__A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_40 vpwr vgnd scs8hd_fill_2
Xmem_right_track_16.LATCH_3_.latch data_in mem_right_track_16.LATCH_3_.latch/Q _142_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_84 vpwr vgnd scs8hd_fill_2
X_164_ _164_/HI _164_/LO vgnd vpwr scs8hd_conb_1
X_095_ _139_/C _139_/D _046_/Y address[3] _095_/X vgnd vpwr scs8hd_or4_4
XFILLER_27_7 vgnd vpwr scs8hd_fill_1
XFILLER_37_116 vpwr vgnd scs8hd_fill_2
XANTENNA__111__A _064_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[4] mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_28_127 vpwr vgnd scs8hd_fill_2
XFILLER_10_75 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_119 vgnd vpwr scs8hd_decap_4
Xmux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_62 vgnd vpwr scs8hd_fill_1
XFILLER_35_94 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_147_ _126_/A _152_/B _147_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__106__A _116_/A vgnd vpwr scs8hd_diode_2
X_078_ _116_/A _081_/B _078_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_18_160 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_218 vpwr vgnd scs8hd_fill_2
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_30 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_track_16.LATCH_3_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mem_left_track_1.LATCH_2_.latch_SLEEPB _120_/Y vgnd vpwr scs8hd_diode_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_15_163 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_2_.latch/Q mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_1.INVTX1_8_.scs8hd_inv_1 left_top_grid_pin_10_ mux_left_track_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_177 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_104 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_left_track_17.LATCH_3_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__103__B _095_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_269 vgnd vpwr scs8hd_decap_8
XFILLER_35_236 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_16.LATCH_2_.latch_SLEEPB _143_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_26_258 vgnd vpwr scs8hd_decap_12
XANTENNA__204__A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_32_228 vgnd vpwr scs8hd_decap_4
XFILLER_32_206 vpwr vgnd scs8hd_fill_2
XFILLER_27_62 vpwr vgnd scs8hd_fill_2
XFILLER_27_40 vpwr vgnd scs8hd_fill_2
XFILLER_17_214 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.INVTX1_2_.scs8hd_inv_1 chany_top_in[7] mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__114__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_4_77 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.INVTX1_3_.scs8hd_inv_1 chanx_right_in[2] mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_2_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_31_272 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_206 vgnd vpwr scs8hd_decap_6
XFILLER_14_228 vgnd vpwr scs8hd_decap_4
X_180_ _180_/A chanx_left_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_53 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__109__A _059_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_210 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A _163_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_209 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_094_ _094_/A _094_/B _094_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_40_84 vgnd vpwr scs8hd_decap_8
XFILLER_40_73 vgnd vpwr scs8hd_decap_8
XFILLER_40_62 vgnd vpwr scs8hd_decap_8
X_163_ _163_/HI _163_/LO vgnd vpwr scs8hd_conb_1
XFILLER_6_213 vgnd vpwr scs8hd_fill_1
XFILLER_6_246 vgnd vpwr scs8hd_decap_12
XANTENNA__111__B _104_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_0.LATCH_2_.latch data_in mem_right_track_0.LATCH_2_.latch/Q _082_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB _159_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.LATCH_2_.latch data_in mem_top_track_8.LATCH_2_.latch/Q _073_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_28_106 vgnd vpwr scs8hd_decap_8
XFILLER_36_150 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_32 vgnd vpwr scs8hd_decap_3
XFILLER_10_87 vgnd vpwr scs8hd_decap_4
XFILLER_19_30 vpwr vgnd scs8hd_fill_2
XFILLER_35_40 vpwr vgnd scs8hd_fill_2
XFILLER_27_172 vgnd vpwr scs8hd_decap_4
Xmux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_96 vgnd vpwr scs8hd_fill_1
XFILLER_19_106 vpwr vgnd scs8hd_fill_2
XFILLER_35_62 vgnd vpwr scs8hd_decap_4
XANTENNA__122__A _094_/A vgnd vpwr scs8hd_diode_2
X_146_ address[4] address[3] _139_/C _114_/D _152_/B vgnd vpwr scs8hd_or4_4
XANTENNA__106__B _104_/X vgnd vpwr scs8hd_diode_2
X_077_ _124_/A _081_/B _077_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_32_6 vgnd vpwr scs8hd_decap_4
Xmux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__207__A _207_/A vgnd vpwr scs8hd_diode_2
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_75 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_15_120 vpwr vgnd scs8hd_fill_2
XFILLER_15_131 vpwr vgnd scs8hd_fill_2
XFILLER_15_175 vpwr vgnd scs8hd_fill_2
XFILLER_30_167 vgnd vpwr scs8hd_decap_8
XANTENNA__117__A _126_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_11 vgnd vpwr scs8hd_decap_4
X_129_ _092_/A _129_/B _129_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_21_145 vgnd vpwr scs8hd_decap_3
XFILLER_21_123 vgnd vpwr scs8hd_decap_3
XFILLER_21_112 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_track_9.LATCH_4_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_234 vpwr vgnd scs8hd_fill_2
XFILLER_29_212 vgnd vpwr scs8hd_decap_3
Xmux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_2_.latch/Q mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_42 vpwr vgnd scs8hd_fill_2
XFILLER_16_86 vpwr vgnd scs8hd_fill_2
XFILLER_32_85 vgnd vpwr scs8hd_decap_4
XFILLER_32_41 vgnd vpwr scs8hd_decap_3
Xmux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_2_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_top_track_0.LATCH_7_.latch data_in mem_top_track_0.LATCH_7_.latch/Q _052_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmem_bottom_track_9.LATCH_4_.latch data_in mem_bottom_track_9.LATCH_4_.latch/Q _108_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_27_96 vpwr vgnd scs8hd_fill_2
XFILLER_17_259 vpwr vgnd scs8hd_fill_2
XANTENNA__114__B _139_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__130__A _064_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_7_.latch_SLEEPB _087_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_174 vgnd vpwr scs8hd_decap_12
XFILLER_4_163 vpwr vgnd scs8hd_fill_2
XFILLER_4_45 vgnd vpwr scs8hd_decap_4
XFILLER_16_270 vgnd vpwr scs8hd_decap_4
Xmem_left_track_9.LATCH_3_.latch data_in mem_left_track_9.LATCH_3_.latch/Q _128_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__109__B _104_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_233 vgnd vpwr scs8hd_decap_8
XANTENNA__125__A _116_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_6_.scs8hd_inv_1 chanx_left_in[3] mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB _111_/Y vgnd vpwr scs8hd_diode_2
XFILLER_39_192 vgnd vpwr scs8hd_decap_12
XFILLER_39_181 vpwr vgnd scs8hd_fill_2
XFILLER_39_170 vgnd vpwr scs8hd_decap_8
Xmux_left_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_3_.latch/Q mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_53 vpwr vgnd scs8hd_fill_2
X_162_ _162_/HI _162_/LO vgnd vpwr scs8hd_conb_1
XFILLER_10_210 vgnd vpwr scs8hd_decap_4
X_093_ _064_/B _094_/B _093_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_258 vgnd vpwr scs8hd_decap_12
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
Xmem_top_track_16.LATCH_4_.latch data_in mem_top_track_16.LATCH_4_.latch/Q _134_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_68 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_195 vgnd vpwr scs8hd_fill_1
XFILLER_10_11 vgnd vpwr scs8hd_decap_3
XFILLER_19_42 vpwr vgnd scs8hd_fill_2
XFILLER_19_53 vpwr vgnd scs8hd_fill_2
XFILLER_19_118 vpwr vgnd scs8hd_fill_2
XFILLER_27_184 vgnd vpwr scs8hd_decap_3
XFILLER_27_162 vgnd vpwr scs8hd_fill_1
XFILLER_42_187 vgnd vpwr scs8hd_decap_12
X_145_ _094_/A _143_/B _145_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_track_0.LATCH_5_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__122__B _121_/B vgnd vpwr scs8hd_diode_2
X_076_ _046_/Y _139_/B _139_/C _051_/D _081_/B vgnd vpwr scs8hd_or4_4
XFILLER_33_198 vpwr vgnd scs8hd_fill_2
XFILLER_33_176 vgnd vpwr scs8hd_decap_4
XFILLER_18_173 vgnd vpwr scs8hd_decap_8
XFILLER_18_184 vgnd vpwr scs8hd_decap_6
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_121 vpwr vgnd scs8hd_fill_2
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_187 vgnd vpwr scs8hd_fill_1
XFILLER_24_154 vgnd vpwr scs8hd_decap_3
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_54 vgnd vpwr scs8hd_decap_4
XFILLER_30_102 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_0.LATCH_3_.latch_SLEEPB _081_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_7 vgnd vpwr scs8hd_decap_3
X_128_ _059_/X _129_/B _128_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__117__B _121_/B vgnd vpwr scs8hd_diode_2
XANTENNA__133__A _126_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_202 vgnd vpwr scs8hd_fill_1
X_059_ address[2] _059_/B _063_/C _059_/X vgnd vpwr scs8hd_or3_4
Xmux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_38_213 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_8.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__043__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_16_32 vgnd vpwr scs8hd_fill_1
XFILLER_16_65 vpwr vgnd scs8hd_fill_2
XFILLER_12_168 vgnd vpwr scs8hd_decap_3
XFILLER_20_190 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_1.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA__128__A _059_/X vgnd vpwr scs8hd_diode_2
XFILLER_11_190 vpwr vgnd scs8hd_fill_2
XFILLER_41_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_271 vgnd vpwr scs8hd_decap_4
XFILLER_5_109 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_5_.latch_SLEEPB _070_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_27_75 vpwr vgnd scs8hd_fill_2
XFILLER_27_53 vpwr vgnd scs8hd_fill_2
XFILLER_17_227 vgnd vpwr scs8hd_decap_4
XFILLER_17_249 vgnd vpwr scs8hd_decap_6
XFILLER_40_241 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.INVTX1_7_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__114__C _139_/C vgnd vpwr scs8hd_diode_2
XANTENNA__130__B _129_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_186 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_bottom_track_17.LATCH_4_.latch data_in mem_bottom_track_17.LATCH_4_.latch/Q _148_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_31_230 vpwr vgnd scs8hd_fill_2
XFILLER_22_274 vgnd vpwr scs8hd_fill_1
XFILLER_13_11 vpwr vgnd scs8hd_fill_2
XFILLER_13_77 vpwr vgnd scs8hd_fill_2
XFILLER_38_52 vgnd vpwr scs8hd_decap_8
XFILLER_38_41 vgnd vpwr scs8hd_decap_8
XFILLER_1_112 vgnd vpwr scs8hd_decap_8
XFILLER_1_145 vgnd vpwr scs8hd_decap_12
XFILLER_38_85 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__125__B _129_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_245 vgnd vpwr scs8hd_decap_12
XFILLER_13_252 vgnd vpwr scs8hd_decap_12
XANTENNA__141__A _118_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 _168_/HI mem_right_track_8.LATCH_7_.latch/Q
+ mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__051__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_24_76 vpwr vgnd scs8hd_fill_2
XFILLER_24_10 vpwr vgnd scs8hd_fill_2
XFILLER_6_215 vgnd vpwr scs8hd_decap_12
X_161_ _161_/HI _161_/LO vgnd vpwr scs8hd_conb_1
X_092_ _092_/A _094_/B _092_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_2_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_right_track_8.LATCH_3_.latch data_in mem_right_track_8.LATCH_3_.latch/Q _091_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__136__A _092_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_163 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__046__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_10_23 vpwr vgnd scs8hd_fill_2
XFILLER_10_56 vgnd vpwr scs8hd_decap_3
XFILLER_19_87 vgnd vpwr scs8hd_decap_3
XFILLER_42_111 vgnd vpwr scs8hd_decap_12
XFILLER_42_100 vgnd vpwr scs8hd_decap_8
XFILLER_35_53 vpwr vgnd scs8hd_fill_2
XFILLER_27_141 vgnd vpwr scs8hd_decap_3
XFILLER_42_199 vgnd vpwr scs8hd_decap_12
X_144_ _064_/B _143_/B _144_/Y vgnd vpwr scs8hd_nor2_4
X_075_ _094_/A _067_/X _075_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_7 vgnd vpwr scs8hd_decap_4
XFILLER_2_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_111 vpwr vgnd scs8hd_fill_2
XFILLER_18_6 vpwr vgnd scs8hd_fill_2
XFILLER_18_130 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB _064_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_2_.scs8hd_inv_1 chany_top_in[8] mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_166 vgnd vpwr scs8hd_decap_8
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_9.INVTX1_5_.scs8hd_inv_1 bottom_left_grid_pin_13_ mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_99 vpwr vgnd scs8hd_fill_2
XFILLER_30_125 vpwr vgnd scs8hd_fill_2
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_15_144 vgnd vpwr scs8hd_decap_4
XFILLER_15_199 vpwr vgnd scs8hd_fill_2
X_058_ _064_/A _118_/A _058_/Y vgnd vpwr scs8hd_nor2_4
X_127_ _118_/A _129_/B _127_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_bottom_track_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_46 vgnd vpwr scs8hd_decap_4
XANTENNA__133__B _134_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _198_/A vgnd vpwr scs8hd_inv_1
XFILLER_21_169 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.INVTX1_6_.scs8hd_inv_1 chanx_left_in[5] mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_8_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_6_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_12_125 vgnd vpwr scs8hd_fill_1
XFILLER_12_147 vgnd vpwr scs8hd_fill_1
XFILLER_32_76 vgnd vpwr scs8hd_fill_1
XFILLER_32_54 vgnd vpwr scs8hd_fill_1
XFILLER_8_129 vgnd vpwr scs8hd_decap_4
XFILLER_20_180 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_228 vpwr vgnd scs8hd_fill_2
XANTENNA__128__B _129_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_140 vpwr vgnd scs8hd_fill_2
XFILLER_11_180 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__144__A _064_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_195 vpwr vgnd scs8hd_fill_2
XFILLER_26_228 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_3_.latch/Q mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_left_track_9.LATCH_3_.latch_SLEEPB _128_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__054__A _064_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_21 vpwr vgnd scs8hd_fill_2
XFILLER_40_253 vpwr vgnd scs8hd_fill_2
XANTENNA__114__D _114_/D vgnd vpwr scs8hd_diode_2
XFILLER_4_143 vgnd vpwr scs8hd_decap_8
XFILLER_4_58 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 _169_/HI mem_top_track_0.LATCH_7_.latch/Q
+ mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__139__A address[4] vgnd vpwr scs8hd_diode_2
XANTENNA__049__A _053_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_45 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.INVTX1_2_.scs8hd_inv_1 chanx_right_in[5] mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_38_64 vpwr vgnd scs8hd_fill_2
XFILLER_1_157 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_257 vgnd vpwr scs8hd_decap_12
XFILLER_13_264 vgnd vpwr scs8hd_decap_12
XANTENNA__141__B _143_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__051__B address[3] vgnd vpwr scs8hd_diode_2
XFILLER_5_90 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A _169_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.INVTX1_3_.scs8hd_inv_1 right_bottom_grid_pin_12_ mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_091_ _059_/X _094_/B _091_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_24_88 vpwr vgnd scs8hd_fill_2
X_160_ _160_/HI _160_/LO vgnd vpwr scs8hd_conb_1
XFILLER_6_205 vgnd vpwr scs8hd_decap_8
XFILLER_6_227 vgnd vpwr scs8hd_decap_12
XFILLER_37_109 vgnd vpwr scs8hd_decap_4
XFILLER_1_15 vgnd vpwr scs8hd_decap_12
XANTENNA__136__B _134_/B vgnd vpwr scs8hd_diode_2
XANTENNA__152__A _094_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_142 vgnd vpwr scs8hd_decap_8
XANTENNA__062__A _064_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_208 vgnd vpwr scs8hd_decap_12
XFILLER_10_68 vgnd vpwr scs8hd_decap_4
XFILLER_10_79 vpwr vgnd scs8hd_fill_2
XFILLER_19_66 vpwr vgnd scs8hd_fill_2
XFILLER_42_156 vgnd vpwr scs8hd_decap_12
XFILLER_42_123 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_1.LATCH_5_.latch_SLEEPB _098_/Y vgnd vpwr scs8hd_diode_2
X_143_ _092_/A _143_/B _143_/Y vgnd vpwr scs8hd_nor2_4
X_074_ _064_/B _067_/X _074_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_134 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_33_156 vgnd vpwr scs8hd_decap_4
XANTENNA__147__A _126_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_3_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_2_91 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[2] mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__057__A _053_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_145 vgnd vpwr scs8hd_decap_4
XFILLER_24_134 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.INVTX1_8_.scs8hd_inv_1 chanx_left_in[7] mux_bottom_track_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_34 vpwr vgnd scs8hd_fill_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_15_123 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_17.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_167 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_16.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_126_ _126_/A _129_/B _126_/Y vgnd vpwr scs8hd_nor2_4
X_057_ _053_/A address[1] address[0] _118_/A vgnd vpwr scs8hd_or3_4
XFILLER_7_58 vgnd vpwr scs8hd_fill_1
Xmux_top_track_8.INVTX1_7_.scs8hd_inv_1 chanx_left_in[6] mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_38_215 vgnd vpwr scs8hd_decap_12
XFILLER_30_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.INVTX1_8_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_2_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_21_137 vpwr vgnd scs8hd_fill_2
XFILLER_29_259 vpwr vgnd scs8hd_fill_2
XFILLER_29_248 vpwr vgnd scs8hd_fill_2
XFILLER_29_226 vpwr vgnd scs8hd_fill_2
XFILLER_16_12 vpwr vgnd scs8hd_fill_2
XFILLER_16_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A _166_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_108 vpwr vgnd scs8hd_fill_2
XFILLER_12_104 vpwr vgnd scs8hd_fill_2
XFILLER_12_115 vpwr vgnd scs8hd_fill_2
XFILLER_16_78 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_207 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__144__B _143_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_163 vpwr vgnd scs8hd_fill_2
X_109_ _059_/X _104_/X _109_/Y vgnd vpwr scs8hd_nor2_4
Xmux_left_track_17.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__054__B _116_/A vgnd vpwr scs8hd_diode_2
XANTENNA__070__A _126_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
XFILLER_4_122 vpwr vgnd scs8hd_fill_2
XFILLER_4_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_276 vgnd vpwr scs8hd_fill_1
XANTENNA__139__B _139_/B vgnd vpwr scs8hd_diode_2
XANTENNA__155__A _118_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__049__B _059_/B vgnd vpwr scs8hd_diode_2
XANTENNA__065__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_13_57 vgnd vpwr scs8hd_fill_1
XFILLER_1_169 vgnd vpwr scs8hd_decap_12
XFILLER_9_214 vpwr vgnd scs8hd_fill_2
XFILLER_13_276 vgnd vpwr scs8hd_fill_1
XFILLER_9_269 vgnd vpwr scs8hd_decap_8
XANTENNA__051__C _139_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_23 vpwr vgnd scs8hd_fill_2
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
X_090_ _118_/A _094_/B _090_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_239 vgnd vpwr scs8hd_decap_4
XFILLER_10_224 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[7] mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_3 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_27 vgnd vpwr scs8hd_decap_12
XANTENNA__152__B _152_/B vgnd vpwr scs8hd_diode_2
XFILLER_36_198 vpwr vgnd scs8hd_fill_2
XFILLER_36_121 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__062__B _092_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_12 vpwr vgnd scs8hd_fill_2
XFILLER_35_11 vpwr vgnd scs8hd_fill_2
XFILLER_27_176 vgnd vpwr scs8hd_fill_1
XFILLER_27_132 vgnd vpwr scs8hd_decap_3
Xmux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_34 vpwr vgnd scs8hd_fill_2
XFILLER_42_168 vgnd vpwr scs8hd_decap_12
XFILLER_35_99 vpwr vgnd scs8hd_fill_2
XFILLER_35_77 vpwr vgnd scs8hd_fill_2
X_142_ _059_/X _143_/B _142_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_073_ _092_/A _067_/X _073_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__147__B _152_/B vgnd vpwr scs8hd_diode_2
XFILLER_18_154 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_0.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_102 vpwr vgnd scs8hd_fill_2
XFILLER_2_81 vpwr vgnd scs8hd_fill_2
XANTENNA__057__B address[1] vgnd vpwr scs8hd_diode_2
XFILLER_24_113 vgnd vpwr scs8hd_decap_8
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_79 vpwr vgnd scs8hd_fill_2
XFILLER_21_13 vpwr vgnd scs8hd_fill_2
XANTENNA__073__A _092_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_113 vgnd vpwr scs8hd_decap_4
X_125_ _116_/A _129_/B _125_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_30_138 vgnd vpwr scs8hd_decap_12
XFILLER_7_15 vgnd vpwr scs8hd_fill_1
XFILLER_15_179 vpwr vgnd scs8hd_fill_2
X_056_ _064_/A _126_/A _056_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_38_227 vgnd vpwr scs8hd_decap_12
XFILLER_38_205 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_116 vgnd vpwr scs8hd_fill_1
XANTENNA__158__A _064_/B vgnd vpwr scs8hd_diode_2
XFILLER_14_190 vgnd vpwr scs8hd_decap_3
XFILLER_29_238 vgnd vpwr scs8hd_decap_6
XANTENNA__068__A _124_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_46 vpwr vgnd scs8hd_fill_2
XFILLER_32_89 vgnd vpwr scs8hd_fill_1
XFILLER_32_23 vgnd vpwr scs8hd_decap_4
XFILLER_32_12 vpwr vgnd scs8hd_fill_2
Xmem_top_track_0.LATCH_2_.latch data_in mem_top_track_0.LATCH_2_.latch/Q _062_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_7_175 vpwr vgnd scs8hd_fill_2
X_108_ _118_/A _104_/X _108_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_21_3 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_16.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_4_.latch_SLEEPB _090_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.tap_buf4_0_.scs8hd_inv_1 mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _203_/A vgnd vpwr scs8hd_inv_1
XFILLER_8_91 vgnd vpwr scs8hd_fill_1
XANTENNA__070__B _067_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_263 vgnd vpwr scs8hd_decap_12
XFILLER_25_252 vpwr vgnd scs8hd_fill_2
Xmem_left_track_17.LATCH_5_.latch data_in mem_left_track_17.LATCH_5_.latch/Q _154_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_167 vgnd vpwr scs8hd_decap_4
XFILLER_4_27 vgnd vpwr scs8hd_decap_4
XANTENNA__139__C _139_/C vgnd vpwr scs8hd_diode_2
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__155__B _153_/X vgnd vpwr scs8hd_diode_2
XFILLER_16_274 vgnd vpwr scs8hd_fill_1
XANTENNA__049__C _063_/C vgnd vpwr scs8hd_diode_2
XFILLER_22_211 vgnd vpwr scs8hd_fill_1
XANTENNA__065__B address[1] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_3_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_right_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__081__A _059_/X vgnd vpwr scs8hd_diode_2
XFILLER_1_104 vpwr vgnd scs8hd_fill_2
XFILLER_1_126 vpwr vgnd scs8hd_fill_2
XFILLER_1_137 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_7_.latch_SLEEPB _115_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_181 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__051__D _051_/D vgnd vpwr scs8hd_diode_2
XFILLER_5_70 vpwr vgnd scs8hd_fill_2
XFILLER_24_57 vpwr vgnd scs8hd_fill_2
XANTENNA__076__A _046_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_56 vgnd vpwr scs8hd_decap_3
XFILLER_10_236 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_1_39 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_1.LATCH_4_.latch data_in mem_bottom_track_1.LATCH_4_.latch/Q _099_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_37 vgnd vpwr scs8hd_decap_3
XFILLER_42_136 vgnd vpwr scs8hd_decap_8
XFILLER_42_125 vpwr vgnd scs8hd_fill_2
XFILLER_35_34 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.INVTX1_3_.scs8hd_inv_1_A right_bottom_grid_pin_12_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_27_155 vgnd vpwr scs8hd_decap_4
XFILLER_19_57 vpwr vgnd scs8hd_fill_2
XFILLER_42_147 vgnd vpwr scs8hd_decap_8
X_141_ _118_/A _143_/B _141_/Y vgnd vpwr scs8hd_nor2_4
X_072_ _059_/X _067_/X _072_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_16.INVTX1_7_.scs8hd_inv_1 chanx_left_in[6] mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
Xmux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_8.LATCH_4_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_18_100 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB _084_/Y vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_3_.latch data_in mem_left_track_1.LATCH_3_.latch/Q _119_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_93 vpwr vgnd scs8hd_fill_2
XANTENNA__057__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_32_191 vpwr vgnd scs8hd_fill_2
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_58 vgnd vpwr scs8hd_fill_1
XANTENNA__073__B _067_/X vgnd vpwr scs8hd_diode_2
X_124_ _124_/A _129_/B _124_/Y vgnd vpwr scs8hd_nor2_4
X_055_ _053_/A address[1] _063_/C _126_/A vgnd vpwr scs8hd_or3_4
XFILLER_23_180 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_17.INVTX1_7_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_7_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_239 vgnd vpwr scs8hd_decap_12
XANTENNA__158__B _153_/X vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ mem_bottom_track_17.LATCH_5_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_right_track_16.LATCH_4_.latch data_in mem_right_track_16.LATCH_4_.latch/Q _141_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__174__A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__068__B _067_/X vgnd vpwr scs8hd_diode_2
XFILLER_32_68 vpwr vgnd scs8hd_fill_2
XFILLER_32_46 vpwr vgnd scs8hd_fill_2
XANTENNA__084__A _094_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_139 vgnd vpwr scs8hd_decap_8
XFILLER_20_150 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_28_272 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_17.LATCH_5_.latch_SLEEPB _154_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_2_.latch_SLEEPB _073_/Y vgnd vpwr scs8hd_diode_2
X_107_ _126_/A _104_/X _107_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_161 vpwr vgnd scs8hd_fill_2
XFILLER_11_172 vpwr vgnd scs8hd_fill_2
XFILLER_27_57 vpwr vgnd scs8hd_fill_2
XANTENNA__079__A _126_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_79 vpwr vgnd scs8hd_fill_2
XFILLER_25_275 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_4_102 vgnd vpwr scs8hd_decap_12
XANTENNA__139__D _139_/D vgnd vpwr scs8hd_diode_2
XFILLER_17_90 vpwr vgnd scs8hd_fill_2
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_234 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__065__C address[0] vgnd vpwr scs8hd_diode_2
XANTENNA__081__B _081_/B vgnd vpwr scs8hd_diode_2
XFILLER_13_26 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_212 vgnd vpwr scs8hd_decap_3
XFILLER_13_234 vpwr vgnd scs8hd_fill_2
XFILLER_0_160 vgnd vpwr scs8hd_fill_1
XFILLER_8_260 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr
+ scs8hd_diode_2
XANTENNA__182__A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_39_153 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_36 vpwr vgnd scs8hd_fill_2
XFILLER_10_248 vgnd vpwr scs8hd_decap_12
XANTENNA__076__B _139_/B vgnd vpwr scs8hd_diode_2
XANTENNA__092__A _092_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_263 vgnd vpwr scs8hd_decap_12
XFILLER_36_167 vgnd vpwr scs8hd_decap_12
XANTENNA__177__A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_10_27 vpwr vgnd scs8hd_fill_2
XFILLER_35_57 vpwr vgnd scs8hd_fill_2
XFILLER_27_189 vpwr vgnd scs8hd_fill_2
XANTENNA__087__A _124_/A vgnd vpwr scs8hd_diode_2
X_140_ _126_/A _143_/B _140_/Y vgnd vpwr scs8hd_nor2_4
X_071_ _118_/A _067_/X _071_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_16.LATCH_4_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_bottom_track_9.INVTX1_2_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_134 vpwr vgnd scs8hd_fill_2
XFILLER_18_145 vgnd vpwr scs8hd_decap_8
XFILLER_41_181 vpwr vgnd scs8hd_fill_2
XFILLER_33_115 vgnd vpwr scs8hd_decap_4
XFILLER_25_90 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_107 vgnd vpwr scs8hd_decap_3
XFILLER_23_170 vgnd vpwr scs8hd_decap_4
Xmux_top_track_16.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[2] mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_left_track_17.LATCH_4_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_054_ _064_/A _116_/A _054_/Y vgnd vpwr scs8hd_nor2_4
X_123_ _046_/Y address[3] _139_/C _114_/D _129_/B vgnd vpwr scs8hd_or4_4
XANTENNA__190__A _190_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_6_.latch_SLEEPB _106_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_0.LATCH_3_.latch data_in mem_right_track_0.LATCH_3_.latch/Q _081_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_top_track_8.LATCH_3_.latch data_in mem_top_track_8.LATCH_3_.latch/Q _072_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__084__B _081_/B vgnd vpwr scs8hd_diode_2
XFILLER_20_140 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_111 vpwr vgnd scs8hd_fill_2
XFILLER_7_144 vpwr vgnd scs8hd_fill_2
XFILLER_7_199 vpwr vgnd scs8hd_fill_2
XFILLER_11_184 vgnd vpwr scs8hd_decap_4
X_106_ _116_/A _104_/X _106_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_3_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XANTENNA__185__A _185_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_82 vgnd vpwr scs8hd_fill_1
XFILLER_27_36 vpwr vgnd scs8hd_fill_2
XANTENNA__079__B _081_/B vgnd vpwr scs8hd_diode_2
XFILLER_40_235 vgnd vpwr scs8hd_decap_3
XFILLER_40_213 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_9.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__095__A _139_/C vgnd vpwr scs8hd_diode_2
XFILLER_4_114 vgnd vpwr scs8hd_decap_4
XFILLER_31_213 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_246 vgnd vpwr scs8hd_decap_12
XFILLER_22_235 vgnd vpwr scs8hd_decap_8
XFILLER_22_224 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_49 vpwr vgnd scs8hd_fill_2
XFILLER_38_68 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_272 vgnd vpwr scs8hd_decap_3
XFILLER_39_132 vpwr vgnd scs8hd_fill_2
XANTENNA__092__B _094_/B vgnd vpwr scs8hd_diode_2
XANTENNA__076__C _139_/C vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_2_.latch/Q mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_17.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_242 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_9.LATCH_5_.latch data_in mem_bottom_track_9.LATCH_5_.latch/Q _107_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_39_6 vpwr vgnd scs8hd_fill_2
XFILLER_5_275 vpwr vgnd scs8hd_fill_2
XFILLER_36_179 vgnd vpwr scs8hd_fill_1
XFILLER_36_102 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_2_.latch_SLEEPB _101_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__193__A chany_top_in[4] vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_2_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_2_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__087__B _094_/B vgnd vpwr scs8hd_diode_2
XFILLER_27_179 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_2_.latch/Q mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_070_ _126_/A _067_/X _070_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_4_3 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.INVTX1_2_.scs8hd_inv_1 chany_top_in[4] mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_bottom_track_1.INVTX1_5_.scs8hd_inv_1 bottom_right_grid_pin_11_ mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_track_8.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_113 vgnd vpwr scs8hd_decap_8
XPHY_80 vgnd vpwr scs8hd_decap_3
XFILLER_33_138 vpwr vgnd scs8hd_fill_2
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_199_ _199_/A chany_top_out[8] vgnd vpwr scs8hd_buf_2
Xmem_left_track_9.LATCH_4_.latch data_in mem_left_track_9.LATCH_4_.latch/Q _127_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_16.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__188__A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_24_138 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ mem_bottom_track_9.LATCH_5_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_171 vgnd vpwr scs8hd_decap_4
XFILLER_21_38 vgnd vpwr scs8hd_decap_3
Xmux_top_track_8.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[1] mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__098__A _126_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_105 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_127 vpwr vgnd scs8hd_fill_2
X_053_ _053_/A _059_/B address[0] _116_/A vgnd vpwr scs8hd_or3_4
Xmux_top_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_3_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_122_ _094_/A _121_/B _122_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB _134_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_119 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A _162_/HI vgnd vpwr
+ scs8hd_diode_2
Xmem_top_track_16.LATCH_5_.latch data_in mem_top_track_16.LATCH_5_.latch/Q _133_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_37_263 vgnd vpwr scs8hd_decap_12
XFILLER_29_208 vpwr vgnd scs8hd_fill_2
XFILLER_16_16 vpwr vgnd scs8hd_fill_2
XFILLER_12_108 vgnd vpwr scs8hd_decap_4
XFILLER_12_119 vgnd vpwr scs8hd_decap_6
XFILLER_16_27 vpwr vgnd scs8hd_fill_2
XFILLER_20_163 vgnd vpwr scs8hd_decap_8
XFILLER_28_252 vgnd vpwr scs8hd_decap_12
XFILLER_28_241 vgnd vpwr scs8hd_decap_8
XFILLER_28_230 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_123 vgnd vpwr scs8hd_decap_4
XFILLER_11_130 vgnd vpwr scs8hd_decap_3
X_105_ _124_/A _104_/X _105_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_167 vgnd vpwr scs8hd_decap_3
XFILLER_19_230 vpwr vgnd scs8hd_fill_2
XFILLER_8_61 vgnd vpwr scs8hd_fill_1
XANTENNA__095__B _139_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_126 vpwr vgnd scs8hd_fill_2
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_211 vgnd vpwr scs8hd_fill_1
XFILLER_17_81 vpwr vgnd scs8hd_fill_2
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_top_track_0.LATCH_6_.latch_SLEEPB _054_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__196__A chany_top_in[1] vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_7_.scs8hd_inv_1 chany_bottom_in[4] mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_22_258 vgnd vpwr scs8hd_decap_12
XFILLER_22_203 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_left_track_17.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_229 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_80 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_17.LATCH_3_.latch_SLEEPB _149_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_195 vgnd vpwr scs8hd_fill_1
Xmux_right_track_0.INVTX1_3_.scs8hd_inv_1 right_top_grid_pin_10_ mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_39_166 vpwr vgnd scs8hd_fill_2
XFILLER_39_188 vpwr vgnd scs8hd_fill_2
XFILLER_24_27 vpwr vgnd scs8hd_fill_2
XANTENNA__076__D _051_/D vgnd vpwr scs8hd_diode_2
XFILLER_40_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_71 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_8_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_6_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_210 vgnd vpwr scs8hd_decap_12
XFILLER_14_93 vgnd vpwr scs8hd_fill_1
XFILLER_39_90 vgnd vpwr scs8hd_decap_4
XFILLER_36_125 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_2_.latch/Q mux_bottom_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_17.LATCH_5_.latch data_in mem_bottom_track_17.LATCH_5_.latch/Q _147_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_35_15 vpwr vgnd scs8hd_fill_2
XFILLER_27_114 vpwr vgnd scs8hd_fill_2
XFILLER_19_16 vgnd vpwr scs8hd_decap_3
XFILLER_19_38 vpwr vgnd scs8hd_fill_2
XFILLER_41_161 vgnd vpwr scs8hd_decap_12
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_198_ _198_/A chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_2_85 vgnd vpwr scs8hd_decap_6
XFILLER_32_150 vgnd vpwr scs8hd_fill_1
XFILLER_24_106 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.INVTX1_7_.scs8hd_inv_1 chanx_left_in[3] mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_17 vpwr vgnd scs8hd_fill_2
XANTENNA__098__B _095_/X vgnd vpwr scs8hd_diode_2
XFILLER_15_117 vgnd vpwr scs8hd_fill_1
X_121_ _064_/B _121_/B _121_/Y vgnd vpwr scs8hd_nor2_4
X_052_ _124_/A _064_/A _052_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_72 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_14_172 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__199__A _199_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_275 vpwr vgnd scs8hd_fill_2
XFILLER_37_253 vpwr vgnd scs8hd_fill_2
Xmem_right_track_8.LATCH_4_.latch data_in mem_right_track_8.LATCH_4_.latch/Q _090_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_8.INVTX1_8_.scs8hd_inv_1 chanx_left_in[5] mux_right_track_8.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_0.INVTX1_8_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_20_186 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB _093_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_264 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_9.INVTX1_8_.scs8hd_inv_1_A left_bottom_grid_pin_12_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_179 vpwr vgnd scs8hd_fill_2
Xmem_left_track_17.LATCH_0_.latch data_in mem_left_track_17.LATCH_0_.latch/Q _159_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_104_ _046_/Y _139_/B _139_/C _139_/D _104_/X vgnd vpwr scs8hd_or4_4
XANTENNA_mem_left_track_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_6 vpwr vgnd scs8hd_fill_2
XFILLER_40_215 vgnd vpwr scs8hd_decap_12
XFILLER_25_234 vpwr vgnd scs8hd_fill_2
XFILLER_25_212 vpwr vgnd scs8hd_fill_2
XANTENNA__095__C _046_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_259 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_248 vgnd vpwr scs8hd_decap_12
XFILLER_31_226 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_4_.latch_SLEEPB _118_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_171 vpwr vgnd scs8hd_fill_2
XFILLER_3_160 vpwr vgnd scs8hd_fill_2
XFILLER_1_108 vpwr vgnd scs8hd_fill_2
XFILLER_38_15 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_3_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_248 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_152 vgnd vpwr scs8hd_decap_3
XFILLER_0_185 vgnd vpwr scs8hd_fill_1
XFILLER_12_270 vgnd vpwr scs8hd_decap_4
XFILLER_5_85 vgnd vpwr scs8hd_decap_3
XFILLER_5_52 vgnd vpwr scs8hd_decap_4
XFILLER_39_178 vgnd vpwr scs8hd_fill_1
XFILLER_39_101 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_4_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_27 vgnd vpwr scs8hd_decap_4
XFILLER_14_50 vpwr vgnd scs8hd_fill_2
XFILLER_5_222 vgnd vpwr scs8hd_decap_12
XFILLER_39_80 vgnd vpwr scs8hd_fill_1
Xmux_right_track_16.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[6] mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[1] mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_159 vgnd vpwr scs8hd_fill_1
XFILLER_27_137 vpwr vgnd scs8hd_fill_2
XFILLER_42_129 vgnd vpwr scs8hd_decap_4
XFILLER_35_192 vpwr vgnd scs8hd_fill_2
XFILLER_35_170 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_41_184 vgnd vpwr scs8hd_decap_12
XFILLER_41_173 vgnd vpwr scs8hd_decap_8
X_197_ chany_top_in[0] chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.tap_buf4_0_.scs8hd_inv_1 mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _199_/A vgnd vpwr scs8hd_inv_1
XFILLER_2_97 vpwr vgnd scs8hd_fill_2
XFILLER_2_64 vpwr vgnd scs8hd_fill_2
XFILLER_32_184 vgnd vpwr scs8hd_decap_4
Xmux_left_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 _163_/HI mem_left_track_1.LATCH_7_.latch/Q
+ mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_23_140 vpwr vgnd scs8hd_fill_2
X_120_ _092_/A _121_/B _120_/Y vgnd vpwr scs8hd_nor2_4
X_051_ address[4] address[3] _139_/C _051_/D _064_/A vgnd vpwr scs8hd_or4_4
XFILLER_23_184 vpwr vgnd scs8hd_fill_2
XFILLER_11_62 vgnd vpwr scs8hd_fill_1
XFILLER_11_95 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_70 vgnd vpwr scs8hd_decap_3
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.LATCH_2_.latch_SLEEPB _157_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_243 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
XFILLER_11_110 vpwr vgnd scs8hd_fill_2
XFILLER_22_61 vgnd vpwr scs8hd_fill_1
XFILLER_11_165 vpwr vgnd scs8hd_fill_2
XFILLER_11_176 vgnd vpwr scs8hd_decap_4
X_103_ _094_/A _095_/X _103_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_34_235 vgnd vpwr scs8hd_decap_12
XFILLER_34_224 vgnd vpwr scs8hd_decap_8
XFILLER_34_213 vgnd vpwr scs8hd_fill_1
XFILLER_19_254 vgnd vpwr scs8hd_fill_1
XFILLER_8_41 vpwr vgnd scs8hd_fill_2
XFILLER_8_85 vgnd vpwr scs8hd_decap_6
XFILLER_6_180 vgnd vpwr scs8hd_decap_4
XFILLER_27_17 vpwr vgnd scs8hd_fill_2
XFILLER_40_227 vgnd vpwr scs8hd_decap_8
XANTENNA__095__D address[3] vgnd vpwr scs8hd_diode_2
XFILLER_4_139 vpwr vgnd scs8hd_fill_2
XFILLER_16_224 vgnd vpwr scs8hd_decap_8
XFILLER_16_235 vgnd vpwr scs8hd_decap_8
XFILLER_16_246 vgnd vpwr scs8hd_decap_12
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_238 vgnd vpwr scs8hd_decap_6
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_13_238 vgnd vpwr scs8hd_decap_6
Xmux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_60 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.tap_buf4_0_.scs8hd_inv_1 mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _185_/A vgnd vpwr scs8hd_inv_1
XFILLER_14_84 vpwr vgnd scs8hd_fill_2
XFILLER_30_72 vpwr vgnd scs8hd_fill_2
XFILLER_5_245 vpwr vgnd scs8hd_fill_2
XFILLER_5_234 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_2_.latch/Q mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_138 vpwr vgnd scs8hd_fill_2
XANTENNA__101__A _092_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_35_182 vgnd vpwr scs8hd_fill_1
XFILLER_35_28 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_215 vgnd vpwr scs8hd_decap_12
XFILLER_18_138 vgnd vpwr scs8hd_decap_4
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XFILLER_33_119 vgnd vpwr scs8hd_fill_1
XPHY_61 vgnd vpwr scs8hd_decap_3
XFILLER_26_182 vpwr vgnd scs8hd_fill_2
XFILLER_26_171 vgnd vpwr scs8hd_decap_4
XFILLER_25_50 vpwr vgnd scs8hd_fill_2
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_196 vgnd vpwr scs8hd_decap_12
X_196_ chany_top_in[1] chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_2_32 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.INVTX1_0_.scs8hd_inv_1 chanx_right_in[0] mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_17_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_050_ address[5] address[6] _051_/D vgnd vpwr scs8hd_or2_4
XANTENNA_mem_bottom_track_9.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_3_.latch_SLEEPB _109_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_3 vgnd vpwr scs8hd_decap_12
XFILLER_11_52 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_141 vgnd vpwr scs8hd_decap_8
XFILLER_14_163 vgnd vpwr scs8hd_decap_3
XFILLER_14_185 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_179_ chanx_right_in[0] chanx_left_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_35_3 vpwr vgnd scs8hd_fill_2
XFILLER_32_29 vpwr vgnd scs8hd_fill_2
XFILLER_20_122 vgnd vpwr scs8hd_decap_4
XFILLER_20_144 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_211 vgnd vpwr scs8hd_fill_1
XFILLER_11_144 vpwr vgnd scs8hd_fill_2
XFILLER_22_84 vpwr vgnd scs8hd_fill_2
XFILLER_22_73 vpwr vgnd scs8hd_fill_2
X_102_ _064_/B _095_/X _102_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_115 vpwr vgnd scs8hd_fill_2
XFILLER_7_159 vpwr vgnd scs8hd_fill_2
XFILLER_34_247 vgnd vpwr scs8hd_decap_8
XFILLER_8_53 vgnd vpwr scs8hd_decap_8
XFILLER_8_64 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.INVTX1_8_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_118 vgnd vpwr scs8hd_fill_1
XFILLER_16_203 vgnd vpwr scs8hd_decap_8
XFILLER_16_258 vgnd vpwr scs8hd_decap_12
XFILLER_17_40 vpwr vgnd scs8hd_fill_2
XFILLER_17_73 vpwr vgnd scs8hd_fill_2
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_94 vpwr vgnd scs8hd_fill_2
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_184 vgnd vpwr scs8hd_decap_12
XANTENNA__104__A _046_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_5_.latch_SLEEPB _079_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_272 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_217 vgnd vpwr scs8hd_decap_3
XFILLER_0_132 vgnd vpwr scs8hd_decap_12
XFILLER_0_165 vpwr vgnd scs8hd_fill_2
XFILLER_0_187 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_8.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_top_track_0.LATCH_3_.latch data_in mem_top_track_0.LATCH_3_.latch/Q _060_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
XFILLER_39_114 vpwr vgnd scs8hd_fill_2
XFILLER_5_65 vgnd vpwr scs8hd_decap_3
Xmem_bottom_track_9.LATCH_0_.latch data_in mem_bottom_track_9.LATCH_0_.latch/Q _112_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_39_136 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_8.LATCH_7_.latch_SLEEPB _068_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_84 vpwr vgnd scs8hd_fill_2
XFILLER_36_106 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__101__B _095_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_2_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__202__A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_227 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.INVTX1_1_.scs8hd_inv_1 chanx_right_in[2] mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_95 vgnd vpwr scs8hd_decap_3
XFILLER_25_73 vpwr vgnd scs8hd_fill_2
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
X_195_ chany_top_in[2] chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_37_7 vpwr vgnd scs8hd_fill_2
XFILLER_2_77 vpwr vgnd scs8hd_fill_2
XFILLER_2_44 vgnd vpwr scs8hd_decap_12
XANTENNA__112__A _094_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_131 vpwr vgnd scs8hd_fill_2
XFILLER_17_161 vpwr vgnd scs8hd_fill_2
XFILLER_32_142 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB _137_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_197 vpwr vgnd scs8hd_fill_2
XFILLER_23_153 vpwr vgnd scs8hd_fill_2
XFILLER_15_109 vpwr vgnd scs8hd_fill_2
Xmem_top_track_16.LATCH_0_.latch data_in mem_top_track_16.LATCH_0_.latch/Q _138_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_31 vpwr vgnd scs8hd_fill_2
XFILLER_14_120 vgnd vpwr scs8hd_decap_8
XANTENNA__107__A _126_/A vgnd vpwr scs8hd_diode_2
X_178_ chanx_right_in[1] chanx_left_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_245 vgnd vpwr scs8hd_decap_8
XFILLER_37_223 vpwr vgnd scs8hd_fill_2
XFILLER_37_212 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_16.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr
+ scs8hd_diode_2
Xmem_bottom_track_1.LATCH_5_.latch data_in mem_bottom_track_1.LATCH_5_.latch/Q _098_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_41 vgnd vpwr scs8hd_decap_3
X_101_ _092_/A _095_/X _101_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_123 vgnd vpwr scs8hd_decap_4
XFILLER_19_234 vpwr vgnd scs8hd_fill_2
XFILLER_34_259 vgnd vpwr scs8hd_decap_12
XFILLER_8_10 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_248 vpwr vgnd scs8hd_fill_2
XFILLER_40_207 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB _060_/Y vgnd vpwr scs8hd_diode_2
XFILLER_25_259 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.INVTX1_4_.scs8hd_inv_1 chanx_right_in[5] mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_left_track_1.LATCH_4_.latch data_in mem_left_track_1.LATCH_4_.latch/Q _118_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_7_.scs8hd_inv_1 chanx_left_in[6] mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_73 vgnd vpwr scs8hd_decap_4
XFILLER_33_40 vpwr vgnd scs8hd_fill_2
XFILLER_3_196 vgnd vpwr scs8hd_decap_12
XANTENNA__104__B _139_/B vgnd vpwr scs8hd_diode_2
XANTENNA__120__A _092_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_6 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_track_9.LATCH_4_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB _152_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_right_track_16.LATCH_5_.latch data_in mem_right_track_16.LATCH_5_.latch/Q _140_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_229 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.INVTX1_2_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA__205__A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_0_144 vgnd vpwr scs8hd_decap_8
XANTENNA__115__A _124_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_3 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_17.LATCH_0_.latch data_in mem_bottom_track_17.LATCH_0_.latch/Q _152_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_left_track_9.LATCH_5_.latch_SLEEPB _126_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_41 vgnd vpwr scs8hd_decap_3
Xmux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_8.LATCH_5_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_39_72 vgnd vpwr scs8hd_decap_8
Xmux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_118 vpwr vgnd scs8hd_fill_2
XFILLER_35_184 vgnd vpwr scs8hd_fill_1
XFILLER_35_151 vpwr vgnd scs8hd_fill_2
XFILLER_2_239 vgnd vpwr scs8hd_decap_12
XFILLER_2_206 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[0] mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_25_30 vpwr vgnd scs8hd_fill_2
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_110 vgnd vpwr scs8hd_fill_1
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_41 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
X_194_ _194_/A chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_56 vgnd vpwr scs8hd_decap_8
XANTENNA__112__B _104_/X vgnd vpwr scs8hd_diode_2
XFILLER_32_154 vpwr vgnd scs8hd_fill_2
XFILLER_17_140 vpwr vgnd scs8hd_fill_2
XFILLER_23_176 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_11_76 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[3] mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_36_84 vpwr vgnd scs8hd_fill_2
XFILLER_36_51 vgnd vpwr scs8hd_fill_1
X_177_ chanx_right_in[2] chanx_left_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA__107__B _104_/X vgnd vpwr scs8hd_diode_2
XANTENNA__123__A _046_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_191 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1_A bottom_left_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_53 vpwr vgnd scs8hd_fill_2
X_100_ _059_/X _095_/X _100_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_19_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_7_.latch_SLEEPB _096_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_213 vpwr vgnd scs8hd_fill_2
XANTENNA__118__A _118_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_6_150 vgnd vpwr scs8hd_decap_3
XFILLER_40_3 vgnd vpwr scs8hd_decap_12
XFILLER_25_238 vgnd vpwr scs8hd_decap_6
XFILLER_25_216 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB _121_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.INVTX1_7_.scs8hd_inv_1 chany_bottom_in[8] mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_2_.latch/Q mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_271 vgnd vpwr scs8hd_decap_4
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_53 vpwr vgnd scs8hd_fill_2
XFILLER_17_86 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_175 vpwr vgnd scs8hd_fill_2
XFILLER_3_164 vgnd vpwr scs8hd_decap_4
XFILLER_3_153 vpwr vgnd scs8hd_fill_2
XFILLER_3_142 vpwr vgnd scs8hd_fill_2
XANTENNA__104__C _139_/C vgnd vpwr scs8hd_diode_2
XANTENNA__120__B _121_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_252 vgnd vpwr scs8hd_decap_12
XFILLER_30_241 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr
+ scs8hd_diode_2
XFILLER_38_19 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_263 vgnd vpwr scs8hd_decap_12
XFILLER_21_252 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB _144_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_156 vgnd vpwr scs8hd_decap_4
Xmux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_2_.latch/Q mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_85 vgnd vpwr scs8hd_decap_4
Xmem_right_track_0.LATCH_4_.latch data_in mem_right_track_0.LATCH_4_.latch/Q _080_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_top_track_8.LATCH_4_.latch data_in mem_top_track_8.LATCH_4_.latch/Q _071_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_274 vgnd vpwr scs8hd_fill_1
XANTENNA__115__B _121_/B vgnd vpwr scs8hd_diode_2
XFILLER_39_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__131__A _094_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_171 vgnd vpwr scs8hd_decap_3
Xmux_right_track_16.INVTX1_1_.scs8hd_inv_1 chany_top_in[5] mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.INVTX1_2_.scs8hd_inv_1 chany_top_in[7] mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_10 vpwr vgnd scs8hd_fill_2
XFILLER_14_32 vpwr vgnd scs8hd_fill_2
XFILLER_14_54 vpwr vgnd scs8hd_fill_2
XFILLER_30_53 vgnd vpwr scs8hd_decap_4
XFILLER_5_259 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ mem_top_track_16.LATCH_5_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_39_62 vpwr vgnd scs8hd_fill_2
XFILLER_29_193 vpwr vgnd scs8hd_fill_2
XFILLER_29_182 vgnd vpwr scs8hd_fill_1
XANTENNA__126__A _126_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_130 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_100 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
Xmux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_left_track_17.LATCH_5_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XFILLER_41_74 vgnd vpwr scs8hd_decap_8
X_193_ chany_top_in[4] chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
XPHY_75 vgnd vpwr scs8hd_decap_3
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_96 vpwr vgnd scs8hd_fill_2
XFILLER_41_85 vpwr vgnd scs8hd_fill_2
XFILLER_32_188 vgnd vpwr scs8hd_fill_1
XFILLER_17_174 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_166 vpwr vgnd scs8hd_fill_2
XFILLER_23_144 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_track_1.LATCH_4_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_63 vgnd vpwr scs8hd_decap_4
Xmux_right_track_0.INVTX1_8_.scs8hd_inv_1 chanx_left_in[4] mux_right_track_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_176_ _176_/A chanx_left_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__123__B address[3] vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_9.LATCH_6_.latch data_in mem_bottom_track_9.LATCH_6_.latch/Q _106_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_203 vpwr vgnd scs8hd_fill_2
XFILLER_11_114 vgnd vpwr scs8hd_decap_8
XFILLER_22_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_3 vgnd vpwr scs8hd_decap_12
XFILLER_34_206 vgnd vpwr scs8hd_fill_1
XFILLER_19_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_261 vgnd vpwr scs8hd_decap_12
XANTENNA__118__B _121_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_23 vgnd vpwr scs8hd_decap_8
XFILLER_8_45 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_78 vgnd vpwr scs8hd_decap_4
X_159_ _094_/A _153_/X _159_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__134__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_3 vgnd vpwr scs8hd_decap_4
Xmem_left_track_9.LATCH_5_.latch data_in mem_left_track_9.LATCH_5_.latch/Q _126_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__044__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _164_/HI vgnd vpwr
+ scs8hd_diode_2
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_53 vpwr vgnd scs8hd_fill_2
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_209 vpwr vgnd scs8hd_fill_2
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_121 vgnd vpwr scs8hd_fill_1
XANTENNA__104__D _139_/D vgnd vpwr scs8hd_diode_2
XANTENNA__129__A _092_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_264 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_275 vpwr vgnd scs8hd_fill_2
XFILLER_0_102 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_64 vgnd vpwr scs8hd_fill_1
XFILLER_8_202 vpwr vgnd scs8hd_fill_2
XFILLER_8_224 vgnd vpwr scs8hd_decap_12
XANTENNA__131__B _129_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_35 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_3_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_194 vgnd vpwr scs8hd_decap_8
XFILLER_38_183 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_8.LATCH_6_.latch_SLEEPB _088_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_88 vpwr vgnd scs8hd_fill_2
XFILLER_30_76 vgnd vpwr scs8hd_decap_3
XFILLER_30_10 vpwr vgnd scs8hd_fill_2
XFILLER_5_249 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__126__B _129_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_5_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__142__A _059_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_120 vpwr vgnd scs8hd_fill_2
XFILLER_27_109 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_8_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_6_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_16.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__052__A _124_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_5_.scs8hd_inv_1 chanx_left_in[0] mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_41_145 vpwr vgnd scs8hd_fill_2
XFILLER_41_134 vpwr vgnd scs8hd_fill_2
XFILLER_41_123 vpwr vgnd scs8hd_fill_2
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XFILLER_26_186 vgnd vpwr scs8hd_fill_1
XPHY_54 vgnd vpwr scs8hd_decap_3
XFILLER_25_54 vgnd vpwr scs8hd_decap_4
XPHY_43 vgnd vpwr scs8hd_decap_3
XPHY_10 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
X_192_ chany_top_in[5] chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_1_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_167 vpwr vgnd scs8hd_fill_2
XFILLER_32_112 vgnd vpwr scs8hd_decap_8
XANTENNA__137__A _064_/B vgnd vpwr scs8hd_diode_2
XFILLER_17_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_123 vpwr vgnd scs8hd_fill_2
XFILLER_23_112 vpwr vgnd scs8hd_fill_2
XANTENNA__047__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_56 vgnd vpwr scs8hd_decap_3
XFILLER_11_89 vgnd vpwr scs8hd_decap_4
X_175_ chanx_right_in[4] chanx_left_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA__123__C _139_/C vgnd vpwr scs8hd_diode_2
XFILLER_35_7 vpwr vgnd scs8hd_fill_2
XFILLER_28_6 vpwr vgnd scs8hd_fill_2
XFILLER_37_259 vpwr vgnd scs8hd_fill_2
XFILLER_9_182 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_215 vpwr vgnd scs8hd_fill_2
XFILLER_22_88 vpwr vgnd scs8hd_fill_2
XFILLER_22_77 vpwr vgnd scs8hd_fill_2
XFILLER_7_119 vgnd vpwr scs8hd_decap_3
XFILLER_11_148 vpwr vgnd scs8hd_fill_2
XFILLER_19_226 vpwr vgnd scs8hd_fill_2
XFILLER_19_248 vgnd vpwr scs8hd_decap_6
XFILLER_42_273 vgnd vpwr scs8hd_decap_4
X_089_ _126_/A _094_/B _089_/Y vgnd vpwr scs8hd_nor2_4
X_158_ _064_/B _153_/X _158_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_163 vgnd vpwr scs8hd_decap_8
XFILLER_10_181 vgnd vpwr scs8hd_decap_8
XANTENNA__134__B _134_/B vgnd vpwr scs8hd_diode_2
XANTENNA__150__A _092_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_229 vgnd vpwr scs8hd_decap_3
XFILLER_18_270 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_0.LATCH_2_.latch_SLEEPB _082_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__060__A _064_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_77 vpwr vgnd scs8hd_fill_2
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_98 vpwr vgnd scs8hd_fill_2
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_251 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__129__B _129_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XANTENNA__145__A _094_/A vgnd vpwr scs8hd_diode_2
XANTENNA__055__A _053_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_243 vgnd vpwr scs8hd_fill_1
Xmem_right_track_8.LATCH_5_.latch data_in mem_right_track_8.LATCH_5_.latch/Q _089_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_28_43 vpwr vgnd scs8hd_fill_2
XFILLER_28_10 vpwr vgnd scs8hd_fill_2
XFILLER_0_169 vgnd vpwr scs8hd_decap_12
XFILLER_28_76 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 _166_/HI mem_right_track_0.LATCH_7_.latch/Q
+ mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_8_236 vgnd vpwr scs8hd_decap_12
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
XFILLER_5_58 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_8.LATCH_4_.latch_SLEEPB _071_/Y vgnd vpwr scs8hd_diode_2
XFILLER_39_118 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_3_.latch/Q mux_bottom_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_left_track_17.LATCH_1_.latch data_in mem_left_track_17.LATCH_1_.latch/Q _158_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_23 vpwr vgnd scs8hd_fill_2
XFILLER_14_67 vpwr vgnd scs8hd_fill_2
XFILLER_30_88 vpwr vgnd scs8hd_fill_2
XFILLER_39_97 vpwr vgnd scs8hd_fill_2
XFILLER_39_86 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_184 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _167_/HI mem_right_track_16.LATCH_2_.latch/Q
+ mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__142__B _143_/B vgnd vpwr scs8hd_diode_2
XANTENNA__052__B _064_/A vgnd vpwr scs8hd_diode_2
XFILLER_41_157 vpwr vgnd scs8hd_fill_2
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_198 vpwr vgnd scs8hd_fill_2
XFILLER_26_154 vpwr vgnd scs8hd_fill_2
XFILLER_25_77 vpwr vgnd scs8hd_fill_2
XPHY_44 vgnd vpwr scs8hd_decap_3
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
X_191_ chany_top_in[6] chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_track_1.INVTX1_7_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_2_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_275 vpwr vgnd scs8hd_fill_2
XFILLER_1_253 vpwr vgnd scs8hd_fill_2
XFILLER_32_102 vpwr vgnd scs8hd_fill_2
XFILLER_32_146 vgnd vpwr scs8hd_decap_4
XFILLER_32_135 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__137__B _134_/B vgnd vpwr scs8hd_diode_2
XANTENNA__153__A _046_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__063__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_11_35 vgnd vpwr scs8hd_decap_4
XFILLER_36_43 vgnd vpwr scs8hd_decap_6
Xmem_bottom_track_1.LATCH_0_.latch data_in mem_bottom_track_1.LATCH_0_.latch/Q _103_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_168 vpwr vgnd scs8hd_fill_2
XANTENNA__123__D _114_/D vgnd vpwr scs8hd_diode_2
X_174_ chanx_right_in[5] chanx_left_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_37_227 vgnd vpwr scs8hd_decap_12
XFILLER_20_105 vpwr vgnd scs8hd_fill_2
XANTENNA__148__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_150 vpwr vgnd scs8hd_fill_2
XFILLER_36_260 vgnd vpwr scs8hd_decap_12
XANTENNA__058__A _064_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_23 vpwr vgnd scs8hd_fill_2
XFILLER_11_127 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB _066_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_238 vgnd vpwr scs8hd_decap_6
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.INVTX1_4_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_9.INVTX1_1_.scs8hd_inv_1 chany_top_in[6] mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_131 vgnd vpwr scs8hd_decap_3
X_157_ _092_/A _153_/X _157_/Y vgnd vpwr scs8hd_nor2_4
X_088_ _116_/A _094_/B _088_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_186 vpwr vgnd scs8hd_fill_2
XFILLER_6_197 vgnd vpwr scs8hd_decap_6
XANTENNA__150__B _152_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__060__B _059_/X vgnd vpwr scs8hd_diode_2
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_241 vgnd vpwr scs8hd_decap_8
XFILLER_17_23 vpwr vgnd scs8hd_fill_2
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_right_track_16.LATCH_0_.latch data_in mem_right_track_16.LATCH_0_.latch/Q _145_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_123 vgnd vpwr scs8hd_decap_4
Xmux_top_track_16.INVTX1_5_.scs8hd_inv_1 chanx_left_in[1] mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_263 vgnd vpwr scs8hd_decap_12
XANTENNA__145__B _143_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__055__B address[1] vgnd vpwr scs8hd_diode_2
XFILLER_21_233 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__071__A _118_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_28_55 vgnd vpwr scs8hd_decap_3
XFILLER_5_15 vgnd vpwr scs8hd_decap_12
XFILLER_8_248 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.LATCH_2_.latch_SLEEPB _129_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_7 vpwr vgnd scs8hd_fill_2
XANTENNA__156__A _059_/X vgnd vpwr scs8hd_diode_2
XFILLER_38_163 vgnd vpwr scs8hd_decap_8
XANTENNA__066__A _064_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A _165_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_23 vpwr vgnd scs8hd_fill_2
XFILLER_39_10 vgnd vpwr scs8hd_decap_12
XFILLER_29_174 vpwr vgnd scs8hd_fill_2
XFILLER_29_163 vpwr vgnd scs8hd_fill_2
XFILLER_4_251 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_188 vpwr vgnd scs8hd_fill_2
XFILLER_35_155 vpwr vgnd scs8hd_fill_2
XFILLER_35_144 vgnd vpwr scs8hd_decap_4
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_41_114 vpwr vgnd scs8hd_fill_2
X_190_ _190_/A chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XFILLER_25_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XFILLER_2_27 vgnd vpwr scs8hd_decap_4
XFILLER_17_144 vpwr vgnd scs8hd_fill_2
XANTENNA__153__B _139_/B vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.INVTX1_2_.scs8hd_inv_1 chany_top_in[4] mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__063__B address[1] vgnd vpwr scs8hd_diode_2
XFILLER_11_14 vpwr vgnd scs8hd_fill_2
XFILLER_36_88 vgnd vpwr scs8hd_decap_4
XFILLER_36_11 vgnd vpwr scs8hd_fill_1
XFILLER_14_103 vpwr vgnd scs8hd_fill_2
XFILLER_22_180 vgnd vpwr scs8hd_decap_8
X_173_ chanx_right_in[6] chanx_left_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_37_239 vgnd vpwr scs8hd_decap_4
Xmux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_128 vgnd vpwr scs8hd_decap_3
XANTENNA__148__B _152_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_4_.latch_SLEEPB _099_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_195 vpwr vgnd scs8hd_fill_2
XFILLER_3_70 vpwr vgnd scs8hd_fill_2
XFILLER_36_272 vgnd vpwr scs8hd_decap_3
XANTENNA__058__B _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_57 vpwr vgnd scs8hd_fill_2
XFILLER_22_46 vgnd vpwr scs8hd_decap_3
XFILLER_11_106 vpwr vgnd scs8hd_fill_2
XANTENNA__074__A _064_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_42_242 vgnd vpwr scs8hd_decap_6
XFILLER_34_209 vgnd vpwr scs8hd_decap_4
X_087_ _124_/A _094_/B _087_/Y vgnd vpwr scs8hd_nor2_4
Xmux_left_track_1.INVTX1_4_.scs8hd_inv_1 chanx_right_in[4] mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_156_ _059_/X _153_/X _156_/Y vgnd vpwr scs8hd_nor2_4
Xmux_bottom_track_1.INVTX1_7_.scs8hd_inv_1 chanx_left_in[5] mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_10_150 vgnd vpwr scs8hd_fill_1
XFILLER_33_220 vpwr vgnd scs8hd_fill_2
XANTENNA__159__A _094_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_253 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__069__A _116_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_6_.scs8hd_inv_1 chanx_left_in[2] mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_23 vpwr vgnd scs8hd_fill_2
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_57 vpwr vgnd scs8hd_fill_2
XFILLER_3_102 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_179 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_231 vpwr vgnd scs8hd_fill_2
XFILLER_15_253 vpwr vgnd scs8hd_fill_2
XFILLER_15_275 vpwr vgnd scs8hd_fill_2
X_139_ address[4] _139_/B _139_/C _139_/D _143_/B vgnd vpwr scs8hd_or4_4
XFILLER_31_3 vgnd vpwr scs8hd_decap_3
XFILLER_21_212 vpwr vgnd scs8hd_fill_2
XFILLER_0_71 vgnd vpwr scs8hd_decap_8
XANTENNA__055__C _063_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__071__B _067_/X vgnd vpwr scs8hd_diode_2
XFILLER_28_89 vgnd vpwr scs8hd_fill_1
XFILLER_28_23 vpwr vgnd scs8hd_fill_2
XFILLER_12_201 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_27 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__172__A _172_/A vgnd vpwr scs8hd_diode_2
XANTENNA__156__B _153_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_8_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_38_131 vgnd vpwr scs8hd_decap_4
XANTENNA__066__B _094_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_36 vgnd vpwr scs8hd_decap_3
XFILLER_30_46 vgnd vpwr scs8hd_decap_3
XANTENNA__082__A _092_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_33 vgnd vpwr scs8hd_decap_8
XFILLER_39_22 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_263 vgnd vpwr scs8hd_decap_12
XFILLER_35_112 vpwr vgnd scs8hd_fill_2
XFILLER_35_178 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_41_104 vgnd vpwr scs8hd_decap_4
XFILLER_26_178 vpwr vgnd scs8hd_fill_2
XFILLER_26_167 vpwr vgnd scs8hd_fill_2
XFILLER_26_145 vgnd vpwr scs8hd_decap_6
XFILLER_26_134 vpwr vgnd scs8hd_fill_2
XFILLER_25_13 vpwr vgnd scs8hd_fill_2
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XANTENNA__077__A _124_/A vgnd vpwr scs8hd_diode_2
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_25_46 vpwr vgnd scs8hd_fill_2
XFILLER_41_89 vgnd vpwr scs8hd_decap_4
XFILLER_1_200 vpwr vgnd scs8hd_fill_2
XFILLER_9_3 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_8.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_17_123 vgnd vpwr scs8hd_decap_4
XANTENNA__153__C _139_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_5_.latch_SLEEPB _147_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[5] mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_31_192 vgnd vpwr scs8hd_decap_4
XFILLER_31_181 vpwr vgnd scs8hd_fill_2
Xmem_top_track_0.LATCH_4_.latch data_in mem_top_track_0.LATCH_4_.latch/Q _058_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__063__C _063_/C vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_track_8.LATCH_4_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_bottom_track_9.LATCH_1_.latch data_in mem_bottom_track_9.LATCH_1_.latch/Q _111_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_36_67 vgnd vpwr scs8hd_fill_1
XFILLER_36_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_137 vpwr vgnd scs8hd_fill_2
X_172_ _172_/A chanx_left_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_9_141 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__180__A _180_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_163 vpwr vgnd scs8hd_fill_2
XFILLER_9_174 vpwr vgnd scs8hd_fill_2
XFILLER_28_207 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__074__B _067_/X vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.LATCH_0_.latch data_in mem_left_track_9.LATCH_0_.latch/Q _131_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__090__A _118_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_240 vgnd vpwr scs8hd_decap_4
XFILLER_8_16 vgnd vpwr scs8hd_decap_4
XFILLER_8_49 vgnd vpwr scs8hd_fill_1
X_086_ address[4] address[3] _139_/C _139_/D _094_/B vgnd vpwr scs8hd_or4_4
X_155_ _118_/A _153_/X _155_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_111 vgnd vpwr scs8hd_decap_8
XFILLER_6_122 vpwr vgnd scs8hd_fill_2
XFILLER_10_162 vgnd vpwr scs8hd_decap_6
XFILLER_33_7 vgnd vpwr scs8hd_fill_1
XFILLER_26_6 vpwr vgnd scs8hd_fill_2
XFILLER_33_243 vgnd vpwr scs8hd_fill_1
XANTENNA__159__B _153_/X vgnd vpwr scs8hd_diode_2
XANTENNA__175__A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__069__B _067_/X vgnd vpwr scs8hd_diode_2
XFILLER_17_36 vpwr vgnd scs8hd_fill_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_57 vpwr vgnd scs8hd_fill_2
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
XANTENNA__085__A address[5] vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_2_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_33_79 vpwr vgnd scs8hd_fill_2
XFILLER_3_114 vgnd vpwr scs8hd_decap_4
XFILLER_15_243 vgnd vpwr scs8hd_fill_1
Xmem_top_track_16.LATCH_1_.latch data_in mem_top_track_16.LATCH_1_.latch/Q _137_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_207_ _207_/A chany_top_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_30_224 vpwr vgnd scs8hd_fill_2
X_138_ _094_/A _134_/B _138_/Y vgnd vpwr scs8hd_nor2_4
X_069_ _116_/A _067_/X _069_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_bottom_track_17.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_61 vgnd vpwr scs8hd_fill_1
XFILLER_0_94 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_16.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_106 vgnd vpwr scs8hd_decap_12
XFILLER_0_128 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_2_.latch/Q mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_8_206 vgnd vpwr scs8hd_decap_6
XFILLER_12_224 vpwr vgnd scs8hd_fill_2
XFILLER_12_235 vgnd vpwr scs8hd_decap_8
XFILLER_12_246 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_8.LATCH_3_.latch_SLEEPB _091_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_39 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_1.LATCH_6_.latch data_in mem_bottom_track_1.LATCH_6_.latch/Q _097_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_110 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__082__B _081_/B vgnd vpwr scs8hd_diode_2
XFILLER_39_45 vpwr vgnd scs8hd_fill_2
XFILLER_29_143 vpwr vgnd scs8hd_fill_2
XFILLER_29_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_5_.latch data_in mem_left_track_1.LATCH_5_.latch/Q _117_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_17.INVTX1_2_.scs8hd_inv_1 chanx_right_in[2] mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_track_16.LATCH_3_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__183__A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_6_.latch_SLEEPB _116_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_0.LATCH_4_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_93 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.tap_buf4_0_.scs8hd_inv_1 mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _207_/A vgnd vpwr scs8hd_inv_1
XFILLER_41_138 vgnd vpwr scs8hd_decap_4
Xmux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_26_102 vpwr vgnd scs8hd_fill_2
XFILLER_25_58 vgnd vpwr scs8hd_fill_1
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XANTENNA__077__B _081_/B vgnd vpwr scs8hd_diode_2
XPHY_36 vgnd vpwr scs8hd_decap_3
XFILLER_41_149 vpwr vgnd scs8hd_fill_2
XANTENNA__093__A _064_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_245 vgnd vpwr scs8hd_decap_8
XFILLER_1_212 vgnd vpwr scs8hd_decap_12
XFILLER_17_113 vgnd vpwr scs8hd_decap_3
XFILLER_40_171 vgnd vpwr scs8hd_decap_8
XFILLER_17_157 vpwr vgnd scs8hd_fill_2
XFILLER_17_179 vpwr vgnd scs8hd_fill_2
XFILLER_31_90 vgnd vpwr scs8hd_decap_3
XANTENNA__153__D _114_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_23_127 vpwr vgnd scs8hd_fill_2
XFILLER_23_116 vgnd vpwr scs8hd_decap_4
XANTENNA__178__A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_23_149 vpwr vgnd scs8hd_fill_2
XANTENNA__088__A _116_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_171_ _171_/HI _171_/LO vgnd vpwr scs8hd_conb_1
Xmem_bottom_track_17.LATCH_1_.latch data_in mem_bottom_track_17.LATCH_1_.latch/Q _151_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_120 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.INVTX1_6_.scs8hd_inv_1 chanx_left_in[2] mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_28_219 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.INVTX1_7_.scs8hd_inv_1 chany_bottom_in[7] mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__090__B _094_/B vgnd vpwr scs8hd_diode_2
XFILLER_42_211 vgnd vpwr scs8hd_decap_6
XFILLER_27_252 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_17.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_154_ _126_/A _153_/X _154_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_145 vgnd vpwr scs8hd_decap_3
X_085_ address[5] _045_/Y _139_/D vgnd vpwr scs8hd_nand2_4
Xmux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_left_track_9.LATCH_5_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_33_233 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_274 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__191__A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_3_.scs8hd_inv_1_A right_top_grid_pin_10_ vgnd vpwr
+ scs8hd_diode_2
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_36 vpwr vgnd scs8hd_fill_2
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__085__B _045_/Y vgnd vpwr scs8hd_diode_2
Xmem_right_track_8.LATCH_0_.latch data_in mem_right_track_8.LATCH_0_.latch/Q _094_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_206_ chany_bottom_in[0] chany_top_out[1] vgnd vpwr scs8hd_buf_2
Xmux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_137_ _064_/B _134_/B _137_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_170 vgnd vpwr scs8hd_decap_12
X_068_ _124_/A _067_/X _068_/Y vgnd vpwr scs8hd_nor2_4
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_2_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_3 vgnd vpwr scs8hd_decap_4
XANTENNA__186__A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB _074_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_4_.latch_SLEEPB _155_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.tap_buf4_0_.scs8hd_inv_1 mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _172_/A vgnd vpwr scs8hd_inv_1
XFILLER_9_82 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_28_47 vpwr vgnd scs8hd_fill_2
XFILLER_0_118 vgnd vpwr scs8hd_decap_6
XANTENNA__096__A _124_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_258 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_8_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_6_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_27 vpwr vgnd scs8hd_fill_2
XFILLER_30_59 vpwr vgnd scs8hd_fill_2
XFILLER_39_68 vpwr vgnd scs8hd_fill_2
XFILLER_39_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A _171_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XFILLER_20_81 vgnd vpwr scs8hd_decap_4
Xmux_left_track_9.tap_buf4_0_.scs8hd_inv_1 mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _176_/A vgnd vpwr scs8hd_inv_1
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_25_26 vpwr vgnd scs8hd_fill_2
XPHY_48 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_37 vgnd vpwr scs8hd_decap_3
XANTENNA__093__B _094_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_224 vgnd vpwr scs8hd_decap_12
XFILLER_40_183 vgnd vpwr scs8hd_decap_12
XFILLER_32_106 vgnd vpwr scs8hd_decap_4
XFILLER_15_92 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__194__A _194_/A vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.LATCH_5_.latch data_in mem_top_track_8.LATCH_5_.latch/Q _070_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_16_180 vgnd vpwr scs8hd_decap_4
Xmem_right_track_0.LATCH_5_.latch data_in mem_right_track_0.LATCH_5_.latch/Q _079_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA__088__B _094_/B vgnd vpwr scs8hd_diode_2
X_170_ _170_/HI _170_/LO vgnd vpwr scs8hd_conb_1
Xmux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_2_.latch/Q mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_132 vgnd vpwr scs8hd_decap_3
XFILLER_9_187 vpwr vgnd scs8hd_fill_2
XFILLER_13_161 vpwr vgnd scs8hd_fill_2
XFILLER_20_109 vgnd vpwr scs8hd_decap_4
XFILLER_3_40 vgnd vpwr scs8hd_decap_8
XFILLER_3_62 vgnd vpwr scs8hd_fill_1
XFILLER_3_51 vpwr vgnd scs8hd_fill_2
XANTENNA__189__A _189_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_1_.scs8hd_inv_1 chany_top_in[5] mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_27 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_3_.latch/Q mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__099__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_209 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A _168_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_131 vpwr vgnd scs8hd_fill_2
X_153_ _046_/Y _139_/B _139_/C _114_/D _153_/X vgnd vpwr scs8hd_or4_4
X_084_ _094_/A _081_/B _084_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_33_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_16.INVTX1_2_.scs8hd_inv_1 chanx_right_in[4] mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_190 vgnd vpwr scs8hd_fill_1
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _167_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_149 vpwr vgnd scs8hd_fill_2
XFILLER_3_138 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_3_.latch/Q mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_9.LATCH_5_.latch_SLEEPB _107_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_245 vgnd vpwr scs8hd_decap_8
X_205_ chany_bottom_in[1] chany_top_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_136_ _092_/A _134_/B _136_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_182 vgnd vpwr scs8hd_decap_12
X_067_ address[4] _139_/B _139_/C _051_/D _067_/X vgnd vpwr scs8hd_or4_4
XFILLER_0_41 vgnd vpwr scs8hd_decap_12
XFILLER_0_85 vpwr vgnd scs8hd_fill_2
XFILLER_21_259 vpwr vgnd scs8hd_fill_2
XFILLER_21_248 vpwr vgnd scs8hd_fill_2
XFILLER_21_237 vgnd vpwr scs8hd_decap_6
XANTENNA__096__B _095_/X vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_9.LATCH_7_.latch data_in mem_bottom_track_9.LATCH_7_.latch/Q _105_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_119_ _059_/X _121_/B _119_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_241 vgnd vpwr scs8hd_decap_3
XFILLER_38_145 vpwr vgnd scs8hd_fill_2
XANTENNA__197__A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_30_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_29_189 vpwr vgnd scs8hd_fill_2
XFILLER_29_178 vpwr vgnd scs8hd_fill_2
XFILLER_29_167 vpwr vgnd scs8hd_fill_2
XFILLER_29_112 vpwr vgnd scs8hd_fill_2
Xmem_left_track_9.LATCH_6_.latch data_in mem_left_track_9.LATCH_6_.latch/Q _125_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_60 vpwr vgnd scs8hd_fill_2
XFILLER_20_93 vgnd vpwr scs8hd_fill_1
XFILLER_35_148 vgnd vpwr scs8hd_fill_1
XFILLER_35_126 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_7_.latch_SLEEPB _077_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_84 vgnd vpwr scs8hd_decap_8
XFILLER_41_118 vpwr vgnd scs8hd_fill_2
XPHY_49 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_236 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ mem_bottom_track_1.LATCH_5_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_40_195 vgnd vpwr scs8hd_decap_12
XFILLER_40_162 vgnd vpwr scs8hd_decap_4
XFILLER_40_140 vgnd vpwr scs8hd_fill_1
XFILLER_15_71 vpwr vgnd scs8hd_fill_2
XFILLER_31_184 vgnd vpwr scs8hd_fill_1
XFILLER_31_173 vpwr vgnd scs8hd_fill_2
XFILLER_31_162 vpwr vgnd scs8hd_fill_2
XFILLER_11_18 vpwr vgnd scs8hd_fill_2
XFILLER_39_240 vgnd vpwr scs8hd_decap_4
XFILLER_14_107 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB _102_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_3 vpwr vgnd scs8hd_fill_2
XFILLER_13_140 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_195 vpwr vgnd scs8hd_fill_2
XFILLER_3_74 vpwr vgnd scs8hd_fill_2
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_85 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.INVTX1_4_.scs8hd_inv_1 chanx_right_in[7] mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__099__B _095_/X vgnd vpwr scs8hd_diode_2
XFILLER_27_276 vgnd vpwr scs8hd_fill_1
X_152_ _094_/A _152_/B _152_/Y vgnd vpwr scs8hd_nor2_4
X_083_ _064_/B _081_/B _083_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_110 vgnd vpwr scs8hd_decap_8
XFILLER_10_154 vpwr vgnd scs8hd_fill_2
XFILLER_10_198 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.INVTX1_3_.scs8hd_inv_1 chanx_right_in[8] mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_12_50 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_33_202 vgnd vpwr scs8hd_decap_3
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_257 vgnd vpwr scs8hd_decap_12
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_224 vpwr vgnd scs8hd_fill_2
XFILLER_24_202 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB _135_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_106 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_204_ chany_bottom_in[2] chany_top_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_15_235 vgnd vpwr scs8hd_decap_8
X_066_ _064_/A _094_/A _066_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_top_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_135_ _059_/X _134_/B _135_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_24_6 vpwr vgnd scs8hd_fill_2
XFILLER_2_194 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_17.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_0_53 vgnd vpwr scs8hd_decap_8
XFILLER_21_216 vpwr vgnd scs8hd_fill_2
XFILLER_9_95 vpwr vgnd scs8hd_fill_2
XFILLER_28_27 vpwr vgnd scs8hd_fill_2
XFILLER_12_205 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_271 vgnd vpwr scs8hd_decap_4
XFILLER_18_82 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
X_118_ _118_/A _121_/B _118_/Y vgnd vpwr scs8hd_nor2_4
X_049_ _053_/A _059_/B _063_/C _124_/A vgnd vpwr scs8hd_or3_4
XFILLER_38_135 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 _162_/HI mem_bottom_track_9.LATCH_7_.latch/Q
+ mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_2_.latch/Q mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB _056_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[3] mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_29_92 vpwr vgnd scs8hd_fill_2
XFILLER_35_116 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_39 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_17.LATCH_2_.latch_SLEEPB _150_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_2_.scs8hd_inv_1 chany_top_in[8] mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_259 vpwr vgnd scs8hd_fill_2
XFILLER_25_193 vpwr vgnd scs8hd_fill_2
XFILLER_25_171 vgnd vpwr scs8hd_decap_4
XFILLER_25_160 vpwr vgnd scs8hd_fill_2
XFILLER_17_105 vpwr vgnd scs8hd_fill_2
Xmem_right_track_8.LATCH_6_.latch data_in mem_right_track_8.LATCH_6_.latch/Q _088_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_39_263 vgnd vpwr scs8hd_decap_12
XFILLER_36_27 vpwr vgnd scs8hd_fill_2
XFILLER_22_163 vgnd vpwr scs8hd_decap_8
XFILLER_22_130 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_17.LATCH_2_.latch data_in mem_left_track_17.LATCH_2_.latch/Q _157_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_left_track_9.LATCH_7_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_112 vpwr vgnd scs8hd_fill_2
XFILLER_13_130 vgnd vpwr scs8hd_fill_1
XFILLER_9_167 vpwr vgnd scs8hd_fill_2
XFILLER_9_178 vpwr vgnd scs8hd_fill_2
XFILLER_36_211 vgnd vpwr scs8hd_decap_3
X_151_ _064_/B _152_/B _151_/Y vgnd vpwr scs8hd_nor2_4
X_082_ _092_/A _081_/B _082_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_126 vgnd vpwr scs8hd_decap_3
XFILLER_10_144 vgnd vpwr scs8hd_decap_6
XFILLER_12_73 vpwr vgnd scs8hd_fill_2
XFILLER_12_84 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.INVTX1_6_.scs8hd_inv_1 chanx_left_in[0] mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _170_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_92 vgnd vpwr scs8hd_decap_4
XFILLER_33_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_8.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_118 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_214 vpwr vgnd scs8hd_fill_2
XFILLER_30_228 vgnd vpwr scs8hd_decap_4
XFILLER_30_206 vgnd vpwr scs8hd_decap_6
X_203_ _203_/A chany_top_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_065_ address[2] address[1] address[0] _094_/A vgnd vpwr scs8hd_or3_4
Xmux_right_track_8.INVTX1_7_.scs8hd_inv_1 chanx_left_in[1] mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_23_83 vgnd vpwr scs8hd_decap_3
X_134_ _118_/A _134_/B _134_/Y vgnd vpwr scs8hd_nor2_4
Xmem_bottom_track_1.LATCH_1_.latch data_in mem_bottom_track_1.LATCH_1_.latch/Q _102_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_2_151 vpwr vgnd scs8hd_fill_2
XFILLER_0_32 vpwr vgnd scs8hd_fill_2
XFILLER_0_98 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB _094_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_52 vgnd vpwr scs8hd_decap_3
XFILLER_12_228 vgnd vpwr scs8hd_decap_4
XFILLER_34_71 vpwr vgnd scs8hd_fill_2
X_117_ _126_/A _121_/B _117_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_221 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_261 vgnd vpwr scs8hd_decap_12
X_048_ enable _139_/C vgnd vpwr scs8hd_inv_8
XFILLER_38_125 vgnd vpwr scs8hd_decap_4
Xmem_left_track_1.LATCH_0_.latch data_in mem_left_track_1.LATCH_0_.latch/Q _122_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_49 vgnd vpwr scs8hd_decap_6
XFILLER_29_136 vpwr vgnd scs8hd_fill_2
XFILLER_37_191 vpwr vgnd scs8hd_fill_2
XFILLER_29_147 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_1.LATCH_3_.latch_SLEEPB _119_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_8_.scs8hd_inv_1_A left_top_grid_pin_10_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_202 vgnd vpwr scs8hd_decap_12
XFILLER_29_71 vpwr vgnd scs8hd_fill_2
Xmem_right_track_16.LATCH_1_.latch data_in mem_right_track_16.LATCH_1_.latch/Q _144_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_6_20 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_97 vgnd vpwr scs8hd_decap_3
XFILLER_34_161 vpwr vgnd scs8hd_fill_2
XFILLER_26_128 vgnd vpwr scs8hd_decap_4
XFILLER_26_106 vgnd vpwr scs8hd_decap_12
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_19_191 vgnd vpwr scs8hd_decap_4
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_3_.latch_SLEEPB _142_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__102__A _064_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_150 vgnd vpwr scs8hd_decap_3
XFILLER_39_275 vpwr vgnd scs8hd_fill_2
XFILLER_22_197 vgnd vpwr scs8hd_decap_4
Xmux_left_track_17.INVTX1_4_.scs8hd_inv_1 chanx_right_in[6] mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[2] mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_83 vpwr vgnd scs8hd_fill_2
XFILLER_26_61 vgnd vpwr scs8hd_decap_4
XFILLER_9_146 vpwr vgnd scs8hd_fill_2
XFILLER_13_175 vpwr vgnd scs8hd_fill_2
XFILLER_27_256 vgnd vpwr scs8hd_decap_12
XFILLER_27_234 vgnd vpwr scs8hd_decap_4
XFILLER_27_223 vpwr vgnd scs8hd_fill_2
X_150_ _092_/A _152_/B _150_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_081_ _059_/X _081_/B _081_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_37_71 vpwr vgnd scs8hd_fill_2
XFILLER_33_237 vgnd vpwr scs8hd_decap_6
XFILLER_17_19 vpwr vgnd scs8hd_fill_2
XFILLER_24_259 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA__200__A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB _158_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_259 vpwr vgnd scs8hd_fill_2
X_202_ chany_bottom_in[4] chany_top_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_23_95 vpwr vgnd scs8hd_fill_2
XFILLER_23_62 vgnd vpwr scs8hd_fill_1
X_133_ _126_/A _134_/B _133_/Y vgnd vpwr scs8hd_nor2_4
X_064_ _064_/A _064_/B _064_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__110__A _092_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_7 vgnd vpwr scs8hd_fill_1
Xmux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_229 vpwr vgnd scs8hd_fill_2
XFILLER_9_31 vpwr vgnd scs8hd_fill_2
XFILLER_9_86 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_40 vpwr vgnd scs8hd_fill_2
XFILLER_34_50 vgnd vpwr scs8hd_fill_1
X_116_ _116_/A _121_/B _116_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_233 vgnd vpwr scs8hd_decap_8
XFILLER_11_273 vgnd vpwr scs8hd_decap_4
XANTENNA__105__A _124_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_047_ address[3] _139_/B vgnd vpwr scs8hd_inv_8
XANTENNA_mem_left_track_1.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_41 vpwr vgnd scs8hd_fill_2
XFILLER_20_85 vgnd vpwr scs8hd_fill_1
XFILLER_6_32 vpwr vgnd scs8hd_fill_2
XFILLER_6_65 vpwr vgnd scs8hd_fill_2
XFILLER_34_151 vpwr vgnd scs8hd_fill_2
XFILLER_26_118 vgnd vpwr scs8hd_fill_1
XPHY_19 vgnd vpwr scs8hd_decap_3
Xmem_right_track_0.LATCH_0_.latch data_in mem_right_track_0.LATCH_0_.latch/Q _084_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_top_track_8.LATCH_0_.latch data_in mem_top_track_8.LATCH_0_.latch/Q _075_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_118 vpwr vgnd scs8hd_fill_2
XFILLER_40_132 vgnd vpwr scs8hd_decap_8
XFILLER_31_95 vpwr vgnd scs8hd_fill_2
XFILLER_31_73 vpwr vgnd scs8hd_fill_2
XFILLER_31_62 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__102__B _095_/X vgnd vpwr scs8hd_diode_2
XFILLER_16_140 vpwr vgnd scs8hd_fill_2
XFILLER_31_143 vpwr vgnd scs8hd_fill_2
XFILLER_31_132 vgnd vpwr scs8hd_decap_8
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_110 vgnd vpwr scs8hd_decap_4
XANTENNA__203__A _203_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_51 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_94 vgnd vpwr scs8hd_decap_3
XFILLER_13_165 vgnd vpwr scs8hd_fill_1
XANTENNA__113__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_36_224 vgnd vpwr scs8hd_decap_12
XFILLER_3_66 vpwr vgnd scs8hd_fill_2
XFILLER_3_55 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_180 vgnd vpwr scs8hd_decap_8
XFILLER_27_268 vgnd vpwr scs8hd_decap_8
Xmux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_2_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_249 vgnd vpwr scs8hd_decap_12
X_080_ _118_/A _081_/B _080_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_5_3 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.tap_buf4_0_.scs8hd_inv_1 mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _189_/A vgnd vpwr scs8hd_inv_1
Xmux_bottom_track_17.INVTX1_7_.scs8hd_inv_1 chanx_left_in[4] mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_224 vpwr vgnd scs8hd_fill_2
XFILLER_33_216 vpwr vgnd scs8hd_fill_2
XFILLER_18_235 vgnd vpwr scs8hd_decap_8
XFILLER_18_246 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_2_.latch_SLEEPB _110_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__108__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_3 vgnd vpwr scs8hd_decap_12
XFILLER_5_194 vpwr vgnd scs8hd_fill_2
XFILLER_33_19 vpwr vgnd scs8hd_fill_2
X_201_ chany_bottom_in[5] chany_top_out[6] vgnd vpwr scs8hd_buf_2
X_063_ address[2] address[1] _063_/C _064_/B vgnd vpwr scs8hd_or3_4
Xmem_top_track_0.LATCH_5_.latch data_in mem_top_track_0.LATCH_5_.latch/Q _056_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_74 vpwr vgnd scs8hd_fill_2
XFILLER_23_41 vgnd vpwr scs8hd_decap_3
X_132_ _046_/Y address[3] _139_/C _051_/D _134_/B vgnd vpwr scs8hd_or4_4
Xmem_bottom_track_9.LATCH_2_.latch data_in mem_bottom_track_9.LATCH_2_.latch/Q _110_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_16.tap_buf4_0_.scs8hd_inv_1 mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _181_/A vgnd vpwr scs8hd_inv_1
XFILLER_0_67 vpwr vgnd scs8hd_fill_2
XANTENNA__110__B _104_/X vgnd vpwr scs8hd_diode_2
XFILLER_0_89 vgnd vpwr scs8hd_decap_4
XFILLER_9_65 vpwr vgnd scs8hd_fill_2
XFILLER_14_271 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_20_241 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_74 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_34_84 vpwr vgnd scs8hd_fill_2
XFILLER_11_241 vgnd vpwr scs8hd_decap_3
XFILLER_18_96 vpwr vgnd scs8hd_fill_2
X_115_ _124_/A _121_/B _115_/Y vgnd vpwr scs8hd_nor2_4
X_046_ address[4] _046_/Y vgnd vpwr scs8hd_inv_8
XFILLER_7_212 vgnd vpwr scs8hd_decap_3
XFILLER_7_245 vgnd vpwr scs8hd_decap_12
XANTENNA__105__B _104_/X vgnd vpwr scs8hd_diode_2
XANTENNA__121__A _064_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.LATCH_1_.latch data_in mem_left_track_9.LATCH_1_.latch/Q _130_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_6 vpwr vgnd scs8hd_fill_2
XFILLER_38_149 vpwr vgnd scs8hd_fill_2
XFILLER_29_116 vgnd vpwr scs8hd_decap_4
XFILLER_29_105 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_0.LATCH_4_.latch_SLEEPB _080_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_182 vgnd vpwr scs8hd_fill_1
XANTENNA__206__A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_4_215 vgnd vpwr scs8hd_decap_12
XFILLER_29_51 vpwr vgnd scs8hd_fill_2
XFILLER_29_40 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_20_64 vpwr vgnd scs8hd_fill_2
XANTENNA__116__A _116_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_2_.latch data_in mem_top_track_16.LATCH_2_.latch/Q _136_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_track_8.LATCH_5_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_141 vpwr vgnd scs8hd_fill_2
XFILLER_40_166 vgnd vpwr scs8hd_fill_1
XFILLER_15_53 vpwr vgnd scs8hd_fill_2
XFILLER_15_75 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_240 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_8.LATCH_6_.latch_SLEEPB _069_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_163 vpwr vgnd scs8hd_fill_2
XFILLER_31_188 vpwr vgnd scs8hd_fill_2
XFILLER_31_177 vpwr vgnd scs8hd_fill_2
XFILLER_31_166 vpwr vgnd scs8hd_fill_2
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_bottom_track_1.LATCH_7_.latch data_in mem_bottom_track_1.LATCH_7_.latch/Q _096_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
.ends

