magic
tech EFS8A
magscale 1 2
timestamp 1602269936
<< locali >>
rect 12759 18785 12794 18819
rect 13771 18785 13806 18819
rect 3985 18071 4019 18309
rect 14841 18071 14875 18241
rect 12943 17697 12978 17731
rect 13277 17119 13311 17221
rect 16347 16609 16382 16643
rect 17359 16609 17394 16643
rect 7021 16439 7055 16609
rect 18003 15997 18130 16031
rect 7199 15895 7233 15963
rect 18337 15895 18371 15997
rect 7199 15861 7205 15895
rect 1771 15657 1777 15691
rect 1771 15589 1805 15657
rect 10344 14841 10412 14875
rect 13838 14841 13908 14875
rect 18463 14433 18498 14467
rect 1771 13719 1805 13787
rect 1771 13685 1777 13719
rect 4019 13345 4146 13379
rect 15209 12631 15243 12937
rect 6279 11305 6285 11339
rect 6279 11237 6313 11305
rect 4537 10659 4571 10761
rect 10051 10217 10057 10251
rect 10051 10149 10085 10217
rect 5273 9979 5307 10149
rect 7199 9367 7233 9435
rect 7199 9333 7205 9367
rect 4439 9129 4445 9163
rect 4439 9061 4473 9129
rect 6469 8415 6503 8585
rect 9315 7191 9349 7259
rect 9315 7157 9321 7191
rect 12081 5083 12115 5321
rect 15019 3927 15053 3995
rect 15019 3893 15025 3927
<< viali >>
rect 13783 19465 13817 19499
rect 10931 19397 10965 19431
rect 4169 19329 4203 19363
rect 9919 19329 9953 19363
rect 1961 19261 1995 19295
rect 2145 19261 2179 19295
rect 4077 19261 4111 19295
rect 4353 19261 4387 19295
rect 4813 19261 4847 19295
rect 5676 19261 5710 19295
rect 6101 19261 6135 19295
rect 6929 19261 6963 19295
rect 7389 19261 7423 19295
rect 9832 19261 9866 19295
rect 10241 19261 10275 19295
rect 10839 19261 10873 19295
rect 12668 19261 12702 19295
rect 13093 19261 13127 19295
rect 13680 19261 13714 19295
rect 14105 19261 14139 19295
rect 3801 19193 3835 19227
rect 5089 19193 5123 19227
rect 11253 19193 11287 19227
rect 2513 19125 2547 19159
rect 3433 19125 3467 19159
rect 5779 19125 5813 19159
rect 6653 19125 6687 19159
rect 7021 19125 7055 19159
rect 8585 19125 8619 19159
rect 12771 19125 12805 19159
rect 10839 18921 10873 18955
rect 2513 18785 2547 18819
rect 4077 18785 4111 18819
rect 4353 18785 4387 18819
rect 5641 18785 5675 18819
rect 5917 18785 5951 18819
rect 7205 18785 7239 18819
rect 7481 18785 7515 18819
rect 10768 18785 10802 18819
rect 11748 18785 11782 18819
rect 12725 18785 12759 18819
rect 13737 18785 13771 18819
rect 1409 18717 1443 18751
rect 3157 18717 3191 18751
rect 4813 18717 4847 18751
rect 5733 18717 5767 18751
rect 6285 18717 6319 18751
rect 7665 18717 7699 18751
rect 9689 18717 9723 18751
rect 4169 18649 4203 18683
rect 7297 18649 7331 18683
rect 11851 18649 11885 18683
rect 13875 18649 13909 18683
rect 1869 18581 1903 18615
rect 7021 18581 7055 18615
rect 8217 18581 8251 18615
rect 12863 18581 12897 18615
rect 1593 18377 1627 18411
rect 5365 18377 5399 18411
rect 5641 18377 5675 18411
rect 6009 18377 6043 18411
rect 6653 18377 6687 18411
rect 7389 18377 7423 18411
rect 8953 18377 8987 18411
rect 18705 18377 18739 18411
rect 3709 18309 3743 18343
rect 3985 18309 4019 18343
rect 4077 18309 4111 18343
rect 4721 18309 4755 18343
rect 8033 18309 8067 18343
rect 1409 18173 1443 18207
rect 2145 18173 2179 18207
rect 2881 18173 2915 18207
rect 3433 18105 3467 18139
rect 10103 18241 10137 18275
rect 10793 18241 10827 18275
rect 14841 18241 14875 18275
rect 4905 18173 4939 18207
rect 7849 18173 7883 18207
rect 7941 18173 7975 18207
rect 8217 18173 8251 18207
rect 9873 18173 9907 18207
rect 10016 18173 10050 18207
rect 11012 18173 11046 18207
rect 12516 18173 12550 18207
rect 13277 18173 13311 18207
rect 13512 18173 13546 18207
rect 14540 18173 14574 18207
rect 8677 18105 8711 18139
rect 12909 18105 12943 18139
rect 14013 18105 14047 18139
rect 14289 18105 14323 18139
rect 15520 18173 15554 18207
rect 15945 18173 15979 18207
rect 18521 18173 18555 18207
rect 19073 18173 19107 18207
rect 15623 18105 15657 18139
rect 2421 18037 2455 18071
rect 3985 18037 4019 18071
rect 6929 18037 6963 18071
rect 11115 18037 11149 18071
rect 11713 18037 11747 18071
rect 12587 18037 12621 18071
rect 13599 18037 13633 18071
rect 14611 18037 14645 18071
rect 14841 18037 14875 18071
rect 15025 18037 15059 18071
rect 4537 17833 4571 17867
rect 1547 17765 1581 17799
rect 2329 17765 2363 17799
rect 4905 17765 4939 17799
rect 8309 17765 8343 17799
rect 1460 17697 1494 17731
rect 2421 17697 2455 17731
rect 2513 17697 2547 17731
rect 2697 17697 2731 17731
rect 4112 17697 4146 17731
rect 5365 17697 5399 17731
rect 5641 17697 5675 17731
rect 5917 17697 5951 17731
rect 7573 17697 7607 17731
rect 7849 17697 7883 17731
rect 9689 17697 9723 17731
rect 10149 17697 10183 17731
rect 11320 17697 11354 17731
rect 12909 17697 12943 17731
rect 13988 17697 14022 17731
rect 15368 17697 15402 17731
rect 16380 17697 16414 17731
rect 3157 17629 3191 17663
rect 6193 17629 6227 17663
rect 10241 17629 10275 17663
rect 1961 17561 1995 17595
rect 7665 17561 7699 17595
rect 8585 17561 8619 17595
rect 14059 17561 14093 17595
rect 4215 17493 4249 17527
rect 7205 17493 7239 17527
rect 10977 17493 11011 17527
rect 11391 17493 11425 17527
rect 13047 17493 13081 17527
rect 15439 17493 15473 17527
rect 16451 17493 16485 17527
rect 1593 17289 1627 17323
rect 14013 17289 14047 17323
rect 17233 17289 17267 17323
rect 13277 17221 13311 17255
rect 15853 17221 15887 17255
rect 2053 17153 2087 17187
rect 5089 17153 5123 17187
rect 13461 17153 13495 17187
rect 16543 17153 16577 17187
rect 1409 17085 1443 17119
rect 2789 17085 2823 17119
rect 3065 17085 3099 17119
rect 4813 17085 4847 17119
rect 4997 17085 5031 17119
rect 6193 17085 6227 17119
rect 7113 17085 7147 17119
rect 7573 17085 7607 17119
rect 8953 17085 8987 17119
rect 9413 17085 9447 17119
rect 9965 17085 9999 17119
rect 10517 17085 10551 17119
rect 10977 17085 11011 17119
rect 12449 17085 12483 17119
rect 12909 17085 12943 17119
rect 13277 17085 13311 17119
rect 15428 17085 15462 17119
rect 16221 17085 16255 17119
rect 16451 17085 16485 17119
rect 3249 17017 3283 17051
rect 5549 17017 5583 17051
rect 6653 17017 6687 17051
rect 8217 17017 8251 17051
rect 10425 17017 10459 17051
rect 15531 17017 15565 17051
rect 16865 17017 16899 17051
rect 2329 16949 2363 16983
rect 3525 16949 3559 16983
rect 4169 16949 4203 16983
rect 7389 16949 7423 16983
rect 8769 16949 8803 16983
rect 9229 16949 9263 16983
rect 10793 16949 10827 16983
rect 11529 16949 11563 16983
rect 12265 16949 12299 16983
rect 12541 16949 12575 16983
rect 14381 16949 14415 16983
rect 8217 16745 8251 16779
rect 9413 16745 9447 16779
rect 10701 16745 10735 16779
rect 11391 16745 11425 16779
rect 2237 16677 2271 16711
rect 2789 16677 2823 16711
rect 7297 16677 7331 16711
rect 7389 16677 7423 16711
rect 12449 16677 12483 16711
rect 17463 16677 17497 16711
rect 4997 16609 5031 16643
rect 5273 16609 5307 16643
rect 5825 16609 5859 16643
rect 7021 16609 7055 16643
rect 7941 16609 7975 16643
rect 9689 16609 9723 16643
rect 10149 16609 10183 16643
rect 11320 16609 11354 16643
rect 12725 16609 12759 16643
rect 13185 16609 13219 16643
rect 15368 16609 15402 16643
rect 16313 16609 16347 16643
rect 17325 16609 17359 16643
rect 18404 16609 18438 16643
rect 2145 16541 2179 16575
rect 3433 16541 3467 16575
rect 4629 16541 4663 16575
rect 5457 16541 5491 16575
rect 6837 16541 6871 16575
rect 1961 16473 1995 16507
rect 10241 16541 10275 16575
rect 13461 16541 13495 16575
rect 3065 16405 3099 16439
rect 7021 16405 7055 16439
rect 9045 16405 9079 16439
rect 14289 16405 14323 16439
rect 15439 16405 15473 16439
rect 16451 16405 16485 16439
rect 18475 16405 18509 16439
rect 4813 16201 4847 16235
rect 8033 16201 8067 16235
rect 11161 16201 11195 16235
rect 16313 16201 16347 16235
rect 18889 16201 18923 16235
rect 2789 16133 2823 16167
rect 14105 16133 14139 16167
rect 19211 16133 19245 16167
rect 2145 16065 2179 16099
rect 3157 16065 3191 16099
rect 5917 16065 5951 16099
rect 6837 16065 6871 16099
rect 11897 16065 11931 16099
rect 15393 16065 15427 16099
rect 18199 16065 18233 16099
rect 3433 15997 3467 16031
rect 4445 15997 4479 16031
rect 5181 15997 5215 16031
rect 5641 15997 5675 16031
rect 8861 15997 8895 16031
rect 9045 15997 9079 16031
rect 9689 15997 9723 16031
rect 12909 15997 12943 16031
rect 13093 15997 13127 16031
rect 14289 15997 14323 16031
rect 14749 15997 14783 16031
rect 15920 15997 15954 16031
rect 16681 15997 16715 16031
rect 16916 15997 16950 16031
rect 17969 15997 18003 16031
rect 18337 15997 18371 16031
rect 19140 15997 19174 16031
rect 19533 15997 19567 16031
rect 1869 15929 1903 15963
rect 1961 15929 1995 15963
rect 3341 15929 3375 15963
rect 9321 15929 9355 15963
rect 10241 15929 10275 15963
rect 10333 15929 10367 15963
rect 10885 15929 10919 15963
rect 13369 15929 13403 15963
rect 13645 15929 13679 15963
rect 15025 15929 15059 15963
rect 17003 15929 17037 15963
rect 17785 15929 17819 15963
rect 1685 15861 1719 15895
rect 6653 15861 6687 15895
rect 7205 15861 7239 15895
rect 7757 15861 7791 15895
rect 8401 15861 8435 15895
rect 12265 15861 12299 15895
rect 15991 15861 16025 15895
rect 17417 15861 17451 15895
rect 18337 15861 18371 15895
rect 18521 15861 18555 15895
rect 1777 15657 1811 15691
rect 2329 15657 2363 15691
rect 3341 15657 3375 15691
rect 4261 15657 4295 15691
rect 4813 15657 4847 15691
rect 5273 15657 5307 15691
rect 7205 15657 7239 15691
rect 8585 15657 8619 15691
rect 9505 15657 9539 15691
rect 10609 15657 10643 15691
rect 11345 15657 11379 15691
rect 13093 15657 13127 15691
rect 19257 15657 19291 15691
rect 2605 15589 2639 15623
rect 5911 15589 5945 15623
rect 7481 15589 7515 15623
rect 8033 15589 8067 15623
rect 10010 15589 10044 15623
rect 11621 15589 11655 15623
rect 13782 15589 13816 15623
rect 15485 15589 15519 15623
rect 16037 15589 16071 15623
rect 4077 15521 4111 15555
rect 5549 15521 5583 15555
rect 9689 15521 9723 15555
rect 13461 15521 13495 15555
rect 14381 15521 14415 15555
rect 16932 15521 16966 15555
rect 17912 15521 17946 15555
rect 19073 15521 19107 15555
rect 1409 15453 1443 15487
rect 6837 15453 6871 15487
rect 7389 15453 7423 15487
rect 11529 15453 11563 15487
rect 12173 15453 12207 15487
rect 15393 15453 15427 15487
rect 18015 15453 18049 15487
rect 2973 15317 3007 15351
rect 6469 15317 6503 15351
rect 10885 15317 10919 15351
rect 12725 15317 12759 15351
rect 17003 15317 17037 15351
rect 1961 15113 1995 15147
rect 7205 15113 7239 15147
rect 9045 15113 9079 15147
rect 9781 15113 9815 15147
rect 10977 15113 11011 15147
rect 11529 15113 11563 15147
rect 15209 15113 15243 15147
rect 16313 15113 16347 15147
rect 17325 15113 17359 15147
rect 17785 15113 17819 15147
rect 3065 15045 3099 15079
rect 3433 15045 3467 15079
rect 5089 15045 5123 15079
rect 19211 15045 19245 15079
rect 1547 14977 1581 15011
rect 2513 14977 2547 15011
rect 8125 14977 8159 15011
rect 10057 14977 10091 15011
rect 12909 14977 12943 15011
rect 13553 14977 13587 15011
rect 15393 14977 15427 15011
rect 16037 14977 16071 15011
rect 1460 14909 1494 14943
rect 4236 14909 4270 14943
rect 5917 14909 5951 14943
rect 12484 14909 12518 14943
rect 16773 14909 16807 14943
rect 16900 14909 16934 14943
rect 18096 14909 18130 14943
rect 18521 14909 18555 14943
rect 19124 14909 19158 14943
rect 19533 14909 19567 14943
rect 2605 14841 2639 14875
rect 4629 14841 4663 14875
rect 5273 14841 5307 14875
rect 5365 14841 5399 14875
rect 6285 14841 6319 14875
rect 7849 14841 7883 14875
rect 7941 14841 7975 14875
rect 10310 14841 10344 14875
rect 13804 14841 13838 14875
rect 15485 14841 15519 14875
rect 2329 14773 2363 14807
rect 4307 14773 4341 14807
rect 6561 14773 6595 14807
rect 7665 14773 7699 14807
rect 9413 14773 9447 14807
rect 11805 14773 11839 14807
rect 12587 14773 12621 14807
rect 13369 14773 13403 14807
rect 14473 14773 14507 14807
rect 14749 14773 14783 14807
rect 17003 14773 17037 14807
rect 18199 14773 18233 14807
rect 19901 14773 19935 14807
rect 1685 14569 1719 14603
rect 4629 14569 4663 14603
rect 6285 14569 6319 14603
rect 7021 14569 7055 14603
rect 8493 14569 8527 14603
rect 9965 14569 9999 14603
rect 10425 14569 10459 14603
rect 13921 14569 13955 14603
rect 16957 14569 16991 14603
rect 2237 14501 2271 14535
rect 2789 14501 2823 14535
rect 5083 14501 5117 14535
rect 7935 14501 7969 14535
rect 11161 14501 11195 14535
rect 12725 14501 12759 14535
rect 13645 14501 13679 14535
rect 15485 14501 15519 14535
rect 16037 14501 16071 14535
rect 18567 14501 18601 14535
rect 5641 14433 5675 14467
rect 6596 14433 6630 14467
rect 7573 14433 7607 14467
rect 14140 14433 14174 14467
rect 17141 14433 17175 14467
rect 17417 14433 17451 14467
rect 18429 14433 18463 14467
rect 19476 14433 19510 14467
rect 2145 14365 2179 14399
rect 3433 14365 3467 14399
rect 4721 14365 4755 14399
rect 11069 14365 11103 14399
rect 11713 14365 11747 14399
rect 12357 14365 12391 14399
rect 12633 14365 12667 14399
rect 13001 14365 13035 14399
rect 15393 14365 15427 14399
rect 6699 14297 6733 14331
rect 8769 14297 8803 14331
rect 14243 14297 14277 14331
rect 19579 14297 19613 14331
rect 3065 14229 3099 14263
rect 5917 14229 5951 14263
rect 7481 14229 7515 14263
rect 15117 14229 15151 14263
rect 2329 14025 2363 14059
rect 2973 14025 3007 14059
rect 4813 14025 4847 14059
rect 6653 14025 6687 14059
rect 8539 14025 8573 14059
rect 9229 14025 9263 14059
rect 9597 14025 9631 14059
rect 11345 14025 11379 14059
rect 11897 14025 11931 14059
rect 14105 14025 14139 14059
rect 18521 14025 18555 14059
rect 19901 14025 19935 14059
rect 8217 13957 8251 13991
rect 12173 13957 12207 13991
rect 13461 13957 13495 13991
rect 15485 13957 15519 13991
rect 17141 13957 17175 13991
rect 18889 13957 18923 13991
rect 1409 13889 1443 13923
rect 6929 13889 6963 13923
rect 9781 13889 9815 13923
rect 12541 13889 12575 13923
rect 13829 13889 13863 13923
rect 14289 13889 14323 13923
rect 16129 13889 16163 13923
rect 19533 13889 19567 13923
rect 2605 13821 2639 13855
rect 3617 13821 3651 13855
rect 4077 13821 4111 13855
rect 5457 13821 5491 13855
rect 5733 13821 5767 13855
rect 6193 13821 6227 13855
rect 7849 13821 7883 13855
rect 8436 13821 8470 13855
rect 18096 13821 18130 13855
rect 19140 13821 19174 13855
rect 4353 13753 4387 13787
rect 5917 13753 5951 13787
rect 7021 13753 7055 13787
rect 7573 13753 7607 13787
rect 8861 13753 8895 13787
rect 10102 13753 10136 13787
rect 12862 13753 12896 13787
rect 14610 13753 14644 13787
rect 16221 13753 16255 13787
rect 16773 13753 16807 13787
rect 1777 13685 1811 13719
rect 3525 13685 3559 13719
rect 10701 13685 10735 13719
rect 11069 13685 11103 13719
rect 15209 13685 15243 13719
rect 15853 13685 15887 13719
rect 17417 13685 17451 13719
rect 18199 13685 18233 13719
rect 19211 13685 19245 13719
rect 1547 13481 1581 13515
rect 2329 13481 2363 13515
rect 3709 13481 3743 13515
rect 10977 13481 11011 13515
rect 12541 13481 12575 13515
rect 14657 13481 14691 13515
rect 16957 13481 16991 13515
rect 18521 13481 18555 13515
rect 3157 13413 3191 13447
rect 4721 13413 4755 13447
rect 5410 13413 5444 13447
rect 7021 13413 7055 13447
rect 10010 13413 10044 13447
rect 11621 13413 11655 13447
rect 14289 13413 14323 13447
rect 15485 13413 15519 13447
rect 1444 13345 1478 13379
rect 2605 13345 2639 13379
rect 2973 13345 3007 13379
rect 3985 13345 4019 13379
rect 6009 13345 6043 13379
rect 8436 13345 8470 13379
rect 9689 13345 9723 13379
rect 13277 13345 13311 13379
rect 13461 13345 13495 13379
rect 16957 13345 16991 13379
rect 17325 13345 17359 13379
rect 18429 13345 18463 13379
rect 18889 13345 18923 13379
rect 1869 13277 1903 13311
rect 5089 13277 5123 13311
rect 6929 13277 6963 13311
rect 11529 13277 11563 13311
rect 13553 13277 13587 13311
rect 15393 13277 15427 13311
rect 15669 13277 15703 13311
rect 4215 13209 4249 13243
rect 6653 13209 6687 13243
rect 7481 13209 7515 13243
rect 10609 13209 10643 13243
rect 12081 13209 12115 13243
rect 16405 13209 16439 13243
rect 6377 13141 6411 13175
rect 8539 13141 8573 13175
rect 15117 13141 15151 13175
rect 2605 12937 2639 12971
rect 3801 12937 3835 12971
rect 5089 12937 5123 12971
rect 6285 12937 6319 12971
rect 10057 12937 10091 12971
rect 11621 12937 11655 12971
rect 13461 12937 13495 12971
rect 15209 12937 15243 12971
rect 15393 12937 15427 12971
rect 17785 12937 17819 12971
rect 2789 12869 2823 12903
rect 7481 12869 7515 12903
rect 5273 12801 5307 12835
rect 6929 12801 6963 12835
rect 7941 12801 7975 12835
rect 9137 12801 9171 12835
rect 10701 12801 10735 12835
rect 12817 12801 12851 12835
rect 13921 12801 13955 12835
rect 14381 12801 14415 12835
rect 15025 12801 15059 12835
rect 1409 12733 1443 12767
rect 2697 12733 2731 12767
rect 2973 12733 3007 12767
rect 8401 12733 8435 12767
rect 8493 12733 8527 12767
rect 8677 12733 8711 12767
rect 2237 12665 2271 12699
rect 3433 12665 3467 12699
rect 5365 12665 5399 12699
rect 5917 12665 5951 12699
rect 6653 12665 6687 12699
rect 7021 12665 7055 12699
rect 10793 12665 10827 12699
rect 11345 12665 11379 12699
rect 12541 12665 12575 12699
rect 12633 12665 12667 12699
rect 14473 12665 14507 12699
rect 19441 12869 19475 12903
rect 15945 12801 15979 12835
rect 16589 12801 16623 12835
rect 18061 12733 18095 12767
rect 18521 12733 18555 12767
rect 19073 12733 19107 12767
rect 19676 12733 19710 12767
rect 15761 12665 15795 12699
rect 16037 12665 16071 12699
rect 19763 12665 19797 12699
rect 1593 12597 1627 12631
rect 4077 12597 4111 12631
rect 4445 12597 4479 12631
rect 8309 12597 8343 12631
rect 9689 12597 9723 12631
rect 10517 12597 10551 12631
rect 12173 12597 12207 12631
rect 15209 12597 15243 12631
rect 16865 12597 16899 12631
rect 17325 12597 17359 12631
rect 18153 12597 18187 12631
rect 20085 12597 20119 12631
rect 3157 12393 3191 12427
rect 3525 12393 3559 12427
rect 5273 12393 5307 12427
rect 5549 12393 5583 12427
rect 7297 12393 7331 12427
rect 8861 12393 8895 12427
rect 10885 12393 10919 12427
rect 11529 12393 11563 12427
rect 13369 12393 13403 12427
rect 14657 12393 14691 12427
rect 15117 12393 15151 12427
rect 16405 12393 16439 12427
rect 16957 12393 16991 12427
rect 18061 12393 18095 12427
rect 18521 12393 18555 12427
rect 2881 12325 2915 12359
rect 6054 12325 6088 12359
rect 7665 12325 7699 12359
rect 8493 12325 8527 12359
rect 10286 12325 10320 12359
rect 11897 12325 11931 12359
rect 13823 12325 13857 12359
rect 15393 12325 15427 12359
rect 15485 12325 15519 12359
rect 1685 12257 1719 12291
rect 2145 12257 2179 12291
rect 2421 12257 2455 12291
rect 2789 12257 2823 12291
rect 4445 12257 4479 12291
rect 4721 12257 4755 12291
rect 6653 12257 6687 12291
rect 9965 12257 9999 12291
rect 17049 12257 17083 12291
rect 17417 12257 17451 12291
rect 18429 12257 18463 12291
rect 18889 12257 18923 12291
rect 4905 12189 4939 12223
rect 5733 12189 5767 12223
rect 7573 12189 7607 12223
rect 11805 12189 11839 12223
rect 12081 12189 12115 12223
rect 13461 12189 13495 12223
rect 15669 12189 15703 12223
rect 8125 12121 8159 12155
rect 12817 12121 12851 12155
rect 14381 12121 14415 12155
rect 7021 12053 7055 12087
rect 5365 11849 5399 11883
rect 6469 11849 6503 11883
rect 7849 11849 7883 11883
rect 8217 11849 8251 11883
rect 8539 11849 8573 11883
rect 11161 11849 11195 11883
rect 11805 11849 11839 11883
rect 12817 11849 12851 11883
rect 13093 11849 13127 11883
rect 14197 11849 14231 11883
rect 14841 11849 14875 11883
rect 16037 11849 16071 11883
rect 5733 11781 5767 11815
rect 6101 11781 6135 11815
rect 9413 11781 9447 11815
rect 12173 11781 12207 11815
rect 19763 11781 19797 11815
rect 2881 11713 2915 11747
rect 3617 11713 3651 11747
rect 6929 11713 6963 11747
rect 13277 11713 13311 11747
rect 15117 11713 15151 11747
rect 15485 11713 15519 11747
rect 1685 11645 1719 11679
rect 2145 11645 2179 11679
rect 2421 11645 2455 11679
rect 2697 11645 2731 11679
rect 5549 11645 5583 11679
rect 8468 11645 8502 11679
rect 9597 11645 9631 11679
rect 10793 11645 10827 11679
rect 11380 11645 11414 11679
rect 11483 11645 11517 11679
rect 16656 11645 16690 11679
rect 17509 11645 17543 11679
rect 18153 11645 18187 11679
rect 19073 11645 19107 11679
rect 19660 11645 19694 11679
rect 20085 11645 20119 11679
rect 4077 11577 4111 11611
rect 4169 11577 4203 11611
rect 4721 11577 4755 11611
rect 7021 11577 7055 11611
rect 7573 11577 7607 11611
rect 9918 11577 9952 11611
rect 13639 11577 13673 11611
rect 15209 11577 15243 11611
rect 16497 11577 16531 11611
rect 18061 11577 18095 11611
rect 3249 11509 3283 11543
rect 5089 11509 5123 11543
rect 8953 11509 8987 11543
rect 10517 11509 10551 11543
rect 14565 11509 14599 11543
rect 16727 11509 16761 11543
rect 17141 11509 17175 11543
rect 17785 11509 17819 11543
rect 1961 11305 1995 11339
rect 3433 11305 3467 11339
rect 3893 11305 3927 11339
rect 5181 11305 5215 11339
rect 5733 11305 5767 11339
rect 6285 11305 6319 11339
rect 6837 11305 6871 11339
rect 7113 11305 7147 11339
rect 8401 11305 8435 11339
rect 12541 11305 12575 11339
rect 15117 11305 15151 11339
rect 15485 11305 15519 11339
rect 17785 11305 17819 11339
rect 18705 11305 18739 11339
rect 19441 11305 19475 11339
rect 4261 11237 4295 11271
rect 7573 11237 7607 11271
rect 9965 11237 9999 11271
rect 11707 11237 11741 11271
rect 13001 11237 13035 11271
rect 13185 11237 13219 11271
rect 13277 11237 13311 11271
rect 16313 11237 16347 11271
rect 1476 11169 1510 11203
rect 2697 11169 2731 11203
rect 2881 11169 2915 11203
rect 7941 11169 7975 11203
rect 8217 11169 8251 11203
rect 17877 11169 17911 11203
rect 18245 11169 18279 11203
rect 19257 11169 19291 11203
rect 3065 11101 3099 11135
rect 4169 11101 4203 11135
rect 5917 11101 5951 11135
rect 9873 11101 9907 11135
rect 11345 11101 11379 11135
rect 13645 11101 13679 11135
rect 16221 11101 16255 11135
rect 4721 11033 4755 11067
rect 8033 11033 8067 11067
rect 10425 11033 10459 11067
rect 12265 11033 12299 11067
rect 16773 11033 16807 11067
rect 1547 10965 1581 10999
rect 2329 10965 2363 10999
rect 9505 10965 9539 10999
rect 3985 10761 4019 10795
rect 4537 10761 4571 10795
rect 6009 10761 6043 10795
rect 6285 10761 6319 10795
rect 7113 10761 7147 10795
rect 8677 10761 8711 10795
rect 10517 10761 10551 10795
rect 10793 10761 10827 10795
rect 12265 10761 12299 10795
rect 13461 10761 13495 10795
rect 13829 10761 13863 10795
rect 15669 10761 15703 10795
rect 16037 10761 16071 10795
rect 20177 10761 20211 10795
rect 4629 10693 4663 10727
rect 9321 10693 9355 10727
rect 13093 10693 13127 10727
rect 17417 10693 17451 10727
rect 17785 10693 17819 10727
rect 3065 10625 3099 10659
rect 4537 10625 4571 10659
rect 7665 10625 7699 10659
rect 9505 10625 9539 10659
rect 11483 10625 11517 10659
rect 14565 10625 14599 10659
rect 15301 10625 15335 10659
rect 16221 10625 16255 10659
rect 19763 10625 19797 10659
rect 1777 10557 1811 10591
rect 2053 10557 2087 10591
rect 2513 10557 2547 10591
rect 4353 10557 4387 10591
rect 4997 10557 5031 10591
rect 5273 10557 5307 10591
rect 11380 10557 11414 10591
rect 11805 10557 11839 10591
rect 14013 10557 14047 10591
rect 14473 10557 14507 10591
rect 18245 10557 18279 10591
rect 18521 10557 18555 10591
rect 19676 10557 19710 10591
rect 2973 10489 3007 10523
rect 3386 10489 3420 10523
rect 7389 10489 7423 10523
rect 7481 10489 7515 10523
rect 9597 10489 9631 10523
rect 10149 10489 10183 10523
rect 12541 10489 12575 10523
rect 12633 10489 12667 10523
rect 16313 10489 16347 10523
rect 16865 10489 16899 10523
rect 1593 10421 1627 10455
rect 4905 10421 4939 10455
rect 8401 10421 8435 10455
rect 11253 10421 11287 10455
rect 18153 10421 18187 10455
rect 19349 10421 19383 10455
rect 2605 10217 2639 10251
rect 3709 10217 3743 10251
rect 4261 10217 4295 10251
rect 5549 10217 5583 10251
rect 6331 10217 6365 10251
rect 6837 10217 6871 10251
rect 10057 10217 10091 10251
rect 10885 10217 10919 10251
rect 12173 10217 12207 10251
rect 16221 10217 16255 10251
rect 16497 10217 16531 10251
rect 16865 10217 16899 10251
rect 18061 10217 18095 10251
rect 18705 10217 18739 10251
rect 1777 10149 1811 10183
rect 4629 10149 4663 10183
rect 5181 10149 5215 10183
rect 5273 10149 5307 10183
rect 7389 10149 7423 10183
rect 13179 10149 13213 10183
rect 15622 10149 15656 10183
rect 17141 10149 17175 10183
rect 17233 10149 17267 10183
rect 2973 10081 3007 10115
rect 1685 10013 1719 10047
rect 4537 10013 4571 10047
rect 6260 10081 6294 10115
rect 9505 10081 9539 10115
rect 10609 10081 10643 10115
rect 11437 10081 11471 10115
rect 18613 10081 18647 10115
rect 19073 10081 19107 10115
rect 7297 10013 7331 10047
rect 7573 10013 7607 10047
rect 9689 10013 9723 10047
rect 12817 10013 12851 10047
rect 15301 10013 15335 10047
rect 17417 10013 17451 10047
rect 2237 9945 2271 9979
rect 5273 9945 5307 9979
rect 3433 9877 3467 9911
rect 5825 9877 5859 9911
rect 8217 9877 8251 9911
rect 11621 9877 11655 9911
rect 12449 9877 12483 9911
rect 13737 9877 13771 9911
rect 14105 9877 14139 9911
rect 18521 9877 18555 9911
rect 2329 9673 2363 9707
rect 2973 9673 3007 9707
rect 4721 9673 4755 9707
rect 4997 9673 5031 9707
rect 5365 9673 5399 9707
rect 8677 9673 8711 9707
rect 9965 9673 9999 9707
rect 10425 9673 10459 9707
rect 11529 9673 11563 9707
rect 14565 9673 14599 9707
rect 14933 9673 14967 9707
rect 16037 9673 16071 9707
rect 16773 9673 16807 9707
rect 19073 9673 19107 9707
rect 11805 9605 11839 9639
rect 12265 9605 12299 9639
rect 17049 9605 17083 9639
rect 3801 9537 3835 9571
rect 6837 9537 6871 9571
rect 9505 9537 9539 9571
rect 10609 9537 10643 9571
rect 13461 9537 13495 9571
rect 13737 9537 13771 9571
rect 16405 9537 16439 9571
rect 19441 9537 19475 9571
rect 1409 9469 1443 9503
rect 5733 9469 5767 9503
rect 9045 9469 9079 9503
rect 9321 9469 9355 9503
rect 15117 9469 15151 9503
rect 16865 9469 16899 9503
rect 17417 9469 17451 9503
rect 18153 9469 18187 9503
rect 19660 9469 19694 9503
rect 20085 9469 20119 9503
rect 1771 9401 1805 9435
rect 3617 9401 3651 9435
rect 4163 9401 4197 9435
rect 10971 9401 11005 9435
rect 13553 9401 13587 9435
rect 15438 9401 15472 9435
rect 19763 9401 19797 9435
rect 2605 9333 2639 9367
rect 6285 9333 6319 9367
rect 6653 9333 6687 9367
rect 7205 9333 7239 9367
rect 7757 9333 7791 9367
rect 8033 9333 8067 9367
rect 12817 9333 12851 9367
rect 13277 9333 13311 9367
rect 17785 9333 17819 9367
rect 18337 9333 18371 9367
rect 1593 9129 1627 9163
rect 2881 9129 2915 9163
rect 3249 9129 3283 9163
rect 3801 9129 3835 9163
rect 4445 9129 4479 9163
rect 7297 9129 7331 9163
rect 8217 9129 8251 9163
rect 9965 9129 9999 9163
rect 12357 9129 12391 9163
rect 13553 9129 13587 9163
rect 15577 9129 15611 9163
rect 6377 9061 6411 9095
rect 11345 9061 11379 9095
rect 12541 9061 12575 9095
rect 12633 9061 12667 9095
rect 16405 9061 16439 9095
rect 1777 8993 1811 9027
rect 2053 8993 2087 9027
rect 6929 8993 6963 9027
rect 7757 8993 7791 9027
rect 8033 8993 8067 9027
rect 10609 8993 10643 9027
rect 11069 8993 11103 9027
rect 14105 8993 14139 9027
rect 17785 8993 17819 9027
rect 17932 8993 17966 9027
rect 19349 8993 19383 9027
rect 4077 8925 4111 8959
rect 6285 8925 6319 8959
rect 12817 8925 12851 8959
rect 16313 8925 16347 8959
rect 16773 8925 16807 8959
rect 17601 8925 17635 8959
rect 18153 8925 18187 8959
rect 7849 8857 7883 8891
rect 17325 8857 17359 8891
rect 2513 8789 2547 8823
rect 4997 8789 5031 8823
rect 8861 8789 8895 8823
rect 14289 8789 14323 8823
rect 18061 8789 18095 8823
rect 18245 8789 18279 8823
rect 18797 8789 18831 8823
rect 19533 8789 19567 8823
rect 1685 8585 1719 8619
rect 2881 8585 2915 8619
rect 3433 8585 3467 8619
rect 5917 8585 5951 8619
rect 6469 8585 6503 8619
rect 6561 8585 6595 8619
rect 7849 8585 7883 8619
rect 8217 8585 8251 8619
rect 10057 8585 10091 8619
rect 11897 8585 11931 8619
rect 13921 8585 13955 8619
rect 15945 8585 15979 8619
rect 17877 8585 17911 8619
rect 19349 8585 19383 8619
rect 4997 8517 5031 8551
rect 5549 8517 5583 8551
rect 2421 8449 2455 8483
rect 3801 8449 3835 8483
rect 6929 8517 6963 8551
rect 15577 8517 15611 8551
rect 8953 8449 8987 8483
rect 10609 8449 10643 8483
rect 12541 8449 12575 8483
rect 13185 8449 13219 8483
rect 14105 8449 14139 8483
rect 14381 8449 14415 8483
rect 16773 8449 16807 8483
rect 18153 8449 18187 8483
rect 18613 8449 18647 8483
rect 6469 8381 6503 8415
rect 6837 8381 6871 8415
rect 7113 8381 7147 8415
rect 7573 8381 7607 8415
rect 8677 8381 8711 8415
rect 8861 8381 8895 8415
rect 11529 8381 11563 8415
rect 12173 8381 12207 8415
rect 19660 8381 19694 8415
rect 20085 8381 20119 8415
rect 1961 8313 1995 8347
rect 2053 8313 2087 8347
rect 4445 8313 4479 8347
rect 4537 8313 4571 8347
rect 6285 8313 6319 8347
rect 10930 8313 10964 8347
rect 12633 8313 12667 8347
rect 14197 8313 14231 8347
rect 16497 8313 16531 8347
rect 16589 8313 16623 8347
rect 18245 8313 18279 8347
rect 19763 8313 19797 8347
rect 4077 8245 4111 8279
rect 9505 8245 9539 8279
rect 10517 8245 10551 8279
rect 13553 8245 13587 8279
rect 16313 8245 16347 8279
rect 17417 8245 17451 8279
rect 3065 8041 3099 8075
rect 3341 8041 3375 8075
rect 4261 8041 4295 8075
rect 5181 8041 5215 8075
rect 8401 8041 8435 8075
rect 8769 8041 8803 8075
rect 10701 8041 10735 8075
rect 12541 8041 12575 8075
rect 12909 8041 12943 8075
rect 14381 8041 14415 8075
rect 16497 8041 16531 8075
rect 18705 8041 18739 8075
rect 1771 7973 1805 8007
rect 3709 7973 3743 8007
rect 6561 7973 6595 8007
rect 11339 7973 11373 8007
rect 13547 7973 13581 8007
rect 15622 7973 15656 8007
rect 17141 7973 17175 8007
rect 17233 7973 17267 8007
rect 1409 7905 1443 7939
rect 4077 7905 4111 7939
rect 5365 7905 5399 7939
rect 5733 7905 5767 7939
rect 6377 7905 6411 7939
rect 7297 7905 7331 7939
rect 7389 7905 7423 7939
rect 10032 7905 10066 7939
rect 10977 7905 11011 7939
rect 15301 7905 15335 7939
rect 18613 7905 18647 7939
rect 19073 7905 19107 7939
rect 4813 7837 4847 7871
rect 7757 7837 7791 7871
rect 8125 7837 8159 7871
rect 13185 7837 13219 7871
rect 17417 7837 17451 7871
rect 18061 7837 18095 7871
rect 7527 7769 7561 7803
rect 11897 7769 11931 7803
rect 16221 7769 16255 7803
rect 2329 7701 2363 7735
rect 2605 7701 2639 7735
rect 6837 7701 6871 7735
rect 7665 7701 7699 7735
rect 10103 7701 10137 7735
rect 14105 7701 14139 7735
rect 18521 7701 18555 7735
rect 4169 7497 4203 7531
rect 5825 7497 5859 7531
rect 8401 7497 8435 7531
rect 10241 7497 10275 7531
rect 15209 7497 15243 7531
rect 17417 7497 17451 7531
rect 17877 7497 17911 7531
rect 19073 7497 19107 7531
rect 7205 7429 7239 7463
rect 7665 7429 7699 7463
rect 8861 7429 8895 7463
rect 12173 7429 12207 7463
rect 14197 7429 14231 7463
rect 14657 7429 14691 7463
rect 16497 7429 16531 7463
rect 17141 7429 17175 7463
rect 18153 7429 18187 7463
rect 1501 7361 1535 7395
rect 2973 7361 3007 7395
rect 4813 7361 4847 7395
rect 5089 7361 5123 7395
rect 6653 7361 6687 7395
rect 7757 7361 7791 7395
rect 8125 7361 8159 7395
rect 10609 7361 10643 7395
rect 13185 7361 13219 7395
rect 13921 7361 13955 7395
rect 19763 7361 19797 7395
rect 3893 7293 3927 7327
rect 4537 7293 4571 7327
rect 7536 7293 7570 7327
rect 8953 7293 8987 7327
rect 10793 7293 10827 7327
rect 11253 7293 11287 7327
rect 14013 7293 14047 7327
rect 15301 7293 15335 7327
rect 16221 7293 16255 7327
rect 18061 7293 18095 7327
rect 18337 7293 18371 7327
rect 19676 7293 19710 7327
rect 1593 7225 1627 7259
rect 2145 7225 2179 7259
rect 3294 7225 3328 7259
rect 4905 7225 4939 7259
rect 7389 7225 7423 7259
rect 11529 7225 11563 7259
rect 12541 7225 12575 7259
rect 12633 7225 12667 7259
rect 15622 7225 15656 7259
rect 18797 7225 18831 7259
rect 2421 7157 2455 7191
rect 2789 7157 2823 7191
rect 6193 7157 6227 7191
rect 9321 7157 9355 7191
rect 9873 7157 9907 7191
rect 11897 7157 11931 7191
rect 13553 7157 13587 7191
rect 19441 7157 19475 7191
rect 20177 7157 20211 7191
rect 1409 6953 1443 6987
rect 2237 6953 2271 6987
rect 6929 6953 6963 6987
rect 7297 6953 7331 6987
rect 9045 6953 9079 6987
rect 9321 6953 9355 6987
rect 10793 6953 10827 6987
rect 11161 6953 11195 6987
rect 14381 6953 14415 6987
rect 15117 6953 15151 6987
rect 15853 6953 15887 6987
rect 17509 6953 17543 6987
rect 18153 6953 18187 6987
rect 4261 6885 4295 6919
rect 9873 6885 9907 6919
rect 10425 6885 10459 6919
rect 11805 6885 11839 6919
rect 13001 6885 13035 6919
rect 13553 6885 13587 6919
rect 16681 6885 16715 6919
rect 17233 6885 17267 6919
rect 2697 6817 2731 6851
rect 2881 6817 2915 6851
rect 5641 6817 5675 6851
rect 5917 6817 5951 6851
rect 7389 6817 7423 6851
rect 7849 6817 7883 6851
rect 8493 6817 8527 6851
rect 14105 6817 14139 6851
rect 15301 6817 15335 6851
rect 18245 6817 18279 6851
rect 18521 6817 18555 6851
rect 19660 6817 19694 6851
rect 3157 6749 3191 6783
rect 3893 6749 3927 6783
rect 4169 6749 4203 6783
rect 6101 6749 6135 6783
rect 7941 6749 7975 6783
rect 9781 6749 9815 6783
rect 11713 6749 11747 6783
rect 12357 6749 12391 6783
rect 13461 6749 13495 6783
rect 16589 6749 16623 6783
rect 4721 6681 4755 6715
rect 5733 6681 5767 6715
rect 12725 6681 12759 6715
rect 15485 6681 15519 6715
rect 1869 6613 1903 6647
rect 5365 6613 5399 6647
rect 16221 6613 16255 6647
rect 19763 6613 19797 6647
rect 3157 6409 3191 6443
rect 3985 6409 4019 6443
rect 5273 6409 5307 6443
rect 5871 6409 5905 6443
rect 13553 6409 13587 6443
rect 15393 6409 15427 6443
rect 16865 6409 16899 6443
rect 17509 6409 17543 6443
rect 19073 6409 19107 6443
rect 20453 6409 20487 6443
rect 2421 6341 2455 6375
rect 7481 6341 7515 6375
rect 9229 6341 9263 6375
rect 9781 6341 9815 6375
rect 16497 6341 16531 6375
rect 1869 6273 1903 6307
rect 4169 6273 4203 6307
rect 4813 6273 4847 6307
rect 6929 6273 6963 6307
rect 7849 6273 7883 6307
rect 8677 6273 8711 6307
rect 12541 6273 12575 6307
rect 12909 6273 12943 6307
rect 14105 6273 14139 6307
rect 19763 6273 19797 6307
rect 2881 6205 2915 6239
rect 5768 6205 5802 6239
rect 6561 6205 6595 6239
rect 10333 6205 10367 6239
rect 18245 6205 18279 6239
rect 18521 6205 18555 6239
rect 19676 6205 19710 6239
rect 20085 6205 20119 6239
rect 1961 6137 1995 6171
rect 3617 6137 3651 6171
rect 4261 6137 4295 6171
rect 6285 6137 6319 6171
rect 7021 6137 7055 6171
rect 8217 6137 8251 6171
rect 8769 6137 8803 6171
rect 10241 6137 10275 6171
rect 10695 6137 10729 6171
rect 12633 6137 12667 6171
rect 14013 6137 14047 6171
rect 14426 6137 14460 6171
rect 15669 6137 15703 6171
rect 15945 6137 15979 6171
rect 16037 6137 16071 6171
rect 17785 6137 17819 6171
rect 1685 6069 1719 6103
rect 5641 6069 5675 6103
rect 11253 6069 11287 6103
rect 11621 6069 11655 6103
rect 12173 6069 12207 6103
rect 15025 6069 15059 6103
rect 18153 6069 18187 6103
rect 2329 5865 2363 5899
rect 3433 5865 3467 5899
rect 4997 5865 5031 5899
rect 5549 5865 5583 5899
rect 7481 5865 7515 5899
rect 9873 5865 9907 5899
rect 11345 5865 11379 5899
rect 11713 5865 11747 5899
rect 18521 5865 18555 5899
rect 1771 5797 1805 5831
rect 2605 5797 2639 5831
rect 4439 5797 4473 5831
rect 6371 5797 6405 5831
rect 8211 5797 8245 5831
rect 10787 5797 10821 5831
rect 12357 5797 12391 5831
rect 13369 5797 13403 5831
rect 15485 5797 15519 5831
rect 16589 5797 16623 5831
rect 17049 5797 17083 5831
rect 3065 5729 3099 5763
rect 4077 5729 4111 5763
rect 7849 5729 7883 5763
rect 14105 5729 14139 5763
rect 18613 5729 18647 5763
rect 18889 5729 18923 5763
rect 1409 5661 1443 5695
rect 6009 5661 6043 5695
rect 10425 5661 10459 5695
rect 12265 5661 12299 5695
rect 12909 5661 12943 5695
rect 15393 5661 15427 5695
rect 16037 5661 16071 5695
rect 16957 5661 16991 5695
rect 17233 5661 17267 5695
rect 10333 5593 10367 5627
rect 3801 5525 3835 5559
rect 5917 5525 5951 5559
rect 6929 5525 6963 5559
rect 8769 5525 8803 5559
rect 9045 5525 9079 5559
rect 14289 5525 14323 5559
rect 15117 5525 15151 5559
rect 18061 5525 18095 5559
rect 3065 5321 3099 5355
rect 4997 5321 5031 5355
rect 6653 5321 6687 5355
rect 7849 5321 7883 5355
rect 9781 5321 9815 5355
rect 11805 5321 11839 5355
rect 12081 5321 12115 5355
rect 12265 5321 12299 5355
rect 13921 5321 13955 5355
rect 14933 5321 14967 5355
rect 15301 5321 15335 5355
rect 19073 5321 19107 5355
rect 2329 5253 2363 5287
rect 3617 5253 3651 5287
rect 10057 5253 10091 5287
rect 1777 5185 1811 5219
rect 7205 5185 7239 5219
rect 8861 5185 8895 5219
rect 10517 5185 10551 5219
rect 3801 5117 3835 5151
rect 5800 5117 5834 5151
rect 10793 5117 10827 5151
rect 11345 5117 11379 5151
rect 16865 5253 16899 5287
rect 19763 5253 19797 5287
rect 12817 5185 12851 5219
rect 13553 5185 13587 5219
rect 14013 5185 14047 5219
rect 16497 5117 16531 5151
rect 18153 5117 18187 5151
rect 19692 5117 19726 5151
rect 20085 5117 20119 5151
rect 1869 5049 1903 5083
rect 4122 5049 4156 5083
rect 6929 5049 6963 5083
rect 7021 5049 7055 5083
rect 8585 5049 8619 5083
rect 8677 5049 8711 5083
rect 11529 5049 11563 5083
rect 12081 5049 12115 5083
rect 12541 5049 12575 5083
rect 12633 5049 12667 5083
rect 14334 5049 14368 5083
rect 15853 5049 15887 5083
rect 15945 5049 15979 5083
rect 18061 5049 18095 5083
rect 2697 4981 2731 5015
rect 4721 4981 4755 5015
rect 5641 4981 5675 5015
rect 5871 4981 5905 5015
rect 6285 4981 6319 5015
rect 8401 4981 8435 5015
rect 17233 4981 17267 5015
rect 17785 4981 17819 5015
rect 19533 4981 19567 5015
rect 3433 4777 3467 4811
rect 7481 4777 7515 4811
rect 7941 4777 7975 4811
rect 9137 4777 9171 4811
rect 10977 4777 11011 4811
rect 12449 4777 12483 4811
rect 12817 4777 12851 4811
rect 15117 4777 15151 4811
rect 16313 4777 16347 4811
rect 16957 4777 16991 4811
rect 18705 4777 18739 4811
rect 1409 4709 1443 4743
rect 3801 4709 3835 4743
rect 4261 4709 4295 4743
rect 4353 4709 4387 4743
rect 4905 4709 4939 4743
rect 6653 4709 6687 4743
rect 7205 4709 7239 4743
rect 8217 4709 8251 4743
rect 11345 4709 11379 4743
rect 11529 4709 11563 4743
rect 11621 4709 11655 4743
rect 13185 4709 13219 4743
rect 15485 4709 15519 4743
rect 18153 4709 18187 4743
rect 2697 4641 2731 4675
rect 2881 4641 2915 4675
rect 3157 4641 3191 4675
rect 9873 4641 9907 4675
rect 10425 4641 10459 4675
rect 17141 4641 17175 4675
rect 17325 4641 17359 4675
rect 18521 4641 18555 4675
rect 6009 4573 6043 4607
rect 6561 4573 6595 4607
rect 8125 4573 8159 4607
rect 10609 4573 10643 4607
rect 12173 4573 12207 4607
rect 13093 4573 13127 4607
rect 13369 4573 13403 4607
rect 14749 4573 14783 4607
rect 15393 4573 15427 4607
rect 2329 4505 2363 4539
rect 6377 4505 6411 4539
rect 8677 4505 8711 4539
rect 15945 4505 15979 4539
rect 1869 4437 1903 4471
rect 14105 4437 14139 4471
rect 16681 4437 16715 4471
rect 1777 4233 1811 4267
rect 2145 4233 2179 4267
rect 3249 4233 3283 4267
rect 4813 4233 4847 4267
rect 8125 4233 8159 4267
rect 9505 4233 9539 4267
rect 9965 4233 9999 4267
rect 13921 4233 13955 4267
rect 19073 4233 19107 4267
rect 4537 4097 4571 4131
rect 5273 4097 5307 4131
rect 5917 4097 5951 4131
rect 12817 4097 12851 4131
rect 16221 4097 16255 4131
rect 16497 4097 16531 4131
rect 19763 4097 19797 4131
rect 2513 4029 2547 4063
rect 2789 4029 2823 4063
rect 5549 4029 5583 4063
rect 6837 4029 6871 4063
rect 8585 4029 8619 4063
rect 10517 4029 10551 4063
rect 11437 4029 11471 4063
rect 12173 4029 12207 4063
rect 14657 4029 14691 4063
rect 15577 4029 15611 4063
rect 18153 4029 18187 4063
rect 18521 4029 18555 4063
rect 19660 4029 19694 4063
rect 20085 4029 20119 4063
rect 2973 3961 3007 3995
rect 3893 3961 3927 3995
rect 3985 3961 4019 3995
rect 5365 3961 5399 3995
rect 6193 3961 6227 3995
rect 7158 3961 7192 3995
rect 8401 3961 8435 3995
rect 8906 3961 8940 3995
rect 10333 3961 10367 3995
rect 10838 3961 10872 3995
rect 12541 3961 12575 3995
rect 12633 3961 12667 3995
rect 15853 3961 15887 3995
rect 16589 3961 16623 3995
rect 17141 3961 17175 3995
rect 3617 3893 3651 3927
rect 6561 3893 6595 3927
rect 7757 3893 7791 3927
rect 11713 3893 11747 3927
rect 13461 3893 13495 3927
rect 14565 3893 14599 3927
rect 15025 3893 15059 3927
rect 17417 3893 17451 3927
rect 17785 3893 17819 3927
rect 18153 3893 18187 3927
rect 1409 3689 1443 3723
rect 5273 3689 5307 3723
rect 7113 3689 7147 3723
rect 7941 3689 7975 3723
rect 9045 3689 9079 3723
rect 9781 3689 9815 3723
rect 13093 3689 13127 3723
rect 14197 3689 14231 3723
rect 15117 3689 15151 3723
rect 16497 3689 16531 3723
rect 18521 3689 18555 3723
rect 2329 3621 2363 3655
rect 3433 3621 3467 3655
rect 4398 3621 4432 3655
rect 6238 3621 6272 3655
rect 8217 3621 8251 3655
rect 9413 3621 9447 3655
rect 11621 3621 11655 3655
rect 12173 3621 12207 3655
rect 12449 3621 12483 3655
rect 13639 3621 13673 3655
rect 14657 3621 14691 3655
rect 15485 3621 15519 3655
rect 2697 3553 2731 3587
rect 2973 3553 3007 3587
rect 3893 3553 3927 3587
rect 4997 3553 5031 3587
rect 9965 3553 9999 3587
rect 10149 3553 10183 3587
rect 13277 3553 13311 3587
rect 17141 3553 17175 3587
rect 17325 3553 17359 3587
rect 18429 3553 18463 3587
rect 18981 3553 19015 3587
rect 3157 3485 3191 3519
rect 4077 3485 4111 3519
rect 5917 3485 5951 3519
rect 8125 3485 8159 3519
rect 8401 3485 8435 3519
rect 11161 3485 11195 3519
rect 11529 3485 11563 3519
rect 15393 3485 15427 3519
rect 17417 3485 17451 3519
rect 1961 3417 1995 3451
rect 6837 3417 6871 3451
rect 15945 3417 15979 3451
rect 5825 3349 5859 3383
rect 7573 3349 7607 3383
rect 10793 3349 10827 3383
rect 18153 3349 18187 3383
rect 2881 3145 2915 3179
rect 8125 3145 8159 3179
rect 8769 3145 8803 3179
rect 11437 3145 11471 3179
rect 13093 3145 13127 3179
rect 14841 3145 14875 3179
rect 15209 3145 15243 3179
rect 15577 3145 15611 3179
rect 17233 3145 17267 3179
rect 19441 3145 19475 3179
rect 4629 3077 4663 3111
rect 6561 3077 6595 3111
rect 12633 3077 12667 3111
rect 16957 3077 16991 3111
rect 5273 3009 5307 3043
rect 6929 3009 6963 3043
rect 8953 3009 8987 3043
rect 9965 3009 9999 3043
rect 10517 3009 10551 3043
rect 11713 3009 11747 3043
rect 15761 3009 15795 3043
rect 16405 3009 16439 3043
rect 19763 3009 19797 3043
rect 1777 2941 1811 2975
rect 2053 2941 2087 2975
rect 2237 2941 2271 2975
rect 3617 2941 3651 2975
rect 4215 2941 4249 2975
rect 12449 2941 12483 2975
rect 13921 2941 13955 2975
rect 18061 2941 18095 2975
rect 18521 2941 18555 2975
rect 19676 2941 19710 2975
rect 20085 2941 20119 2975
rect 4353 2873 4387 2907
rect 5089 2873 5123 2907
rect 5365 2873 5399 2907
rect 5917 2873 5951 2907
rect 7021 2873 7055 2907
rect 7573 2873 7607 2907
rect 9045 2873 9079 2907
rect 9597 2873 9631 2907
rect 10838 2873 10872 2907
rect 13737 2873 13771 2907
rect 14242 2873 14276 2907
rect 15853 2873 15887 2907
rect 19073 2873 19107 2907
rect 2605 2805 2639 2839
rect 3525 2805 3559 2839
rect 6193 2805 6227 2839
rect 10333 2805 10367 2839
rect 12081 2805 12115 2839
rect 13369 2805 13403 2839
rect 17785 2805 17819 2839
rect 18153 2805 18187 2839
rect 1409 2601 1443 2635
rect 3617 2601 3651 2635
rect 6009 2601 6043 2635
rect 7389 2601 7423 2635
rect 7849 2601 7883 2635
rect 8861 2601 8895 2635
rect 9137 2601 9171 2635
rect 10057 2601 10091 2635
rect 11437 2601 11471 2635
rect 14289 2601 14323 2635
rect 16957 2601 16991 2635
rect 18061 2601 18095 2635
rect 18429 2601 18463 2635
rect 2329 2533 2363 2567
rect 3157 2533 3191 2567
rect 4629 2533 4663 2567
rect 5410 2533 5444 2567
rect 8262 2533 8296 2567
rect 10333 2533 10367 2567
rect 10838 2533 10872 2567
rect 13185 2533 13219 2567
rect 13690 2533 13724 2567
rect 14565 2533 14599 2567
rect 15669 2533 15703 2567
rect 16497 2533 16531 2567
rect 19349 2533 19383 2567
rect 1961 2465 1995 2499
rect 2513 2465 2547 2499
rect 2973 2465 3007 2499
rect 4144 2465 4178 2499
rect 5089 2465 5123 2499
rect 6996 2465 7030 2499
rect 10517 2465 10551 2499
rect 11713 2465 11747 2499
rect 12081 2465 12115 2499
rect 12909 2465 12943 2499
rect 13369 2465 13403 2499
rect 17141 2465 17175 2499
rect 17693 2465 17727 2499
rect 18337 2465 18371 2499
rect 18889 2465 18923 2499
rect 7941 2397 7975 2431
rect 9505 2397 9539 2431
rect 15577 2397 15611 2431
rect 15853 2397 15887 2431
rect 4215 2329 4249 2363
rect 6745 2329 6779 2363
rect 17325 2329 17359 2363
rect 4905 2261 4939 2295
rect 6377 2261 6411 2295
rect 7067 2261 7101 2295
rect 15209 2261 15243 2295
<< metal1 >>
rect 1104 19610 20884 19632
rect 1104 19558 4648 19610
rect 4700 19558 4712 19610
rect 4764 19558 4776 19610
rect 4828 19558 4840 19610
rect 4892 19558 11982 19610
rect 12034 19558 12046 19610
rect 12098 19558 12110 19610
rect 12162 19558 12174 19610
rect 12226 19558 19315 19610
rect 19367 19558 19379 19610
rect 19431 19558 19443 19610
rect 19495 19558 19507 19610
rect 19559 19558 20884 19610
rect 1104 19536 20884 19558
rect 4246 19456 4252 19508
rect 4304 19496 4310 19508
rect 13771 19499 13829 19505
rect 13771 19496 13783 19499
rect 4304 19468 13783 19496
rect 4304 19456 4310 19468
rect 13771 19465 13783 19468
rect 13817 19465 13829 19499
rect 13771 19459 13829 19465
rect 6730 19388 6736 19440
rect 6788 19428 6794 19440
rect 10919 19431 10977 19437
rect 10919 19428 10931 19431
rect 6788 19400 10931 19428
rect 6788 19388 6794 19400
rect 10919 19397 10931 19400
rect 10965 19397 10977 19431
rect 10919 19391 10977 19397
rect 4154 19320 4160 19372
rect 4212 19360 4218 19372
rect 5442 19360 5448 19372
rect 4212 19332 5448 19360
rect 4212 19320 4218 19332
rect 5442 19320 5448 19332
rect 5500 19320 5506 19372
rect 7006 19320 7012 19372
rect 7064 19360 7070 19372
rect 9907 19363 9965 19369
rect 9907 19360 9919 19363
rect 7064 19332 9919 19360
rect 7064 19320 7070 19332
rect 9907 19329 9919 19332
rect 9953 19329 9965 19363
rect 9907 19323 9965 19329
rect 1949 19295 2007 19301
rect 1949 19261 1961 19295
rect 1995 19292 2007 19295
rect 2130 19292 2136 19304
rect 1995 19264 2136 19292
rect 1995 19261 2007 19264
rect 1949 19255 2007 19261
rect 2130 19252 2136 19264
rect 2188 19252 2194 19304
rect 4062 19292 4068 19304
rect 4023 19264 4068 19292
rect 4062 19252 4068 19264
rect 4120 19252 4126 19304
rect 4338 19292 4344 19304
rect 4166 19264 4344 19292
rect 2314 19184 2320 19236
rect 2372 19224 2378 19236
rect 3789 19227 3847 19233
rect 3789 19224 3801 19227
rect 2372 19196 3801 19224
rect 2372 19184 2378 19196
rect 3789 19193 3801 19196
rect 3835 19224 3847 19227
rect 4166 19224 4194 19264
rect 4338 19252 4344 19264
rect 4396 19252 4402 19304
rect 4801 19295 4859 19301
rect 4801 19261 4813 19295
rect 4847 19292 4859 19295
rect 4982 19292 4988 19304
rect 4847 19264 4988 19292
rect 4847 19261 4859 19264
rect 4801 19255 4859 19261
rect 4982 19252 4988 19264
rect 5040 19252 5046 19304
rect 5534 19252 5540 19304
rect 5592 19292 5598 19304
rect 5664 19295 5722 19301
rect 5664 19292 5676 19295
rect 5592 19264 5676 19292
rect 5592 19252 5598 19264
rect 5664 19261 5676 19264
rect 5710 19292 5722 19295
rect 6089 19295 6147 19301
rect 6089 19292 6101 19295
rect 5710 19264 6101 19292
rect 5710 19261 5722 19264
rect 5664 19255 5722 19261
rect 6089 19261 6101 19264
rect 6135 19261 6147 19295
rect 6089 19255 6147 19261
rect 6454 19252 6460 19304
rect 6512 19292 6518 19304
rect 6917 19295 6975 19301
rect 6917 19292 6929 19295
rect 6512 19264 6929 19292
rect 6512 19252 6518 19264
rect 6917 19261 6929 19264
rect 6963 19261 6975 19295
rect 6917 19255 6975 19261
rect 7282 19252 7288 19304
rect 7340 19292 7346 19304
rect 7377 19295 7435 19301
rect 7377 19292 7389 19295
rect 7340 19264 7389 19292
rect 7340 19252 7346 19264
rect 7377 19261 7389 19264
rect 7423 19261 7435 19295
rect 7377 19255 7435 19261
rect 9820 19295 9878 19301
rect 9820 19261 9832 19295
rect 9866 19292 9878 19295
rect 10229 19295 10287 19301
rect 10229 19292 10241 19295
rect 9866 19264 10241 19292
rect 9866 19261 9878 19264
rect 9820 19255 9878 19261
rect 10229 19261 10241 19264
rect 10275 19292 10287 19295
rect 10318 19292 10324 19304
rect 10275 19264 10324 19292
rect 10275 19261 10287 19264
rect 10229 19255 10287 19261
rect 10318 19252 10324 19264
rect 10376 19252 10382 19304
rect 10827 19295 10885 19301
rect 10827 19261 10839 19295
rect 10873 19261 10885 19295
rect 10827 19255 10885 19261
rect 5077 19227 5135 19233
rect 5077 19224 5089 19227
rect 3835 19196 4194 19224
rect 4223 19196 5089 19224
rect 3835 19193 3847 19196
rect 3789 19187 3847 19193
rect 2501 19159 2559 19165
rect 2501 19125 2513 19159
rect 2547 19156 2559 19159
rect 2590 19156 2596 19168
rect 2547 19128 2596 19156
rect 2547 19125 2559 19128
rect 2501 19119 2559 19125
rect 2590 19116 2596 19128
rect 2648 19116 2654 19168
rect 2866 19116 2872 19168
rect 2924 19156 2930 19168
rect 3418 19156 3424 19168
rect 2924 19128 3424 19156
rect 2924 19116 2930 19128
rect 3418 19116 3424 19128
rect 3476 19116 3482 19168
rect 4062 19116 4068 19168
rect 4120 19156 4126 19168
rect 4223 19156 4251 19196
rect 5077 19193 5089 19196
rect 5123 19193 5135 19227
rect 5077 19187 5135 19193
rect 6178 19184 6184 19236
rect 6236 19224 6242 19236
rect 6236 19196 6868 19224
rect 6236 19184 6242 19196
rect 4120 19128 4251 19156
rect 4120 19116 4126 19128
rect 5166 19116 5172 19168
rect 5224 19156 5230 19168
rect 5767 19159 5825 19165
rect 5767 19156 5779 19159
rect 5224 19128 5779 19156
rect 5224 19116 5230 19128
rect 5767 19125 5779 19128
rect 5813 19125 5825 19159
rect 5767 19119 5825 19125
rect 6454 19116 6460 19168
rect 6512 19156 6518 19168
rect 6641 19159 6699 19165
rect 6641 19156 6653 19159
rect 6512 19128 6653 19156
rect 6512 19116 6518 19128
rect 6641 19125 6653 19128
rect 6687 19125 6699 19159
rect 6840 19156 6868 19196
rect 7098 19184 7104 19236
rect 7156 19224 7162 19236
rect 10842 19224 10870 19255
rect 11698 19252 11704 19304
rect 11756 19292 11762 19304
rect 12656 19295 12714 19301
rect 12656 19292 12668 19295
rect 11756 19264 12668 19292
rect 11756 19252 11762 19264
rect 12656 19261 12668 19264
rect 12702 19292 12714 19295
rect 13081 19295 13139 19301
rect 13081 19292 13093 19295
rect 12702 19264 13093 19292
rect 12702 19261 12714 19264
rect 12656 19255 12714 19261
rect 13081 19261 13093 19264
rect 13127 19261 13139 19295
rect 13081 19255 13139 19261
rect 13262 19252 13268 19304
rect 13320 19292 13326 19304
rect 13668 19295 13726 19301
rect 13668 19292 13680 19295
rect 13320 19264 13680 19292
rect 13320 19252 13326 19264
rect 13668 19261 13680 19264
rect 13714 19292 13726 19295
rect 14093 19295 14151 19301
rect 14093 19292 14105 19295
rect 13714 19264 14105 19292
rect 13714 19261 13726 19264
rect 13668 19255 13726 19261
rect 14093 19261 14105 19264
rect 14139 19261 14151 19295
rect 14093 19255 14151 19261
rect 11238 19224 11244 19236
rect 7156 19196 11244 19224
rect 7156 19184 7162 19196
rect 11238 19184 11244 19196
rect 11296 19184 11302 19236
rect 7009 19159 7067 19165
rect 7009 19156 7021 19159
rect 6840 19128 7021 19156
rect 6641 19119 6699 19125
rect 7009 19125 7021 19128
rect 7055 19125 7067 19159
rect 7009 19119 7067 19125
rect 8573 19159 8631 19165
rect 8573 19125 8585 19159
rect 8619 19156 8631 19159
rect 8938 19156 8944 19168
rect 8619 19128 8944 19156
rect 8619 19125 8631 19128
rect 8573 19119 8631 19125
rect 8938 19116 8944 19128
rect 8996 19116 9002 19168
rect 9490 19116 9496 19168
rect 9548 19156 9554 19168
rect 12759 19159 12817 19165
rect 12759 19156 12771 19159
rect 9548 19128 12771 19156
rect 9548 19116 9554 19128
rect 12759 19125 12771 19128
rect 12805 19125 12817 19159
rect 12759 19119 12817 19125
rect 1104 19066 20884 19088
rect 1104 19014 8315 19066
rect 8367 19014 8379 19066
rect 8431 19014 8443 19066
rect 8495 19014 8507 19066
rect 8559 19014 15648 19066
rect 15700 19014 15712 19066
rect 15764 19014 15776 19066
rect 15828 19014 15840 19066
rect 15892 19014 20884 19066
rect 1104 18992 20884 19014
rect 5810 18912 5816 18964
rect 5868 18952 5874 18964
rect 10827 18955 10885 18961
rect 10827 18952 10839 18955
rect 5868 18924 10839 18952
rect 5868 18912 5874 18924
rect 10827 18921 10839 18924
rect 10873 18921 10885 18955
rect 10827 18915 10885 18921
rect 11238 18912 11244 18964
rect 11296 18952 11302 18964
rect 19058 18952 19064 18964
rect 11296 18924 19064 18952
rect 11296 18912 11302 18924
rect 19058 18912 19064 18924
rect 19116 18912 19122 18964
rect 5350 18844 5356 18896
rect 5408 18884 5414 18896
rect 5408 18856 7512 18884
rect 5408 18844 5414 18856
rect 2314 18776 2320 18828
rect 2372 18816 2378 18828
rect 2501 18819 2559 18825
rect 2501 18816 2513 18819
rect 2372 18788 2513 18816
rect 2372 18776 2378 18788
rect 2501 18785 2513 18788
rect 2547 18785 2559 18819
rect 2501 18779 2559 18785
rect 4065 18819 4123 18825
rect 4065 18785 4077 18819
rect 4111 18785 4123 18819
rect 4338 18816 4344 18828
rect 4299 18788 4344 18816
rect 4065 18779 4123 18785
rect 1394 18748 1400 18760
rect 1355 18720 1400 18748
rect 1394 18708 1400 18720
rect 1452 18708 1458 18760
rect 3142 18748 3148 18760
rect 3103 18720 3148 18748
rect 3142 18708 3148 18720
rect 3200 18708 3206 18760
rect 4080 18748 4108 18779
rect 4338 18776 4344 18788
rect 4396 18776 4402 18828
rect 5626 18816 5632 18828
rect 4448 18788 5632 18816
rect 4448 18748 4476 18788
rect 5626 18776 5632 18788
rect 5684 18776 5690 18828
rect 5920 18825 5948 18856
rect 7484 18828 7512 18856
rect 5905 18819 5963 18825
rect 5905 18785 5917 18819
rect 5951 18785 5963 18819
rect 5905 18779 5963 18785
rect 6638 18776 6644 18828
rect 6696 18816 6702 18828
rect 7193 18819 7251 18825
rect 7193 18816 7205 18819
rect 6696 18788 7205 18816
rect 6696 18776 6702 18788
rect 7193 18785 7205 18788
rect 7239 18785 7251 18819
rect 7466 18816 7472 18828
rect 7427 18788 7472 18816
rect 7193 18779 7251 18785
rect 7466 18776 7472 18788
rect 7524 18776 7530 18828
rect 10756 18819 10814 18825
rect 10756 18785 10768 18819
rect 10802 18816 10814 18819
rect 11146 18816 11152 18828
rect 10802 18788 11152 18816
rect 10802 18785 10814 18788
rect 10756 18779 10814 18785
rect 11146 18776 11152 18788
rect 11204 18776 11210 18828
rect 11514 18776 11520 18828
rect 11572 18816 11578 18828
rect 11736 18819 11794 18825
rect 11736 18816 11748 18819
rect 11572 18788 11748 18816
rect 11572 18776 11578 18788
rect 11736 18785 11748 18788
rect 11782 18785 11794 18819
rect 11736 18779 11794 18785
rect 12713 18819 12771 18825
rect 12713 18785 12725 18819
rect 12759 18816 12771 18819
rect 12802 18816 12808 18828
rect 12759 18788 12808 18816
rect 12759 18785 12771 18788
rect 12713 18779 12771 18785
rect 12802 18776 12808 18788
rect 12860 18776 12866 18828
rect 13722 18816 13728 18828
rect 13683 18788 13728 18816
rect 13722 18776 13728 18788
rect 13780 18776 13786 18828
rect 4080 18720 4476 18748
rect 4801 18751 4859 18757
rect 4801 18717 4813 18751
rect 4847 18748 4859 18751
rect 5074 18748 5080 18760
rect 4847 18720 5080 18748
rect 4847 18717 4859 18720
rect 4801 18711 4859 18717
rect 5074 18708 5080 18720
rect 5132 18708 5138 18760
rect 5442 18708 5448 18760
rect 5500 18748 5506 18760
rect 5721 18751 5779 18757
rect 5721 18748 5733 18751
rect 5500 18720 5733 18748
rect 5500 18708 5506 18720
rect 5721 18717 5733 18720
rect 5767 18748 5779 18751
rect 5994 18748 6000 18760
rect 5767 18720 6000 18748
rect 5767 18717 5779 18720
rect 5721 18711 5779 18717
rect 5994 18708 6000 18720
rect 6052 18708 6058 18760
rect 6270 18748 6276 18760
rect 6231 18720 6276 18748
rect 6270 18708 6276 18720
rect 6328 18708 6334 18760
rect 6822 18708 6828 18760
rect 6880 18748 6886 18760
rect 7653 18751 7711 18757
rect 7653 18748 7665 18751
rect 6880 18720 7665 18748
rect 6880 18708 6886 18720
rect 7653 18717 7665 18720
rect 7699 18717 7711 18751
rect 7653 18711 7711 18717
rect 9398 18708 9404 18760
rect 9456 18748 9462 18760
rect 9677 18751 9735 18757
rect 9677 18748 9689 18751
rect 9456 18720 9689 18748
rect 9456 18708 9462 18720
rect 9677 18717 9689 18720
rect 9723 18717 9735 18751
rect 9677 18711 9735 18717
rect 4157 18683 4215 18689
rect 4157 18649 4169 18683
rect 4203 18680 4215 18683
rect 4246 18680 4252 18692
rect 4203 18652 4252 18680
rect 4203 18649 4215 18652
rect 4157 18643 4215 18649
rect 4246 18640 4252 18652
rect 4304 18640 4310 18692
rect 6012 18680 6040 18708
rect 7285 18683 7343 18689
rect 7285 18680 7297 18683
rect 6012 18652 7297 18680
rect 7285 18649 7297 18652
rect 7331 18680 7343 18683
rect 7374 18680 7380 18692
rect 7331 18652 7380 18680
rect 7331 18649 7343 18652
rect 7285 18643 7343 18649
rect 7374 18640 7380 18652
rect 7432 18640 7438 18692
rect 10594 18640 10600 18692
rect 10652 18680 10658 18692
rect 11839 18683 11897 18689
rect 11839 18680 11851 18683
rect 10652 18652 11851 18680
rect 10652 18640 10658 18652
rect 11839 18649 11851 18652
rect 11885 18649 11897 18683
rect 13863 18683 13921 18689
rect 13863 18680 13875 18683
rect 11839 18643 11897 18649
rect 11992 18652 13875 18680
rect 1854 18612 1860 18624
rect 1815 18584 1860 18612
rect 1854 18572 1860 18584
rect 1912 18572 1918 18624
rect 7009 18615 7067 18621
rect 7009 18581 7021 18615
rect 7055 18612 7067 18615
rect 7190 18612 7196 18624
rect 7055 18584 7196 18612
rect 7055 18581 7067 18584
rect 7009 18575 7067 18581
rect 7190 18572 7196 18584
rect 7248 18572 7254 18624
rect 8202 18612 8208 18624
rect 8163 18584 8208 18612
rect 8202 18572 8208 18584
rect 8260 18572 8266 18624
rect 9122 18572 9128 18624
rect 9180 18612 9186 18624
rect 11992 18612 12020 18652
rect 13863 18649 13875 18652
rect 13909 18649 13921 18683
rect 13863 18643 13921 18649
rect 9180 18584 12020 18612
rect 9180 18572 9186 18584
rect 12618 18572 12624 18624
rect 12676 18612 12682 18624
rect 12851 18615 12909 18621
rect 12851 18612 12863 18615
rect 12676 18584 12863 18612
rect 12676 18572 12682 18584
rect 12851 18581 12863 18584
rect 12897 18581 12909 18615
rect 12851 18575 12909 18581
rect 1104 18522 20884 18544
rect 1104 18470 4648 18522
rect 4700 18470 4712 18522
rect 4764 18470 4776 18522
rect 4828 18470 4840 18522
rect 4892 18470 11982 18522
rect 12034 18470 12046 18522
rect 12098 18470 12110 18522
rect 12162 18470 12174 18522
rect 12226 18470 19315 18522
rect 19367 18470 19379 18522
rect 19431 18470 19443 18522
rect 19495 18470 19507 18522
rect 19559 18470 20884 18522
rect 1104 18448 20884 18470
rect 1578 18408 1584 18420
rect 1539 18380 1584 18408
rect 1578 18368 1584 18380
rect 1636 18368 1642 18420
rect 3142 18368 3148 18420
rect 3200 18408 3206 18420
rect 5350 18408 5356 18420
rect 3200 18380 5356 18408
rect 3200 18368 3206 18380
rect 5350 18368 5356 18380
rect 5408 18368 5414 18420
rect 5626 18408 5632 18420
rect 5587 18380 5632 18408
rect 5626 18368 5632 18380
rect 5684 18368 5690 18420
rect 5994 18408 6000 18420
rect 5955 18380 6000 18408
rect 5994 18368 6000 18380
rect 6052 18368 6058 18420
rect 6638 18408 6644 18420
rect 6599 18380 6644 18408
rect 6638 18368 6644 18380
rect 6696 18368 6702 18420
rect 7374 18408 7380 18420
rect 7335 18380 7380 18408
rect 7374 18368 7380 18380
rect 7432 18368 7438 18420
rect 7466 18368 7472 18420
rect 7524 18408 7530 18420
rect 8941 18411 8999 18417
rect 8941 18408 8953 18411
rect 7524 18380 8953 18408
rect 7524 18368 7530 18380
rect 8941 18377 8953 18380
rect 8987 18377 8999 18411
rect 8941 18371 8999 18377
rect 18693 18411 18751 18417
rect 18693 18377 18705 18411
rect 18739 18408 18751 18411
rect 19702 18408 19708 18420
rect 18739 18380 19708 18408
rect 18739 18377 18751 18380
rect 18693 18371 18751 18377
rect 19702 18368 19708 18380
rect 19760 18368 19766 18420
rect 2038 18300 2044 18352
rect 2096 18340 2102 18352
rect 2682 18340 2688 18352
rect 2096 18312 2688 18340
rect 2096 18300 2102 18312
rect 2682 18300 2688 18312
rect 2740 18340 2746 18352
rect 3697 18343 3755 18349
rect 3697 18340 3709 18343
rect 2740 18312 3709 18340
rect 2740 18300 2746 18312
rect 3697 18309 3709 18312
rect 3743 18340 3755 18343
rect 3973 18343 4031 18349
rect 3973 18340 3985 18343
rect 3743 18312 3985 18340
rect 3743 18309 3755 18312
rect 3697 18303 3755 18309
rect 3973 18309 3985 18312
rect 4019 18340 4031 18343
rect 4065 18343 4123 18349
rect 4065 18340 4077 18343
rect 4019 18312 4077 18340
rect 4019 18309 4031 18312
rect 3973 18303 4031 18309
rect 4065 18309 4077 18312
rect 4111 18309 4123 18343
rect 4706 18340 4712 18352
rect 4619 18312 4712 18340
rect 4065 18303 4123 18309
rect 4706 18300 4712 18312
rect 4764 18340 4770 18352
rect 6656 18340 6684 18368
rect 4764 18312 6684 18340
rect 4764 18300 4770 18312
rect 7558 18300 7564 18352
rect 7616 18340 7622 18352
rect 8021 18343 8079 18349
rect 8021 18340 8033 18343
rect 7616 18312 8033 18340
rect 7616 18300 7622 18312
rect 8021 18309 8033 18312
rect 8067 18309 8079 18343
rect 8021 18303 8079 18309
rect 106 18232 112 18284
rect 164 18272 170 18284
rect 10091 18275 10149 18281
rect 10091 18272 10103 18275
rect 164 18244 10103 18272
rect 164 18232 170 18244
rect 10091 18241 10103 18244
rect 10137 18241 10149 18275
rect 10091 18235 10149 18241
rect 10781 18275 10839 18281
rect 10781 18241 10793 18275
rect 10827 18272 10839 18275
rect 11146 18272 11152 18284
rect 10827 18244 11152 18272
rect 10827 18241 10839 18244
rect 10781 18235 10839 18241
rect 11146 18232 11152 18244
rect 11204 18232 11210 18284
rect 13078 18232 13084 18284
rect 13136 18272 13142 18284
rect 13722 18272 13728 18284
rect 13136 18244 13728 18272
rect 13136 18232 13142 18244
rect 1397 18207 1455 18213
rect 1397 18173 1409 18207
rect 1443 18204 1455 18207
rect 1486 18204 1492 18216
rect 1443 18176 1492 18204
rect 1443 18173 1455 18176
rect 1397 18167 1455 18173
rect 1486 18164 1492 18176
rect 1544 18164 1550 18216
rect 2133 18207 2191 18213
rect 2133 18173 2145 18207
rect 2179 18204 2191 18207
rect 2866 18204 2872 18216
rect 2179 18176 2872 18204
rect 2179 18173 2191 18176
rect 2133 18167 2191 18173
rect 2866 18164 2872 18176
rect 2924 18164 2930 18216
rect 3602 18164 3608 18216
rect 3660 18204 3666 18216
rect 4062 18204 4068 18216
rect 3660 18176 4068 18204
rect 3660 18164 3666 18176
rect 4062 18164 4068 18176
rect 4120 18204 4126 18216
rect 4706 18204 4712 18216
rect 4120 18176 4712 18204
rect 4120 18164 4126 18176
rect 4706 18164 4712 18176
rect 4764 18164 4770 18216
rect 4893 18207 4951 18213
rect 4893 18173 4905 18207
rect 4939 18204 4951 18207
rect 5626 18204 5632 18216
rect 4939 18176 5632 18204
rect 4939 18173 4951 18176
rect 4893 18167 4951 18173
rect 3421 18139 3479 18145
rect 3421 18105 3433 18139
rect 3467 18136 3479 18139
rect 4246 18136 4252 18148
rect 3467 18108 4252 18136
rect 3467 18105 3479 18108
rect 3421 18099 3479 18105
rect 4246 18096 4252 18108
rect 4304 18096 4310 18148
rect 4908 18136 4936 18167
rect 5626 18164 5632 18176
rect 5684 18164 5690 18216
rect 7837 18207 7895 18213
rect 7837 18173 7849 18207
rect 7883 18204 7895 18207
rect 7926 18204 7932 18216
rect 7883 18176 7932 18204
rect 7883 18173 7895 18176
rect 7837 18167 7895 18173
rect 7926 18164 7932 18176
rect 7984 18164 7990 18216
rect 8202 18204 8208 18216
rect 8163 18176 8208 18204
rect 8202 18164 8208 18176
rect 8260 18164 8266 18216
rect 9861 18207 9919 18213
rect 9861 18173 9873 18207
rect 9907 18204 9919 18207
rect 10004 18207 10062 18213
rect 10004 18204 10016 18207
rect 9907 18176 10016 18204
rect 9907 18173 9919 18176
rect 9861 18167 9919 18173
rect 10004 18173 10016 18176
rect 10050 18204 10062 18207
rect 10502 18204 10508 18216
rect 10050 18176 10508 18204
rect 10050 18173 10062 18176
rect 10004 18167 10062 18173
rect 10502 18164 10508 18176
rect 10560 18164 10566 18216
rect 10686 18164 10692 18216
rect 10744 18204 10750 18216
rect 13515 18213 13543 18244
rect 13722 18232 13728 18244
rect 13780 18272 13786 18284
rect 14829 18275 14887 18281
rect 14829 18272 14841 18275
rect 13780 18244 14044 18272
rect 13780 18232 13786 18244
rect 11000 18207 11058 18213
rect 11000 18204 11012 18207
rect 10744 18176 11012 18204
rect 10744 18164 10750 18176
rect 11000 18173 11012 18176
rect 11046 18173 11058 18207
rect 11000 18167 11058 18173
rect 12504 18207 12562 18213
rect 12504 18173 12516 18207
rect 12550 18204 12562 18207
rect 13265 18207 13323 18213
rect 13265 18204 13277 18207
rect 12550 18176 13277 18204
rect 12550 18173 12562 18176
rect 12504 18167 12562 18173
rect 13265 18173 13277 18176
rect 13311 18173 13323 18207
rect 13500 18207 13558 18213
rect 13500 18204 13512 18207
rect 13478 18176 13512 18204
rect 13265 18167 13323 18173
rect 13500 18173 13512 18176
rect 13546 18173 13558 18207
rect 13500 18167 13558 18173
rect 4448 18108 4936 18136
rect 8665 18139 8723 18145
rect 2314 18028 2320 18080
rect 2372 18068 2378 18080
rect 2409 18071 2467 18077
rect 2409 18068 2421 18071
rect 2372 18040 2421 18068
rect 2372 18028 2378 18040
rect 2409 18037 2421 18040
rect 2455 18037 2467 18071
rect 2409 18031 2467 18037
rect 3973 18071 4031 18077
rect 3973 18037 3985 18071
rect 4019 18068 4031 18071
rect 4448 18068 4476 18108
rect 8665 18105 8677 18139
rect 8711 18136 8723 18139
rect 9674 18136 9680 18148
rect 8711 18108 9680 18136
rect 8711 18105 8723 18108
rect 8665 18099 8723 18105
rect 9674 18096 9680 18108
rect 9732 18096 9738 18148
rect 12802 18136 12808 18148
rect 10289 18108 12808 18136
rect 6914 18068 6920 18080
rect 4019 18040 4476 18068
rect 6875 18040 6920 18068
rect 4019 18037 4031 18040
rect 3973 18031 4031 18037
rect 6914 18028 6920 18040
rect 6972 18028 6978 18080
rect 9858 18028 9864 18080
rect 9916 18068 9922 18080
rect 10289 18068 10317 18108
rect 12802 18096 12808 18108
rect 12860 18136 12866 18148
rect 12897 18139 12955 18145
rect 12897 18136 12909 18139
rect 12860 18108 12909 18136
rect 12860 18096 12866 18108
rect 12897 18105 12909 18108
rect 12943 18105 12955 18139
rect 13280 18136 13308 18167
rect 13722 18136 13728 18148
rect 13280 18108 13728 18136
rect 12897 18099 12955 18105
rect 13722 18096 13728 18108
rect 13780 18096 13786 18148
rect 14016 18145 14044 18244
rect 14614 18244 14841 18272
rect 14614 18216 14642 18244
rect 14829 18241 14841 18244
rect 14875 18241 14887 18275
rect 14829 18235 14887 18241
rect 14550 18213 14556 18216
rect 14528 18207 14556 18213
rect 14528 18173 14540 18207
rect 14608 18204 14642 18216
rect 14608 18176 14701 18204
rect 14528 18167 14556 18173
rect 14550 18164 14556 18167
rect 14608 18164 14614 18176
rect 14734 18164 14740 18216
rect 14792 18204 14798 18216
rect 15508 18207 15566 18213
rect 15508 18204 15520 18207
rect 14792 18176 15520 18204
rect 14792 18164 14798 18176
rect 15508 18173 15520 18176
rect 15554 18204 15566 18207
rect 15933 18207 15991 18213
rect 15933 18204 15945 18207
rect 15554 18176 15945 18204
rect 15554 18173 15566 18176
rect 15508 18167 15566 18173
rect 15933 18173 15945 18176
rect 15979 18173 15991 18207
rect 15933 18167 15991 18173
rect 18414 18164 18420 18216
rect 18472 18204 18478 18216
rect 18509 18207 18567 18213
rect 18509 18204 18521 18207
rect 18472 18176 18521 18204
rect 18472 18164 18478 18176
rect 18509 18173 18521 18176
rect 18555 18204 18567 18207
rect 19061 18207 19119 18213
rect 19061 18204 19073 18207
rect 18555 18176 19073 18204
rect 18555 18173 18567 18176
rect 18509 18167 18567 18173
rect 19061 18173 19073 18176
rect 19107 18173 19119 18207
rect 19061 18167 19119 18173
rect 14001 18139 14059 18145
rect 14001 18105 14013 18139
rect 14047 18136 14059 18139
rect 14277 18139 14335 18145
rect 14277 18136 14289 18139
rect 14047 18108 14289 18136
rect 14047 18105 14059 18108
rect 14001 18099 14059 18105
rect 14277 18105 14289 18108
rect 14323 18105 14335 18139
rect 14277 18099 14335 18105
rect 14366 18096 14372 18148
rect 14424 18136 14430 18148
rect 15611 18139 15669 18145
rect 15611 18136 15623 18139
rect 14424 18108 15623 18136
rect 14424 18096 14430 18108
rect 15611 18105 15623 18108
rect 15657 18105 15669 18139
rect 15611 18099 15669 18105
rect 9916 18040 10317 18068
rect 9916 18028 9922 18040
rect 10870 18028 10876 18080
rect 10928 18068 10934 18080
rect 11103 18071 11161 18077
rect 11103 18068 11115 18071
rect 10928 18040 11115 18068
rect 10928 18028 10934 18040
rect 11103 18037 11115 18040
rect 11149 18037 11161 18071
rect 11103 18031 11161 18037
rect 11514 18028 11520 18080
rect 11572 18068 11578 18080
rect 11701 18071 11759 18077
rect 11701 18068 11713 18071
rect 11572 18040 11713 18068
rect 11572 18028 11578 18040
rect 11701 18037 11713 18040
rect 11747 18037 11759 18071
rect 11701 18031 11759 18037
rect 12434 18028 12440 18080
rect 12492 18068 12498 18080
rect 12575 18071 12633 18077
rect 12575 18068 12587 18071
rect 12492 18040 12587 18068
rect 12492 18028 12498 18040
rect 12575 18037 12587 18040
rect 12621 18037 12633 18071
rect 12575 18031 12633 18037
rect 12710 18028 12716 18080
rect 12768 18068 12774 18080
rect 13587 18071 13645 18077
rect 13587 18068 13599 18071
rect 12768 18040 13599 18068
rect 12768 18028 12774 18040
rect 13587 18037 13599 18040
rect 13633 18037 13645 18071
rect 13587 18031 13645 18037
rect 14182 18028 14188 18080
rect 14240 18068 14246 18080
rect 14599 18071 14657 18077
rect 14599 18068 14611 18071
rect 14240 18040 14611 18068
rect 14240 18028 14246 18040
rect 14599 18037 14611 18040
rect 14645 18037 14657 18071
rect 14599 18031 14657 18037
rect 14829 18071 14887 18077
rect 14829 18037 14841 18071
rect 14875 18068 14887 18071
rect 15013 18071 15071 18077
rect 15013 18068 15025 18071
rect 14875 18040 15025 18068
rect 14875 18037 14887 18040
rect 14829 18031 14887 18037
rect 15013 18037 15025 18040
rect 15059 18068 15071 18071
rect 16758 18068 16764 18080
rect 15059 18040 16764 18068
rect 15059 18037 15071 18040
rect 15013 18031 15071 18037
rect 16758 18028 16764 18040
rect 16816 18028 16822 18080
rect 1104 17978 20884 18000
rect 1104 17926 8315 17978
rect 8367 17926 8379 17978
rect 8431 17926 8443 17978
rect 8495 17926 8507 17978
rect 8559 17926 15648 17978
rect 15700 17926 15712 17978
rect 15764 17926 15776 17978
rect 15828 17926 15840 17978
rect 15892 17926 20884 17978
rect 1104 17904 20884 17926
rect 4338 17824 4344 17876
rect 4396 17864 4402 17876
rect 4525 17867 4583 17873
rect 4525 17864 4537 17867
rect 4396 17836 4537 17864
rect 4396 17824 4402 17836
rect 4525 17833 4537 17836
rect 4571 17833 4583 17867
rect 4525 17827 4583 17833
rect 5994 17824 6000 17876
rect 6052 17864 6058 17876
rect 12526 17864 12532 17876
rect 6052 17836 12532 17864
rect 6052 17824 6058 17836
rect 12526 17824 12532 17836
rect 12584 17824 12590 17876
rect 1302 17756 1308 17808
rect 1360 17796 1366 17808
rect 1535 17799 1593 17805
rect 1535 17796 1547 17799
rect 1360 17768 1547 17796
rect 1360 17756 1366 17768
rect 1535 17765 1547 17768
rect 1581 17765 1593 17799
rect 1535 17759 1593 17765
rect 2317 17799 2375 17805
rect 2317 17765 2329 17799
rect 2363 17796 2375 17799
rect 4246 17796 4252 17808
rect 2363 17768 4252 17796
rect 2363 17765 2375 17768
rect 2317 17759 2375 17765
rect 1448 17731 1506 17737
rect 1448 17697 1460 17731
rect 1494 17728 1506 17731
rect 1854 17728 1860 17740
rect 1494 17700 1860 17728
rect 1494 17697 1506 17700
rect 1448 17691 1506 17697
rect 1854 17688 1860 17700
rect 1912 17688 1918 17740
rect 2406 17728 2412 17740
rect 2367 17700 2412 17728
rect 2406 17688 2412 17700
rect 2464 17688 2470 17740
rect 2516 17737 2544 17768
rect 4246 17756 4252 17768
rect 4304 17796 4310 17808
rect 4893 17799 4951 17805
rect 4893 17796 4905 17799
rect 4304 17768 4905 17796
rect 4304 17756 4310 17768
rect 4893 17765 4905 17768
rect 4939 17765 4951 17799
rect 4893 17759 4951 17765
rect 8297 17799 8355 17805
rect 8297 17765 8309 17799
rect 8343 17796 8355 17799
rect 10410 17796 10416 17808
rect 8343 17768 10416 17796
rect 8343 17765 8355 17768
rect 8297 17759 8355 17765
rect 10410 17756 10416 17768
rect 10468 17756 10474 17808
rect 2501 17731 2559 17737
rect 2501 17697 2513 17731
rect 2547 17697 2559 17731
rect 2501 17691 2559 17697
rect 2685 17731 2743 17737
rect 2685 17697 2697 17731
rect 2731 17697 2743 17731
rect 2685 17691 2743 17697
rect 2314 17620 2320 17672
rect 2372 17660 2378 17672
rect 2700 17660 2728 17691
rect 3970 17688 3976 17740
rect 4028 17728 4034 17740
rect 4100 17731 4158 17737
rect 4100 17728 4112 17731
rect 4028 17700 4112 17728
rect 4028 17688 4034 17700
rect 4100 17697 4112 17700
rect 4146 17697 4158 17731
rect 4100 17691 4158 17697
rect 4982 17688 4988 17740
rect 5040 17728 5046 17740
rect 5353 17731 5411 17737
rect 5353 17728 5365 17731
rect 5040 17700 5365 17728
rect 5040 17688 5046 17700
rect 5353 17697 5365 17700
rect 5399 17728 5411 17731
rect 5626 17728 5632 17740
rect 5399 17700 5632 17728
rect 5399 17697 5411 17700
rect 5353 17691 5411 17697
rect 5626 17688 5632 17700
rect 5684 17688 5690 17740
rect 5902 17728 5908 17740
rect 5863 17700 5908 17728
rect 5902 17688 5908 17700
rect 5960 17688 5966 17740
rect 7561 17731 7619 17737
rect 7561 17697 7573 17731
rect 7607 17728 7619 17731
rect 7650 17728 7656 17740
rect 7607 17700 7656 17728
rect 7607 17697 7619 17700
rect 7561 17691 7619 17697
rect 7650 17688 7656 17700
rect 7708 17688 7714 17740
rect 7837 17731 7895 17737
rect 7837 17697 7849 17731
rect 7883 17728 7895 17731
rect 8202 17728 8208 17740
rect 7883 17700 8208 17728
rect 7883 17697 7895 17700
rect 7837 17691 7895 17697
rect 8202 17688 8208 17700
rect 8260 17688 8266 17740
rect 9306 17688 9312 17740
rect 9364 17728 9370 17740
rect 9677 17731 9735 17737
rect 9677 17728 9689 17731
rect 9364 17700 9689 17728
rect 9364 17688 9370 17700
rect 9677 17697 9689 17700
rect 9723 17697 9735 17731
rect 10134 17728 10140 17740
rect 10095 17700 10140 17728
rect 9677 17691 9735 17697
rect 10134 17688 10140 17700
rect 10192 17688 10198 17740
rect 11308 17731 11366 17737
rect 11308 17697 11320 17731
rect 11354 17728 11366 17731
rect 11514 17728 11520 17740
rect 11354 17700 11520 17728
rect 11354 17697 11366 17700
rect 11308 17691 11366 17697
rect 11514 17688 11520 17700
rect 11572 17688 11578 17740
rect 12897 17731 12955 17737
rect 12897 17697 12909 17731
rect 12943 17728 12955 17731
rect 12986 17728 12992 17740
rect 12943 17700 12992 17728
rect 12943 17697 12955 17700
rect 12897 17691 12955 17697
rect 12986 17688 12992 17700
rect 13044 17688 13050 17740
rect 13976 17731 14034 17737
rect 13976 17697 13988 17731
rect 14022 17728 14034 17731
rect 14090 17728 14096 17740
rect 14022 17700 14096 17728
rect 14022 17697 14034 17700
rect 13976 17691 14034 17697
rect 14090 17688 14096 17700
rect 14148 17688 14154 17740
rect 15356 17731 15414 17737
rect 15356 17697 15368 17731
rect 15402 17728 15414 17731
rect 15470 17728 15476 17740
rect 15402 17700 15476 17728
rect 15402 17697 15414 17700
rect 15356 17691 15414 17697
rect 15470 17688 15476 17700
rect 15528 17688 15534 17740
rect 16368 17731 16426 17737
rect 16368 17697 16380 17731
rect 16414 17728 16426 17731
rect 17218 17728 17224 17740
rect 16414 17700 17224 17728
rect 16414 17697 16426 17700
rect 16368 17691 16426 17697
rect 17218 17688 17224 17700
rect 17276 17688 17282 17740
rect 2372 17632 2728 17660
rect 3145 17663 3203 17669
rect 2372 17620 2378 17632
rect 3145 17629 3157 17663
rect 3191 17660 3203 17663
rect 4430 17660 4436 17672
rect 3191 17632 4436 17660
rect 3191 17629 3203 17632
rect 3145 17623 3203 17629
rect 4430 17620 4436 17632
rect 4488 17620 4494 17672
rect 6181 17663 6239 17669
rect 6181 17629 6193 17663
rect 6227 17660 6239 17663
rect 6730 17660 6736 17672
rect 6227 17632 6736 17660
rect 6227 17629 6239 17632
rect 6181 17623 6239 17629
rect 6730 17620 6736 17632
rect 6788 17620 6794 17672
rect 10042 17620 10048 17672
rect 10100 17660 10106 17672
rect 10229 17663 10287 17669
rect 10229 17660 10241 17663
rect 10100 17632 10241 17660
rect 10100 17620 10106 17632
rect 10229 17629 10241 17632
rect 10275 17629 10287 17663
rect 10229 17623 10287 17629
rect 1486 17552 1492 17604
rect 1544 17592 1550 17604
rect 1949 17595 2007 17601
rect 1949 17592 1961 17595
rect 1544 17564 1961 17592
rect 1544 17552 1550 17564
rect 1949 17561 1961 17564
rect 1995 17592 2007 17595
rect 4062 17592 4068 17604
rect 1995 17564 4068 17592
rect 1995 17561 2007 17564
rect 1949 17555 2007 17561
rect 4062 17552 4068 17564
rect 4120 17592 4126 17604
rect 7098 17592 7104 17604
rect 4120 17564 7104 17592
rect 4120 17552 4126 17564
rect 7098 17552 7104 17564
rect 7156 17552 7162 17604
rect 7558 17552 7564 17604
rect 7616 17592 7622 17604
rect 7653 17595 7711 17601
rect 7653 17592 7665 17595
rect 7616 17564 7665 17592
rect 7616 17552 7622 17564
rect 7653 17561 7665 17564
rect 7699 17592 7711 17595
rect 8573 17595 8631 17601
rect 8573 17592 8585 17595
rect 7699 17564 8585 17592
rect 7699 17561 7711 17564
rect 7653 17555 7711 17561
rect 8573 17561 8585 17564
rect 8619 17561 8631 17595
rect 8573 17555 8631 17561
rect 9030 17552 9036 17604
rect 9088 17592 9094 17604
rect 14047 17595 14105 17601
rect 14047 17592 14059 17595
rect 9088 17564 14059 17592
rect 9088 17552 9094 17564
rect 14047 17561 14059 17564
rect 14093 17561 14105 17595
rect 14047 17555 14105 17561
rect 3878 17484 3884 17536
rect 3936 17524 3942 17536
rect 4203 17527 4261 17533
rect 4203 17524 4215 17527
rect 3936 17496 4215 17524
rect 3936 17484 3942 17496
rect 4203 17493 4215 17496
rect 4249 17493 4261 17527
rect 7190 17524 7196 17536
rect 7151 17496 7196 17524
rect 4203 17487 4261 17493
rect 7190 17484 7196 17496
rect 7248 17484 7254 17536
rect 10686 17484 10692 17536
rect 10744 17524 10750 17536
rect 10965 17527 11023 17533
rect 10965 17524 10977 17527
rect 10744 17496 10977 17524
rect 10744 17484 10750 17496
rect 10965 17493 10977 17496
rect 11011 17493 11023 17527
rect 10965 17487 11023 17493
rect 11054 17484 11060 17536
rect 11112 17524 11118 17536
rect 11379 17527 11437 17533
rect 11379 17524 11391 17527
rect 11112 17496 11391 17524
rect 11112 17484 11118 17496
rect 11379 17493 11391 17496
rect 11425 17493 11437 17527
rect 11379 17487 11437 17493
rect 13035 17527 13093 17533
rect 13035 17493 13047 17527
rect 13081 17524 13093 17527
rect 13814 17524 13820 17536
rect 13081 17496 13820 17524
rect 13081 17493 13093 17496
rect 13035 17487 13093 17493
rect 13814 17484 13820 17496
rect 13872 17484 13878 17536
rect 14182 17484 14188 17536
rect 14240 17524 14246 17536
rect 15427 17527 15485 17533
rect 15427 17524 15439 17527
rect 14240 17496 15439 17524
rect 14240 17484 14246 17496
rect 15427 17493 15439 17496
rect 15473 17493 15485 17527
rect 15427 17487 15485 17493
rect 16114 17484 16120 17536
rect 16172 17524 16178 17536
rect 16439 17527 16497 17533
rect 16439 17524 16451 17527
rect 16172 17496 16451 17524
rect 16172 17484 16178 17496
rect 16439 17493 16451 17496
rect 16485 17493 16497 17527
rect 16439 17487 16497 17493
rect 1104 17434 20884 17456
rect 1104 17382 4648 17434
rect 4700 17382 4712 17434
rect 4764 17382 4776 17434
rect 4828 17382 4840 17434
rect 4892 17382 11982 17434
rect 12034 17382 12046 17434
rect 12098 17382 12110 17434
rect 12162 17382 12174 17434
rect 12226 17382 19315 17434
rect 19367 17382 19379 17434
rect 19431 17382 19443 17434
rect 19495 17382 19507 17434
rect 19559 17382 20884 17434
rect 1104 17360 20884 17382
rect 1578 17320 1584 17332
rect 1539 17292 1584 17320
rect 1578 17280 1584 17292
rect 1636 17280 1642 17332
rect 6362 17280 6368 17332
rect 6420 17320 6426 17332
rect 12710 17320 12716 17332
rect 6420 17292 12716 17320
rect 6420 17280 6426 17292
rect 12710 17280 12716 17292
rect 12768 17280 12774 17332
rect 13906 17320 13912 17332
rect 13464 17292 13912 17320
rect 5626 17252 5632 17264
rect 4816 17224 5632 17252
rect 2041 17187 2099 17193
rect 2041 17153 2053 17187
rect 2087 17184 2099 17187
rect 3970 17184 3976 17196
rect 2087 17156 3976 17184
rect 2087 17153 2099 17156
rect 2041 17147 2099 17153
rect 1397 17119 1455 17125
rect 1397 17085 1409 17119
rect 1443 17116 1455 17119
rect 2056 17116 2084 17147
rect 3970 17144 3976 17156
rect 4028 17144 4034 17196
rect 2774 17116 2780 17128
rect 1443 17088 2084 17116
rect 2735 17088 2780 17116
rect 1443 17085 1455 17088
rect 1397 17079 1455 17085
rect 2774 17076 2780 17088
rect 2832 17076 2838 17128
rect 4816 17125 4844 17224
rect 5626 17212 5632 17224
rect 5684 17212 5690 17264
rect 6822 17212 6828 17264
rect 6880 17252 6886 17264
rect 6880 17224 10133 17252
rect 6880 17212 6886 17224
rect 5074 17184 5080 17196
rect 5035 17156 5080 17184
rect 5074 17144 5080 17156
rect 5132 17144 5138 17196
rect 9766 17184 9772 17196
rect 5460 17156 7236 17184
rect 3053 17119 3111 17125
rect 3053 17085 3065 17119
rect 3099 17116 3111 17119
rect 4801 17119 4859 17125
rect 3099 17088 4154 17116
rect 3099 17085 3111 17088
rect 3053 17079 3111 17085
rect 3234 17048 3240 17060
rect 3195 17020 3240 17048
rect 3234 17008 3240 17020
rect 3292 17008 3298 17060
rect 3344 16992 3372 17088
rect 4126 17048 4154 17088
rect 4801 17085 4813 17119
rect 4847 17085 4859 17119
rect 4801 17079 4859 17085
rect 4985 17119 5043 17125
rect 4985 17085 4997 17119
rect 5031 17116 5043 17119
rect 5258 17116 5264 17128
rect 5031 17088 5264 17116
rect 5031 17085 5043 17088
rect 4985 17079 5043 17085
rect 5258 17076 5264 17088
rect 5316 17116 5322 17128
rect 5460 17116 5488 17156
rect 7208 17128 7236 17156
rect 8956 17156 9772 17184
rect 5316 17088 5488 17116
rect 5316 17076 5322 17088
rect 5718 17076 5724 17128
rect 5776 17116 5782 17128
rect 6181 17119 6239 17125
rect 6181 17116 6193 17119
rect 5776 17088 6193 17116
rect 5776 17076 5782 17088
rect 6181 17085 6193 17088
rect 6227 17116 6239 17119
rect 6822 17116 6828 17128
rect 6227 17088 6828 17116
rect 6227 17085 6239 17088
rect 6181 17079 6239 17085
rect 6822 17076 6828 17088
rect 6880 17116 6886 17128
rect 7101 17119 7159 17125
rect 7101 17116 7113 17119
rect 6880 17088 7113 17116
rect 6880 17076 6886 17088
rect 7101 17085 7113 17088
rect 7147 17085 7159 17119
rect 7101 17079 7159 17085
rect 7190 17076 7196 17128
rect 7248 17116 7254 17128
rect 8956 17125 8984 17156
rect 9766 17144 9772 17156
rect 9824 17144 9830 17196
rect 10105 17184 10133 17224
rect 10686 17212 10692 17264
rect 10744 17252 10750 17264
rect 13265 17255 13323 17261
rect 13265 17252 13277 17255
rect 10744 17224 13277 17252
rect 10744 17212 10750 17224
rect 13265 17221 13277 17224
rect 13311 17221 13323 17255
rect 13265 17215 13323 17221
rect 10226 17184 10232 17196
rect 10105 17156 10232 17184
rect 10226 17144 10232 17156
rect 10284 17184 10290 17196
rect 10284 17156 10548 17184
rect 10284 17144 10290 17156
rect 7561 17119 7619 17125
rect 7561 17116 7573 17119
rect 7248 17088 7573 17116
rect 7248 17076 7254 17088
rect 7561 17085 7573 17088
rect 7607 17085 7619 17119
rect 7561 17079 7619 17085
rect 8941 17119 8999 17125
rect 8941 17085 8953 17119
rect 8987 17085 8999 17119
rect 9401 17119 9459 17125
rect 9401 17116 9413 17119
rect 8941 17079 8999 17085
rect 9048 17088 9413 17116
rect 5537 17051 5595 17057
rect 5537 17048 5549 17051
rect 4126 17020 5549 17048
rect 5537 17017 5549 17020
rect 5583 17048 5595 17051
rect 5902 17048 5908 17060
rect 5583 17020 5908 17048
rect 5583 17017 5595 17020
rect 5537 17011 5595 17017
rect 5902 17008 5908 17020
rect 5960 17008 5966 17060
rect 6641 17051 6699 17057
rect 6641 17017 6653 17051
rect 6687 17048 6699 17051
rect 7650 17048 7656 17060
rect 6687 17020 7656 17048
rect 6687 17017 6699 17020
rect 6641 17011 6699 17017
rect 7650 17008 7656 17020
rect 7708 17008 7714 17060
rect 8202 17048 8208 17060
rect 8115 17020 8208 17048
rect 8202 17008 8208 17020
rect 8260 17048 8266 17060
rect 8846 17048 8852 17060
rect 8260 17020 8852 17048
rect 8260 17008 8266 17020
rect 8846 17008 8852 17020
rect 8904 17008 8910 17060
rect 2314 16980 2320 16992
rect 2275 16952 2320 16980
rect 2314 16940 2320 16952
rect 2372 16940 2378 16992
rect 3326 16940 3332 16992
rect 3384 16980 3390 16992
rect 3513 16983 3571 16989
rect 3513 16980 3525 16983
rect 3384 16952 3525 16980
rect 3384 16940 3390 16952
rect 3513 16949 3525 16952
rect 3559 16949 3571 16983
rect 3513 16943 3571 16949
rect 3970 16940 3976 16992
rect 4028 16980 4034 16992
rect 4157 16983 4215 16989
rect 4157 16980 4169 16983
rect 4028 16952 4169 16980
rect 4028 16940 4034 16952
rect 4157 16949 4169 16952
rect 4203 16980 4215 16983
rect 6086 16980 6092 16992
rect 4203 16952 6092 16980
rect 4203 16949 4215 16952
rect 4157 16943 4215 16949
rect 6086 16940 6092 16952
rect 6144 16940 6150 16992
rect 7374 16980 7380 16992
rect 7335 16952 7380 16980
rect 7374 16940 7380 16952
rect 7432 16940 7438 16992
rect 8754 16980 8760 16992
rect 8715 16952 8760 16980
rect 8754 16940 8760 16952
rect 8812 16980 8818 16992
rect 9048 16980 9076 17088
rect 9401 17085 9413 17088
rect 9447 17116 9459 17119
rect 9953 17119 10011 17125
rect 9953 17116 9965 17119
rect 9447 17088 9965 17116
rect 9447 17085 9459 17088
rect 9401 17079 9459 17085
rect 9953 17085 9965 17088
rect 9999 17116 10011 17119
rect 10134 17116 10140 17128
rect 9999 17088 10140 17116
rect 9999 17085 10011 17088
rect 9953 17079 10011 17085
rect 10134 17076 10140 17088
rect 10192 17076 10198 17128
rect 10520 17125 10548 17156
rect 11330 17144 11336 17196
rect 11388 17184 11394 17196
rect 12986 17184 12992 17196
rect 11388 17156 12992 17184
rect 11388 17144 11394 17156
rect 12986 17144 12992 17156
rect 13044 17184 13050 17196
rect 13464 17193 13492 17292
rect 13906 17280 13912 17292
rect 13964 17280 13970 17332
rect 14001 17323 14059 17329
rect 14001 17289 14013 17323
rect 14047 17320 14059 17323
rect 14090 17320 14096 17332
rect 14047 17292 14096 17320
rect 14047 17289 14059 17292
rect 14001 17283 14059 17289
rect 14090 17280 14096 17292
rect 14148 17280 14154 17332
rect 17218 17320 17224 17332
rect 17179 17292 17224 17320
rect 17218 17280 17224 17292
rect 17276 17320 17282 17332
rect 18782 17320 18788 17332
rect 17276 17292 18788 17320
rect 17276 17280 17282 17292
rect 18782 17280 18788 17292
rect 18840 17280 18846 17332
rect 15470 17212 15476 17264
rect 15528 17252 15534 17264
rect 15841 17255 15899 17261
rect 15841 17252 15853 17255
rect 15528 17224 15853 17252
rect 15528 17212 15534 17224
rect 15841 17221 15853 17224
rect 15887 17221 15899 17255
rect 15841 17215 15899 17221
rect 13449 17187 13507 17193
rect 13449 17184 13461 17187
rect 13044 17156 13461 17184
rect 13044 17144 13050 17156
rect 13449 17153 13461 17156
rect 13495 17153 13507 17187
rect 13449 17147 13507 17153
rect 13630 17144 13636 17196
rect 13688 17184 13694 17196
rect 16531 17187 16589 17193
rect 16531 17184 16543 17187
rect 13688 17156 16543 17184
rect 13688 17144 13694 17156
rect 16531 17153 16543 17156
rect 16577 17153 16589 17187
rect 16531 17147 16589 17153
rect 10505 17119 10563 17125
rect 10505 17085 10517 17119
rect 10551 17085 10563 17119
rect 10505 17079 10563 17085
rect 10965 17119 11023 17125
rect 10965 17085 10977 17119
rect 11011 17085 11023 17119
rect 10965 17079 11023 17085
rect 10410 17048 10416 17060
rect 10371 17020 10416 17048
rect 10410 17008 10416 17020
rect 10468 17048 10474 17060
rect 10980 17048 11008 17079
rect 12250 17076 12256 17128
rect 12308 17116 12314 17128
rect 12437 17119 12495 17125
rect 12437 17116 12449 17119
rect 12308 17088 12449 17116
rect 12308 17076 12314 17088
rect 12437 17085 12449 17088
rect 12483 17085 12495 17119
rect 12437 17079 12495 17085
rect 12897 17119 12955 17125
rect 12897 17085 12909 17119
rect 12943 17085 12955 17119
rect 12897 17079 12955 17085
rect 13265 17119 13323 17125
rect 13265 17085 13277 17119
rect 13311 17116 13323 17119
rect 15416 17119 15474 17125
rect 15416 17116 15428 17119
rect 13311 17088 15428 17116
rect 13311 17085 13323 17088
rect 13265 17079 13323 17085
rect 15416 17085 15428 17088
rect 15462 17116 15474 17119
rect 16209 17119 16267 17125
rect 16209 17116 16221 17119
rect 15462 17088 16221 17116
rect 15462 17085 15474 17088
rect 15416 17079 15474 17085
rect 16209 17085 16221 17088
rect 16255 17085 16267 17119
rect 16209 17079 16267 17085
rect 16439 17119 16497 17125
rect 16439 17085 16451 17119
rect 16485 17085 16497 17119
rect 16439 17079 16497 17085
rect 12912 17048 12940 17079
rect 14090 17048 14096 17060
rect 10468 17020 11008 17048
rect 12360 17020 12940 17048
rect 12979 17020 14096 17048
rect 10468 17008 10474 17020
rect 12360 16992 12388 17020
rect 9214 16980 9220 16992
rect 8812 16952 9076 16980
rect 9175 16952 9220 16980
rect 8812 16940 8818 16952
rect 9214 16940 9220 16952
rect 9272 16940 9278 16992
rect 10778 16980 10784 16992
rect 10739 16952 10784 16980
rect 10778 16940 10784 16952
rect 10836 16940 10842 16992
rect 11514 16980 11520 16992
rect 11475 16952 11520 16980
rect 11514 16940 11520 16952
rect 11572 16940 11578 16992
rect 12253 16983 12311 16989
rect 12253 16949 12265 16983
rect 12299 16980 12311 16983
rect 12342 16980 12348 16992
rect 12299 16952 12348 16980
rect 12299 16949 12311 16952
rect 12253 16943 12311 16949
rect 12342 16940 12348 16952
rect 12400 16940 12406 16992
rect 12526 16980 12532 16992
rect 12487 16952 12532 16980
rect 12526 16940 12532 16952
rect 12584 16940 12590 16992
rect 12802 16940 12808 16992
rect 12860 16980 12866 16992
rect 12979 16980 13007 17020
rect 14090 17008 14096 17020
rect 14148 17008 14154 17060
rect 15519 17051 15577 17057
rect 15519 17048 15531 17051
rect 14292 17020 15531 17048
rect 12860 16952 13007 16980
rect 12860 16940 12866 16952
rect 13998 16940 14004 16992
rect 14056 16980 14062 16992
rect 14292 16980 14320 17020
rect 15519 17017 15531 17020
rect 15565 17017 15577 17051
rect 15519 17011 15577 17017
rect 16022 17008 16028 17060
rect 16080 17048 16086 17060
rect 16454 17048 16482 17079
rect 16853 17051 16911 17057
rect 16853 17048 16865 17051
rect 16080 17020 16865 17048
rect 16080 17008 16086 17020
rect 16853 17017 16865 17020
rect 16899 17048 16911 17051
rect 18322 17048 18328 17060
rect 16899 17020 18328 17048
rect 16899 17017 16911 17020
rect 16853 17011 16911 17017
rect 18322 17008 18328 17020
rect 18380 17008 18386 17060
rect 14056 16952 14320 16980
rect 14369 16983 14427 16989
rect 14056 16940 14062 16952
rect 14369 16949 14381 16983
rect 14415 16980 14427 16983
rect 15378 16980 15384 16992
rect 14415 16952 15384 16980
rect 14415 16949 14427 16952
rect 14369 16943 14427 16949
rect 15378 16940 15384 16952
rect 15436 16940 15442 16992
rect 1104 16890 20884 16912
rect 1104 16838 8315 16890
rect 8367 16838 8379 16890
rect 8431 16838 8443 16890
rect 8495 16838 8507 16890
rect 8559 16838 15648 16890
rect 15700 16838 15712 16890
rect 15764 16838 15776 16890
rect 15828 16838 15840 16890
rect 15892 16838 20884 16890
rect 1104 16816 20884 16838
rect 1854 16736 1860 16788
rect 1912 16776 1918 16788
rect 1912 16748 2820 16776
rect 1912 16736 1918 16748
rect 2222 16708 2228 16720
rect 2183 16680 2228 16708
rect 2222 16668 2228 16680
rect 2280 16668 2286 16720
rect 2792 16717 2820 16748
rect 6546 16736 6552 16788
rect 6604 16776 6610 16788
rect 7558 16776 7564 16788
rect 6604 16748 7564 16776
rect 6604 16736 6610 16748
rect 7558 16736 7564 16748
rect 7616 16776 7622 16788
rect 8205 16779 8263 16785
rect 8205 16776 8217 16779
rect 7616 16748 8217 16776
rect 7616 16736 7622 16748
rect 8205 16745 8217 16748
rect 8251 16745 8263 16779
rect 8205 16739 8263 16745
rect 9306 16736 9312 16788
rect 9364 16776 9370 16788
rect 9401 16779 9459 16785
rect 9401 16776 9413 16779
rect 9364 16748 9413 16776
rect 9364 16736 9370 16748
rect 9401 16745 9413 16748
rect 9447 16776 9459 16779
rect 9582 16776 9588 16788
rect 9447 16748 9588 16776
rect 9447 16745 9459 16748
rect 9401 16739 9459 16745
rect 9582 16736 9588 16748
rect 9640 16736 9646 16788
rect 10226 16736 10232 16788
rect 10284 16776 10290 16788
rect 10689 16779 10747 16785
rect 10689 16776 10701 16779
rect 10284 16748 10701 16776
rect 10284 16736 10290 16748
rect 10689 16745 10701 16748
rect 10735 16745 10747 16779
rect 10689 16739 10747 16745
rect 11379 16779 11437 16785
rect 11379 16745 11391 16779
rect 11425 16776 11437 16779
rect 16206 16776 16212 16788
rect 11425 16748 16212 16776
rect 11425 16745 11437 16748
rect 11379 16739 11437 16745
rect 2777 16711 2835 16717
rect 2777 16677 2789 16711
rect 2823 16677 2835 16711
rect 2777 16671 2835 16677
rect 6914 16668 6920 16720
rect 6972 16708 6978 16720
rect 7285 16711 7343 16717
rect 7285 16708 7297 16711
rect 6972 16680 7297 16708
rect 6972 16668 6978 16680
rect 7285 16677 7297 16680
rect 7331 16677 7343 16711
rect 7285 16671 7343 16677
rect 7377 16711 7435 16717
rect 7377 16677 7389 16711
rect 7423 16708 7435 16711
rect 7742 16708 7748 16720
rect 7423 16680 7748 16708
rect 7423 16677 7435 16680
rect 7377 16671 7435 16677
rect 7742 16668 7748 16680
rect 7800 16668 7806 16720
rect 10704 16708 10732 16739
rect 16206 16736 16212 16748
rect 16264 16736 16270 16788
rect 12250 16708 12256 16720
rect 10704 16680 12256 16708
rect 12250 16668 12256 16680
rect 12308 16708 12314 16720
rect 12437 16711 12495 16717
rect 12437 16708 12449 16711
rect 12308 16680 12449 16708
rect 12308 16668 12314 16680
rect 12437 16677 12449 16680
rect 12483 16708 12495 16711
rect 12483 16680 13308 16708
rect 12483 16677 12495 16680
rect 12437 16671 12495 16677
rect 4982 16640 4988 16652
rect 4943 16612 4988 16640
rect 4982 16600 4988 16612
rect 5040 16600 5046 16652
rect 5258 16640 5264 16652
rect 5219 16612 5264 16640
rect 5258 16600 5264 16612
rect 5316 16600 5322 16652
rect 5626 16600 5632 16652
rect 5684 16640 5690 16652
rect 5813 16643 5871 16649
rect 5813 16640 5825 16643
rect 5684 16612 5825 16640
rect 5684 16600 5690 16612
rect 5813 16609 5825 16612
rect 5859 16640 5871 16643
rect 7009 16643 7067 16649
rect 7009 16640 7021 16643
rect 5859 16612 7021 16640
rect 5859 16609 5871 16612
rect 5813 16603 5871 16609
rect 7009 16609 7021 16612
rect 7055 16609 7067 16643
rect 7009 16603 7067 16609
rect 7929 16643 7987 16649
rect 7929 16609 7941 16643
rect 7975 16640 7987 16643
rect 8018 16640 8024 16652
rect 7975 16612 8024 16640
rect 7975 16609 7987 16612
rect 7929 16603 7987 16609
rect 8018 16600 8024 16612
rect 8076 16600 8082 16652
rect 8110 16600 8116 16652
rect 8168 16640 8174 16652
rect 9677 16643 9735 16649
rect 9677 16640 9689 16643
rect 8168 16612 9689 16640
rect 8168 16600 8174 16612
rect 9677 16609 9689 16612
rect 9723 16640 9735 16643
rect 9950 16640 9956 16652
rect 9723 16612 9956 16640
rect 9723 16609 9735 16612
rect 9677 16603 9735 16609
rect 9950 16600 9956 16612
rect 10008 16600 10014 16652
rect 10134 16640 10140 16652
rect 10095 16612 10140 16640
rect 10134 16600 10140 16612
rect 10192 16600 10198 16652
rect 11308 16643 11366 16649
rect 11308 16609 11320 16643
rect 11354 16640 11366 16643
rect 11422 16640 11428 16652
rect 11354 16612 11428 16640
rect 11354 16609 11366 16612
rect 11308 16603 11366 16609
rect 11422 16600 11428 16612
rect 11480 16600 11486 16652
rect 12710 16640 12716 16652
rect 12671 16612 12716 16640
rect 12710 16600 12716 16612
rect 12768 16600 12774 16652
rect 13170 16640 13176 16652
rect 13131 16612 13176 16640
rect 13170 16600 13176 16612
rect 13228 16600 13234 16652
rect 13280 16640 13308 16680
rect 13354 16668 13360 16720
rect 13412 16708 13418 16720
rect 17451 16711 17509 16717
rect 17451 16708 17463 16711
rect 13412 16680 17463 16708
rect 13412 16668 13418 16680
rect 17451 16677 17463 16680
rect 17497 16677 17509 16711
rect 17451 16671 17509 16677
rect 15356 16643 15414 16649
rect 13280 16612 13814 16640
rect 2133 16575 2191 16581
rect 2133 16541 2145 16575
rect 2179 16572 2191 16575
rect 3050 16572 3056 16584
rect 2179 16544 3056 16572
rect 2179 16541 2191 16544
rect 2133 16535 2191 16541
rect 3050 16532 3056 16544
rect 3108 16572 3114 16584
rect 3421 16575 3479 16581
rect 3421 16572 3433 16575
rect 3108 16544 3433 16572
rect 3108 16532 3114 16544
rect 3421 16541 3433 16544
rect 3467 16541 3479 16575
rect 3421 16535 3479 16541
rect 4617 16575 4675 16581
rect 4617 16541 4629 16575
rect 4663 16572 4675 16575
rect 5276 16572 5304 16600
rect 5442 16572 5448 16584
rect 4663 16544 5304 16572
rect 5403 16544 5448 16572
rect 4663 16541 4675 16544
rect 4617 16535 4675 16541
rect 5442 16532 5448 16544
rect 5500 16532 5506 16584
rect 6822 16572 6828 16584
rect 6783 16544 6828 16572
rect 6822 16532 6828 16544
rect 6880 16532 6886 16584
rect 10226 16572 10232 16584
rect 10187 16544 10232 16572
rect 10226 16532 10232 16544
rect 10284 16532 10290 16584
rect 13449 16575 13507 16581
rect 13449 16541 13461 16575
rect 13495 16572 13507 16575
rect 13538 16572 13544 16584
rect 13495 16544 13544 16572
rect 13495 16541 13507 16544
rect 13449 16535 13507 16541
rect 13538 16532 13544 16544
rect 13596 16532 13602 16584
rect 13786 16572 13814 16612
rect 15356 16609 15368 16643
rect 15402 16640 15414 16643
rect 15470 16640 15476 16652
rect 15402 16612 15476 16640
rect 15402 16609 15414 16612
rect 15356 16603 15414 16609
rect 15470 16600 15476 16612
rect 15528 16600 15534 16652
rect 16298 16640 16304 16652
rect 16259 16612 16304 16640
rect 16298 16600 16304 16612
rect 16356 16600 16362 16652
rect 17310 16640 17316 16652
rect 17271 16612 17316 16640
rect 17310 16600 17316 16612
rect 17368 16600 17374 16652
rect 18392 16643 18450 16649
rect 18392 16609 18404 16643
rect 18438 16640 18450 16643
rect 18506 16640 18512 16652
rect 18438 16612 18512 16640
rect 18438 16609 18450 16612
rect 18392 16603 18450 16609
rect 18506 16600 18512 16612
rect 18564 16600 18570 16652
rect 18230 16572 18236 16584
rect 13786 16544 18236 16572
rect 18230 16532 18236 16544
rect 18288 16532 18294 16584
rect 1949 16507 2007 16513
rect 1949 16473 1961 16507
rect 1995 16504 2007 16507
rect 2774 16504 2780 16516
rect 1995 16476 2780 16504
rect 1995 16473 2007 16476
rect 1949 16467 2007 16473
rect 2774 16464 2780 16476
rect 2832 16504 2838 16516
rect 3142 16504 3148 16516
rect 2832 16476 3148 16504
rect 2832 16464 2838 16476
rect 3142 16464 3148 16476
rect 3200 16464 3206 16516
rect 6086 16464 6092 16516
rect 6144 16504 6150 16516
rect 16022 16504 16028 16516
rect 6144 16476 16028 16504
rect 6144 16464 6150 16476
rect 16022 16464 16028 16476
rect 16080 16464 16086 16516
rect 2406 16396 2412 16448
rect 2464 16436 2470 16448
rect 3053 16439 3111 16445
rect 3053 16436 3065 16439
rect 2464 16408 3065 16436
rect 2464 16396 2470 16408
rect 3053 16405 3065 16408
rect 3099 16436 3111 16439
rect 3602 16436 3608 16448
rect 3099 16408 3608 16436
rect 3099 16405 3111 16408
rect 3053 16399 3111 16405
rect 3602 16396 3608 16408
rect 3660 16396 3666 16448
rect 7009 16439 7067 16445
rect 7009 16405 7021 16439
rect 7055 16436 7067 16439
rect 9033 16439 9091 16445
rect 9033 16436 9045 16439
rect 7055 16408 9045 16436
rect 7055 16405 7067 16408
rect 7009 16399 7067 16405
rect 9033 16405 9045 16408
rect 9079 16436 9091 16439
rect 9766 16436 9772 16448
rect 9079 16408 9772 16436
rect 9079 16405 9091 16408
rect 9033 16399 9091 16405
rect 9766 16396 9772 16408
rect 9824 16396 9830 16448
rect 14274 16436 14280 16448
rect 14235 16408 14280 16436
rect 14274 16396 14280 16408
rect 14332 16396 14338 16448
rect 15102 16396 15108 16448
rect 15160 16436 15166 16448
rect 15427 16439 15485 16445
rect 15427 16436 15439 16439
rect 15160 16408 15439 16436
rect 15160 16396 15166 16408
rect 15427 16405 15439 16408
rect 15473 16405 15485 16439
rect 15427 16399 15485 16405
rect 15930 16396 15936 16448
rect 15988 16436 15994 16448
rect 16439 16439 16497 16445
rect 16439 16436 16451 16439
rect 15988 16408 16451 16436
rect 15988 16396 15994 16408
rect 16439 16405 16451 16408
rect 16485 16405 16497 16439
rect 16439 16399 16497 16405
rect 17126 16396 17132 16448
rect 17184 16436 17190 16448
rect 18463 16439 18521 16445
rect 18463 16436 18475 16439
rect 17184 16408 18475 16436
rect 17184 16396 17190 16408
rect 18463 16405 18475 16408
rect 18509 16405 18521 16439
rect 18463 16399 18521 16405
rect 1104 16346 20884 16368
rect 1104 16294 4648 16346
rect 4700 16294 4712 16346
rect 4764 16294 4776 16346
rect 4828 16294 4840 16346
rect 4892 16294 11982 16346
rect 12034 16294 12046 16346
rect 12098 16294 12110 16346
rect 12162 16294 12174 16346
rect 12226 16294 19315 16346
rect 19367 16294 19379 16346
rect 19431 16294 19443 16346
rect 19495 16294 19507 16346
rect 19559 16294 20884 16346
rect 1104 16272 20884 16294
rect 4801 16235 4859 16241
rect 4801 16201 4813 16235
rect 4847 16232 4859 16235
rect 5258 16232 5264 16244
rect 4847 16204 5264 16232
rect 4847 16201 4859 16204
rect 4801 16195 4859 16201
rect 5258 16192 5264 16204
rect 5316 16192 5322 16244
rect 6914 16192 6920 16244
rect 6972 16232 6978 16244
rect 8021 16235 8079 16241
rect 8021 16232 8033 16235
rect 6972 16204 8033 16232
rect 6972 16192 6978 16204
rect 8021 16201 8033 16204
rect 8067 16201 8079 16235
rect 8021 16195 8079 16201
rect 9950 16192 9956 16244
rect 10008 16232 10014 16244
rect 11149 16235 11207 16241
rect 11149 16232 11161 16235
rect 10008 16204 11161 16232
rect 10008 16192 10014 16204
rect 11149 16201 11161 16204
rect 11195 16232 11207 16235
rect 12710 16232 12716 16244
rect 11195 16204 12716 16232
rect 11195 16201 11207 16204
rect 11149 16195 11207 16201
rect 12710 16192 12716 16204
rect 12768 16192 12774 16244
rect 13906 16192 13912 16244
rect 13964 16232 13970 16244
rect 16298 16232 16304 16244
rect 13964 16204 16304 16232
rect 13964 16192 13970 16204
rect 16298 16192 16304 16204
rect 16356 16192 16362 16244
rect 17402 16232 17408 16244
rect 16960 16204 17408 16232
rect 2777 16167 2835 16173
rect 2777 16164 2789 16167
rect 1688 16136 2789 16164
rect 1394 15920 1400 15972
rect 1452 15960 1458 15972
rect 1688 15960 1716 16136
rect 2777 16133 2789 16136
rect 2823 16133 2835 16167
rect 2777 16127 2835 16133
rect 9674 16124 9680 16176
rect 9732 16164 9738 16176
rect 13630 16164 13636 16176
rect 9732 16136 13636 16164
rect 9732 16124 9738 16136
rect 13630 16124 13636 16136
rect 13688 16124 13694 16176
rect 14090 16164 14096 16176
rect 14051 16136 14096 16164
rect 14090 16124 14096 16136
rect 14148 16164 14154 16176
rect 16960 16164 16988 16204
rect 17402 16192 17408 16204
rect 17460 16192 17466 16244
rect 17954 16192 17960 16244
rect 18012 16232 18018 16244
rect 18877 16235 18935 16241
rect 18877 16232 18889 16235
rect 18012 16204 18889 16232
rect 18012 16192 18018 16204
rect 18877 16201 18889 16204
rect 18923 16201 18935 16235
rect 18877 16195 18935 16201
rect 14148 16136 16988 16164
rect 14148 16124 14154 16136
rect 1854 16056 1860 16108
rect 1912 16096 1918 16108
rect 2133 16099 2191 16105
rect 2133 16096 2145 16099
rect 1912 16068 2145 16096
rect 1912 16056 1918 16068
rect 2133 16065 2145 16068
rect 2179 16065 2191 16099
rect 2133 16059 2191 16065
rect 2222 16056 2228 16108
rect 2280 16096 2286 16108
rect 3145 16099 3203 16105
rect 3145 16096 3157 16099
rect 2280 16068 3157 16096
rect 2280 16056 2286 16068
rect 3145 16065 3157 16068
rect 3191 16096 3203 16099
rect 5905 16099 5963 16105
rect 3191 16068 3464 16096
rect 3191 16065 3203 16068
rect 3145 16059 3203 16065
rect 3436 16037 3464 16068
rect 5905 16065 5917 16099
rect 5951 16096 5963 16099
rect 6822 16096 6828 16108
rect 5951 16068 6828 16096
rect 5951 16065 5963 16068
rect 5905 16059 5963 16065
rect 6822 16056 6828 16068
rect 6880 16056 6886 16108
rect 11885 16099 11943 16105
rect 11885 16096 11897 16099
rect 8864 16068 11897 16096
rect 3421 16031 3479 16037
rect 3421 15997 3433 16031
rect 3467 15997 3479 16031
rect 4430 16028 4436 16040
rect 4343 16000 4436 16028
rect 3421 15991 3479 15997
rect 4430 15988 4436 16000
rect 4488 16028 4494 16040
rect 5169 16031 5227 16037
rect 5169 16028 5181 16031
rect 4488 16000 5181 16028
rect 4488 15988 4494 16000
rect 5169 15997 5181 16000
rect 5215 15997 5227 16031
rect 5169 15991 5227 15997
rect 1857 15963 1915 15969
rect 1857 15960 1869 15963
rect 1452 15932 1869 15960
rect 1452 15920 1458 15932
rect 1857 15929 1869 15932
rect 1903 15929 1915 15963
rect 1857 15923 1915 15929
rect 1949 15963 2007 15969
rect 1949 15929 1961 15963
rect 1995 15929 2007 15963
rect 3329 15963 3387 15969
rect 3329 15960 3341 15963
rect 1949 15923 2007 15929
rect 2608 15932 3341 15960
rect 1673 15895 1731 15901
rect 1673 15861 1685 15895
rect 1719 15892 1731 15895
rect 1964 15892 1992 15923
rect 2608 15892 2636 15932
rect 3329 15929 3341 15932
rect 3375 15929 3387 15963
rect 5184 15960 5212 15991
rect 5258 15988 5264 16040
rect 5316 16028 5322 16040
rect 5629 16031 5687 16037
rect 5629 16028 5641 16031
rect 5316 16000 5641 16028
rect 5316 15988 5322 16000
rect 5629 15997 5641 16000
rect 5675 15997 5687 16031
rect 5629 15991 5687 15997
rect 8202 15988 8208 16040
rect 8260 16028 8266 16040
rect 8864 16037 8892 16068
rect 11885 16065 11897 16068
rect 11931 16096 11943 16099
rect 14642 16096 14648 16108
rect 11931 16068 14648 16096
rect 11931 16065 11943 16068
rect 11885 16059 11943 16065
rect 12912 16037 12940 16068
rect 14642 16056 14648 16068
rect 14700 16056 14706 16108
rect 8849 16031 8907 16037
rect 8849 16028 8861 16031
rect 8260 16000 8861 16028
rect 8260 15988 8266 16000
rect 8849 15997 8861 16000
rect 8895 15997 8907 16031
rect 8849 15991 8907 15997
rect 9033 16031 9091 16037
rect 9033 15997 9045 16031
rect 9079 16028 9091 16031
rect 9677 16031 9735 16037
rect 9677 16028 9689 16031
rect 9079 16000 9689 16028
rect 9079 15997 9091 16000
rect 9033 15991 9091 15997
rect 9677 15997 9689 16000
rect 9723 15997 9735 16031
rect 9677 15991 9735 15997
rect 12897 16031 12955 16037
rect 12897 15997 12909 16031
rect 12943 15997 12955 16031
rect 12897 15991 12955 15997
rect 13081 16031 13139 16037
rect 13081 15997 13093 16031
rect 13127 16028 13139 16031
rect 13170 16028 13176 16040
rect 13127 16000 13176 16028
rect 13127 15997 13139 16000
rect 13081 15991 13139 15997
rect 6454 15960 6460 15972
rect 5184 15932 6460 15960
rect 3329 15923 3387 15929
rect 6454 15920 6460 15932
rect 6512 15960 6518 15972
rect 8220 15960 8248 15988
rect 8754 15960 8760 15972
rect 6512 15932 8248 15960
rect 8404 15932 8760 15960
rect 6512 15920 6518 15932
rect 1719 15864 2636 15892
rect 6641 15895 6699 15901
rect 1719 15861 1731 15864
rect 1673 15855 1731 15861
rect 6641 15861 6653 15895
rect 6687 15892 6699 15895
rect 7098 15892 7104 15904
rect 6687 15864 7104 15892
rect 6687 15861 6699 15864
rect 6641 15855 6699 15861
rect 7098 15852 7104 15864
rect 7156 15892 7162 15904
rect 7193 15895 7251 15901
rect 7193 15892 7205 15895
rect 7156 15864 7205 15892
rect 7156 15852 7162 15864
rect 7193 15861 7205 15864
rect 7239 15861 7251 15895
rect 7742 15892 7748 15904
rect 7703 15864 7748 15892
rect 7193 15855 7251 15861
rect 7742 15852 7748 15864
rect 7800 15852 7806 15904
rect 8110 15852 8116 15904
rect 8168 15892 8174 15904
rect 8404 15901 8432 15932
rect 8754 15920 8760 15932
rect 8812 15960 8818 15972
rect 9048 15960 9076 15991
rect 9306 15960 9312 15972
rect 8812 15932 9076 15960
rect 9267 15932 9312 15960
rect 8812 15920 8818 15932
rect 9306 15920 9312 15932
rect 9364 15920 9370 15972
rect 9950 15920 9956 15972
rect 10008 15960 10014 15972
rect 10229 15963 10287 15969
rect 10229 15960 10241 15963
rect 10008 15932 10241 15960
rect 10008 15920 10014 15932
rect 10229 15929 10241 15932
rect 10275 15929 10287 15963
rect 10229 15923 10287 15929
rect 10318 15920 10324 15972
rect 10376 15960 10382 15972
rect 10376 15932 10421 15960
rect 10376 15920 10382 15932
rect 10502 15920 10508 15972
rect 10560 15960 10566 15972
rect 10873 15963 10931 15969
rect 10873 15960 10885 15963
rect 10560 15932 10885 15960
rect 10560 15920 10566 15932
rect 10873 15929 10885 15932
rect 10919 15960 10931 15963
rect 12158 15960 12164 15972
rect 10919 15932 12164 15960
rect 10919 15929 10931 15932
rect 10873 15923 10931 15929
rect 12158 15920 12164 15932
rect 12216 15920 12222 15972
rect 13096 15960 13124 15991
rect 13170 15988 13176 16000
rect 13228 15988 13234 16040
rect 14274 16028 14280 16040
rect 14235 16000 14280 16028
rect 14274 15988 14280 16000
rect 14332 15988 14338 16040
rect 14752 16037 14780 16136
rect 17034 16124 17040 16176
rect 17092 16164 17098 16176
rect 19199 16167 19257 16173
rect 19199 16164 19211 16167
rect 17092 16136 19211 16164
rect 17092 16124 17098 16136
rect 19199 16133 19211 16136
rect 19245 16133 19257 16167
rect 19199 16127 19257 16133
rect 15381 16099 15439 16105
rect 15381 16065 15393 16099
rect 15427 16096 15439 16099
rect 15470 16096 15476 16108
rect 15427 16068 15476 16096
rect 15427 16065 15439 16068
rect 15381 16059 15439 16065
rect 15470 16056 15476 16068
rect 15528 16096 15534 16108
rect 16298 16096 16304 16108
rect 15528 16068 16304 16096
rect 15528 16056 15534 16068
rect 16298 16056 16304 16068
rect 16356 16056 16362 16108
rect 16574 16056 16580 16108
rect 16632 16096 16638 16108
rect 18187 16099 18245 16105
rect 18187 16096 18199 16099
rect 16632 16068 18199 16096
rect 16632 16056 16638 16068
rect 18187 16065 18199 16068
rect 18233 16065 18245 16099
rect 18187 16059 18245 16065
rect 14737 16031 14795 16037
rect 14737 15997 14749 16031
rect 14783 15997 14795 16031
rect 14737 15991 14795 15997
rect 15908 16031 15966 16037
rect 15908 15997 15920 16031
rect 15954 16028 15966 16031
rect 16022 16028 16028 16040
rect 15954 16000 16028 16028
rect 15954 15997 15966 16000
rect 15908 15991 15966 15997
rect 16022 15988 16028 16000
rect 16080 16028 16086 16040
rect 16669 16031 16727 16037
rect 16669 16028 16681 16031
rect 16080 16000 16681 16028
rect 16080 15988 16086 16000
rect 16669 15997 16681 16000
rect 16715 15997 16727 16031
rect 16669 15991 16727 15997
rect 16904 16031 16962 16037
rect 16904 15997 16916 16031
rect 16950 16028 16962 16031
rect 17954 16028 17960 16040
rect 16950 16000 17816 16028
rect 17915 16000 17960 16028
rect 16950 15997 16962 16000
rect 16904 15991 16962 15997
rect 12360 15932 13124 15960
rect 13357 15963 13415 15969
rect 12360 15904 12388 15932
rect 13357 15929 13369 15963
rect 13403 15960 13415 15963
rect 13446 15960 13452 15972
rect 13403 15932 13452 15960
rect 13403 15929 13415 15932
rect 13357 15923 13415 15929
rect 13446 15920 13452 15932
rect 13504 15960 13510 15972
rect 13633 15963 13691 15969
rect 13633 15960 13645 15963
rect 13504 15932 13645 15960
rect 13504 15920 13510 15932
rect 13633 15929 13645 15932
rect 13679 15929 13691 15963
rect 13633 15923 13691 15929
rect 14918 15920 14924 15972
rect 14976 15960 14982 15972
rect 15013 15963 15071 15969
rect 15013 15960 15025 15963
rect 14976 15932 15025 15960
rect 14976 15920 14982 15932
rect 15013 15929 15025 15932
rect 15059 15929 15071 15963
rect 15013 15923 15071 15929
rect 16206 15920 16212 15972
rect 16264 15960 16270 15972
rect 17788 15969 17816 16000
rect 17954 15988 17960 16000
rect 18012 15988 18018 16040
rect 19150 16037 19156 16040
rect 18325 16031 18383 16037
rect 18325 15997 18337 16031
rect 18371 16028 18383 16031
rect 19128 16031 19156 16037
rect 19128 16028 19140 16031
rect 18371 16000 19140 16028
rect 18371 15997 18383 16000
rect 18325 15991 18383 15997
rect 19128 15997 19140 16000
rect 19208 16028 19214 16040
rect 19521 16031 19579 16037
rect 19521 16028 19533 16031
rect 19208 16000 19533 16028
rect 19128 15991 19156 15997
rect 19150 15988 19156 15991
rect 19208 15988 19214 16000
rect 19521 15997 19533 16000
rect 19567 15997 19579 16031
rect 19521 15991 19579 15997
rect 16991 15963 17049 15969
rect 16991 15960 17003 15963
rect 16264 15932 17003 15960
rect 16264 15920 16270 15932
rect 16991 15929 17003 15932
rect 17037 15929 17049 15963
rect 16991 15923 17049 15929
rect 17773 15963 17831 15969
rect 17773 15929 17785 15963
rect 17819 15960 17831 15963
rect 18966 15960 18972 15972
rect 17819 15932 18972 15960
rect 17819 15929 17831 15932
rect 17773 15923 17831 15929
rect 18966 15920 18972 15932
rect 19024 15920 19030 15972
rect 8389 15895 8447 15901
rect 8389 15892 8401 15895
rect 8168 15864 8401 15892
rect 8168 15852 8174 15864
rect 8389 15861 8401 15864
rect 8435 15861 8447 15895
rect 8389 15855 8447 15861
rect 12253 15895 12311 15901
rect 12253 15861 12265 15895
rect 12299 15892 12311 15895
rect 12342 15892 12348 15904
rect 12299 15864 12348 15892
rect 12299 15861 12311 15864
rect 12253 15855 12311 15861
rect 12342 15852 12348 15864
rect 12400 15852 12406 15904
rect 15979 15895 16037 15901
rect 15979 15861 15991 15895
rect 16025 15892 16037 15895
rect 16390 15892 16396 15904
rect 16025 15864 16396 15892
rect 16025 15861 16037 15864
rect 15979 15855 16037 15861
rect 16390 15852 16396 15864
rect 16448 15852 16454 15904
rect 17310 15852 17316 15904
rect 17368 15892 17374 15904
rect 17405 15895 17463 15901
rect 17405 15892 17417 15895
rect 17368 15864 17417 15892
rect 17368 15852 17374 15864
rect 17405 15861 17417 15864
rect 17451 15892 17463 15895
rect 18325 15895 18383 15901
rect 18325 15892 18337 15895
rect 17451 15864 18337 15892
rect 17451 15861 17463 15864
rect 17405 15855 17463 15861
rect 18325 15861 18337 15864
rect 18371 15861 18383 15895
rect 18506 15892 18512 15904
rect 18467 15864 18512 15892
rect 18325 15855 18383 15861
rect 18506 15852 18512 15864
rect 18564 15852 18570 15904
rect 1104 15802 20884 15824
rect 1104 15750 8315 15802
rect 8367 15750 8379 15802
rect 8431 15750 8443 15802
rect 8495 15750 8507 15802
rect 8559 15750 15648 15802
rect 15700 15750 15712 15802
rect 15764 15750 15776 15802
rect 15828 15750 15840 15802
rect 15892 15750 20884 15802
rect 1104 15728 20884 15750
rect 1670 15648 1676 15700
rect 1728 15688 1734 15700
rect 1765 15691 1823 15697
rect 1765 15688 1777 15691
rect 1728 15660 1777 15688
rect 1728 15648 1734 15660
rect 1765 15657 1777 15660
rect 1811 15657 1823 15691
rect 1765 15651 1823 15657
rect 2222 15648 2228 15700
rect 2280 15688 2286 15700
rect 2317 15691 2375 15697
rect 2317 15688 2329 15691
rect 2280 15660 2329 15688
rect 2280 15648 2286 15660
rect 2317 15657 2329 15660
rect 2363 15688 2375 15691
rect 3329 15691 3387 15697
rect 3329 15688 3341 15691
rect 2363 15660 3341 15688
rect 2363 15657 2375 15660
rect 2317 15651 2375 15657
rect 3329 15657 3341 15660
rect 3375 15657 3387 15691
rect 4246 15688 4252 15700
rect 4207 15660 4252 15688
rect 3329 15651 3387 15657
rect 4246 15648 4252 15660
rect 4304 15648 4310 15700
rect 4801 15691 4859 15697
rect 4801 15657 4813 15691
rect 4847 15688 4859 15691
rect 4982 15688 4988 15700
rect 4847 15660 4988 15688
rect 4847 15657 4859 15660
rect 4801 15651 4859 15657
rect 4982 15648 4988 15660
rect 5040 15648 5046 15700
rect 5258 15688 5264 15700
rect 5219 15660 5264 15688
rect 5258 15648 5264 15660
rect 5316 15648 5322 15700
rect 7193 15691 7251 15697
rect 7193 15657 7205 15691
rect 7239 15688 7251 15691
rect 7742 15688 7748 15700
rect 7239 15660 7748 15688
rect 7239 15657 7251 15660
rect 7193 15651 7251 15657
rect 7742 15648 7748 15660
rect 7800 15648 7806 15700
rect 8202 15648 8208 15700
rect 8260 15688 8266 15700
rect 8573 15691 8631 15697
rect 8573 15688 8585 15691
rect 8260 15660 8585 15688
rect 8260 15648 8266 15660
rect 8573 15657 8585 15660
rect 8619 15657 8631 15691
rect 8573 15651 8631 15657
rect 9493 15691 9551 15697
rect 9493 15657 9505 15691
rect 9539 15688 9551 15691
rect 10318 15688 10324 15700
rect 9539 15660 10324 15688
rect 9539 15657 9551 15660
rect 9493 15651 9551 15657
rect 10318 15648 10324 15660
rect 10376 15688 10382 15700
rect 10597 15691 10655 15697
rect 10597 15688 10609 15691
rect 10376 15660 10609 15688
rect 10376 15648 10382 15660
rect 10597 15657 10609 15660
rect 10643 15657 10655 15691
rect 10597 15651 10655 15657
rect 11333 15691 11391 15697
rect 11333 15657 11345 15691
rect 11379 15688 11391 15691
rect 11422 15688 11428 15700
rect 11379 15660 11428 15688
rect 11379 15657 11391 15660
rect 11333 15651 11391 15657
rect 2590 15620 2596 15632
rect 2551 15592 2596 15620
rect 2590 15580 2596 15592
rect 2648 15580 2654 15632
rect 5899 15623 5957 15629
rect 5899 15589 5911 15623
rect 5945 15620 5957 15623
rect 7098 15620 7104 15632
rect 5945 15592 7104 15620
rect 5945 15589 5957 15592
rect 5899 15583 5957 15589
rect 7098 15580 7104 15592
rect 7156 15580 7162 15632
rect 7466 15620 7472 15632
rect 7427 15592 7472 15620
rect 7466 15580 7472 15592
rect 7524 15580 7530 15632
rect 8018 15620 8024 15632
rect 7979 15592 8024 15620
rect 8018 15580 8024 15592
rect 8076 15580 8082 15632
rect 9766 15580 9772 15632
rect 9824 15620 9830 15632
rect 9998 15623 10056 15629
rect 9998 15620 10010 15623
rect 9824 15592 10010 15620
rect 9824 15580 9830 15592
rect 9998 15589 10010 15592
rect 10044 15589 10056 15623
rect 9998 15583 10056 15589
rect 3970 15512 3976 15564
rect 4028 15552 4034 15564
rect 4065 15555 4123 15561
rect 4065 15552 4077 15555
rect 4028 15524 4077 15552
rect 4028 15512 4034 15524
rect 4065 15521 4077 15524
rect 4111 15521 4123 15555
rect 4065 15515 4123 15521
rect 5442 15512 5448 15564
rect 5500 15552 5506 15564
rect 5537 15555 5595 15561
rect 5537 15552 5549 15555
rect 5500 15524 5549 15552
rect 5500 15512 5506 15524
rect 5537 15521 5549 15524
rect 5583 15521 5595 15555
rect 5537 15515 5595 15521
rect 9306 15512 9312 15564
rect 9364 15552 9370 15564
rect 9677 15555 9735 15561
rect 9677 15552 9689 15555
rect 9364 15524 9689 15552
rect 9364 15512 9370 15524
rect 9677 15521 9689 15524
rect 9723 15521 9735 15555
rect 9677 15515 9735 15521
rect 1397 15487 1455 15493
rect 1397 15453 1409 15487
rect 1443 15484 1455 15487
rect 2866 15484 2872 15496
rect 1443 15456 2872 15484
rect 1443 15453 1455 15456
rect 1397 15447 1455 15453
rect 2866 15444 2872 15456
rect 2924 15484 2930 15496
rect 3418 15484 3424 15496
rect 2924 15456 3424 15484
rect 2924 15444 2930 15456
rect 3418 15444 3424 15456
rect 3476 15444 3482 15496
rect 6825 15487 6883 15493
rect 6825 15453 6837 15487
rect 6871 15484 6883 15487
rect 7377 15487 7435 15493
rect 7377 15484 7389 15487
rect 6871 15456 7389 15484
rect 6871 15453 6883 15456
rect 6825 15447 6883 15453
rect 7377 15453 7389 15456
rect 7423 15484 7435 15487
rect 7558 15484 7564 15496
rect 7423 15456 7564 15484
rect 7423 15453 7435 15456
rect 7377 15447 7435 15453
rect 7558 15444 7564 15456
rect 7616 15444 7622 15496
rect 8018 15444 8024 15496
rect 8076 15484 8082 15496
rect 11348 15484 11376 15651
rect 11422 15648 11428 15660
rect 11480 15648 11486 15700
rect 12710 15648 12716 15700
rect 12768 15688 12774 15700
rect 13081 15691 13139 15697
rect 13081 15688 13093 15691
rect 12768 15660 13093 15688
rect 12768 15648 12774 15660
rect 13081 15657 13093 15660
rect 13127 15688 13139 15691
rect 18046 15688 18052 15700
rect 13127 15660 18052 15688
rect 13127 15657 13139 15660
rect 13081 15651 13139 15657
rect 18046 15648 18052 15660
rect 18104 15648 18110 15700
rect 19245 15691 19303 15697
rect 19245 15657 19257 15691
rect 19291 15688 19303 15691
rect 19610 15688 19616 15700
rect 19291 15660 19616 15688
rect 19291 15657 19303 15660
rect 19245 15651 19303 15657
rect 19610 15648 19616 15660
rect 19668 15648 19674 15700
rect 11606 15620 11612 15632
rect 11567 15592 11612 15620
rect 11606 15580 11612 15592
rect 11664 15580 11670 15632
rect 13262 15580 13268 15632
rect 13320 15620 13326 15632
rect 13770 15623 13828 15629
rect 13770 15620 13782 15623
rect 13320 15592 13782 15620
rect 13320 15580 13326 15592
rect 13770 15589 13782 15592
rect 13816 15589 13828 15623
rect 15470 15620 15476 15632
rect 13770 15583 13828 15589
rect 14384 15592 15476 15620
rect 13446 15552 13452 15564
rect 13407 15524 13452 15552
rect 13446 15512 13452 15524
rect 13504 15512 13510 15564
rect 14384 15561 14412 15592
rect 15470 15580 15476 15592
rect 15528 15580 15534 15632
rect 16022 15620 16028 15632
rect 15983 15592 16028 15620
rect 16022 15580 16028 15592
rect 16080 15580 16086 15632
rect 14369 15555 14427 15561
rect 14369 15521 14381 15555
rect 14415 15521 14427 15555
rect 14369 15515 14427 15521
rect 16920 15555 16978 15561
rect 16920 15521 16932 15555
rect 16966 15552 16978 15555
rect 17310 15552 17316 15564
rect 16966 15524 17316 15552
rect 16966 15521 16978 15524
rect 16920 15515 16978 15521
rect 17310 15512 17316 15524
rect 17368 15512 17374 15564
rect 17770 15512 17776 15564
rect 17828 15552 17834 15564
rect 17900 15555 17958 15561
rect 17900 15552 17912 15555
rect 17828 15524 17912 15552
rect 17828 15512 17834 15524
rect 17900 15521 17912 15524
rect 17946 15521 17958 15555
rect 17900 15515 17958 15521
rect 18598 15512 18604 15564
rect 18656 15552 18662 15564
rect 19061 15555 19119 15561
rect 19061 15552 19073 15555
rect 18656 15524 19073 15552
rect 18656 15512 18662 15524
rect 19061 15521 19073 15524
rect 19107 15521 19119 15555
rect 19061 15515 19119 15521
rect 8076 15456 11376 15484
rect 11517 15487 11575 15493
rect 8076 15444 8082 15456
rect 11517 15453 11529 15487
rect 11563 15484 11575 15487
rect 11790 15484 11796 15496
rect 11563 15456 11796 15484
rect 11563 15453 11575 15456
rect 11517 15447 11575 15453
rect 11790 15444 11796 15456
rect 11848 15444 11854 15496
rect 12158 15484 12164 15496
rect 12071 15456 12164 15484
rect 12158 15444 12164 15456
rect 12216 15484 12222 15496
rect 12986 15484 12992 15496
rect 12216 15456 12992 15484
rect 12216 15444 12222 15456
rect 12986 15444 12992 15456
rect 13044 15444 13050 15496
rect 15378 15484 15384 15496
rect 15339 15456 15384 15484
rect 15378 15444 15384 15456
rect 15436 15444 15442 15496
rect 18003 15487 18061 15493
rect 18003 15484 18015 15487
rect 15539 15456 18015 15484
rect 3786 15376 3792 15428
rect 3844 15416 3850 15428
rect 5258 15416 5264 15428
rect 3844 15388 5264 15416
rect 3844 15376 3850 15388
rect 5258 15376 5264 15388
rect 5316 15376 5322 15428
rect 6086 15376 6092 15428
rect 6144 15416 6150 15428
rect 12618 15416 12624 15428
rect 6144 15388 12624 15416
rect 6144 15376 6150 15388
rect 12618 15376 12624 15388
rect 12676 15376 12682 15428
rect 13630 15376 13636 15428
rect 13688 15416 13694 15428
rect 15539 15416 15567 15456
rect 18003 15453 18015 15456
rect 18049 15453 18061 15487
rect 18003 15447 18061 15453
rect 13688 15388 15567 15416
rect 13688 15376 13694 15388
rect 2958 15348 2964 15360
rect 2919 15320 2964 15348
rect 2958 15308 2964 15320
rect 3016 15308 3022 15360
rect 6454 15348 6460 15360
rect 6415 15320 6460 15348
rect 6454 15308 6460 15320
rect 6512 15308 6518 15360
rect 9950 15308 9956 15360
rect 10008 15348 10014 15360
rect 10873 15351 10931 15357
rect 10873 15348 10885 15351
rect 10008 15320 10885 15348
rect 10008 15308 10014 15320
rect 10873 15317 10885 15320
rect 10919 15317 10931 15351
rect 10873 15311 10931 15317
rect 12342 15308 12348 15360
rect 12400 15348 12406 15360
rect 12713 15351 12771 15357
rect 12713 15348 12725 15351
rect 12400 15320 12725 15348
rect 12400 15308 12406 15320
rect 12713 15317 12725 15320
rect 12759 15317 12771 15351
rect 12713 15311 12771 15317
rect 16482 15308 16488 15360
rect 16540 15348 16546 15360
rect 16991 15351 17049 15357
rect 16991 15348 17003 15351
rect 16540 15320 17003 15348
rect 16540 15308 16546 15320
rect 16991 15317 17003 15320
rect 17037 15317 17049 15351
rect 16991 15311 17049 15317
rect 1104 15258 20884 15280
rect 1104 15206 4648 15258
rect 4700 15206 4712 15258
rect 4764 15206 4776 15258
rect 4828 15206 4840 15258
rect 4892 15206 11982 15258
rect 12034 15206 12046 15258
rect 12098 15206 12110 15258
rect 12162 15206 12174 15258
rect 12226 15206 19315 15258
rect 19367 15206 19379 15258
rect 19431 15206 19443 15258
rect 19495 15206 19507 15258
rect 19559 15206 20884 15258
rect 1104 15184 20884 15206
rect 1949 15147 2007 15153
rect 1949 15113 1961 15147
rect 1995 15144 2007 15147
rect 5902 15144 5908 15156
rect 1995 15116 5908 15144
rect 1995 15113 2007 15116
rect 1949 15107 2007 15113
rect 1964 15076 1992 15107
rect 5902 15104 5908 15116
rect 5960 15104 5966 15156
rect 6454 15104 6460 15156
rect 6512 15144 6518 15156
rect 7193 15147 7251 15153
rect 7193 15144 7205 15147
rect 6512 15116 7205 15144
rect 6512 15104 6518 15116
rect 7193 15113 7205 15116
rect 7239 15144 7251 15147
rect 7466 15144 7472 15156
rect 7239 15116 7472 15144
rect 7239 15113 7251 15116
rect 7193 15107 7251 15113
rect 7466 15104 7472 15116
rect 7524 15104 7530 15156
rect 9033 15147 9091 15153
rect 9033 15113 9045 15147
rect 9079 15144 9091 15147
rect 9306 15144 9312 15156
rect 9079 15116 9312 15144
rect 9079 15113 9091 15116
rect 9033 15107 9091 15113
rect 9306 15104 9312 15116
rect 9364 15104 9370 15156
rect 9766 15144 9772 15156
rect 9727 15116 9772 15144
rect 9766 15104 9772 15116
rect 9824 15104 9830 15156
rect 10965 15147 11023 15153
rect 10965 15113 10977 15147
rect 11011 15144 11023 15147
rect 11517 15147 11575 15153
rect 11517 15144 11529 15147
rect 11011 15116 11529 15144
rect 11011 15113 11023 15116
rect 10965 15107 11023 15113
rect 11517 15113 11529 15116
rect 11563 15144 11575 15147
rect 11606 15144 11612 15156
rect 11563 15116 11612 15144
rect 11563 15113 11575 15116
rect 11517 15107 11575 15113
rect 11606 15104 11612 15116
rect 11664 15104 11670 15156
rect 15197 15147 15255 15153
rect 15197 15113 15209 15147
rect 15243 15144 15255 15147
rect 15378 15144 15384 15156
rect 15243 15116 15384 15144
rect 15243 15113 15255 15116
rect 15197 15107 15255 15113
rect 15378 15104 15384 15116
rect 15436 15104 15442 15156
rect 15470 15104 15476 15156
rect 15528 15144 15534 15156
rect 16301 15147 16359 15153
rect 16301 15144 16313 15147
rect 15528 15116 16313 15144
rect 15528 15104 15534 15116
rect 16301 15113 16313 15116
rect 16347 15113 16359 15147
rect 17310 15144 17316 15156
rect 17271 15116 17316 15144
rect 16301 15107 16359 15113
rect 17310 15104 17316 15116
rect 17368 15104 17374 15156
rect 17770 15144 17776 15156
rect 17731 15116 17776 15144
rect 17770 15104 17776 15116
rect 17828 15104 17834 15156
rect 3050 15076 3056 15088
rect 1479 15048 1992 15076
rect 3011 15048 3056 15076
rect 1479 14949 1507 15048
rect 3050 15036 3056 15048
rect 3108 15036 3114 15088
rect 3418 15076 3424 15088
rect 3379 15048 3424 15076
rect 3418 15036 3424 15048
rect 3476 15036 3482 15088
rect 5077 15079 5135 15085
rect 5077 15045 5089 15079
rect 5123 15076 5135 15079
rect 11146 15076 11152 15088
rect 5123 15048 11152 15076
rect 5123 15045 5135 15048
rect 5077 15039 5135 15045
rect 1535 15011 1593 15017
rect 1535 14977 1547 15011
rect 1581 15008 1593 15011
rect 2501 15011 2559 15017
rect 2501 15008 2513 15011
rect 1581 14980 2513 15008
rect 1581 14977 1593 14980
rect 1535 14971 1593 14977
rect 2501 14977 2513 14980
rect 2547 15008 2559 15011
rect 2958 15008 2964 15020
rect 2547 14980 2964 15008
rect 2547 14977 2559 14980
rect 2501 14971 2559 14977
rect 2958 14968 2964 14980
rect 3016 14968 3022 15020
rect 1448 14943 1507 14949
rect 1448 14909 1460 14943
rect 1494 14912 1507 14943
rect 1494 14909 1506 14912
rect 1448 14903 1506 14909
rect 3510 14900 3516 14952
rect 3568 14940 3574 14952
rect 4224 14943 4282 14949
rect 4224 14940 4236 14943
rect 3568 14912 4236 14940
rect 3568 14900 3574 14912
rect 4224 14909 4236 14912
rect 4270 14940 4282 14943
rect 5092 14940 5120 15039
rect 11146 15036 11152 15048
rect 11204 15036 11210 15088
rect 12618 15036 12624 15088
rect 12676 15076 12682 15088
rect 19199 15079 19257 15085
rect 19199 15076 19211 15079
rect 12676 15048 19211 15076
rect 12676 15036 12682 15048
rect 19199 15045 19211 15048
rect 19245 15045 19257 15079
rect 19199 15039 19257 15045
rect 8018 14968 8024 15020
rect 8076 15008 8082 15020
rect 8113 15011 8171 15017
rect 8113 15008 8125 15011
rect 8076 14980 8125 15008
rect 8076 14968 8082 14980
rect 8113 14977 8125 14980
rect 8159 14977 8171 15011
rect 8113 14971 8171 14977
rect 10045 15011 10103 15017
rect 10045 14977 10057 15011
rect 10091 15008 10103 15011
rect 10226 15008 10232 15020
rect 10091 14980 10232 15008
rect 10091 14977 10103 14980
rect 10045 14971 10103 14977
rect 10226 14968 10232 14980
rect 10284 14968 10290 15020
rect 10410 14968 10416 15020
rect 10468 15008 10474 15020
rect 11238 15008 11244 15020
rect 10468 14980 11244 15008
rect 10468 14968 10474 14980
rect 11238 14968 11244 14980
rect 11296 15008 11302 15020
rect 12897 15011 12955 15017
rect 12897 15008 12909 15011
rect 11296 14980 12909 15008
rect 11296 14968 11302 14980
rect 4270 14912 5120 14940
rect 5905 14943 5963 14949
rect 4270 14909 4282 14912
rect 4224 14903 4282 14909
rect 5905 14909 5917 14943
rect 5951 14940 5963 14943
rect 7558 14940 7564 14952
rect 5951 14912 7564 14940
rect 5951 14909 5963 14912
rect 5905 14903 5963 14909
rect 7558 14900 7564 14912
rect 7616 14900 7622 14952
rect 11698 14940 11704 14952
rect 10105 14912 11704 14940
rect 2590 14872 2596 14884
rect 2551 14844 2596 14872
rect 2590 14832 2596 14844
rect 2648 14832 2654 14884
rect 4617 14875 4675 14881
rect 4617 14872 4629 14875
rect 4126 14844 4629 14872
rect 1670 14764 1676 14816
rect 1728 14804 1734 14816
rect 2317 14807 2375 14813
rect 2317 14804 2329 14807
rect 1728 14776 2329 14804
rect 1728 14764 1734 14776
rect 2317 14773 2329 14776
rect 2363 14804 2375 14807
rect 3694 14804 3700 14816
rect 2363 14776 3700 14804
rect 2363 14773 2375 14776
rect 2317 14767 2375 14773
rect 3694 14764 3700 14776
rect 3752 14764 3758 14816
rect 3970 14764 3976 14816
rect 4028 14804 4034 14816
rect 4126 14804 4154 14844
rect 4617 14841 4629 14844
rect 4663 14841 4675 14875
rect 5258 14872 5264 14884
rect 4617 14835 4675 14841
rect 4724 14844 5264 14872
rect 4028 14776 4154 14804
rect 4295 14807 4353 14813
rect 4028 14764 4034 14776
rect 4295 14773 4307 14807
rect 4341 14804 4353 14807
rect 4724 14804 4752 14844
rect 5258 14832 5264 14844
rect 5316 14832 5322 14884
rect 5353 14875 5411 14881
rect 5353 14841 5365 14875
rect 5399 14872 5411 14875
rect 5626 14872 5632 14884
rect 5399 14844 5632 14872
rect 5399 14841 5411 14844
rect 5353 14835 5411 14841
rect 5626 14832 5632 14844
rect 5684 14832 5690 14884
rect 6273 14875 6331 14881
rect 6273 14841 6285 14875
rect 6319 14872 6331 14875
rect 7098 14872 7104 14884
rect 6319 14844 7104 14872
rect 6319 14841 6331 14844
rect 6273 14835 6331 14841
rect 7098 14832 7104 14844
rect 7156 14832 7162 14884
rect 7190 14832 7196 14884
rect 7248 14872 7254 14884
rect 7837 14875 7895 14881
rect 7837 14872 7849 14875
rect 7248 14844 7849 14872
rect 7248 14832 7254 14844
rect 7837 14841 7849 14844
rect 7883 14841 7895 14875
rect 7837 14835 7895 14841
rect 7929 14875 7987 14881
rect 7929 14841 7941 14875
rect 7975 14841 7987 14875
rect 7929 14835 7987 14841
rect 4341 14776 4752 14804
rect 5644 14804 5672 14832
rect 6549 14807 6607 14813
rect 6549 14804 6561 14807
rect 5644 14776 6561 14804
rect 4341 14773 4353 14776
rect 4295 14767 4353 14773
rect 6549 14773 6561 14776
rect 6595 14804 6607 14807
rect 7006 14804 7012 14816
rect 6595 14776 7012 14804
rect 6595 14773 6607 14776
rect 6549 14767 6607 14773
rect 7006 14764 7012 14776
rect 7064 14764 7070 14816
rect 7653 14807 7711 14813
rect 7653 14773 7665 14807
rect 7699 14804 7711 14807
rect 7944 14804 7972 14835
rect 8018 14832 8024 14884
rect 8076 14872 8082 14884
rect 10105 14872 10133 14912
rect 11698 14900 11704 14912
rect 11756 14900 11762 14952
rect 12487 14949 12515 14980
rect 12897 14977 12909 14980
rect 12943 14977 12955 15011
rect 13538 15008 13544 15020
rect 13499 14980 13544 15008
rect 12897 14971 12955 14977
rect 12472 14943 12530 14949
rect 12472 14909 12484 14943
rect 12518 14909 12530 14943
rect 12912 14940 12940 14971
rect 13538 14968 13544 14980
rect 13596 14968 13602 15020
rect 15381 15011 15439 15017
rect 15381 14977 15393 15011
rect 15427 15008 15439 15011
rect 15470 15008 15476 15020
rect 15427 14980 15476 15008
rect 15427 14977 15439 14980
rect 15381 14971 15439 14977
rect 15470 14968 15476 14980
rect 15528 14968 15534 15020
rect 16022 15008 16028 15020
rect 15983 14980 16028 15008
rect 16022 14968 16028 14980
rect 16080 14968 16086 15020
rect 17310 14968 17316 15020
rect 17368 15008 17374 15020
rect 18690 15008 18696 15020
rect 17368 14980 18696 15008
rect 17368 14968 17374 14980
rect 18690 14968 18696 14980
rect 18748 15008 18754 15020
rect 18748 14980 19155 15008
rect 18748 14968 18754 14980
rect 15194 14940 15200 14952
rect 12912 14912 15200 14940
rect 12472 14903 12530 14909
rect 15194 14900 15200 14912
rect 15252 14900 15258 14952
rect 16758 14940 16764 14952
rect 16719 14912 16764 14940
rect 16758 14900 16764 14912
rect 16816 14940 16822 14952
rect 16888 14943 16946 14949
rect 16888 14940 16900 14943
rect 16816 14912 16900 14940
rect 16816 14900 16822 14912
rect 16888 14909 16900 14912
rect 16934 14909 16946 14943
rect 18084 14943 18142 14949
rect 18084 14940 18096 14943
rect 16888 14903 16946 14909
rect 17604 14912 18096 14940
rect 10298 14875 10356 14881
rect 10298 14872 10310 14875
rect 8076 14844 10133 14872
rect 8076 14832 8082 14844
rect 10289 14841 10310 14872
rect 10344 14841 10356 14875
rect 13792 14875 13850 14881
rect 13792 14872 13804 14875
rect 10289 14835 10356 14841
rect 13372 14844 13804 14872
rect 8202 14804 8208 14816
rect 7699 14776 8208 14804
rect 7699 14773 7711 14776
rect 7653 14767 7711 14773
rect 8202 14764 8208 14776
rect 8260 14764 8266 14816
rect 9401 14807 9459 14813
rect 9401 14773 9413 14807
rect 9447 14804 9459 14807
rect 9490 14804 9496 14816
rect 9447 14776 9496 14804
rect 9447 14773 9459 14776
rect 9401 14767 9459 14773
rect 9490 14764 9496 14776
rect 9548 14804 9554 14816
rect 9766 14804 9772 14816
rect 9548 14776 9772 14804
rect 9548 14764 9554 14776
rect 9766 14764 9772 14776
rect 9824 14804 9830 14816
rect 10134 14804 10140 14816
rect 9824 14776 10140 14804
rect 9824 14764 9830 14776
rect 10134 14764 10140 14776
rect 10192 14804 10198 14816
rect 10289 14804 10317 14835
rect 11790 14804 11796 14816
rect 10192 14776 10317 14804
rect 11751 14776 11796 14804
rect 10192 14764 10198 14776
rect 11790 14764 11796 14776
rect 11848 14764 11854 14816
rect 11882 14764 11888 14816
rect 11940 14804 11946 14816
rect 12575 14807 12633 14813
rect 12575 14804 12587 14807
rect 11940 14776 12587 14804
rect 11940 14764 11946 14776
rect 12575 14773 12587 14776
rect 12621 14773 12633 14807
rect 12575 14767 12633 14773
rect 12894 14764 12900 14816
rect 12952 14804 12958 14816
rect 13262 14804 13268 14816
rect 12952 14776 13268 14804
rect 12952 14764 12958 14776
rect 13262 14764 13268 14776
rect 13320 14804 13326 14816
rect 13372 14813 13400 14844
rect 13792 14841 13804 14844
rect 13838 14841 13850 14875
rect 15473 14875 15531 14881
rect 13792 14835 13850 14841
rect 14752 14844 15332 14872
rect 14752 14813 14780 14844
rect 13357 14807 13415 14813
rect 13357 14804 13369 14807
rect 13320 14776 13369 14804
rect 13320 14764 13326 14776
rect 13357 14773 13369 14776
rect 13403 14773 13415 14807
rect 13357 14767 13415 14773
rect 14461 14807 14519 14813
rect 14461 14773 14473 14807
rect 14507 14804 14519 14807
rect 14737 14807 14795 14813
rect 14737 14804 14749 14807
rect 14507 14776 14749 14804
rect 14507 14773 14519 14776
rect 14461 14767 14519 14773
rect 14737 14773 14749 14776
rect 14783 14773 14795 14807
rect 15304 14804 15332 14844
rect 15473 14841 15485 14875
rect 15519 14841 15531 14875
rect 15473 14835 15531 14841
rect 15488 14804 15516 14835
rect 17604 14816 17632 14912
rect 18084 14909 18096 14912
rect 18130 14940 18142 14943
rect 18414 14940 18420 14952
rect 18130 14912 18420 14940
rect 18130 14909 18142 14912
rect 18084 14903 18142 14909
rect 18414 14900 18420 14912
rect 18472 14940 18478 14952
rect 19127 14949 19155 14980
rect 18509 14943 18567 14949
rect 18509 14940 18521 14943
rect 18472 14912 18521 14940
rect 18472 14900 18478 14912
rect 18509 14909 18521 14912
rect 18555 14909 18567 14943
rect 18509 14903 18567 14909
rect 19112 14943 19170 14949
rect 19112 14909 19124 14943
rect 19158 14940 19170 14943
rect 19521 14943 19579 14949
rect 19521 14940 19533 14943
rect 19158 14912 19533 14940
rect 19158 14909 19170 14912
rect 19112 14903 19170 14909
rect 19521 14909 19533 14912
rect 19567 14909 19579 14943
rect 19521 14903 19579 14909
rect 15304 14776 15516 14804
rect 14737 14767 14795 14773
rect 16850 14764 16856 14816
rect 16908 14804 16914 14816
rect 16991 14807 17049 14813
rect 16991 14804 17003 14807
rect 16908 14776 17003 14804
rect 16908 14764 16914 14776
rect 16991 14773 17003 14776
rect 17037 14773 17049 14807
rect 16991 14767 17049 14773
rect 17586 14764 17592 14816
rect 17644 14764 17650 14816
rect 17678 14764 17684 14816
rect 17736 14804 17742 14816
rect 18187 14807 18245 14813
rect 18187 14804 18199 14807
rect 17736 14776 18199 14804
rect 17736 14764 17742 14776
rect 18187 14773 18199 14776
rect 18233 14773 18245 14807
rect 18187 14767 18245 14773
rect 18598 14764 18604 14816
rect 18656 14804 18662 14816
rect 19889 14807 19947 14813
rect 19889 14804 19901 14807
rect 18656 14776 19901 14804
rect 18656 14764 18662 14776
rect 19889 14773 19901 14776
rect 19935 14773 19947 14807
rect 19889 14767 19947 14773
rect 1104 14714 20884 14736
rect 1104 14662 8315 14714
rect 8367 14662 8379 14714
rect 8431 14662 8443 14714
rect 8495 14662 8507 14714
rect 8559 14662 15648 14714
rect 15700 14662 15712 14714
rect 15764 14662 15776 14714
rect 15828 14662 15840 14714
rect 15892 14662 20884 14714
rect 1104 14640 20884 14662
rect 1670 14600 1676 14612
rect 1631 14572 1676 14600
rect 1670 14560 1676 14572
rect 1728 14560 1734 14612
rect 2958 14560 2964 14612
rect 3016 14600 3022 14612
rect 4430 14600 4436 14612
rect 3016 14572 4436 14600
rect 3016 14560 3022 14572
rect 4430 14560 4436 14572
rect 4488 14560 4494 14612
rect 4617 14603 4675 14609
rect 4617 14569 4629 14603
rect 4663 14600 4675 14603
rect 5258 14600 5264 14612
rect 4663 14572 5264 14600
rect 4663 14569 4675 14572
rect 4617 14563 4675 14569
rect 5258 14560 5264 14572
rect 5316 14560 5322 14612
rect 5442 14560 5448 14612
rect 5500 14600 5506 14612
rect 6273 14603 6331 14609
rect 6273 14600 6285 14603
rect 5500 14572 6285 14600
rect 5500 14560 5506 14572
rect 6273 14569 6285 14572
rect 6319 14569 6331 14603
rect 7006 14600 7012 14612
rect 6967 14572 7012 14600
rect 6273 14563 6331 14569
rect 7006 14560 7012 14572
rect 7064 14560 7070 14612
rect 8202 14560 8208 14612
rect 8260 14600 8266 14612
rect 8481 14603 8539 14609
rect 8481 14600 8493 14603
rect 8260 14572 8493 14600
rect 8260 14560 8266 14572
rect 8481 14569 8493 14572
rect 8527 14569 8539 14603
rect 9950 14600 9956 14612
rect 9911 14572 9956 14600
rect 8481 14563 8539 14569
rect 9950 14560 9956 14572
rect 10008 14560 10014 14612
rect 10226 14560 10232 14612
rect 10284 14600 10290 14612
rect 10413 14603 10471 14609
rect 10413 14600 10425 14603
rect 10284 14572 10425 14600
rect 10284 14560 10290 14572
rect 10413 14569 10425 14572
rect 10459 14569 10471 14603
rect 10413 14563 10471 14569
rect 13538 14560 13544 14612
rect 13596 14600 13602 14612
rect 13909 14603 13967 14609
rect 13909 14600 13921 14603
rect 13596 14572 13921 14600
rect 13596 14560 13602 14572
rect 13909 14569 13921 14572
rect 13955 14569 13967 14603
rect 13909 14563 13967 14569
rect 15286 14560 15292 14612
rect 15344 14600 15350 14612
rect 15344 14572 16160 14600
rect 15344 14560 15350 14572
rect 2130 14492 2136 14544
rect 2188 14532 2194 14544
rect 2225 14535 2283 14541
rect 2225 14532 2237 14535
rect 2188 14504 2237 14532
rect 2188 14492 2194 14504
rect 2225 14501 2237 14504
rect 2271 14501 2283 14535
rect 2225 14495 2283 14501
rect 2777 14535 2835 14541
rect 2777 14501 2789 14535
rect 2823 14532 2835 14535
rect 3050 14532 3056 14544
rect 2823 14504 3056 14532
rect 2823 14501 2835 14504
rect 2777 14495 2835 14501
rect 3050 14492 3056 14504
rect 3108 14492 3114 14544
rect 3326 14492 3332 14544
rect 3384 14532 3390 14544
rect 3602 14532 3608 14544
rect 3384 14504 3608 14532
rect 3384 14492 3390 14504
rect 3602 14492 3608 14504
rect 3660 14492 3666 14544
rect 5071 14535 5129 14541
rect 5071 14501 5083 14535
rect 5117 14532 5129 14535
rect 7098 14532 7104 14544
rect 5117 14504 7104 14532
rect 5117 14501 5129 14504
rect 5071 14495 5129 14501
rect 5276 14476 5304 14504
rect 7098 14492 7104 14504
rect 7156 14532 7162 14544
rect 7923 14535 7981 14541
rect 7923 14532 7935 14535
rect 7156 14504 7935 14532
rect 7156 14492 7162 14504
rect 7923 14501 7935 14504
rect 7969 14532 7981 14535
rect 8294 14532 8300 14544
rect 7969 14504 8300 14532
rect 7969 14501 7981 14504
rect 7923 14495 7981 14501
rect 8294 14492 8300 14504
rect 8352 14532 8358 14544
rect 9490 14532 9496 14544
rect 8352 14504 9496 14532
rect 8352 14492 8358 14504
rect 9490 14492 9496 14504
rect 9548 14492 9554 14544
rect 11146 14532 11152 14544
rect 11107 14504 11152 14532
rect 11146 14492 11152 14504
rect 11204 14492 11210 14544
rect 12710 14532 12716 14544
rect 12671 14504 12716 14532
rect 12710 14492 12716 14504
rect 12768 14492 12774 14544
rect 12894 14492 12900 14544
rect 12952 14532 12958 14544
rect 13633 14535 13691 14541
rect 13633 14532 13645 14535
rect 12952 14504 13645 14532
rect 12952 14492 12958 14504
rect 13633 14501 13645 14504
rect 13679 14501 13691 14535
rect 13633 14495 13691 14501
rect 15378 14492 15384 14544
rect 15436 14532 15442 14544
rect 15473 14535 15531 14541
rect 15473 14532 15485 14535
rect 15436 14504 15485 14532
rect 15436 14492 15442 14504
rect 15473 14501 15485 14504
rect 15519 14501 15531 14535
rect 16022 14532 16028 14544
rect 15983 14504 16028 14532
rect 15473 14495 15531 14501
rect 16022 14492 16028 14504
rect 16080 14492 16086 14544
rect 16132 14532 16160 14572
rect 16666 14560 16672 14612
rect 16724 14600 16730 14612
rect 16945 14603 17003 14609
rect 16945 14600 16957 14603
rect 16724 14572 16957 14600
rect 16724 14560 16730 14572
rect 16945 14569 16957 14572
rect 16991 14569 17003 14603
rect 16945 14563 17003 14569
rect 18555 14535 18613 14541
rect 18555 14532 18567 14535
rect 16132 14504 18567 14532
rect 18555 14501 18567 14504
rect 18601 14501 18613 14535
rect 18555 14495 18613 14501
rect 5258 14424 5264 14476
rect 5316 14424 5322 14476
rect 5626 14464 5632 14476
rect 5587 14436 5632 14464
rect 5626 14424 5632 14436
rect 5684 14424 5690 14476
rect 5902 14424 5908 14476
rect 5960 14464 5966 14476
rect 6638 14473 6644 14476
rect 6584 14467 6644 14473
rect 6584 14464 6596 14467
rect 5960 14436 6596 14464
rect 5960 14424 5966 14436
rect 6584 14433 6596 14436
rect 6630 14433 6644 14467
rect 6584 14427 6644 14433
rect 6638 14424 6644 14427
rect 6696 14424 6702 14476
rect 7374 14424 7380 14476
rect 7432 14464 7438 14476
rect 7561 14467 7619 14473
rect 7561 14464 7573 14467
rect 7432 14436 7573 14464
rect 7432 14424 7438 14436
rect 7561 14433 7573 14436
rect 7607 14464 7619 14467
rect 8202 14464 8208 14476
rect 7607 14436 8208 14464
rect 7607 14433 7619 14436
rect 7561 14427 7619 14433
rect 8202 14424 8208 14436
rect 8260 14424 8266 14476
rect 13262 14424 13268 14476
rect 13320 14464 13326 14476
rect 13722 14464 13728 14476
rect 13320 14436 13728 14464
rect 13320 14424 13326 14436
rect 13722 14424 13728 14436
rect 13780 14464 13786 14476
rect 14090 14464 14096 14476
rect 14148 14473 14154 14476
rect 14148 14467 14186 14473
rect 13780 14436 14096 14464
rect 13780 14424 13786 14436
rect 14090 14424 14096 14436
rect 14174 14433 14186 14467
rect 14148 14427 14186 14433
rect 17129 14467 17187 14473
rect 17129 14433 17141 14467
rect 17175 14464 17187 14467
rect 17218 14464 17224 14476
rect 17175 14436 17224 14464
rect 17175 14433 17187 14436
rect 17129 14427 17187 14433
rect 14148 14424 14154 14427
rect 17218 14424 17224 14436
rect 17276 14424 17282 14476
rect 17402 14464 17408 14476
rect 17363 14436 17408 14464
rect 17402 14424 17408 14436
rect 17460 14424 17466 14476
rect 18414 14464 18420 14476
rect 18375 14436 18420 14464
rect 18414 14424 18420 14436
rect 18472 14424 18478 14476
rect 19058 14424 19064 14476
rect 19116 14464 19122 14476
rect 19464 14467 19522 14473
rect 19464 14464 19476 14467
rect 19116 14436 19476 14464
rect 19116 14424 19122 14436
rect 19464 14433 19476 14436
rect 19510 14464 19522 14467
rect 19886 14464 19892 14476
rect 19510 14436 19892 14464
rect 19510 14433 19522 14436
rect 19464 14427 19522 14433
rect 19886 14424 19892 14436
rect 19944 14424 19950 14476
rect 1670 14356 1676 14408
rect 1728 14396 1734 14408
rect 2133 14399 2191 14405
rect 2133 14396 2145 14399
rect 1728 14368 2145 14396
rect 1728 14356 1734 14368
rect 2133 14365 2145 14368
rect 2179 14396 2191 14399
rect 3421 14399 3479 14405
rect 3421 14396 3433 14399
rect 2179 14368 3433 14396
rect 2179 14365 2191 14368
rect 2133 14359 2191 14365
rect 3421 14365 3433 14368
rect 3467 14365 3479 14399
rect 3421 14359 3479 14365
rect 4522 14356 4528 14408
rect 4580 14396 4586 14408
rect 4709 14399 4767 14405
rect 4709 14396 4721 14399
rect 4580 14368 4721 14396
rect 4580 14356 4586 14368
rect 4709 14365 4721 14368
rect 4755 14365 4767 14399
rect 4709 14359 4767 14365
rect 7466 14356 7472 14408
rect 7524 14396 7530 14408
rect 9674 14396 9680 14408
rect 7524 14368 9680 14396
rect 7524 14356 7530 14368
rect 9674 14356 9680 14368
rect 9732 14356 9738 14408
rect 10042 14356 10048 14408
rect 10100 14396 10106 14408
rect 10686 14396 10692 14408
rect 10100 14368 10692 14396
rect 10100 14356 10106 14368
rect 10686 14356 10692 14368
rect 10744 14356 10750 14408
rect 11054 14396 11060 14408
rect 11015 14368 11060 14396
rect 11054 14356 11060 14368
rect 11112 14356 11118 14408
rect 11698 14396 11704 14408
rect 11659 14368 11704 14396
rect 11698 14356 11704 14368
rect 11756 14396 11762 14408
rect 12345 14399 12403 14405
rect 12345 14396 12357 14399
rect 11756 14368 12357 14396
rect 11756 14356 11762 14368
rect 12345 14365 12357 14368
rect 12391 14396 12403 14399
rect 12621 14399 12679 14405
rect 12621 14396 12633 14399
rect 12391 14368 12633 14396
rect 12391 14365 12403 14368
rect 12345 14359 12403 14365
rect 12621 14365 12633 14368
rect 12667 14365 12679 14399
rect 12986 14396 12992 14408
rect 12947 14368 12992 14396
rect 12621 14359 12679 14365
rect 12986 14356 12992 14368
rect 13044 14356 13050 14408
rect 13446 14356 13452 14408
rect 13504 14396 13510 14408
rect 13504 14368 14642 14396
rect 13504 14356 13510 14368
rect 6687 14331 6745 14337
rect 6687 14297 6699 14331
rect 6733 14328 6745 14331
rect 6914 14328 6920 14340
rect 6733 14300 6920 14328
rect 6733 14297 6745 14300
rect 6687 14291 6745 14297
rect 6914 14288 6920 14300
rect 6972 14288 6978 14340
rect 7190 14288 7196 14340
rect 7248 14328 7254 14340
rect 8757 14331 8815 14337
rect 8757 14328 8769 14331
rect 7248 14300 8769 14328
rect 7248 14288 7254 14300
rect 8757 14297 8769 14300
rect 8803 14297 8815 14331
rect 14231 14331 14289 14337
rect 14231 14328 14243 14331
rect 8757 14291 8815 14297
rect 13280 14300 14243 14328
rect 3050 14260 3056 14272
rect 3011 14232 3056 14260
rect 3050 14220 3056 14232
rect 3108 14220 3114 14272
rect 5718 14220 5724 14272
rect 5776 14260 5782 14272
rect 5905 14263 5963 14269
rect 5905 14260 5917 14263
rect 5776 14232 5917 14260
rect 5776 14220 5782 14232
rect 5905 14229 5917 14232
rect 5951 14229 5963 14263
rect 7466 14260 7472 14272
rect 7427 14232 7472 14260
rect 5905 14223 5963 14229
rect 7466 14220 7472 14232
rect 7524 14220 7530 14272
rect 10962 14220 10968 14272
rect 11020 14260 11026 14272
rect 13280 14260 13308 14300
rect 14231 14297 14243 14300
rect 14277 14297 14289 14331
rect 14614 14328 14642 14368
rect 15010 14356 15016 14408
rect 15068 14396 15074 14408
rect 15381 14399 15439 14405
rect 15381 14396 15393 14399
rect 15068 14368 15393 14396
rect 15068 14356 15074 14368
rect 15381 14365 15393 14368
rect 15427 14365 15439 14399
rect 15381 14359 15439 14365
rect 16758 14356 16764 14408
rect 16816 14396 16822 14408
rect 17770 14396 17776 14408
rect 16816 14368 17776 14396
rect 16816 14356 16822 14368
rect 17770 14356 17776 14368
rect 17828 14356 17834 14408
rect 19567 14331 19625 14337
rect 19567 14328 19579 14331
rect 14614 14300 19579 14328
rect 14231 14291 14289 14297
rect 19567 14297 19579 14300
rect 19613 14297 19625 14331
rect 19567 14291 19625 14297
rect 11020 14232 13308 14260
rect 15105 14263 15163 14269
rect 11020 14220 11026 14232
rect 15105 14229 15117 14263
rect 15151 14260 15163 14263
rect 15470 14260 15476 14272
rect 15151 14232 15476 14260
rect 15151 14229 15163 14232
rect 15105 14223 15163 14229
rect 15470 14220 15476 14232
rect 15528 14220 15534 14272
rect 1104 14170 20884 14192
rect 1104 14118 4648 14170
rect 4700 14118 4712 14170
rect 4764 14118 4776 14170
rect 4828 14118 4840 14170
rect 4892 14118 11982 14170
rect 12034 14118 12046 14170
rect 12098 14118 12110 14170
rect 12162 14118 12174 14170
rect 12226 14118 19315 14170
rect 19367 14118 19379 14170
rect 19431 14118 19443 14170
rect 19495 14118 19507 14170
rect 19559 14118 20884 14170
rect 1104 14096 20884 14118
rect 2130 14016 2136 14068
rect 2188 14056 2194 14068
rect 2317 14059 2375 14065
rect 2317 14056 2329 14059
rect 2188 14028 2329 14056
rect 2188 14016 2194 14028
rect 2317 14025 2329 14028
rect 2363 14056 2375 14059
rect 2961 14059 3019 14065
rect 2961 14056 2973 14059
rect 2363 14028 2973 14056
rect 2363 14025 2375 14028
rect 2317 14019 2375 14025
rect 2961 14025 2973 14028
rect 3007 14025 3019 14059
rect 4801 14059 4859 14065
rect 4801 14056 4813 14059
rect 2961 14019 3019 14025
rect 4126 14028 4813 14056
rect 2590 13948 2596 14000
rect 2648 13988 2654 14000
rect 2648 13960 3648 13988
rect 2648 13948 2654 13960
rect 1397 13923 1455 13929
rect 1397 13889 1409 13923
rect 1443 13920 1455 13923
rect 3050 13920 3056 13932
rect 1443 13892 3056 13920
rect 1443 13889 1455 13892
rect 1397 13883 1455 13889
rect 3050 13880 3056 13892
rect 3108 13880 3114 13932
rect 3620 13920 3648 13960
rect 3694 13948 3700 14000
rect 3752 13988 3758 14000
rect 4126 13988 4154 14028
rect 4801 14025 4813 14028
rect 4847 14056 4859 14059
rect 5258 14056 5264 14068
rect 4847 14028 5264 14056
rect 4847 14025 4859 14028
rect 4801 14019 4859 14025
rect 5258 14016 5264 14028
rect 5316 14016 5322 14068
rect 5350 14016 5356 14068
rect 5408 14056 5414 14068
rect 6086 14056 6092 14068
rect 5408 14028 6092 14056
rect 5408 14016 5414 14028
rect 6086 14016 6092 14028
rect 6144 14016 6150 14068
rect 6638 14056 6644 14068
rect 6599 14028 6644 14056
rect 6638 14016 6644 14028
rect 6696 14016 6702 14068
rect 7466 14016 7472 14068
rect 7524 14056 7530 14068
rect 8527 14059 8585 14065
rect 8527 14056 8539 14059
rect 7524 14028 8539 14056
rect 7524 14016 7530 14028
rect 8527 14025 8539 14028
rect 8573 14025 8585 14059
rect 9214 14056 9220 14068
rect 9175 14028 9220 14056
rect 8527 14019 8585 14025
rect 9214 14016 9220 14028
rect 9272 14016 9278 14068
rect 9490 14016 9496 14068
rect 9548 14056 9554 14068
rect 9585 14059 9643 14065
rect 9585 14056 9597 14059
rect 9548 14028 9597 14056
rect 9548 14016 9554 14028
rect 9585 14025 9597 14028
rect 9631 14056 9643 14059
rect 9858 14056 9864 14068
rect 9631 14028 9864 14056
rect 9631 14025 9643 14028
rect 9585 14019 9643 14025
rect 9858 14016 9864 14028
rect 9916 14016 9922 14068
rect 11054 14016 11060 14068
rect 11112 14056 11118 14068
rect 11333 14059 11391 14065
rect 11333 14056 11345 14059
rect 11112 14028 11345 14056
rect 11112 14016 11118 14028
rect 11333 14025 11345 14028
rect 11379 14025 11391 14059
rect 11333 14019 11391 14025
rect 11422 14016 11428 14068
rect 11480 14056 11486 14068
rect 11885 14059 11943 14065
rect 11885 14056 11897 14059
rect 11480 14028 11897 14056
rect 11480 14016 11486 14028
rect 11885 14025 11897 14028
rect 11931 14056 11943 14059
rect 12710 14056 12716 14068
rect 11931 14028 12716 14056
rect 11931 14025 11943 14028
rect 11885 14019 11943 14025
rect 12710 14016 12716 14028
rect 12768 14016 12774 14068
rect 14090 14056 14096 14068
rect 14051 14028 14096 14056
rect 14090 14016 14096 14028
rect 14148 14016 14154 14068
rect 15194 14016 15200 14068
rect 15252 14056 15258 14068
rect 18509 14059 18567 14065
rect 18509 14056 18521 14059
rect 15252 14028 18521 14056
rect 15252 14016 15258 14028
rect 3752 13960 4154 13988
rect 3752 13948 3758 13960
rect 6270 13920 6276 13932
rect 3620 13892 6276 13920
rect 2590 13852 2596 13864
rect 2551 13824 2596 13852
rect 2590 13812 2596 13824
rect 2648 13812 2654 13864
rect 3620 13861 3648 13892
rect 6270 13880 6276 13892
rect 6328 13880 6334 13932
rect 6638 13920 6644 13932
rect 6472 13892 6644 13920
rect 3605 13855 3663 13861
rect 3605 13821 3617 13855
rect 3651 13852 3663 13855
rect 3694 13852 3700 13864
rect 3651 13824 3700 13852
rect 3651 13821 3663 13824
rect 3605 13815 3663 13821
rect 3694 13812 3700 13824
rect 3752 13812 3758 13864
rect 4065 13855 4123 13861
rect 4065 13821 4077 13855
rect 4111 13821 4123 13855
rect 4065 13815 4123 13821
rect 5445 13855 5503 13861
rect 5445 13821 5457 13855
rect 5491 13852 5503 13855
rect 5626 13852 5632 13864
rect 5491 13824 5632 13852
rect 5491 13821 5503 13824
rect 5445 13815 5503 13821
rect 1762 13716 1768 13728
rect 1723 13688 1768 13716
rect 1762 13676 1768 13688
rect 1820 13676 1826 13728
rect 3418 13676 3424 13728
rect 3476 13716 3482 13728
rect 3513 13719 3571 13725
rect 3513 13716 3525 13719
rect 3476 13688 3525 13716
rect 3476 13676 3482 13688
rect 3513 13685 3525 13688
rect 3559 13716 3571 13719
rect 3602 13716 3608 13728
rect 3559 13688 3608 13716
rect 3559 13685 3571 13688
rect 3513 13679 3571 13685
rect 3602 13676 3608 13688
rect 3660 13716 3666 13728
rect 4080 13716 4108 13815
rect 5626 13812 5632 13824
rect 5684 13812 5690 13864
rect 5721 13855 5779 13861
rect 5721 13821 5733 13855
rect 5767 13852 5779 13855
rect 6181 13855 6239 13861
rect 6181 13852 6193 13855
rect 5767 13824 6193 13852
rect 5767 13821 5779 13824
rect 5721 13815 5779 13821
rect 6181 13821 6193 13824
rect 6227 13852 6239 13855
rect 6472 13852 6500 13892
rect 6638 13880 6644 13892
rect 6696 13880 6702 13932
rect 6917 13923 6975 13929
rect 6917 13889 6929 13923
rect 6963 13920 6975 13923
rect 7484 13920 7512 14016
rect 7742 13948 7748 14000
rect 7800 13988 7806 14000
rect 7926 13988 7932 14000
rect 7800 13960 7932 13988
rect 7800 13948 7806 13960
rect 7926 13948 7932 13960
rect 7984 13948 7990 14000
rect 8202 13988 8208 14000
rect 8163 13960 8208 13988
rect 8202 13948 8208 13960
rect 8260 13948 8266 14000
rect 6963 13892 7512 13920
rect 9232 13920 9260 14016
rect 10134 13948 10140 14000
rect 10192 13988 10198 14000
rect 12161 13991 12219 13997
rect 12161 13988 12173 13991
rect 10192 13960 12173 13988
rect 10192 13948 10198 13960
rect 12161 13957 12173 13960
rect 12207 13957 12219 13991
rect 12161 13951 12219 13957
rect 13449 13991 13507 13997
rect 13449 13957 13461 13991
rect 13495 13988 13507 13991
rect 15378 13988 15384 14000
rect 13495 13960 15384 13988
rect 13495 13957 13507 13960
rect 13449 13951 13507 13957
rect 9769 13923 9827 13929
rect 9769 13920 9781 13923
rect 9232 13892 9781 13920
rect 6963 13889 6975 13892
rect 6917 13883 6975 13889
rect 9769 13889 9781 13892
rect 9815 13889 9827 13923
rect 9769 13883 9827 13889
rect 6227 13824 6500 13852
rect 7837 13855 7895 13861
rect 6227 13821 6239 13824
rect 6181 13815 6239 13821
rect 7837 13821 7849 13855
rect 7883 13852 7895 13855
rect 8294 13852 8300 13864
rect 7883 13824 8300 13852
rect 7883 13821 7895 13824
rect 7837 13815 7895 13821
rect 8294 13812 8300 13824
rect 8352 13812 8358 13864
rect 8424 13855 8482 13861
rect 8424 13821 8436 13855
rect 8470 13821 8482 13855
rect 8424 13815 8482 13821
rect 4338 13784 4344 13796
rect 4299 13756 4344 13784
rect 4338 13744 4344 13756
rect 4396 13744 4402 13796
rect 5905 13787 5963 13793
rect 5905 13753 5917 13787
rect 5951 13784 5963 13787
rect 7006 13784 7012 13796
rect 5951 13756 6361 13784
rect 6967 13756 7012 13784
rect 5951 13753 5963 13756
rect 5905 13747 5963 13753
rect 3660 13688 4108 13716
rect 6333 13716 6361 13756
rect 7006 13744 7012 13756
rect 7064 13744 7070 13796
rect 7190 13744 7196 13796
rect 7248 13784 7254 13796
rect 7558 13784 7564 13796
rect 7248 13756 7564 13784
rect 7248 13744 7254 13756
rect 7558 13744 7564 13756
rect 7616 13744 7622 13796
rect 8202 13744 8208 13796
rect 8260 13784 8266 13796
rect 8439 13784 8467 13815
rect 8849 13787 8907 13793
rect 8849 13784 8861 13787
rect 8260 13756 8861 13784
rect 8260 13744 8266 13756
rect 8849 13753 8861 13756
rect 8895 13784 8907 13787
rect 9030 13784 9036 13796
rect 8895 13756 9036 13784
rect 8895 13753 8907 13756
rect 8849 13747 8907 13753
rect 9030 13744 9036 13756
rect 9088 13744 9094 13796
rect 9858 13744 9864 13796
rect 9916 13784 9922 13796
rect 10090 13787 10148 13793
rect 10090 13784 10102 13787
rect 9916 13756 10102 13784
rect 9916 13744 9922 13756
rect 10090 13753 10102 13756
rect 10136 13753 10148 13787
rect 10090 13747 10148 13753
rect 11330 13744 11336 13796
rect 11388 13784 11394 13796
rect 11974 13784 11980 13796
rect 11388 13756 11980 13784
rect 11388 13744 11394 13756
rect 11974 13744 11980 13756
rect 12032 13744 12038 13796
rect 12176 13784 12204 13951
rect 15378 13948 15384 13960
rect 15436 13988 15442 14000
rect 15473 13991 15531 13997
rect 15473 13988 15485 13991
rect 15436 13960 15485 13988
rect 15436 13948 15442 13960
rect 15473 13957 15485 13960
rect 15519 13957 15531 13991
rect 16942 13988 16948 14000
rect 15473 13951 15531 13957
rect 15923 13960 16948 13988
rect 12526 13920 12532 13932
rect 12487 13892 12532 13920
rect 12526 13880 12532 13892
rect 12584 13880 12590 13932
rect 13817 13923 13875 13929
rect 13817 13889 13829 13923
rect 13863 13920 13875 13923
rect 14277 13923 14335 13929
rect 14277 13920 14289 13923
rect 13863 13892 14289 13920
rect 13863 13889 13875 13892
rect 13817 13883 13875 13889
rect 14277 13889 14289 13892
rect 14323 13920 14335 13923
rect 15923 13920 15951 13960
rect 16942 13948 16948 13960
rect 17000 13948 17006 14000
rect 17129 13991 17187 13997
rect 17129 13957 17141 13991
rect 17175 13988 17187 13991
rect 17402 13988 17408 14000
rect 17175 13960 17408 13988
rect 17175 13957 17187 13960
rect 17129 13951 17187 13957
rect 17402 13948 17408 13960
rect 17460 13948 17466 14000
rect 14323 13892 15951 13920
rect 16117 13923 16175 13929
rect 14323 13889 14335 13892
rect 14277 13883 14335 13889
rect 16117 13889 16129 13923
rect 16163 13920 16175 13923
rect 16390 13920 16396 13932
rect 16163 13892 16396 13920
rect 16163 13889 16175 13892
rect 16117 13883 16175 13889
rect 16390 13880 16396 13892
rect 16448 13880 16454 13932
rect 18099 13861 18127 14028
rect 18509 14025 18521 14028
rect 18555 14056 18567 14059
rect 18598 14056 18604 14068
rect 18555 14028 18604 14056
rect 18555 14025 18567 14028
rect 18509 14019 18567 14025
rect 18598 14016 18604 14028
rect 18656 14016 18662 14068
rect 19886 14056 19892 14068
rect 19847 14028 19892 14056
rect 19886 14016 19892 14028
rect 19944 14016 19950 14068
rect 18414 13948 18420 14000
rect 18472 13988 18478 14000
rect 18877 13991 18935 13997
rect 18877 13988 18889 13991
rect 18472 13960 18889 13988
rect 18472 13948 18478 13960
rect 18877 13957 18889 13960
rect 18923 13957 18935 13991
rect 18877 13951 18935 13957
rect 19076 13960 19334 13988
rect 18322 13880 18328 13932
rect 18380 13920 18386 13932
rect 19076 13920 19104 13960
rect 18380 13892 19104 13920
rect 19306 13920 19334 13960
rect 19521 13923 19579 13929
rect 19521 13920 19533 13923
rect 19306 13892 19533 13920
rect 18380 13880 18386 13892
rect 18084 13855 18142 13861
rect 18084 13821 18096 13855
rect 18130 13821 18142 13855
rect 18084 13815 18142 13821
rect 19128 13855 19186 13861
rect 19128 13821 19140 13855
rect 19174 13852 19186 13855
rect 19306 13852 19334 13892
rect 19521 13889 19533 13892
rect 19567 13889 19579 13923
rect 19521 13883 19579 13889
rect 19174 13824 19334 13852
rect 19174 13821 19186 13824
rect 19128 13815 19186 13821
rect 12894 13793 12900 13796
rect 12850 13787 12900 13793
rect 12850 13784 12862 13787
rect 12176 13756 12862 13784
rect 12850 13753 12862 13756
rect 12896 13753 12900 13787
rect 12850 13747 12900 13753
rect 12894 13744 12900 13747
rect 12952 13784 12958 13796
rect 14090 13784 14096 13796
rect 12952 13756 14096 13784
rect 12952 13744 12958 13756
rect 14090 13744 14096 13756
rect 14148 13784 14154 13796
rect 14598 13787 14656 13793
rect 14598 13784 14610 13787
rect 14148 13756 14610 13784
rect 14148 13744 14154 13756
rect 14598 13753 14610 13756
rect 14644 13753 14656 13787
rect 16209 13787 16267 13793
rect 16209 13784 16221 13787
rect 14598 13747 14656 13753
rect 15856 13756 16221 13784
rect 9674 13716 9680 13728
rect 6333 13688 9680 13716
rect 3660 13676 3666 13688
rect 9674 13676 9680 13688
rect 9732 13676 9738 13728
rect 10689 13719 10747 13725
rect 10689 13685 10701 13719
rect 10735 13716 10747 13719
rect 11057 13719 11115 13725
rect 11057 13716 11069 13719
rect 10735 13688 11069 13716
rect 10735 13685 10747 13688
rect 10689 13679 10747 13685
rect 11057 13685 11069 13688
rect 11103 13716 11115 13719
rect 11146 13716 11152 13728
rect 11103 13688 11152 13716
rect 11103 13685 11115 13688
rect 11057 13679 11115 13685
rect 11146 13676 11152 13688
rect 11204 13716 11210 13728
rect 11606 13716 11612 13728
rect 11204 13688 11612 13716
rect 11204 13676 11210 13688
rect 11606 13676 11612 13688
rect 11664 13676 11670 13728
rect 15197 13719 15255 13725
rect 15197 13685 15209 13719
rect 15243 13716 15255 13719
rect 15378 13716 15384 13728
rect 15243 13688 15384 13716
rect 15243 13685 15255 13688
rect 15197 13679 15255 13685
rect 15378 13676 15384 13688
rect 15436 13716 15442 13728
rect 15856 13725 15884 13756
rect 16209 13753 16221 13756
rect 16255 13753 16267 13787
rect 16758 13784 16764 13796
rect 16719 13756 16764 13784
rect 16209 13747 16267 13753
rect 16758 13744 16764 13756
rect 16816 13744 16822 13796
rect 15841 13719 15899 13725
rect 15841 13716 15853 13719
rect 15436 13688 15853 13716
rect 15436 13676 15442 13688
rect 15841 13685 15853 13688
rect 15887 13685 15899 13719
rect 15841 13679 15899 13685
rect 16666 13676 16672 13728
rect 16724 13716 16730 13728
rect 17034 13716 17040 13728
rect 16724 13688 17040 13716
rect 16724 13676 16730 13688
rect 17034 13676 17040 13688
rect 17092 13676 17098 13728
rect 17218 13676 17224 13728
rect 17276 13716 17282 13728
rect 17405 13719 17463 13725
rect 17405 13716 17417 13719
rect 17276 13688 17417 13716
rect 17276 13676 17282 13688
rect 17405 13685 17417 13688
rect 17451 13685 17463 13719
rect 17405 13679 17463 13685
rect 17494 13676 17500 13728
rect 17552 13716 17558 13728
rect 18187 13719 18245 13725
rect 18187 13716 18199 13719
rect 17552 13688 18199 13716
rect 17552 13676 17558 13688
rect 18187 13685 18199 13688
rect 18233 13685 18245 13719
rect 18187 13679 18245 13685
rect 18598 13676 18604 13728
rect 18656 13716 18662 13728
rect 19199 13719 19257 13725
rect 19199 13716 19211 13719
rect 18656 13688 19211 13716
rect 18656 13676 18662 13688
rect 19199 13685 19211 13688
rect 19245 13685 19257 13719
rect 19199 13679 19257 13685
rect 1104 13626 20884 13648
rect 1104 13574 8315 13626
rect 8367 13574 8379 13626
rect 8431 13574 8443 13626
rect 8495 13574 8507 13626
rect 8559 13574 15648 13626
rect 15700 13574 15712 13626
rect 15764 13574 15776 13626
rect 15828 13574 15840 13626
rect 15892 13574 20884 13626
rect 1104 13552 20884 13574
rect 1535 13515 1593 13521
rect 1535 13481 1547 13515
rect 1581 13512 1593 13515
rect 1670 13512 1676 13524
rect 1581 13484 1676 13512
rect 1581 13481 1593 13484
rect 1535 13475 1593 13481
rect 1670 13472 1676 13484
rect 1728 13472 1734 13524
rect 2314 13512 2320 13524
rect 2227 13484 2320 13512
rect 2314 13472 2320 13484
rect 2372 13512 2378 13524
rect 3510 13512 3516 13524
rect 2372 13484 3516 13512
rect 2372 13472 2378 13484
rect 3510 13472 3516 13484
rect 3568 13472 3574 13524
rect 3694 13512 3700 13524
rect 3655 13484 3700 13512
rect 3694 13472 3700 13484
rect 3752 13472 3758 13524
rect 8202 13512 8208 13524
rect 4908 13484 8208 13512
rect 3145 13447 3203 13453
rect 3145 13413 3157 13447
rect 3191 13444 3203 13447
rect 4522 13444 4528 13456
rect 3191 13416 4528 13444
rect 3191 13413 3203 13416
rect 3145 13407 3203 13413
rect 4522 13404 4528 13416
rect 4580 13444 4586 13456
rect 4709 13447 4767 13453
rect 4709 13444 4721 13447
rect 4580 13416 4721 13444
rect 4580 13404 4586 13416
rect 4709 13413 4721 13416
rect 4755 13413 4767 13447
rect 4709 13407 4767 13413
rect 1302 13336 1308 13388
rect 1360 13376 1366 13388
rect 1432 13379 1490 13385
rect 1432 13376 1444 13379
rect 1360 13348 1444 13376
rect 1360 13336 1366 13348
rect 1432 13345 1444 13348
rect 1478 13345 1490 13379
rect 1432 13339 1490 13345
rect 1447 13308 1475 13339
rect 1762 13336 1768 13388
rect 1820 13376 1826 13388
rect 2590 13376 2596 13388
rect 1820 13348 2596 13376
rect 1820 13336 1826 13348
rect 2590 13336 2596 13348
rect 2648 13336 2654 13388
rect 2961 13379 3019 13385
rect 2961 13345 2973 13379
rect 3007 13376 3019 13379
rect 3786 13376 3792 13388
rect 3007 13348 3792 13376
rect 3007 13345 3019 13348
rect 2961 13339 3019 13345
rect 3786 13336 3792 13348
rect 3844 13336 3850 13388
rect 3973 13379 4031 13385
rect 3973 13345 3985 13379
rect 4019 13376 4031 13379
rect 4062 13376 4068 13388
rect 4019 13348 4068 13376
rect 4019 13345 4031 13348
rect 3973 13339 4031 13345
rect 4062 13336 4068 13348
rect 4120 13336 4126 13388
rect 1857 13311 1915 13317
rect 1857 13308 1869 13311
rect 1447 13280 1869 13308
rect 1857 13277 1869 13280
rect 1903 13308 1915 13311
rect 4908 13308 4936 13484
rect 8202 13472 8208 13484
rect 8260 13472 8266 13524
rect 10962 13512 10968 13524
rect 10923 13484 10968 13512
rect 10962 13472 10968 13484
rect 11020 13472 11026 13524
rect 11146 13472 11152 13524
rect 11204 13512 11210 13524
rect 11514 13512 11520 13524
rect 11204 13484 11520 13512
rect 11204 13472 11210 13484
rect 11514 13472 11520 13484
rect 11572 13472 11578 13524
rect 12526 13512 12532 13524
rect 12487 13484 12532 13512
rect 12526 13472 12532 13484
rect 12584 13472 12590 13524
rect 13906 13472 13912 13524
rect 13964 13512 13970 13524
rect 14366 13512 14372 13524
rect 13964 13484 14372 13512
rect 13964 13472 13970 13484
rect 14366 13472 14372 13484
rect 14424 13512 14430 13524
rect 14645 13515 14703 13521
rect 14645 13512 14657 13515
rect 14424 13484 14657 13512
rect 14424 13472 14430 13484
rect 14645 13481 14657 13484
rect 14691 13481 14703 13515
rect 16942 13512 16948 13524
rect 16903 13484 16948 13512
rect 14645 13475 14703 13481
rect 16942 13472 16948 13484
rect 17000 13472 17006 13524
rect 18509 13515 18567 13521
rect 18509 13512 18521 13515
rect 17788 13484 18521 13512
rect 5258 13404 5264 13456
rect 5316 13444 5322 13456
rect 5398 13447 5456 13453
rect 5398 13444 5410 13447
rect 5316 13416 5410 13444
rect 5316 13404 5322 13416
rect 5398 13413 5410 13416
rect 5444 13413 5456 13447
rect 6270 13444 6276 13456
rect 5398 13407 5456 13413
rect 6012 13416 6276 13444
rect 6012 13385 6040 13416
rect 6270 13404 6276 13416
rect 6328 13444 6334 13456
rect 7009 13447 7067 13453
rect 7009 13444 7021 13447
rect 6328 13416 7021 13444
rect 6328 13404 6334 13416
rect 7009 13413 7021 13416
rect 7055 13413 7067 13447
rect 7009 13407 7067 13413
rect 9858 13404 9864 13456
rect 9916 13444 9922 13456
rect 9998 13447 10056 13453
rect 9998 13444 10010 13447
rect 9916 13416 10010 13444
rect 9916 13404 9922 13416
rect 9998 13413 10010 13416
rect 10044 13413 10056 13447
rect 11606 13444 11612 13456
rect 11567 13416 11612 13444
rect 9998 13407 10056 13413
rect 11606 13404 11612 13416
rect 11664 13404 11670 13456
rect 13722 13444 13728 13456
rect 13280 13416 13728 13444
rect 5997 13379 6055 13385
rect 5997 13345 6009 13379
rect 6043 13345 6055 13379
rect 5997 13339 6055 13345
rect 7926 13336 7932 13388
rect 7984 13376 7990 13388
rect 8424 13379 8482 13385
rect 8424 13376 8436 13379
rect 7984 13348 8436 13376
rect 7984 13336 7990 13348
rect 8424 13345 8436 13348
rect 8470 13345 8482 13379
rect 9674 13376 9680 13388
rect 9635 13348 9680 13376
rect 8424 13339 8482 13345
rect 9674 13336 9680 13348
rect 9732 13336 9738 13388
rect 13280 13385 13308 13416
rect 13722 13404 13728 13416
rect 13780 13444 13786 13456
rect 13780 13416 13952 13444
rect 13780 13404 13786 13416
rect 13924 13388 13952 13416
rect 14090 13404 14096 13456
rect 14148 13444 14154 13456
rect 14277 13447 14335 13453
rect 14277 13444 14289 13447
rect 14148 13416 14289 13444
rect 14148 13404 14154 13416
rect 14277 13413 14289 13416
rect 14323 13413 14335 13447
rect 14277 13407 14335 13413
rect 15378 13404 15384 13456
rect 15436 13444 15442 13456
rect 15473 13447 15531 13453
rect 15473 13444 15485 13447
rect 15436 13416 15485 13444
rect 15436 13404 15442 13416
rect 15473 13413 15485 13416
rect 15519 13413 15531 13447
rect 17218 13444 17224 13456
rect 15473 13407 15531 13413
rect 16960 13416 17224 13444
rect 13265 13379 13323 13385
rect 13265 13345 13277 13379
rect 13311 13345 13323 13379
rect 13446 13376 13452 13388
rect 13407 13348 13452 13376
rect 13265 13339 13323 13345
rect 13446 13336 13452 13348
rect 13504 13336 13510 13388
rect 13906 13336 13912 13388
rect 13964 13336 13970 13388
rect 16960 13385 16988 13416
rect 17218 13404 17224 13416
rect 17276 13404 17282 13456
rect 16945 13379 17003 13385
rect 16945 13345 16957 13379
rect 16991 13345 17003 13379
rect 16945 13339 17003 13345
rect 17034 13336 17040 13388
rect 17092 13376 17098 13388
rect 17313 13379 17371 13385
rect 17313 13376 17325 13379
rect 17092 13348 17325 13376
rect 17092 13336 17098 13348
rect 17313 13345 17325 13348
rect 17359 13345 17371 13379
rect 17788 13376 17816 13484
rect 18509 13481 18521 13484
rect 18555 13481 18567 13515
rect 18509 13475 18567 13481
rect 18782 13472 18788 13524
rect 18840 13512 18846 13524
rect 20162 13512 20168 13524
rect 18840 13484 20168 13512
rect 18840 13472 18846 13484
rect 20162 13472 20168 13484
rect 20220 13472 20226 13524
rect 17313 13339 17371 13345
rect 17420 13348 17816 13376
rect 5074 13308 5080 13320
rect 1903 13280 4936 13308
rect 4987 13280 5080 13308
rect 1903 13277 1915 13280
rect 1857 13271 1915 13277
rect 5074 13268 5080 13280
rect 5132 13308 5138 13320
rect 5534 13308 5540 13320
rect 5132 13280 5540 13308
rect 5132 13268 5138 13280
rect 5534 13268 5540 13280
rect 5592 13268 5598 13320
rect 6917 13311 6975 13317
rect 6917 13308 6929 13311
rect 6656 13280 6929 13308
rect 6656 13249 6684 13280
rect 6917 13277 6929 13280
rect 6963 13277 6975 13311
rect 11514 13308 11520 13320
rect 11427 13280 11520 13308
rect 6917 13271 6975 13277
rect 11514 13268 11520 13280
rect 11572 13308 11578 13320
rect 11882 13308 11888 13320
rect 11572 13280 11888 13308
rect 11572 13268 11578 13280
rect 11882 13268 11888 13280
rect 11940 13268 11946 13320
rect 13538 13308 13544 13320
rect 13499 13280 13544 13308
rect 13538 13268 13544 13280
rect 13596 13268 13602 13320
rect 15194 13268 15200 13320
rect 15252 13308 15258 13320
rect 15381 13311 15439 13317
rect 15381 13308 15393 13311
rect 15252 13280 15393 13308
rect 15252 13268 15258 13280
rect 15381 13277 15393 13280
rect 15427 13277 15439 13311
rect 15381 13271 15439 13277
rect 15470 13268 15476 13320
rect 15528 13308 15534 13320
rect 15657 13311 15715 13317
rect 15657 13308 15669 13311
rect 15528 13280 15669 13308
rect 15528 13268 15534 13280
rect 15657 13277 15669 13280
rect 15703 13277 15715 13311
rect 17420 13308 17448 13348
rect 18230 13336 18236 13388
rect 18288 13376 18294 13388
rect 18417 13379 18475 13385
rect 18417 13376 18429 13379
rect 18288 13348 18429 13376
rect 18288 13336 18294 13348
rect 18417 13345 18429 13348
rect 18463 13345 18475 13379
rect 18874 13376 18880 13388
rect 18835 13348 18880 13376
rect 18417 13339 18475 13345
rect 18874 13336 18880 13348
rect 18932 13336 18938 13388
rect 15657 13271 15715 13277
rect 15856 13280 17448 13308
rect 4203 13243 4261 13249
rect 4203 13209 4215 13243
rect 4249 13240 4261 13243
rect 6641 13243 6699 13249
rect 6641 13240 6653 13243
rect 4249 13212 6653 13240
rect 4249 13209 4261 13212
rect 4203 13203 4261 13209
rect 6641 13209 6653 13212
rect 6687 13209 6699 13243
rect 7466 13240 7472 13252
rect 7427 13212 7472 13240
rect 6641 13203 6699 13209
rect 7466 13200 7472 13212
rect 7524 13200 7530 13252
rect 10597 13243 10655 13249
rect 10597 13209 10609 13243
rect 10643 13240 10655 13243
rect 11422 13240 11428 13252
rect 10643 13212 11428 13240
rect 10643 13209 10655 13212
rect 10597 13203 10655 13209
rect 11422 13200 11428 13212
rect 11480 13200 11486 13252
rect 12069 13243 12127 13249
rect 12069 13209 12081 13243
rect 12115 13209 12127 13243
rect 12069 13203 12127 13209
rect 2590 13132 2596 13184
rect 2648 13172 2654 13184
rect 2958 13172 2964 13184
rect 2648 13144 2964 13172
rect 2648 13132 2654 13144
rect 2958 13132 2964 13144
rect 3016 13132 3022 13184
rect 6086 13132 6092 13184
rect 6144 13172 6150 13184
rect 6365 13175 6423 13181
rect 6365 13172 6377 13175
rect 6144 13144 6377 13172
rect 6144 13132 6150 13144
rect 6365 13141 6377 13144
rect 6411 13172 6423 13175
rect 8527 13175 8585 13181
rect 8527 13172 8539 13175
rect 6411 13144 8539 13172
rect 6411 13141 6423 13144
rect 6365 13135 6423 13141
rect 8527 13141 8539 13144
rect 8573 13141 8585 13175
rect 8527 13135 8585 13141
rect 10410 13132 10416 13184
rect 10468 13172 10474 13184
rect 11790 13172 11796 13184
rect 10468 13144 11796 13172
rect 10468 13132 10474 13144
rect 11790 13132 11796 13144
rect 11848 13172 11854 13184
rect 12084 13172 12112 13203
rect 12894 13200 12900 13252
rect 12952 13240 12958 13252
rect 15856 13240 15884 13280
rect 16390 13240 16396 13252
rect 12952 13212 15884 13240
rect 16303 13212 16396 13240
rect 12952 13200 12958 13212
rect 16390 13200 16396 13212
rect 16448 13240 16454 13252
rect 18598 13240 18604 13252
rect 16448 13212 18604 13240
rect 16448 13200 16454 13212
rect 18598 13200 18604 13212
rect 18656 13200 18662 13252
rect 12802 13172 12808 13184
rect 11848 13144 12808 13172
rect 11848 13132 11854 13144
rect 12802 13132 12808 13144
rect 12860 13132 12866 13184
rect 15010 13132 15016 13184
rect 15068 13172 15074 13184
rect 15105 13175 15163 13181
rect 15105 13172 15117 13175
rect 15068 13144 15117 13172
rect 15068 13132 15074 13144
rect 15105 13141 15117 13144
rect 15151 13172 15163 13175
rect 16758 13172 16764 13184
rect 15151 13144 16764 13172
rect 15151 13141 15163 13144
rect 15105 13135 15163 13141
rect 16758 13132 16764 13144
rect 16816 13132 16822 13184
rect 1104 13082 20884 13104
rect 1104 13030 4648 13082
rect 4700 13030 4712 13082
rect 4764 13030 4776 13082
rect 4828 13030 4840 13082
rect 4892 13030 11982 13082
rect 12034 13030 12046 13082
rect 12098 13030 12110 13082
rect 12162 13030 12174 13082
rect 12226 13030 19315 13082
rect 19367 13030 19379 13082
rect 19431 13030 19443 13082
rect 19495 13030 19507 13082
rect 19559 13030 20884 13082
rect 1104 13008 20884 13030
rect 2593 12971 2651 12977
rect 2593 12937 2605 12971
rect 2639 12968 2651 12971
rect 2682 12968 2688 12980
rect 2639 12940 2688 12968
rect 2639 12937 2651 12940
rect 2593 12931 2651 12937
rect 2682 12928 2688 12940
rect 2740 12928 2746 12980
rect 3786 12968 3792 12980
rect 3747 12940 3792 12968
rect 3786 12928 3792 12940
rect 3844 12928 3850 12980
rect 5077 12971 5135 12977
rect 5077 12937 5089 12971
rect 5123 12968 5135 12971
rect 5258 12968 5264 12980
rect 5123 12940 5264 12968
rect 5123 12937 5135 12940
rect 5077 12931 5135 12937
rect 5258 12928 5264 12940
rect 5316 12968 5322 12980
rect 5718 12968 5724 12980
rect 5316 12940 5724 12968
rect 5316 12928 5322 12940
rect 5718 12928 5724 12940
rect 5776 12928 5782 12980
rect 6270 12968 6276 12980
rect 6231 12940 6276 12968
rect 6270 12928 6276 12940
rect 6328 12928 6334 12980
rect 9674 12928 9680 12980
rect 9732 12968 9738 12980
rect 10045 12971 10103 12977
rect 10045 12968 10057 12971
rect 9732 12940 10057 12968
rect 9732 12928 9738 12940
rect 10045 12937 10057 12940
rect 10091 12937 10103 12971
rect 11606 12968 11612 12980
rect 11567 12940 11612 12968
rect 10045 12931 10103 12937
rect 11606 12928 11612 12940
rect 11664 12928 11670 12980
rect 12342 12968 12348 12980
rect 11716 12940 12348 12968
rect 2774 12900 2780 12912
rect 2735 12872 2780 12900
rect 2774 12860 2780 12872
rect 2832 12860 2838 12912
rect 7466 12900 7472 12912
rect 7427 12872 7472 12900
rect 7466 12860 7472 12872
rect 7524 12860 7530 12912
rect 9582 12860 9588 12912
rect 9640 12900 9646 12912
rect 9858 12900 9864 12912
rect 9640 12872 9864 12900
rect 9640 12860 9646 12872
rect 9858 12860 9864 12872
rect 9916 12860 9922 12912
rect 11716 12900 11744 12940
rect 12342 12928 12348 12940
rect 12400 12968 12406 12980
rect 13446 12968 13452 12980
rect 12400 12940 13452 12968
rect 12400 12928 12406 12940
rect 13446 12928 13452 12940
rect 13504 12968 13510 12980
rect 13722 12968 13728 12980
rect 13504 12940 13728 12968
rect 13504 12928 13510 12940
rect 13722 12928 13728 12940
rect 13780 12968 13786 12980
rect 15197 12971 15255 12977
rect 15197 12968 15209 12971
rect 13780 12940 15209 12968
rect 13780 12928 13786 12940
rect 15197 12937 15209 12940
rect 15243 12937 15255 12971
rect 15378 12968 15384 12980
rect 15339 12940 15384 12968
rect 15197 12931 15255 12937
rect 15378 12928 15384 12940
rect 15436 12928 15442 12980
rect 17402 12928 17408 12980
rect 17460 12968 17466 12980
rect 17773 12971 17831 12977
rect 17773 12968 17785 12971
rect 17460 12940 17785 12968
rect 17460 12928 17466 12940
rect 17773 12937 17785 12940
rect 17819 12937 17831 12971
rect 17773 12931 17831 12937
rect 10105 12872 11744 12900
rect 5261 12835 5319 12841
rect 5261 12801 5273 12835
rect 5307 12832 5319 12835
rect 6086 12832 6092 12844
rect 5307 12804 6092 12832
rect 5307 12801 5319 12804
rect 5261 12795 5319 12801
rect 6086 12792 6092 12804
rect 6144 12792 6150 12844
rect 6914 12832 6920 12844
rect 6875 12804 6920 12832
rect 6914 12792 6920 12804
rect 6972 12792 6978 12844
rect 7929 12835 7987 12841
rect 7929 12801 7941 12835
rect 7975 12832 7987 12835
rect 9125 12835 9183 12841
rect 7975 12804 8708 12832
rect 7975 12801 7987 12804
rect 7929 12795 7987 12801
rect 106 12724 112 12776
rect 164 12764 170 12776
rect 1397 12767 1455 12773
rect 1397 12764 1409 12767
rect 164 12736 1409 12764
rect 164 12724 170 12736
rect 1397 12733 1409 12736
rect 1443 12764 1455 12767
rect 2314 12764 2320 12776
rect 1443 12736 2320 12764
rect 1443 12733 1455 12736
rect 1397 12727 1455 12733
rect 2314 12724 2320 12736
rect 2372 12724 2378 12776
rect 2682 12764 2688 12776
rect 2643 12736 2688 12764
rect 2682 12724 2688 12736
rect 2740 12724 2746 12776
rect 2958 12764 2964 12776
rect 2919 12736 2964 12764
rect 2958 12724 2964 12736
rect 3016 12724 3022 12776
rect 7742 12724 7748 12776
rect 7800 12764 7806 12776
rect 8202 12764 8208 12776
rect 7800 12736 8208 12764
rect 7800 12724 7806 12736
rect 8202 12724 8208 12736
rect 8260 12764 8266 12776
rect 8680 12773 8708 12804
rect 9125 12801 9137 12835
rect 9171 12832 9183 12835
rect 10105 12832 10133 12872
rect 11790 12860 11796 12912
rect 11848 12900 11854 12912
rect 17494 12900 17500 12912
rect 11848 12872 17500 12900
rect 11848 12860 11854 12872
rect 17494 12860 17500 12872
rect 17552 12860 17558 12912
rect 9171 12804 10133 12832
rect 10689 12835 10747 12841
rect 9171 12801 9183 12804
rect 9125 12795 9183 12801
rect 10689 12801 10701 12835
rect 10735 12832 10747 12835
rect 10962 12832 10968 12844
rect 10735 12804 10968 12832
rect 10735 12801 10747 12804
rect 10689 12795 10747 12801
rect 10962 12792 10968 12804
rect 11020 12792 11026 12844
rect 12802 12832 12808 12844
rect 12763 12804 12808 12832
rect 12802 12792 12808 12804
rect 12860 12792 12866 12844
rect 13906 12832 13912 12844
rect 13867 12804 13912 12832
rect 13906 12792 13912 12804
rect 13964 12792 13970 12844
rect 14366 12832 14372 12844
rect 14327 12804 14372 12832
rect 14366 12792 14372 12804
rect 14424 12792 14430 12844
rect 15010 12832 15016 12844
rect 14971 12804 15016 12832
rect 15010 12792 15016 12804
rect 15068 12792 15074 12844
rect 15933 12835 15991 12841
rect 15933 12801 15945 12835
rect 15979 12832 15991 12835
rect 16390 12832 16396 12844
rect 15979 12804 16396 12832
rect 15979 12801 15991 12804
rect 15933 12795 15991 12801
rect 16390 12792 16396 12804
rect 16448 12792 16454 12844
rect 16577 12835 16635 12841
rect 16577 12801 16589 12835
rect 16623 12832 16635 12835
rect 16758 12832 16764 12844
rect 16623 12804 16764 12832
rect 16623 12801 16635 12804
rect 16577 12795 16635 12801
rect 16758 12792 16764 12804
rect 16816 12792 16822 12844
rect 17788 12832 17816 12931
rect 18230 12860 18236 12912
rect 18288 12900 18294 12912
rect 19429 12903 19487 12909
rect 19429 12900 19441 12903
rect 18288 12872 19441 12900
rect 18288 12860 18294 12872
rect 19429 12869 19441 12872
rect 19475 12869 19487 12903
rect 19429 12863 19487 12869
rect 17788 12804 18552 12832
rect 8389 12767 8447 12773
rect 8389 12764 8401 12767
rect 8260 12736 8401 12764
rect 8260 12724 8266 12736
rect 8389 12733 8401 12736
rect 8435 12733 8447 12767
rect 8389 12727 8447 12733
rect 8481 12767 8539 12773
rect 8481 12733 8493 12767
rect 8527 12733 8539 12767
rect 8481 12727 8539 12733
rect 8665 12767 8723 12773
rect 8665 12733 8677 12767
rect 8711 12764 8723 12767
rect 9582 12764 9588 12776
rect 8711 12736 9588 12764
rect 8711 12733 8723 12736
rect 8665 12727 8723 12733
rect 2225 12699 2283 12705
rect 2225 12665 2237 12699
rect 2271 12696 2283 12699
rect 2406 12696 2412 12708
rect 2271 12668 2412 12696
rect 2271 12665 2283 12668
rect 2225 12659 2283 12665
rect 2406 12656 2412 12668
rect 2464 12696 2470 12708
rect 2976 12696 3004 12724
rect 2464 12668 3004 12696
rect 2464 12656 2470 12668
rect 3142 12656 3148 12708
rect 3200 12696 3206 12708
rect 3421 12699 3479 12705
rect 3421 12696 3433 12699
rect 3200 12668 3433 12696
rect 3200 12656 3206 12668
rect 3421 12665 3433 12668
rect 3467 12696 3479 12699
rect 3510 12696 3516 12708
rect 3467 12668 3516 12696
rect 3467 12665 3479 12668
rect 3421 12659 3479 12665
rect 3510 12656 3516 12668
rect 3568 12656 3574 12708
rect 3786 12656 3792 12708
rect 3844 12696 3850 12708
rect 5074 12696 5080 12708
rect 3844 12668 5080 12696
rect 3844 12656 3850 12668
rect 5074 12656 5080 12668
rect 5132 12656 5138 12708
rect 5353 12699 5411 12705
rect 5353 12665 5365 12699
rect 5399 12665 5411 12699
rect 5902 12696 5908 12708
rect 5863 12668 5908 12696
rect 5353 12659 5411 12665
rect 14 12588 20 12640
rect 72 12628 78 12640
rect 1581 12631 1639 12637
rect 1581 12628 1593 12631
rect 72 12600 1593 12628
rect 72 12588 78 12600
rect 1581 12597 1593 12600
rect 1627 12597 1639 12631
rect 1581 12591 1639 12597
rect 1946 12588 1952 12640
rect 2004 12628 2010 12640
rect 4062 12628 4068 12640
rect 2004 12600 4068 12628
rect 2004 12588 2010 12600
rect 4062 12588 4068 12600
rect 4120 12588 4126 12640
rect 4246 12588 4252 12640
rect 4304 12628 4310 12640
rect 4433 12631 4491 12637
rect 4433 12628 4445 12631
rect 4304 12600 4445 12628
rect 4304 12588 4310 12600
rect 4433 12597 4445 12600
rect 4479 12597 4491 12631
rect 4433 12591 4491 12597
rect 5258 12588 5264 12640
rect 5316 12628 5322 12640
rect 5368 12628 5396 12659
rect 5902 12656 5908 12668
rect 5960 12656 5966 12708
rect 6641 12699 6699 12705
rect 6641 12665 6653 12699
rect 6687 12696 6699 12699
rect 7006 12696 7012 12708
rect 6687 12668 7012 12696
rect 6687 12665 6699 12668
rect 6641 12659 6699 12665
rect 7006 12656 7012 12668
rect 7064 12656 7070 12708
rect 6270 12628 6276 12640
rect 5316 12600 6276 12628
rect 5316 12588 5322 12600
rect 6270 12588 6276 12600
rect 6328 12588 6334 12640
rect 8297 12631 8355 12637
rect 8297 12597 8309 12631
rect 8343 12628 8355 12631
rect 8496 12628 8524 12727
rect 9582 12724 9588 12736
rect 9640 12724 9646 12776
rect 11606 12724 11612 12776
rect 11664 12764 11670 12776
rect 11882 12764 11888 12776
rect 11664 12736 11888 12764
rect 11664 12724 11670 12736
rect 11882 12724 11888 12736
rect 11940 12724 11946 12776
rect 18046 12764 18052 12776
rect 18007 12736 18052 12764
rect 18046 12724 18052 12736
rect 18104 12724 18110 12776
rect 18524 12773 18552 12804
rect 18966 12792 18972 12844
rect 19024 12832 19030 12844
rect 19024 12804 19707 12832
rect 19024 12792 19030 12804
rect 18509 12767 18567 12773
rect 18509 12733 18521 12767
rect 18555 12764 18567 12767
rect 18874 12764 18880 12776
rect 18555 12736 18880 12764
rect 18555 12733 18567 12736
rect 18509 12727 18567 12733
rect 18874 12724 18880 12736
rect 18932 12764 18938 12776
rect 19679 12773 19707 12804
rect 19061 12767 19119 12773
rect 19061 12764 19073 12767
rect 18932 12736 19073 12764
rect 18932 12724 18938 12736
rect 19061 12733 19073 12736
rect 19107 12733 19119 12767
rect 19061 12727 19119 12733
rect 19664 12767 19722 12773
rect 19664 12733 19676 12767
rect 19710 12764 19722 12767
rect 19710 12736 20116 12764
rect 19710 12733 19722 12736
rect 19664 12727 19722 12733
rect 10781 12699 10839 12705
rect 10781 12665 10793 12699
rect 10827 12665 10839 12699
rect 10781 12659 10839 12665
rect 11333 12699 11391 12705
rect 11333 12665 11345 12699
rect 11379 12696 11391 12699
rect 11698 12696 11704 12708
rect 11379 12668 11704 12696
rect 11379 12665 11391 12668
rect 11333 12659 11391 12665
rect 8662 12628 8668 12640
rect 8343 12600 8668 12628
rect 8343 12597 8355 12600
rect 8297 12591 8355 12597
rect 8662 12588 8668 12600
rect 8720 12588 8726 12640
rect 9674 12628 9680 12640
rect 9635 12600 9680 12628
rect 9674 12588 9680 12600
rect 9732 12588 9738 12640
rect 10502 12628 10508 12640
rect 10463 12600 10508 12628
rect 10502 12588 10508 12600
rect 10560 12628 10566 12640
rect 10796 12628 10824 12659
rect 11698 12656 11704 12668
rect 11756 12696 11762 12708
rect 12066 12696 12072 12708
rect 11756 12668 12072 12696
rect 11756 12656 11762 12668
rect 12066 12656 12072 12668
rect 12124 12656 12130 12708
rect 12526 12696 12532 12708
rect 12487 12668 12532 12696
rect 12526 12656 12532 12668
rect 12584 12656 12590 12708
rect 12621 12699 12679 12705
rect 12621 12665 12633 12699
rect 12667 12665 12679 12699
rect 14458 12696 14464 12708
rect 14419 12668 14464 12696
rect 12621 12659 12679 12665
rect 10560 12600 10824 12628
rect 10560 12588 10566 12600
rect 11882 12588 11888 12640
rect 11940 12628 11946 12640
rect 12161 12631 12219 12637
rect 12161 12628 12173 12631
rect 11940 12600 12173 12628
rect 11940 12588 11946 12600
rect 12161 12597 12173 12600
rect 12207 12628 12219 12631
rect 12636 12628 12664 12659
rect 14458 12656 14464 12668
rect 14516 12656 14522 12708
rect 15749 12699 15807 12705
rect 15749 12665 15761 12699
rect 15795 12696 15807 12699
rect 16022 12696 16028 12708
rect 15795 12668 16028 12696
rect 15795 12665 15807 12668
rect 15749 12659 15807 12665
rect 16022 12656 16028 12668
rect 16080 12656 16086 12708
rect 18414 12656 18420 12708
rect 18472 12696 18478 12708
rect 19751 12699 19809 12705
rect 19751 12696 19763 12699
rect 18472 12668 19763 12696
rect 18472 12656 18478 12668
rect 19751 12665 19763 12668
rect 19797 12665 19809 12699
rect 19751 12659 19809 12665
rect 20088 12640 20116 12736
rect 12207 12600 12664 12628
rect 15197 12631 15255 12637
rect 12207 12597 12219 12600
rect 12161 12591 12219 12597
rect 15197 12597 15209 12631
rect 15243 12628 15255 12631
rect 16853 12631 16911 12637
rect 16853 12628 16865 12631
rect 15243 12600 16865 12628
rect 15243 12597 15255 12600
rect 15197 12591 15255 12597
rect 16853 12597 16865 12600
rect 16899 12628 16911 12631
rect 17034 12628 17040 12640
rect 16899 12600 17040 12628
rect 16899 12597 16911 12600
rect 16853 12591 16911 12597
rect 17034 12588 17040 12600
rect 17092 12588 17098 12640
rect 17310 12628 17316 12640
rect 17271 12600 17316 12628
rect 17310 12588 17316 12600
rect 17368 12588 17374 12640
rect 18138 12628 18144 12640
rect 18099 12600 18144 12628
rect 18138 12588 18144 12600
rect 18196 12588 18202 12640
rect 20070 12628 20076 12640
rect 20031 12600 20076 12628
rect 20070 12588 20076 12600
rect 20128 12588 20134 12640
rect 1104 12538 20884 12560
rect 1104 12486 8315 12538
rect 8367 12486 8379 12538
rect 8431 12486 8443 12538
rect 8495 12486 8507 12538
rect 8559 12486 15648 12538
rect 15700 12486 15712 12538
rect 15764 12486 15776 12538
rect 15828 12486 15840 12538
rect 15892 12486 20884 12538
rect 1104 12464 20884 12486
rect 2774 12384 2780 12436
rect 2832 12424 2838 12436
rect 3145 12427 3203 12433
rect 3145 12424 3157 12427
rect 2832 12396 3157 12424
rect 2832 12384 2838 12396
rect 3145 12393 3157 12396
rect 3191 12393 3203 12427
rect 3145 12387 3203 12393
rect 3326 12384 3332 12436
rect 3384 12424 3390 12436
rect 3513 12427 3571 12433
rect 3513 12424 3525 12427
rect 3384 12396 3525 12424
rect 3384 12384 3390 12396
rect 3513 12393 3525 12396
rect 3559 12393 3571 12427
rect 5258 12424 5264 12436
rect 5219 12396 5264 12424
rect 3513 12387 3571 12393
rect 5258 12384 5264 12396
rect 5316 12384 5322 12436
rect 5534 12424 5540 12436
rect 5495 12396 5540 12424
rect 5534 12384 5540 12396
rect 5592 12384 5598 12436
rect 6914 12384 6920 12436
rect 6972 12424 6978 12436
rect 7285 12427 7343 12433
rect 7285 12424 7297 12427
rect 6972 12396 7297 12424
rect 6972 12384 6978 12396
rect 7285 12393 7297 12396
rect 7331 12393 7343 12427
rect 7285 12387 7343 12393
rect 7466 12384 7472 12436
rect 7524 12424 7530 12436
rect 8202 12424 8208 12436
rect 7524 12396 8208 12424
rect 7524 12384 7530 12396
rect 8202 12384 8208 12396
rect 8260 12424 8266 12436
rect 8849 12427 8907 12433
rect 8849 12424 8861 12427
rect 8260 12396 8861 12424
rect 8260 12384 8266 12396
rect 8849 12393 8861 12396
rect 8895 12393 8907 12427
rect 8849 12387 8907 12393
rect 10873 12427 10931 12433
rect 10873 12393 10885 12427
rect 10919 12424 10931 12427
rect 11514 12424 11520 12436
rect 10919 12396 11370 12424
rect 11475 12396 11520 12424
rect 10919 12393 10931 12396
rect 10873 12387 10931 12393
rect 2866 12356 2872 12368
rect 2827 12328 2872 12356
rect 2866 12316 2872 12328
rect 2924 12316 2930 12368
rect 1670 12288 1676 12300
rect 1631 12260 1676 12288
rect 1670 12248 1676 12260
rect 1728 12248 1734 12300
rect 2130 12288 2136 12300
rect 2091 12260 2136 12288
rect 2130 12248 2136 12260
rect 2188 12248 2194 12300
rect 2406 12288 2412 12300
rect 2367 12260 2412 12288
rect 2406 12248 2412 12260
rect 2464 12248 2470 12300
rect 2777 12291 2835 12297
rect 2777 12257 2789 12291
rect 2823 12288 2835 12291
rect 3344 12288 3372 12384
rect 5718 12316 5724 12368
rect 5776 12356 5782 12368
rect 6042 12359 6100 12365
rect 6042 12356 6054 12359
rect 5776 12328 6054 12356
rect 5776 12316 5782 12328
rect 6042 12325 6054 12328
rect 6088 12356 6100 12359
rect 6270 12356 6276 12368
rect 6088 12328 6276 12356
rect 6088 12325 6100 12328
rect 6042 12319 6100 12325
rect 6270 12316 6276 12328
rect 6328 12316 6334 12368
rect 7006 12356 7012 12368
rect 6656 12328 7012 12356
rect 2823 12260 3372 12288
rect 2823 12257 2835 12260
rect 2777 12251 2835 12257
rect 3510 12248 3516 12300
rect 3568 12288 3574 12300
rect 4430 12288 4436 12300
rect 3568 12260 4436 12288
rect 3568 12248 3574 12260
rect 4430 12248 4436 12260
rect 4488 12248 4494 12300
rect 4709 12291 4767 12297
rect 4709 12257 4721 12291
rect 4755 12288 4767 12291
rect 5074 12288 5080 12300
rect 4755 12260 5080 12288
rect 4755 12257 4767 12260
rect 4709 12251 4767 12257
rect 5074 12248 5080 12260
rect 5132 12248 5138 12300
rect 6656 12297 6684 12328
rect 7006 12316 7012 12328
rect 7064 12356 7070 12368
rect 7653 12359 7711 12365
rect 7653 12356 7665 12359
rect 7064 12328 7665 12356
rect 7064 12316 7070 12328
rect 7653 12325 7665 12328
rect 7699 12356 7711 12359
rect 7834 12356 7840 12368
rect 7699 12328 7840 12356
rect 7699 12325 7711 12328
rect 7653 12319 7711 12325
rect 7834 12316 7840 12328
rect 7892 12316 7898 12368
rect 7926 12316 7932 12368
rect 7984 12356 7990 12368
rect 8481 12359 8539 12365
rect 8481 12356 8493 12359
rect 7984 12328 8493 12356
rect 7984 12316 7990 12328
rect 8481 12325 8493 12328
rect 8527 12325 8539 12359
rect 8481 12319 8539 12325
rect 6641 12291 6699 12297
rect 6641 12257 6653 12291
rect 6687 12257 6699 12291
rect 6641 12251 6699 12257
rect 4893 12223 4951 12229
rect 4893 12189 4905 12223
rect 4939 12220 4951 12223
rect 5718 12220 5724 12232
rect 4939 12192 5724 12220
rect 4939 12189 4951 12192
rect 4893 12183 4951 12189
rect 5718 12180 5724 12192
rect 5776 12180 5782 12232
rect 7561 12223 7619 12229
rect 7561 12189 7573 12223
rect 7607 12220 7619 12223
rect 8202 12220 8208 12232
rect 7607 12192 8208 12220
rect 7607 12189 7619 12192
rect 7561 12183 7619 12189
rect 8202 12180 8208 12192
rect 8260 12180 8266 12232
rect 8496 12220 8524 12319
rect 9674 12316 9680 12368
rect 9732 12356 9738 12368
rect 10274 12359 10332 12365
rect 10274 12356 10286 12359
rect 9732 12328 10286 12356
rect 9732 12316 9738 12328
rect 10274 12325 10286 12328
rect 10320 12325 10332 12359
rect 11342 12356 11370 12396
rect 11514 12384 11520 12396
rect 11572 12384 11578 12436
rect 13357 12427 13415 12433
rect 13357 12393 13369 12427
rect 13403 12424 13415 12427
rect 13538 12424 13544 12436
rect 13403 12396 13544 12424
rect 13403 12393 13415 12396
rect 13357 12387 13415 12393
rect 13538 12384 13544 12396
rect 13596 12384 13602 12436
rect 14458 12384 14464 12436
rect 14516 12424 14522 12436
rect 14645 12427 14703 12433
rect 14645 12424 14657 12427
rect 14516 12396 14657 12424
rect 14516 12384 14522 12396
rect 14645 12393 14657 12396
rect 14691 12393 14703 12427
rect 14645 12387 14703 12393
rect 15105 12427 15163 12433
rect 15105 12393 15117 12427
rect 15151 12424 15163 12427
rect 15194 12424 15200 12436
rect 15151 12396 15200 12424
rect 15151 12393 15163 12396
rect 15105 12387 15163 12393
rect 15194 12384 15200 12396
rect 15252 12384 15258 12436
rect 15286 12384 15292 12436
rect 15344 12424 15350 12436
rect 16393 12427 16451 12433
rect 15344 12396 15424 12424
rect 15344 12384 15350 12396
rect 11882 12356 11888 12368
rect 11342 12328 11888 12356
rect 10274 12319 10332 12325
rect 11882 12316 11888 12328
rect 11940 12316 11946 12368
rect 13811 12359 13869 12365
rect 13811 12325 13823 12359
rect 13857 12356 13869 12359
rect 14090 12356 14096 12368
rect 13857 12328 14096 12356
rect 13857 12325 13869 12328
rect 13811 12319 13869 12325
rect 14090 12316 14096 12328
rect 14148 12316 14154 12368
rect 15396 12365 15424 12396
rect 16393 12393 16405 12427
rect 16439 12424 16451 12427
rect 16482 12424 16488 12436
rect 16439 12396 16488 12424
rect 16439 12393 16451 12396
rect 16393 12387 16451 12393
rect 16482 12384 16488 12396
rect 16540 12384 16546 12436
rect 16574 12384 16580 12436
rect 16632 12424 16638 12436
rect 16945 12427 17003 12433
rect 16945 12424 16957 12427
rect 16632 12396 16957 12424
rect 16632 12384 16638 12396
rect 16945 12393 16957 12396
rect 16991 12393 17003 12427
rect 18046 12424 18052 12436
rect 18007 12396 18052 12424
rect 16945 12387 17003 12393
rect 18046 12384 18052 12396
rect 18104 12384 18110 12436
rect 18506 12424 18512 12436
rect 18467 12396 18512 12424
rect 18506 12384 18512 12396
rect 18564 12384 18570 12436
rect 15381 12359 15439 12365
rect 15381 12325 15393 12359
rect 15427 12325 15439 12359
rect 15381 12319 15439 12325
rect 15473 12359 15531 12365
rect 15473 12325 15485 12359
rect 15519 12356 15531 12359
rect 16022 12356 16028 12368
rect 15519 12328 16028 12356
rect 15519 12325 15531 12328
rect 15473 12319 15531 12325
rect 16022 12316 16028 12328
rect 16080 12316 16086 12368
rect 17052 12328 18460 12356
rect 17052 12300 17080 12328
rect 9950 12288 9956 12300
rect 9911 12260 9956 12288
rect 9950 12248 9956 12260
rect 10008 12248 10014 12300
rect 17034 12288 17040 12300
rect 16995 12260 17040 12288
rect 17034 12248 17040 12260
rect 17092 12248 17098 12300
rect 17405 12291 17463 12297
rect 17405 12257 17417 12291
rect 17451 12288 17463 12291
rect 17494 12288 17500 12300
rect 17451 12260 17500 12288
rect 17451 12257 17463 12260
rect 17405 12251 17463 12257
rect 17494 12248 17500 12260
rect 17552 12248 17558 12300
rect 18432 12297 18460 12328
rect 18417 12291 18475 12297
rect 18417 12257 18429 12291
rect 18463 12288 18475 12291
rect 18690 12288 18696 12300
rect 18463 12260 18696 12288
rect 18463 12257 18475 12260
rect 18417 12251 18475 12257
rect 18690 12248 18696 12260
rect 18748 12248 18754 12300
rect 18874 12288 18880 12300
rect 18835 12260 18880 12288
rect 18874 12248 18880 12260
rect 18932 12248 18938 12300
rect 11606 12220 11612 12232
rect 8496 12192 11612 12220
rect 11606 12180 11612 12192
rect 11664 12180 11670 12232
rect 11790 12220 11796 12232
rect 11751 12192 11796 12220
rect 11790 12180 11796 12192
rect 11848 12180 11854 12232
rect 12066 12220 12072 12232
rect 12027 12192 12072 12220
rect 12066 12180 12072 12192
rect 12124 12180 12130 12232
rect 13449 12223 13507 12229
rect 13449 12189 13461 12223
rect 13495 12220 13507 12223
rect 14550 12220 14556 12232
rect 13495 12192 14556 12220
rect 13495 12189 13507 12192
rect 13449 12183 13507 12189
rect 14550 12180 14556 12192
rect 14608 12180 14614 12232
rect 15470 12180 15476 12232
rect 15528 12220 15534 12232
rect 15657 12223 15715 12229
rect 15657 12220 15669 12223
rect 15528 12192 15669 12220
rect 15528 12180 15534 12192
rect 15657 12189 15669 12192
rect 15703 12189 15715 12223
rect 15657 12183 15715 12189
rect 5902 12112 5908 12164
rect 5960 12152 5966 12164
rect 8113 12155 8171 12161
rect 8113 12152 8125 12155
rect 5960 12124 8125 12152
rect 5960 12112 5966 12124
rect 7576 12096 7604 12124
rect 8113 12121 8125 12124
rect 8159 12121 8171 12155
rect 8113 12115 8171 12121
rect 12526 12112 12532 12164
rect 12584 12152 12590 12164
rect 12805 12155 12863 12161
rect 12805 12152 12817 12155
rect 12584 12124 12817 12152
rect 12584 12112 12590 12124
rect 12805 12121 12817 12124
rect 12851 12152 12863 12155
rect 14369 12155 14427 12161
rect 12851 12124 13814 12152
rect 12851 12121 12863 12124
rect 12805 12115 12863 12121
rect 7006 12084 7012 12096
rect 6967 12056 7012 12084
rect 7006 12044 7012 12056
rect 7064 12044 7070 12096
rect 7558 12044 7564 12096
rect 7616 12044 7622 12096
rect 9214 12044 9220 12096
rect 9272 12084 9278 12096
rect 12618 12084 12624 12096
rect 9272 12056 12624 12084
rect 9272 12044 9278 12056
rect 12618 12044 12624 12056
rect 12676 12044 12682 12096
rect 13786 12084 13814 12124
rect 14369 12121 14381 12155
rect 14415 12152 14427 12155
rect 16022 12152 16028 12164
rect 14415 12124 16028 12152
rect 14415 12121 14427 12124
rect 14369 12115 14427 12121
rect 16022 12112 16028 12124
rect 16080 12112 16086 12164
rect 14918 12084 14924 12096
rect 13786 12056 14924 12084
rect 14918 12044 14924 12056
rect 14976 12044 14982 12096
rect 1104 11994 20884 12016
rect 1104 11942 4648 11994
rect 4700 11942 4712 11994
rect 4764 11942 4776 11994
rect 4828 11942 4840 11994
rect 4892 11942 11982 11994
rect 12034 11942 12046 11994
rect 12098 11942 12110 11994
rect 12162 11942 12174 11994
rect 12226 11942 19315 11994
rect 19367 11942 19379 11994
rect 19431 11942 19443 11994
rect 19495 11942 19507 11994
rect 19559 11942 20884 11994
rect 1104 11920 20884 11942
rect 106 11840 112 11892
rect 164 11880 170 11892
rect 164 11852 4251 11880
rect 164 11840 170 11852
rect 4223 11812 4251 11852
rect 4430 11840 4436 11892
rect 4488 11880 4494 11892
rect 5353 11883 5411 11889
rect 5353 11880 5365 11883
rect 4488 11852 5365 11880
rect 4488 11840 4494 11852
rect 5353 11849 5365 11852
rect 5399 11849 5411 11883
rect 5353 11843 5411 11849
rect 6270 11840 6276 11892
rect 6328 11880 6334 11892
rect 6457 11883 6515 11889
rect 6457 11880 6469 11883
rect 6328 11852 6469 11880
rect 6328 11840 6334 11852
rect 6457 11849 6469 11852
rect 6503 11849 6515 11883
rect 7834 11880 7840 11892
rect 7795 11852 7840 11880
rect 6457 11843 6515 11849
rect 5721 11815 5779 11821
rect 5721 11812 5733 11815
rect 4223 11784 5733 11812
rect 5721 11781 5733 11784
rect 5767 11781 5779 11815
rect 6086 11812 6092 11824
rect 6047 11784 6092 11812
rect 5721 11775 5779 11781
rect 6086 11772 6092 11784
rect 6144 11772 6150 11824
rect 6472 11812 6500 11843
rect 7834 11840 7840 11852
rect 7892 11840 7898 11892
rect 8202 11880 8208 11892
rect 8163 11852 8208 11880
rect 8202 11840 8208 11852
rect 8260 11880 8266 11892
rect 8527 11883 8585 11889
rect 8527 11880 8539 11883
rect 8260 11852 8539 11880
rect 8260 11840 8266 11852
rect 8527 11849 8539 11852
rect 8573 11849 8585 11883
rect 8527 11843 8585 11849
rect 9950 11840 9956 11892
rect 10008 11880 10014 11892
rect 11149 11883 11207 11889
rect 11149 11880 11161 11883
rect 10008 11852 11161 11880
rect 10008 11840 10014 11852
rect 11149 11849 11161 11852
rect 11195 11849 11207 11883
rect 11149 11843 11207 11849
rect 11330 11840 11336 11892
rect 11388 11880 11394 11892
rect 11793 11883 11851 11889
rect 11793 11880 11805 11883
rect 11388 11852 11805 11880
rect 11388 11840 11411 11852
rect 11793 11849 11805 11852
rect 11839 11849 11851 11883
rect 11793 11843 11851 11849
rect 12342 11840 12348 11892
rect 12400 11880 12406 11892
rect 12805 11883 12863 11889
rect 12805 11880 12817 11883
rect 12400 11852 12817 11880
rect 12400 11840 12406 11852
rect 12805 11849 12817 11852
rect 12851 11880 12863 11883
rect 13081 11883 13139 11889
rect 13081 11880 13093 11883
rect 12851 11852 13093 11880
rect 12851 11849 12863 11852
rect 12805 11843 12863 11849
rect 13081 11849 13093 11852
rect 13127 11880 13139 11883
rect 14090 11880 14096 11892
rect 13127 11852 14096 11880
rect 13127 11849 13139 11852
rect 13081 11843 13139 11849
rect 14090 11840 14096 11852
rect 14148 11840 14154 11892
rect 14185 11883 14243 11889
rect 14185 11849 14197 11883
rect 14231 11880 14243 11883
rect 14458 11880 14464 11892
rect 14231 11852 14464 11880
rect 14231 11849 14243 11852
rect 14185 11843 14243 11849
rect 14458 11840 14464 11852
rect 14516 11880 14522 11892
rect 14829 11883 14887 11889
rect 14829 11880 14841 11883
rect 14516 11852 14841 11880
rect 14516 11840 14522 11852
rect 14829 11849 14841 11852
rect 14875 11849 14887 11883
rect 16022 11880 16028 11892
rect 15983 11852 16028 11880
rect 14829 11843 14887 11849
rect 9401 11815 9459 11821
rect 9401 11812 9413 11815
rect 6472 11784 9413 11812
rect 9401 11781 9413 11784
rect 9447 11812 9459 11815
rect 9674 11812 9680 11824
rect 9447 11784 9680 11812
rect 9447 11781 9459 11784
rect 9401 11775 9459 11781
rect 9674 11772 9680 11784
rect 9732 11772 9738 11824
rect 2869 11747 2927 11753
rect 2869 11713 2881 11747
rect 2915 11744 2927 11747
rect 3050 11744 3056 11756
rect 2915 11716 3056 11744
rect 2915 11713 2927 11716
rect 2869 11707 2927 11713
rect 3050 11704 3056 11716
rect 3108 11704 3114 11756
rect 3418 11704 3424 11756
rect 3476 11744 3482 11756
rect 3605 11747 3663 11753
rect 3605 11744 3617 11747
rect 3476 11716 3617 11744
rect 3476 11704 3482 11716
rect 3605 11713 3617 11716
rect 3651 11744 3663 11747
rect 4798 11744 4804 11756
rect 3651 11716 4804 11744
rect 3651 11713 3663 11716
rect 3605 11707 3663 11713
rect 4798 11704 4804 11716
rect 4856 11704 4862 11756
rect 1670 11676 1676 11688
rect 1583 11648 1676 11676
rect 1670 11636 1676 11648
rect 1728 11676 1734 11688
rect 2130 11676 2136 11688
rect 1728 11648 1992 11676
rect 2091 11648 2136 11676
rect 1728 11636 1734 11648
rect 1964 11540 1992 11648
rect 2130 11636 2136 11648
rect 2188 11636 2194 11688
rect 2406 11676 2412 11688
rect 2319 11648 2412 11676
rect 2406 11636 2412 11648
rect 2464 11636 2470 11688
rect 2682 11676 2688 11688
rect 2643 11648 2688 11676
rect 2682 11636 2688 11648
rect 2740 11636 2746 11688
rect 3326 11636 3332 11688
rect 3384 11676 3390 11688
rect 3878 11676 3884 11688
rect 3384 11648 3884 11676
rect 3384 11636 3390 11648
rect 3878 11636 3884 11648
rect 3936 11636 3942 11688
rect 5537 11679 5595 11685
rect 5537 11645 5549 11679
rect 5583 11676 5595 11679
rect 5626 11676 5632 11688
rect 5583 11648 5632 11676
rect 5583 11645 5595 11648
rect 5537 11639 5595 11645
rect 5626 11636 5632 11648
rect 5684 11676 5690 11688
rect 6104 11676 6132 11772
rect 6546 11704 6552 11756
rect 6604 11744 6610 11756
rect 6917 11747 6975 11753
rect 6917 11744 6929 11747
rect 6604 11716 6929 11744
rect 6604 11704 6610 11716
rect 6917 11713 6929 11716
rect 6963 11744 6975 11747
rect 7098 11744 7104 11756
rect 6963 11716 7104 11744
rect 6963 11713 6975 11716
rect 6917 11707 6975 11713
rect 7098 11704 7104 11716
rect 7156 11704 7162 11756
rect 5684 11648 6132 11676
rect 8456 11679 8514 11685
rect 5684 11636 5690 11648
rect 8456 11645 8468 11679
rect 8502 11676 8514 11679
rect 8502 11648 8984 11676
rect 8502 11645 8514 11648
rect 8456 11639 8514 11645
rect 2424 11608 2452 11636
rect 3418 11608 3424 11620
rect 2424 11580 3424 11608
rect 3418 11568 3424 11580
rect 3476 11568 3482 11620
rect 4062 11608 4068 11620
rect 4023 11580 4068 11608
rect 4062 11568 4068 11580
rect 4120 11568 4126 11620
rect 4157 11611 4215 11617
rect 4157 11577 4169 11611
rect 4203 11608 4215 11611
rect 4246 11608 4252 11620
rect 4203 11580 4252 11608
rect 4203 11577 4215 11580
rect 4157 11571 4215 11577
rect 4246 11568 4252 11580
rect 4304 11568 4310 11620
rect 4709 11611 4767 11617
rect 4709 11577 4721 11611
rect 4755 11608 4767 11611
rect 4755 11580 6592 11608
rect 4755 11577 4767 11580
rect 4709 11571 4767 11577
rect 3237 11543 3295 11549
rect 3237 11540 3249 11543
rect 1964 11512 3249 11540
rect 3237 11509 3249 11512
rect 3283 11540 3295 11543
rect 3694 11540 3700 11552
rect 3283 11512 3700 11540
rect 3283 11509 3295 11512
rect 3237 11503 3295 11509
rect 3694 11500 3700 11512
rect 3752 11500 3758 11552
rect 5074 11540 5080 11552
rect 5035 11512 5080 11540
rect 5074 11500 5080 11512
rect 5132 11500 5138 11552
rect 6564 11540 6592 11580
rect 7006 11568 7012 11620
rect 7064 11608 7070 11620
rect 7561 11611 7619 11617
rect 7561 11608 7573 11611
rect 7064 11580 7109 11608
rect 7392 11580 7573 11608
rect 7064 11568 7070 11580
rect 6914 11540 6920 11552
rect 6564 11512 6920 11540
rect 6914 11500 6920 11512
rect 6972 11540 6978 11552
rect 7392 11540 7420 11580
rect 7561 11577 7573 11580
rect 7607 11577 7619 11611
rect 7561 11571 7619 11577
rect 8956 11549 8984 11648
rect 9490 11636 9496 11688
rect 9548 11676 9554 11688
rect 9585 11679 9643 11685
rect 9585 11676 9597 11679
rect 9548 11648 9597 11676
rect 9548 11636 9554 11648
rect 9585 11645 9597 11648
rect 9631 11645 9643 11679
rect 10781 11679 10839 11685
rect 10781 11676 10793 11679
rect 9585 11639 9643 11645
rect 9968 11648 10793 11676
rect 9968 11620 9996 11648
rect 10781 11645 10793 11648
rect 10827 11645 10839 11679
rect 10781 11639 10839 11645
rect 10962 11636 10968 11688
rect 11020 11676 11026 11688
rect 11146 11676 11152 11688
rect 11020 11648 11152 11676
rect 11020 11636 11026 11648
rect 11146 11636 11152 11648
rect 11204 11636 11210 11688
rect 11383 11685 11411 11840
rect 11882 11772 11888 11824
rect 11940 11812 11946 11824
rect 12161 11815 12219 11821
rect 12161 11812 12173 11815
rect 11940 11784 12173 11812
rect 11940 11772 11946 11784
rect 12161 11781 12173 11784
rect 12207 11781 12219 11815
rect 12161 11775 12219 11781
rect 13265 11747 13323 11753
rect 13265 11713 13277 11747
rect 13311 11744 13323 11747
rect 13538 11744 13544 11756
rect 13311 11716 13544 11744
rect 13311 11713 13323 11716
rect 13265 11707 13323 11713
rect 13538 11704 13544 11716
rect 13596 11704 13602 11756
rect 11368 11679 11426 11685
rect 11368 11645 11380 11679
rect 11414 11645 11426 11679
rect 11368 11639 11426 11645
rect 11471 11679 11529 11685
rect 11471 11645 11483 11679
rect 11517 11676 11529 11679
rect 13078 11676 13084 11688
rect 11517 11648 13084 11676
rect 11517 11645 11529 11648
rect 11471 11639 11529 11645
rect 13078 11636 13084 11648
rect 13136 11636 13142 11688
rect 13446 11636 13452 11688
rect 13504 11676 13510 11688
rect 14182 11676 14188 11688
rect 13504 11648 14188 11676
rect 13504 11636 13510 11648
rect 14182 11636 14188 11648
rect 14240 11636 14246 11688
rect 9674 11568 9680 11620
rect 9732 11608 9738 11620
rect 9950 11617 9956 11620
rect 9906 11611 9956 11617
rect 9906 11608 9918 11611
rect 9732 11580 9918 11608
rect 9732 11568 9738 11580
rect 9906 11577 9918 11580
rect 9952 11577 9956 11611
rect 9906 11571 9956 11577
rect 9950 11568 9956 11571
rect 10008 11568 10014 11620
rect 10134 11568 10140 11620
rect 10192 11608 10198 11620
rect 13354 11608 13360 11620
rect 10192 11580 13360 11608
rect 10192 11568 10198 11580
rect 13354 11568 13360 11580
rect 13412 11568 13418 11620
rect 13627 11611 13685 11617
rect 13627 11577 13639 11611
rect 13673 11608 13685 11611
rect 14090 11608 14096 11620
rect 13673 11580 14096 11608
rect 13673 11577 13685 11580
rect 13627 11571 13685 11577
rect 14090 11568 14096 11580
rect 14148 11568 14154 11620
rect 14844 11608 14872 11843
rect 16022 11840 16028 11852
rect 16080 11840 16086 11892
rect 16298 11840 16304 11892
rect 16356 11880 16362 11892
rect 21634 11880 21640 11892
rect 16356 11852 21640 11880
rect 16356 11840 16362 11852
rect 21634 11840 21640 11852
rect 21692 11840 21698 11892
rect 14918 11772 14924 11824
rect 14976 11812 14982 11824
rect 19751 11815 19809 11821
rect 19751 11812 19763 11815
rect 14976 11784 19763 11812
rect 14976 11772 14982 11784
rect 19751 11781 19763 11784
rect 19797 11781 19809 11815
rect 19751 11775 19809 11781
rect 15102 11744 15108 11756
rect 15063 11716 15108 11744
rect 15102 11704 15108 11716
rect 15160 11704 15166 11756
rect 15470 11744 15476 11756
rect 15431 11716 15476 11744
rect 15470 11704 15476 11716
rect 15528 11704 15534 11756
rect 17402 11704 17408 11756
rect 17460 11744 17466 11756
rect 17460 11716 19691 11744
rect 17460 11704 17466 11716
rect 16644 11679 16702 11685
rect 16644 11645 16656 11679
rect 16690 11676 16702 11679
rect 17494 11676 17500 11688
rect 16690 11648 17172 11676
rect 17407 11648 17500 11676
rect 16690 11645 16702 11648
rect 16644 11639 16702 11645
rect 15197 11611 15255 11617
rect 15197 11608 15209 11611
rect 14844 11580 15209 11608
rect 15197 11577 15209 11580
rect 15243 11577 15255 11611
rect 15197 11571 15255 11577
rect 16485 11611 16543 11617
rect 16485 11577 16497 11611
rect 16531 11608 16543 11611
rect 17034 11608 17040 11620
rect 16531 11580 17040 11608
rect 16531 11577 16543 11580
rect 16485 11571 16543 11577
rect 6972 11512 7420 11540
rect 8941 11543 8999 11549
rect 6972 11500 6978 11512
rect 8941 11509 8953 11543
rect 8987 11540 8999 11543
rect 9030 11540 9036 11552
rect 8987 11512 9036 11540
rect 8987 11509 8999 11512
rect 8941 11503 8999 11509
rect 9030 11500 9036 11512
rect 9088 11500 9094 11552
rect 10502 11540 10508 11552
rect 10463 11512 10508 11540
rect 10502 11500 10508 11512
rect 10560 11500 10566 11552
rect 14550 11540 14556 11552
rect 14511 11512 14556 11540
rect 14550 11500 14556 11512
rect 14608 11500 14614 11552
rect 14642 11500 14648 11552
rect 14700 11540 14706 11552
rect 16500 11540 16528 11571
rect 17034 11568 17040 11580
rect 17092 11568 17098 11620
rect 14700 11512 16528 11540
rect 16715 11543 16773 11549
rect 14700 11500 14706 11512
rect 16715 11509 16727 11543
rect 16761 11540 16773 11543
rect 16850 11540 16856 11552
rect 16761 11512 16856 11540
rect 16761 11509 16773 11512
rect 16715 11503 16773 11509
rect 16850 11500 16856 11512
rect 16908 11500 16914 11552
rect 17144 11549 17172 11648
rect 17494 11636 17500 11648
rect 17552 11676 17558 11688
rect 17954 11676 17960 11688
rect 17552 11648 17960 11676
rect 17552 11636 17558 11648
rect 17954 11636 17960 11648
rect 18012 11636 18018 11688
rect 18141 11679 18199 11685
rect 18141 11645 18153 11679
rect 18187 11645 18199 11679
rect 18141 11639 18199 11645
rect 17586 11568 17592 11620
rect 17644 11608 17650 11620
rect 18049 11611 18107 11617
rect 18049 11608 18061 11611
rect 17644 11580 18061 11608
rect 17644 11568 17650 11580
rect 18049 11577 18061 11580
rect 18095 11577 18107 11611
rect 18049 11571 18107 11577
rect 17129 11543 17187 11549
rect 17129 11509 17141 11543
rect 17175 11540 17187 11543
rect 17218 11540 17224 11552
rect 17175 11512 17224 11540
rect 17175 11509 17187 11512
rect 17129 11503 17187 11509
rect 17218 11500 17224 11512
rect 17276 11500 17282 11552
rect 17494 11500 17500 11552
rect 17552 11540 17558 11552
rect 17773 11543 17831 11549
rect 17773 11540 17785 11543
rect 17552 11512 17785 11540
rect 17552 11500 17558 11512
rect 17773 11509 17785 11512
rect 17819 11540 17831 11543
rect 18156 11540 18184 11639
rect 18874 11636 18880 11688
rect 18932 11676 18938 11688
rect 19058 11676 19064 11688
rect 18932 11648 19064 11676
rect 18932 11636 18938 11648
rect 19058 11636 19064 11648
rect 19116 11636 19122 11688
rect 19663 11685 19691 11716
rect 19648 11679 19706 11685
rect 19648 11645 19660 11679
rect 19694 11676 19706 11679
rect 20070 11676 20076 11688
rect 19694 11648 20076 11676
rect 19694 11645 19706 11648
rect 19648 11639 19706 11645
rect 20070 11636 20076 11648
rect 20128 11636 20134 11688
rect 17819 11512 18184 11540
rect 17819 11509 17831 11512
rect 17773 11503 17831 11509
rect 1104 11450 20884 11472
rect 1104 11398 8315 11450
rect 8367 11398 8379 11450
rect 8431 11398 8443 11450
rect 8495 11398 8507 11450
rect 8559 11398 15648 11450
rect 15700 11398 15712 11450
rect 15764 11398 15776 11450
rect 15828 11398 15840 11450
rect 15892 11398 20884 11450
rect 1104 11376 20884 11398
rect 1949 11339 2007 11345
rect 1949 11305 1961 11339
rect 1995 11336 2007 11339
rect 2682 11336 2688 11348
rect 1995 11308 2688 11336
rect 1995 11305 2007 11308
rect 1949 11299 2007 11305
rect 2682 11296 2688 11308
rect 2740 11296 2746 11348
rect 3418 11336 3424 11348
rect 3379 11308 3424 11336
rect 3418 11296 3424 11308
rect 3476 11296 3482 11348
rect 3878 11336 3884 11348
rect 3839 11308 3884 11336
rect 3878 11296 3884 11308
rect 3936 11296 3942 11348
rect 4062 11296 4068 11348
rect 4120 11336 4126 11348
rect 5169 11339 5227 11345
rect 5169 11336 5181 11339
rect 4120 11308 5181 11336
rect 4120 11296 4126 11308
rect 5169 11305 5181 11308
rect 5215 11336 5227 11339
rect 5350 11336 5356 11348
rect 5215 11308 5356 11336
rect 5215 11305 5227 11308
rect 5169 11299 5227 11305
rect 5350 11296 5356 11308
rect 5408 11296 5414 11348
rect 5718 11336 5724 11348
rect 5679 11308 5724 11336
rect 5718 11296 5724 11308
rect 5776 11296 5782 11348
rect 6086 11296 6092 11348
rect 6144 11336 6150 11348
rect 6270 11336 6276 11348
rect 6144 11308 6276 11336
rect 6144 11296 6150 11308
rect 6270 11296 6276 11308
rect 6328 11296 6334 11348
rect 6825 11339 6883 11345
rect 6825 11305 6837 11339
rect 6871 11336 6883 11339
rect 7006 11336 7012 11348
rect 6871 11308 7012 11336
rect 6871 11305 6883 11308
rect 6825 11299 6883 11305
rect 7006 11296 7012 11308
rect 7064 11296 7070 11348
rect 7098 11296 7104 11348
rect 7156 11336 7162 11348
rect 7156 11308 7201 11336
rect 7156 11296 7162 11308
rect 8110 11296 8116 11348
rect 8168 11336 8174 11348
rect 8389 11339 8447 11345
rect 8389 11336 8401 11339
rect 8168 11308 8401 11336
rect 8168 11296 8174 11308
rect 8389 11305 8401 11308
rect 8435 11305 8447 11339
rect 10870 11336 10876 11348
rect 8389 11299 8447 11305
rect 8588 11308 10876 11336
rect 3510 11268 3516 11280
rect 2700 11240 3516 11268
rect 2700 11209 2728 11240
rect 3510 11228 3516 11240
rect 3568 11228 3574 11280
rect 4246 11268 4252 11280
rect 4207 11240 4252 11268
rect 4246 11228 4252 11240
rect 4304 11228 4310 11280
rect 7190 11228 7196 11280
rect 7248 11268 7254 11280
rect 7561 11271 7619 11277
rect 7561 11268 7573 11271
rect 7248 11240 7573 11268
rect 7248 11228 7254 11240
rect 7561 11237 7573 11240
rect 7607 11268 7619 11271
rect 8588 11268 8616 11308
rect 10870 11296 10876 11308
rect 10928 11296 10934 11348
rect 11790 11296 11796 11348
rect 11848 11336 11854 11348
rect 12529 11339 12587 11345
rect 12529 11336 12541 11339
rect 11848 11308 12541 11336
rect 11848 11296 11854 11308
rect 12529 11305 12541 11308
rect 12575 11305 12587 11339
rect 13998 11336 14004 11348
rect 12529 11299 12587 11305
rect 13188 11308 14004 11336
rect 7607 11240 8616 11268
rect 9953 11271 10011 11277
rect 7607 11237 7619 11240
rect 7561 11231 7619 11237
rect 9953 11237 9965 11271
rect 9999 11268 10011 11271
rect 10502 11268 10508 11280
rect 9999 11240 10508 11268
rect 9999 11237 10011 11240
rect 9953 11231 10011 11237
rect 10502 11228 10508 11240
rect 10560 11228 10566 11280
rect 11695 11271 11753 11277
rect 11695 11237 11707 11271
rect 11741 11268 11753 11271
rect 12342 11268 12348 11280
rect 11741 11240 12348 11268
rect 11741 11237 11753 11240
rect 11695 11231 11753 11237
rect 12342 11228 12348 11240
rect 12400 11228 12406 11280
rect 13188 11277 13216 11308
rect 13998 11296 14004 11308
rect 14056 11296 14062 11348
rect 15102 11336 15108 11348
rect 15063 11308 15108 11336
rect 15102 11296 15108 11308
rect 15160 11296 15166 11348
rect 15286 11296 15292 11348
rect 15344 11336 15350 11348
rect 15473 11339 15531 11345
rect 15473 11336 15485 11339
rect 15344 11308 15485 11336
rect 15344 11296 15350 11308
rect 15473 11305 15485 11308
rect 15519 11305 15531 11339
rect 15473 11299 15531 11305
rect 16022 11296 16028 11348
rect 16080 11336 16086 11348
rect 17773 11339 17831 11345
rect 17773 11336 17785 11339
rect 16080 11308 17785 11336
rect 16080 11296 16086 11308
rect 17773 11305 17785 11308
rect 17819 11305 17831 11339
rect 18690 11336 18696 11348
rect 18651 11308 18696 11336
rect 17773 11299 17831 11305
rect 18690 11296 18696 11308
rect 18748 11296 18754 11348
rect 19429 11339 19487 11345
rect 19429 11305 19441 11339
rect 19475 11336 19487 11339
rect 19702 11336 19708 11348
rect 19475 11308 19708 11336
rect 19475 11305 19487 11308
rect 19429 11299 19487 11305
rect 19702 11296 19708 11308
rect 19760 11296 19766 11348
rect 12989 11271 13047 11277
rect 12989 11237 13001 11271
rect 13035 11268 13047 11271
rect 13173 11271 13231 11277
rect 13173 11268 13185 11271
rect 13035 11240 13185 11268
rect 13035 11237 13047 11240
rect 12989 11231 13047 11237
rect 13173 11237 13185 11240
rect 13219 11237 13231 11271
rect 13173 11231 13231 11237
rect 13262 11228 13268 11280
rect 13320 11268 13326 11280
rect 16298 11268 16304 11280
rect 13320 11240 13365 11268
rect 16259 11240 16304 11268
rect 13320 11228 13326 11240
rect 16298 11228 16304 11240
rect 16356 11228 16362 11280
rect 17218 11228 17224 11280
rect 17276 11268 17282 11280
rect 18598 11268 18604 11280
rect 17276 11240 18604 11268
rect 17276 11228 17282 11240
rect 18598 11228 18604 11240
rect 18656 11268 18662 11280
rect 18656 11240 19288 11268
rect 18656 11228 18662 11240
rect 1464 11203 1522 11209
rect 1464 11169 1476 11203
rect 1510 11169 1522 11203
rect 1464 11163 1522 11169
rect 2685 11203 2743 11209
rect 2685 11169 2697 11203
rect 2731 11169 2743 11203
rect 2866 11200 2872 11212
rect 2827 11172 2872 11200
rect 2685 11163 2743 11169
rect 1479 11064 1507 11163
rect 2866 11160 2872 11172
rect 2924 11160 2930 11212
rect 4798 11160 4804 11212
rect 4856 11200 4862 11212
rect 7466 11200 7472 11212
rect 4856 11172 7472 11200
rect 4856 11160 4862 11172
rect 7466 11160 7472 11172
rect 7524 11200 7530 11212
rect 7929 11203 7987 11209
rect 7929 11200 7941 11203
rect 7524 11172 7941 11200
rect 7524 11160 7530 11172
rect 7929 11169 7941 11172
rect 7975 11169 7987 11203
rect 8202 11200 8208 11212
rect 8163 11172 8208 11200
rect 7929 11163 7987 11169
rect 8202 11160 8208 11172
rect 8260 11200 8266 11212
rect 8846 11200 8852 11212
rect 8260 11172 8852 11200
rect 8260 11160 8266 11172
rect 8846 11160 8852 11172
rect 8904 11160 8910 11212
rect 17862 11200 17868 11212
rect 17823 11172 17868 11200
rect 17862 11160 17868 11172
rect 17920 11160 17926 11212
rect 17954 11160 17960 11212
rect 18012 11200 18018 11212
rect 18230 11200 18236 11212
rect 18012 11172 18236 11200
rect 18012 11160 18018 11172
rect 18230 11160 18236 11172
rect 18288 11160 18294 11212
rect 19260 11209 19288 11240
rect 19245 11203 19303 11209
rect 19245 11169 19257 11203
rect 19291 11200 19303 11203
rect 19610 11200 19616 11212
rect 19291 11172 19616 11200
rect 19291 11169 19303 11172
rect 19245 11163 19303 11169
rect 19610 11160 19616 11172
rect 19668 11160 19674 11212
rect 3050 11132 3056 11144
rect 3011 11104 3056 11132
rect 3050 11092 3056 11104
rect 3108 11092 3114 11144
rect 4157 11135 4215 11141
rect 4157 11101 4169 11135
rect 4203 11132 4215 11135
rect 4203 11104 4292 11132
rect 4203 11101 4215 11104
rect 4157 11095 4215 11101
rect 4062 11064 4068 11076
rect 1479 11036 4068 11064
rect 4062 11024 4068 11036
rect 4120 11024 4126 11076
rect 106 10956 112 11008
rect 164 10996 170 11008
rect 1535 10999 1593 11005
rect 1535 10996 1547 10999
rect 164 10968 1547 10996
rect 164 10956 170 10968
rect 1535 10965 1547 10968
rect 1581 10965 1593 10999
rect 1535 10959 1593 10965
rect 2317 10999 2375 11005
rect 2317 10965 2329 10999
rect 2363 10996 2375 10999
rect 3694 10996 3700 11008
rect 2363 10968 3700 10996
rect 2363 10965 2375 10968
rect 2317 10959 2375 10965
rect 3694 10956 3700 10968
rect 3752 10956 3758 11008
rect 4264 10996 4292 11104
rect 4338 11092 4344 11144
rect 4396 11132 4402 11144
rect 5905 11135 5963 11141
rect 5905 11132 5917 11135
rect 4396 11104 5917 11132
rect 4396 11092 4402 11104
rect 5905 11101 5917 11104
rect 5951 11132 5963 11135
rect 6270 11132 6276 11144
rect 5951 11104 6276 11132
rect 5951 11101 5963 11104
rect 5905 11095 5963 11101
rect 6270 11092 6276 11104
rect 6328 11092 6334 11144
rect 6638 11092 6644 11144
rect 6696 11132 6702 11144
rect 9861 11135 9919 11141
rect 9861 11132 9873 11135
rect 6696 11104 9873 11132
rect 6696 11092 6702 11104
rect 9861 11101 9873 11104
rect 9907 11132 9919 11135
rect 10686 11132 10692 11144
rect 9907 11104 10692 11132
rect 9907 11101 9919 11104
rect 9861 11095 9919 11101
rect 10686 11092 10692 11104
rect 10744 11092 10750 11144
rect 11330 11132 11336 11144
rect 11291 11104 11336 11132
rect 11330 11092 11336 11104
rect 11388 11092 11394 11144
rect 13630 11132 13636 11144
rect 13591 11104 13636 11132
rect 13630 11092 13636 11104
rect 13688 11092 13694 11144
rect 16209 11135 16267 11141
rect 16209 11101 16221 11135
rect 16255 11132 16267 11135
rect 16482 11132 16488 11144
rect 16255 11104 16488 11132
rect 16255 11101 16267 11104
rect 16209 11095 16267 11101
rect 16482 11092 16488 11104
rect 16540 11132 16546 11144
rect 16540 11104 16947 11132
rect 16540 11092 16546 11104
rect 4522 11024 4528 11076
rect 4580 11064 4586 11076
rect 4709 11067 4767 11073
rect 4709 11064 4721 11067
rect 4580 11036 4721 11064
rect 4580 11024 4586 11036
rect 4709 11033 4721 11036
rect 4755 11033 4767 11067
rect 4709 11027 4767 11033
rect 8021 11067 8079 11073
rect 8021 11033 8033 11067
rect 8067 11064 8079 11067
rect 8662 11064 8668 11076
rect 8067 11036 8668 11064
rect 8067 11033 8079 11036
rect 8021 11027 8079 11033
rect 8662 11024 8668 11036
rect 8720 11024 8726 11076
rect 10410 11064 10416 11076
rect 10371 11036 10416 11064
rect 10410 11024 10416 11036
rect 10468 11024 10474 11076
rect 12253 11067 12311 11073
rect 12253 11033 12265 11067
rect 12299 11064 12311 11067
rect 12618 11064 12624 11076
rect 12299 11036 12624 11064
rect 12299 11033 12311 11036
rect 12253 11027 12311 11033
rect 12618 11024 12624 11036
rect 12676 11064 12682 11076
rect 13262 11064 13268 11076
rect 12676 11036 13268 11064
rect 12676 11024 12682 11036
rect 13262 11024 13268 11036
rect 13320 11024 13326 11076
rect 16758 11064 16764 11076
rect 16719 11036 16764 11064
rect 16758 11024 16764 11036
rect 16816 11024 16822 11076
rect 16919 11064 16947 11104
rect 17678 11064 17684 11076
rect 16919 11036 17684 11064
rect 17678 11024 17684 11036
rect 17736 11024 17742 11076
rect 5810 10996 5816 11008
rect 4264 10968 5816 10996
rect 5810 10956 5816 10968
rect 5868 10956 5874 11008
rect 7650 10956 7656 11008
rect 7708 10996 7714 11008
rect 7834 10996 7840 11008
rect 7708 10968 7840 10996
rect 7708 10956 7714 10968
rect 7834 10956 7840 10968
rect 7892 10956 7898 11008
rect 9490 10996 9496 11008
rect 9451 10968 9496 10996
rect 9490 10956 9496 10968
rect 9548 10956 9554 11008
rect 12710 10956 12716 11008
rect 12768 10996 12774 11008
rect 18138 10996 18144 11008
rect 12768 10968 18144 10996
rect 12768 10956 12774 10968
rect 18138 10956 18144 10968
rect 18196 10956 18202 11008
rect 1104 10906 20884 10928
rect 1104 10854 4648 10906
rect 4700 10854 4712 10906
rect 4764 10854 4776 10906
rect 4828 10854 4840 10906
rect 4892 10854 11982 10906
rect 12034 10854 12046 10906
rect 12098 10854 12110 10906
rect 12162 10854 12174 10906
rect 12226 10854 19315 10906
rect 19367 10854 19379 10906
rect 19431 10854 19443 10906
rect 19495 10854 19507 10906
rect 19559 10854 20884 10906
rect 1104 10832 20884 10854
rect 3973 10795 4031 10801
rect 3973 10761 3985 10795
rect 4019 10792 4031 10795
rect 4246 10792 4252 10804
rect 4019 10764 4252 10792
rect 4019 10761 4031 10764
rect 3973 10755 4031 10761
rect 4246 10752 4252 10764
rect 4304 10752 4310 10804
rect 4525 10795 4583 10801
rect 4525 10761 4537 10795
rect 4571 10792 4583 10795
rect 5997 10795 6055 10801
rect 5997 10792 6009 10795
rect 4571 10764 6009 10792
rect 4571 10761 4583 10764
rect 4525 10755 4583 10761
rect 5997 10761 6009 10764
rect 6043 10792 6055 10795
rect 6086 10792 6092 10804
rect 6043 10764 6092 10792
rect 6043 10761 6055 10764
rect 5997 10755 6055 10761
rect 6086 10752 6092 10764
rect 6144 10752 6150 10804
rect 6270 10792 6276 10804
rect 6231 10764 6276 10792
rect 6270 10752 6276 10764
rect 6328 10752 6334 10804
rect 7006 10752 7012 10804
rect 7064 10792 7070 10804
rect 7101 10795 7159 10801
rect 7101 10792 7113 10795
rect 7064 10764 7113 10792
rect 7064 10752 7070 10764
rect 7101 10761 7113 10764
rect 7147 10761 7159 10795
rect 7101 10755 7159 10761
rect 7466 10752 7472 10804
rect 7524 10792 7530 10804
rect 7742 10792 7748 10804
rect 7524 10764 7748 10792
rect 7524 10752 7530 10764
rect 7742 10752 7748 10764
rect 7800 10792 7806 10804
rect 8665 10795 8723 10801
rect 8665 10792 8677 10795
rect 7800 10764 8677 10792
rect 7800 10752 7806 10764
rect 8665 10761 8677 10764
rect 8711 10761 8723 10795
rect 10502 10792 10508 10804
rect 10463 10764 10508 10792
rect 8665 10755 8723 10761
rect 10502 10752 10508 10764
rect 10560 10752 10566 10804
rect 10686 10752 10692 10804
rect 10744 10792 10750 10804
rect 10781 10795 10839 10801
rect 10781 10792 10793 10795
rect 10744 10764 10793 10792
rect 10744 10752 10750 10764
rect 10781 10761 10793 10764
rect 10827 10761 10839 10795
rect 10781 10755 10839 10761
rect 12253 10795 12311 10801
rect 12253 10761 12265 10795
rect 12299 10792 12311 10795
rect 12342 10792 12348 10804
rect 12299 10764 12348 10792
rect 12299 10761 12311 10764
rect 12253 10755 12311 10761
rect 12342 10752 12348 10764
rect 12400 10752 12406 10804
rect 13262 10752 13268 10804
rect 13320 10792 13326 10804
rect 13449 10795 13507 10801
rect 13449 10792 13461 10795
rect 13320 10764 13461 10792
rect 13320 10752 13326 10764
rect 13449 10761 13461 10764
rect 13495 10761 13507 10795
rect 13449 10755 13507 10761
rect 13722 10752 13728 10804
rect 13780 10792 13786 10804
rect 13817 10795 13875 10801
rect 13817 10792 13829 10795
rect 13780 10764 13829 10792
rect 13780 10752 13786 10764
rect 13817 10761 13829 10764
rect 13863 10761 13875 10795
rect 13817 10755 13875 10761
rect 15657 10795 15715 10801
rect 15657 10761 15669 10795
rect 15703 10792 15715 10795
rect 16025 10795 16083 10801
rect 16025 10792 16037 10795
rect 15703 10764 16037 10792
rect 15703 10761 15715 10764
rect 15657 10755 15715 10761
rect 16025 10761 16037 10764
rect 16071 10792 16083 10795
rect 16298 10792 16304 10804
rect 16071 10764 16304 10792
rect 16071 10761 16083 10764
rect 16025 10755 16083 10761
rect 16298 10752 16304 10764
rect 16356 10752 16362 10804
rect 20162 10792 20168 10804
rect 20123 10764 20168 10792
rect 20162 10752 20168 10764
rect 20220 10752 20226 10804
rect 3602 10724 3608 10736
rect 2516 10696 3608 10724
rect 2516 10597 2544 10696
rect 3602 10684 3608 10696
rect 3660 10724 3666 10736
rect 4617 10727 4675 10733
rect 4617 10724 4629 10727
rect 3660 10696 4629 10724
rect 3660 10684 3666 10696
rect 4617 10693 4629 10696
rect 4663 10693 4675 10727
rect 4617 10687 4675 10693
rect 9309 10727 9367 10733
rect 9309 10693 9321 10727
rect 9355 10724 9367 10727
rect 9398 10724 9404 10736
rect 9355 10696 9404 10724
rect 9355 10693 9367 10696
rect 9309 10687 9367 10693
rect 3053 10659 3111 10665
rect 3053 10625 3065 10659
rect 3099 10656 3111 10659
rect 3234 10656 3240 10668
rect 3099 10628 3240 10656
rect 3099 10625 3111 10628
rect 3053 10619 3111 10625
rect 3234 10616 3240 10628
rect 3292 10616 3298 10668
rect 4525 10659 4583 10665
rect 4525 10656 4537 10659
rect 3620 10628 4537 10656
rect 1765 10591 1823 10597
rect 1765 10557 1777 10591
rect 1811 10557 1823 10591
rect 1765 10551 1823 10557
rect 2041 10591 2099 10597
rect 2041 10557 2053 10591
rect 2087 10588 2099 10591
rect 2501 10591 2559 10597
rect 2501 10588 2513 10591
rect 2087 10560 2513 10588
rect 2087 10557 2099 10560
rect 2041 10551 2099 10557
rect 2501 10557 2513 10560
rect 2547 10557 2559 10591
rect 2501 10551 2559 10557
rect 1780 10520 1808 10551
rect 2590 10520 2596 10532
rect 1780 10492 2596 10520
rect 2590 10480 2596 10492
rect 2648 10480 2654 10532
rect 2961 10523 3019 10529
rect 2961 10489 2973 10523
rect 3007 10520 3019 10523
rect 3374 10523 3432 10529
rect 3374 10520 3386 10523
rect 3007 10492 3386 10520
rect 3007 10489 3019 10492
rect 2961 10483 3019 10489
rect 3374 10489 3386 10492
rect 3420 10520 3432 10523
rect 3620 10520 3648 10628
rect 4525 10625 4537 10628
rect 4571 10625 4583 10659
rect 4632 10656 4660 10687
rect 9398 10684 9404 10696
rect 9456 10724 9462 10736
rect 13081 10727 13139 10733
rect 13081 10724 13093 10727
rect 9456 10696 9536 10724
rect 9456 10684 9462 10696
rect 7466 10656 7472 10668
rect 4632 10628 7472 10656
rect 4525 10619 4583 10625
rect 4341 10591 4399 10597
rect 4341 10557 4353 10591
rect 4387 10588 4399 10591
rect 4982 10588 4988 10600
rect 4387 10560 4988 10588
rect 4387 10557 4399 10560
rect 4341 10551 4399 10557
rect 4982 10548 4988 10560
rect 5040 10548 5046 10600
rect 5276 10597 5304 10628
rect 7466 10616 7472 10628
rect 7524 10616 7530 10668
rect 7558 10616 7564 10668
rect 7616 10656 7622 10668
rect 9508 10665 9536 10696
rect 10152 10696 13093 10724
rect 7653 10659 7711 10665
rect 7653 10656 7665 10659
rect 7616 10628 7665 10656
rect 7616 10616 7622 10628
rect 7653 10625 7665 10628
rect 7699 10625 7711 10659
rect 7653 10619 7711 10625
rect 9493 10659 9551 10665
rect 9493 10625 9505 10659
rect 9539 10625 9551 10659
rect 9493 10619 9551 10625
rect 5261 10591 5319 10597
rect 5261 10557 5273 10591
rect 5307 10557 5319 10591
rect 5261 10551 5319 10557
rect 3420 10492 3648 10520
rect 3420 10489 3432 10492
rect 3374 10483 3432 10489
rect 3786 10480 3792 10532
rect 3844 10520 3850 10532
rect 3844 10492 4936 10520
rect 3844 10480 3850 10492
rect 1578 10452 1584 10464
rect 1539 10424 1584 10452
rect 1578 10412 1584 10424
rect 1636 10412 1642 10464
rect 4908 10461 4936 10492
rect 7190 10480 7196 10532
rect 7248 10520 7254 10532
rect 7377 10523 7435 10529
rect 7377 10520 7389 10523
rect 7248 10492 7389 10520
rect 7248 10480 7254 10492
rect 7377 10489 7389 10492
rect 7423 10489 7435 10523
rect 7377 10483 7435 10489
rect 7469 10523 7527 10529
rect 7469 10489 7481 10523
rect 7515 10489 7527 10523
rect 9582 10520 9588 10532
rect 9543 10492 9588 10520
rect 7469 10483 7527 10489
rect 4893 10455 4951 10461
rect 4893 10421 4905 10455
rect 4939 10421 4951 10455
rect 4893 10415 4951 10421
rect 7006 10412 7012 10464
rect 7064 10452 7070 10464
rect 7484 10452 7512 10483
rect 9582 10480 9588 10492
rect 9640 10480 9646 10532
rect 10152 10529 10180 10696
rect 13081 10693 13093 10696
rect 13127 10724 13139 10727
rect 13538 10724 13544 10736
rect 13127 10696 13544 10724
rect 13127 10693 13139 10696
rect 13081 10687 13139 10693
rect 13538 10684 13544 10696
rect 13596 10684 13602 10736
rect 14366 10684 14372 10736
rect 14424 10724 14430 10736
rect 17405 10727 17463 10733
rect 17405 10724 17417 10727
rect 14424 10696 17417 10724
rect 14424 10684 14430 10696
rect 17405 10693 17417 10696
rect 17451 10724 17463 10727
rect 17773 10727 17831 10733
rect 17773 10724 17785 10727
rect 17451 10696 17785 10724
rect 17451 10693 17463 10696
rect 17405 10687 17463 10693
rect 17773 10693 17785 10696
rect 17819 10724 17831 10727
rect 18230 10724 18236 10736
rect 17819 10696 18236 10724
rect 17819 10693 17831 10696
rect 17773 10687 17831 10693
rect 18230 10684 18236 10696
rect 18288 10724 18294 10736
rect 18506 10724 18512 10736
rect 18288 10696 18512 10724
rect 18288 10684 18294 10696
rect 18506 10684 18512 10696
rect 18564 10684 18570 10736
rect 11471 10659 11529 10665
rect 11471 10625 11483 10659
rect 11517 10656 11529 10659
rect 12986 10656 12992 10668
rect 11517 10628 12992 10656
rect 11517 10625 11529 10628
rect 11471 10619 11529 10625
rect 12986 10616 12992 10628
rect 13044 10616 13050 10668
rect 14090 10656 14096 10668
rect 14016 10628 14096 10656
rect 10686 10548 10692 10600
rect 10744 10588 10750 10600
rect 10962 10588 10968 10600
rect 10744 10560 10968 10588
rect 10744 10548 10750 10560
rect 10962 10548 10968 10560
rect 11020 10588 11026 10600
rect 14016 10597 14044 10628
rect 14090 10616 14096 10628
rect 14148 10616 14154 10668
rect 14550 10656 14556 10668
rect 14511 10628 14556 10656
rect 14550 10616 14556 10628
rect 14608 10616 14614 10668
rect 15289 10659 15347 10665
rect 15289 10625 15301 10659
rect 15335 10656 15347 10659
rect 16209 10659 16267 10665
rect 16209 10656 16221 10659
rect 15335 10628 16221 10656
rect 15335 10625 15347 10628
rect 15289 10619 15347 10625
rect 16209 10625 16221 10628
rect 16255 10656 16267 10659
rect 19751 10659 19809 10665
rect 19751 10656 19763 10659
rect 16255 10628 19763 10656
rect 16255 10625 16267 10628
rect 16209 10619 16267 10625
rect 19751 10625 19763 10628
rect 19797 10625 19809 10659
rect 19751 10619 19809 10625
rect 11368 10591 11426 10597
rect 11368 10588 11380 10591
rect 11020 10560 11380 10588
rect 11020 10548 11026 10560
rect 11368 10557 11380 10560
rect 11414 10588 11426 10591
rect 11793 10591 11851 10597
rect 11793 10588 11805 10591
rect 11414 10560 11805 10588
rect 11414 10557 11426 10560
rect 11368 10551 11426 10557
rect 11793 10557 11805 10560
rect 11839 10557 11851 10591
rect 11793 10551 11851 10557
rect 14001 10591 14059 10597
rect 14001 10557 14013 10591
rect 14047 10557 14059 10591
rect 14461 10591 14519 10597
rect 14461 10588 14473 10591
rect 14001 10551 14059 10557
rect 14108 10560 14473 10588
rect 10137 10523 10195 10529
rect 10137 10489 10149 10523
rect 10183 10489 10195 10523
rect 12526 10520 12532 10532
rect 12487 10492 12532 10520
rect 10137 10483 10195 10489
rect 7064 10424 7512 10452
rect 8389 10455 8447 10461
rect 7064 10412 7070 10424
rect 8389 10421 8401 10455
rect 8435 10452 8447 10455
rect 8662 10452 8668 10464
rect 8435 10424 8668 10452
rect 8435 10421 8447 10424
rect 8389 10415 8447 10421
rect 8662 10412 8668 10424
rect 8720 10412 8726 10464
rect 8754 10412 8760 10464
rect 8812 10452 8818 10464
rect 10152 10452 10180 10483
rect 12526 10480 12532 10492
rect 12584 10480 12590 10532
rect 12621 10523 12679 10529
rect 12621 10489 12633 10523
rect 12667 10489 12679 10523
rect 12621 10483 12679 10489
rect 8812 10424 10180 10452
rect 11241 10455 11299 10461
rect 8812 10412 8818 10424
rect 11241 10421 11253 10455
rect 11287 10452 11299 10455
rect 11330 10452 11336 10464
rect 11287 10424 11336 10452
rect 11287 10421 11299 10424
rect 11241 10415 11299 10421
rect 11330 10412 11336 10424
rect 11388 10412 11394 10464
rect 12434 10412 12440 10464
rect 12492 10452 12498 10464
rect 12636 10452 12664 10483
rect 13722 10480 13728 10532
rect 13780 10520 13786 10532
rect 14108 10520 14136 10560
rect 14461 10557 14473 10560
rect 14507 10557 14519 10591
rect 14461 10551 14519 10557
rect 17310 10548 17316 10600
rect 17368 10588 17374 10600
rect 18230 10588 18236 10600
rect 17368 10560 18236 10588
rect 17368 10548 17374 10560
rect 18230 10548 18236 10560
rect 18288 10548 18294 10600
rect 18506 10588 18512 10600
rect 18467 10560 18512 10588
rect 18506 10548 18512 10560
rect 18564 10548 18570 10600
rect 19664 10591 19722 10597
rect 19664 10557 19676 10591
rect 19710 10588 19722 10591
rect 20162 10588 20168 10600
rect 19710 10560 20168 10588
rect 19710 10557 19722 10560
rect 19664 10551 19722 10557
rect 20162 10548 20168 10560
rect 20220 10548 20226 10600
rect 13780 10492 14136 10520
rect 13780 10480 13786 10492
rect 16298 10480 16304 10532
rect 16356 10520 16362 10532
rect 16853 10523 16911 10529
rect 16356 10492 16401 10520
rect 16356 10480 16362 10492
rect 16853 10489 16865 10523
rect 16899 10489 16911 10523
rect 16853 10483 16911 10489
rect 12492 10424 12664 10452
rect 12492 10412 12498 10424
rect 13814 10412 13820 10464
rect 13872 10452 13878 10464
rect 16868 10452 16896 10483
rect 17310 10452 17316 10464
rect 13872 10424 17316 10452
rect 13872 10412 13878 10424
rect 17310 10412 17316 10424
rect 17368 10412 17374 10464
rect 17862 10412 17868 10464
rect 17920 10452 17926 10464
rect 18141 10455 18199 10461
rect 18141 10452 18153 10455
rect 17920 10424 18153 10452
rect 17920 10412 17926 10424
rect 18141 10421 18153 10424
rect 18187 10421 18199 10455
rect 18141 10415 18199 10421
rect 19337 10455 19395 10461
rect 19337 10421 19349 10455
rect 19383 10452 19395 10455
rect 19610 10452 19616 10464
rect 19383 10424 19616 10452
rect 19383 10421 19395 10424
rect 19337 10415 19395 10421
rect 19610 10412 19616 10424
rect 19668 10412 19674 10464
rect 1104 10362 20884 10384
rect 1104 10310 8315 10362
rect 8367 10310 8379 10362
rect 8431 10310 8443 10362
rect 8495 10310 8507 10362
rect 8559 10310 15648 10362
rect 15700 10310 15712 10362
rect 15764 10310 15776 10362
rect 15828 10310 15840 10362
rect 15892 10310 20884 10362
rect 1104 10288 20884 10310
rect 2130 10208 2136 10260
rect 2188 10248 2194 10260
rect 2593 10251 2651 10257
rect 2593 10248 2605 10251
rect 2188 10220 2605 10248
rect 2188 10208 2194 10220
rect 2593 10217 2605 10220
rect 2639 10217 2651 10251
rect 2593 10211 2651 10217
rect 3234 10208 3240 10260
rect 3292 10248 3298 10260
rect 3697 10251 3755 10257
rect 3697 10248 3709 10251
rect 3292 10220 3709 10248
rect 3292 10208 3298 10220
rect 3697 10217 3709 10220
rect 3743 10217 3755 10251
rect 4246 10248 4252 10260
rect 4207 10220 4252 10248
rect 3697 10211 3755 10217
rect 4246 10208 4252 10220
rect 4304 10208 4310 10260
rect 5537 10251 5595 10257
rect 5537 10217 5549 10251
rect 5583 10248 5595 10251
rect 5810 10248 5816 10260
rect 5583 10220 5816 10248
rect 5583 10217 5595 10220
rect 5537 10211 5595 10217
rect 5810 10208 5816 10220
rect 5868 10208 5874 10260
rect 6319 10251 6377 10257
rect 6319 10217 6331 10251
rect 6365 10248 6377 10251
rect 6638 10248 6644 10260
rect 6365 10220 6644 10248
rect 6365 10217 6377 10220
rect 6319 10211 6377 10217
rect 6638 10208 6644 10220
rect 6696 10208 6702 10260
rect 6730 10208 6736 10260
rect 6788 10248 6794 10260
rect 6825 10251 6883 10257
rect 6825 10248 6837 10251
rect 6788 10220 6837 10248
rect 6788 10208 6794 10220
rect 6825 10217 6837 10220
rect 6871 10217 6883 10251
rect 6825 10211 6883 10217
rect 9950 10208 9956 10260
rect 10008 10248 10014 10260
rect 10045 10251 10103 10257
rect 10045 10248 10057 10251
rect 10008 10220 10057 10248
rect 10008 10208 10014 10220
rect 10045 10217 10057 10220
rect 10091 10248 10103 10251
rect 10226 10248 10232 10260
rect 10091 10220 10232 10248
rect 10091 10217 10103 10220
rect 10045 10211 10103 10217
rect 10226 10208 10232 10220
rect 10284 10208 10290 10260
rect 10778 10208 10784 10260
rect 10836 10248 10842 10260
rect 10873 10251 10931 10257
rect 10873 10248 10885 10251
rect 10836 10220 10885 10248
rect 10836 10208 10842 10220
rect 10873 10217 10885 10220
rect 10919 10217 10931 10251
rect 10873 10211 10931 10217
rect 12161 10251 12219 10257
rect 12161 10217 12173 10251
rect 12207 10248 12219 10251
rect 12526 10248 12532 10260
rect 12207 10220 12532 10248
rect 12207 10217 12219 10220
rect 12161 10211 12219 10217
rect 12526 10208 12532 10220
rect 12584 10208 12590 10260
rect 16209 10251 16267 10257
rect 12636 10220 15976 10248
rect 1765 10183 1823 10189
rect 1765 10149 1777 10183
rect 1811 10180 1823 10183
rect 2314 10180 2320 10192
rect 1811 10152 2320 10180
rect 1811 10149 1823 10152
rect 1765 10143 1823 10149
rect 2314 10140 2320 10152
rect 2372 10140 2378 10192
rect 4522 10140 4528 10192
rect 4580 10180 4586 10192
rect 4617 10183 4675 10189
rect 4617 10180 4629 10183
rect 4580 10152 4629 10180
rect 4580 10140 4586 10152
rect 4617 10149 4629 10152
rect 4663 10149 4675 10183
rect 4617 10143 4675 10149
rect 5169 10183 5227 10189
rect 5169 10149 5181 10183
rect 5215 10180 5227 10183
rect 5261 10183 5319 10189
rect 5261 10180 5273 10183
rect 5215 10152 5273 10180
rect 5215 10149 5227 10152
rect 5169 10143 5227 10149
rect 5261 10149 5273 10152
rect 5307 10180 5319 10183
rect 5442 10180 5448 10192
rect 5307 10152 5448 10180
rect 5307 10149 5319 10152
rect 5261 10143 5319 10149
rect 5442 10140 5448 10152
rect 5500 10140 5506 10192
rect 7377 10183 7435 10189
rect 7377 10149 7389 10183
rect 7423 10180 7435 10183
rect 7650 10180 7656 10192
rect 7423 10152 7656 10180
rect 7423 10149 7435 10152
rect 7377 10143 7435 10149
rect 7650 10140 7656 10152
rect 7708 10140 7714 10192
rect 11146 10140 11152 10192
rect 11204 10180 11210 10192
rect 11204 10152 11468 10180
rect 11204 10140 11210 10152
rect 2590 10072 2596 10124
rect 2648 10112 2654 10124
rect 2961 10115 3019 10121
rect 2961 10112 2973 10115
rect 2648 10084 2973 10112
rect 2648 10072 2654 10084
rect 2961 10081 2973 10084
rect 3007 10081 3019 10115
rect 2961 10075 3019 10081
rect 6248 10115 6306 10121
rect 6248 10081 6260 10115
rect 6294 10112 6306 10115
rect 6546 10112 6552 10124
rect 6294 10084 6552 10112
rect 6294 10081 6306 10084
rect 6248 10075 6306 10081
rect 6546 10072 6552 10084
rect 6604 10072 6610 10124
rect 9493 10115 9551 10121
rect 9493 10081 9505 10115
rect 9539 10112 9551 10115
rect 9582 10112 9588 10124
rect 9539 10084 9588 10112
rect 9539 10081 9551 10084
rect 9493 10075 9551 10081
rect 9582 10072 9588 10084
rect 9640 10112 9646 10124
rect 11440 10121 11468 10152
rect 10597 10115 10655 10121
rect 10597 10112 10609 10115
rect 9640 10084 10609 10112
rect 9640 10072 9646 10084
rect 10597 10081 10609 10084
rect 10643 10081 10655 10115
rect 10597 10075 10655 10081
rect 11425 10115 11483 10121
rect 11425 10081 11437 10115
rect 11471 10081 11483 10115
rect 11425 10075 11483 10081
rect 1394 10004 1400 10056
rect 1452 10044 1458 10056
rect 1673 10047 1731 10053
rect 1673 10044 1685 10047
rect 1452 10016 1685 10044
rect 1452 10004 1458 10016
rect 1673 10013 1685 10016
rect 1719 10013 1731 10047
rect 1673 10007 1731 10013
rect 4525 10047 4583 10053
rect 4525 10013 4537 10047
rect 4571 10044 4583 10047
rect 4614 10044 4620 10056
rect 4571 10016 4620 10044
rect 4571 10013 4583 10016
rect 4525 10007 4583 10013
rect 4614 10004 4620 10016
rect 4672 10044 4678 10056
rect 5350 10044 5356 10056
rect 4672 10016 5356 10044
rect 4672 10004 4678 10016
rect 5350 10004 5356 10016
rect 5408 10004 5414 10056
rect 6822 10004 6828 10056
rect 6880 10044 6886 10056
rect 7282 10044 7288 10056
rect 6880 10016 7288 10044
rect 6880 10004 6886 10016
rect 7282 10004 7288 10016
rect 7340 10004 7346 10056
rect 7558 10044 7564 10056
rect 7471 10016 7564 10044
rect 7558 10004 7564 10016
rect 7616 10004 7622 10056
rect 9677 10047 9735 10053
rect 9677 10013 9689 10047
rect 9723 10044 9735 10047
rect 9950 10044 9956 10056
rect 9723 10016 9956 10044
rect 9723 10013 9735 10016
rect 9677 10007 9735 10013
rect 9950 10004 9956 10016
rect 10008 10044 10014 10056
rect 12636 10044 12664 10220
rect 13167 10183 13225 10189
rect 13167 10149 13179 10183
rect 13213 10180 13225 10183
rect 13262 10180 13268 10192
rect 13213 10152 13268 10180
rect 13213 10149 13225 10152
rect 13167 10143 13225 10149
rect 13262 10140 13268 10152
rect 13320 10180 13326 10192
rect 14550 10180 14556 10192
rect 13320 10152 14556 10180
rect 13320 10140 13326 10152
rect 14550 10140 14556 10152
rect 14608 10180 14614 10192
rect 15610 10183 15668 10189
rect 15610 10180 15622 10183
rect 14608 10152 15622 10180
rect 14608 10140 14614 10152
rect 15610 10149 15622 10152
rect 15656 10149 15668 10183
rect 15948 10180 15976 10220
rect 16209 10217 16221 10251
rect 16255 10248 16267 10251
rect 16298 10248 16304 10260
rect 16255 10220 16304 10248
rect 16255 10217 16267 10220
rect 16209 10211 16267 10217
rect 16298 10208 16304 10220
rect 16356 10208 16362 10260
rect 16482 10248 16488 10260
rect 16443 10220 16488 10248
rect 16482 10208 16488 10220
rect 16540 10208 16546 10260
rect 16850 10248 16856 10260
rect 16811 10220 16856 10248
rect 16850 10208 16856 10220
rect 16908 10208 16914 10260
rect 17954 10208 17960 10260
rect 18012 10248 18018 10260
rect 18049 10251 18107 10257
rect 18049 10248 18061 10251
rect 18012 10220 18061 10248
rect 18012 10208 18018 10220
rect 18049 10217 18061 10220
rect 18095 10217 18107 10251
rect 18690 10248 18696 10260
rect 18651 10220 18696 10248
rect 18049 10211 18107 10217
rect 18690 10208 18696 10220
rect 18748 10208 18754 10260
rect 16574 10180 16580 10192
rect 15948 10152 16580 10180
rect 15610 10143 15668 10149
rect 16574 10140 16580 10152
rect 16632 10140 16638 10192
rect 16868 10180 16896 10208
rect 17129 10183 17187 10189
rect 17129 10180 17141 10183
rect 16868 10152 17141 10180
rect 17129 10149 17141 10152
rect 17175 10149 17187 10183
rect 17129 10143 17187 10149
rect 17218 10140 17224 10192
rect 17276 10180 17282 10192
rect 17276 10152 17321 10180
rect 17276 10140 17282 10152
rect 18506 10140 18512 10192
rect 18564 10180 18570 10192
rect 18966 10180 18972 10192
rect 18564 10152 18972 10180
rect 18564 10140 18570 10152
rect 18966 10140 18972 10152
rect 19024 10180 19030 10192
rect 19024 10152 19104 10180
rect 19024 10140 19030 10152
rect 16022 10112 16028 10124
rect 13786 10084 16028 10112
rect 12802 10044 12808 10056
rect 10008 10016 12664 10044
rect 12763 10016 12808 10044
rect 10008 10004 10014 10016
rect 12802 10004 12808 10016
rect 12860 10044 12866 10056
rect 13786 10044 13814 10084
rect 16022 10072 16028 10084
rect 16080 10072 16086 10124
rect 18598 10112 18604 10124
rect 18559 10084 18604 10112
rect 18598 10072 18604 10084
rect 18656 10072 18662 10124
rect 19076 10121 19104 10152
rect 19061 10115 19119 10121
rect 19061 10081 19073 10115
rect 19107 10081 19119 10115
rect 19061 10075 19119 10081
rect 15286 10044 15292 10056
rect 12860 10016 13814 10044
rect 15247 10016 15292 10044
rect 12860 10004 12866 10016
rect 15286 10004 15292 10016
rect 15344 10004 15350 10056
rect 17310 10004 17316 10056
rect 17368 10044 17374 10056
rect 17405 10047 17463 10053
rect 17405 10044 17417 10047
rect 17368 10016 17417 10044
rect 17368 10004 17374 10016
rect 17405 10013 17417 10016
rect 17451 10013 17463 10047
rect 17405 10007 17463 10013
rect 2225 9979 2283 9985
rect 2225 9945 2237 9979
rect 2271 9976 2283 9979
rect 4982 9976 4988 9988
rect 2271 9948 4988 9976
rect 2271 9945 2283 9948
rect 2225 9939 2283 9945
rect 4982 9936 4988 9948
rect 5040 9976 5046 9988
rect 5261 9979 5319 9985
rect 5261 9976 5273 9979
rect 5040 9948 5273 9976
rect 5040 9936 5046 9948
rect 5261 9945 5273 9948
rect 5307 9945 5319 9979
rect 5368 9976 5396 10004
rect 7576 9976 7604 10004
rect 8754 9976 8760 9988
rect 5368 9948 7604 9976
rect 8036 9948 8760 9976
rect 5261 9939 5319 9945
rect 3421 9911 3479 9917
rect 3421 9877 3433 9911
rect 3467 9908 3479 9911
rect 3510 9908 3516 9920
rect 3467 9880 3516 9908
rect 3467 9877 3479 9880
rect 3421 9871 3479 9877
rect 3510 9868 3516 9880
rect 3568 9868 3574 9920
rect 4062 9868 4068 9920
rect 4120 9908 4126 9920
rect 5813 9911 5871 9917
rect 5813 9908 5825 9911
rect 4120 9880 5825 9908
rect 4120 9868 4126 9880
rect 5813 9877 5825 9880
rect 5859 9908 5871 9911
rect 8036 9908 8064 9948
rect 8754 9936 8760 9948
rect 8812 9936 8818 9988
rect 9398 9936 9404 9988
rect 9456 9976 9462 9988
rect 13446 9976 13452 9988
rect 9456 9948 13452 9976
rect 9456 9936 9462 9948
rect 13446 9936 13452 9948
rect 13504 9936 13510 9988
rect 13630 9936 13636 9988
rect 13688 9976 13694 9988
rect 13814 9976 13820 9988
rect 13688 9948 13820 9976
rect 13688 9936 13694 9948
rect 13814 9936 13820 9948
rect 13872 9936 13878 9988
rect 16482 9936 16488 9988
rect 16540 9976 16546 9988
rect 18322 9976 18328 9988
rect 16540 9948 18328 9976
rect 16540 9936 16546 9948
rect 18322 9936 18328 9948
rect 18380 9936 18386 9988
rect 8202 9908 8208 9920
rect 5859 9880 8064 9908
rect 8163 9880 8208 9908
rect 5859 9877 5871 9880
rect 5813 9871 5871 9877
rect 8202 9868 8208 9880
rect 8260 9868 8266 9920
rect 11609 9911 11667 9917
rect 11609 9877 11621 9911
rect 11655 9908 11667 9911
rect 11790 9908 11796 9920
rect 11655 9880 11796 9908
rect 11655 9877 11667 9880
rect 11609 9871 11667 9877
rect 11790 9868 11796 9880
rect 11848 9868 11854 9920
rect 12434 9908 12440 9920
rect 12395 9880 12440 9908
rect 12434 9868 12440 9880
rect 12492 9868 12498 9920
rect 13722 9908 13728 9920
rect 13683 9880 13728 9908
rect 13722 9868 13728 9880
rect 13780 9868 13786 9920
rect 14090 9908 14096 9920
rect 14051 9880 14096 9908
rect 14090 9868 14096 9880
rect 14148 9868 14154 9920
rect 18230 9868 18236 9920
rect 18288 9908 18294 9920
rect 18509 9911 18567 9917
rect 18509 9908 18521 9911
rect 18288 9880 18521 9908
rect 18288 9868 18294 9880
rect 18509 9877 18521 9880
rect 18555 9908 18567 9911
rect 19702 9908 19708 9920
rect 18555 9880 19708 9908
rect 18555 9877 18567 9880
rect 18509 9871 18567 9877
rect 19702 9868 19708 9880
rect 19760 9868 19766 9920
rect 1104 9818 20884 9840
rect 1104 9766 4648 9818
rect 4700 9766 4712 9818
rect 4764 9766 4776 9818
rect 4828 9766 4840 9818
rect 4892 9766 11982 9818
rect 12034 9766 12046 9818
rect 12098 9766 12110 9818
rect 12162 9766 12174 9818
rect 12226 9766 19315 9818
rect 19367 9766 19379 9818
rect 19431 9766 19443 9818
rect 19495 9766 19507 9818
rect 19559 9766 20884 9818
rect 1104 9744 20884 9766
rect 2314 9704 2320 9716
rect 2275 9676 2320 9704
rect 2314 9664 2320 9676
rect 2372 9664 2378 9716
rect 2866 9664 2872 9716
rect 2924 9704 2930 9716
rect 2961 9707 3019 9713
rect 2961 9704 2973 9707
rect 2924 9676 2973 9704
rect 2924 9664 2930 9676
rect 2961 9673 2973 9676
rect 3007 9673 3019 9707
rect 2961 9667 3019 9673
rect 4522 9664 4528 9716
rect 4580 9704 4586 9716
rect 4709 9707 4767 9713
rect 4709 9704 4721 9707
rect 4580 9676 4721 9704
rect 4580 9664 4586 9676
rect 4709 9673 4721 9676
rect 4755 9704 4767 9707
rect 4985 9707 5043 9713
rect 4985 9704 4997 9707
rect 4755 9676 4997 9704
rect 4755 9673 4767 9676
rect 4709 9667 4767 9673
rect 4985 9673 4997 9676
rect 5031 9673 5043 9707
rect 5350 9704 5356 9716
rect 5311 9676 5356 9704
rect 4985 9667 5043 9673
rect 5350 9664 5356 9676
rect 5408 9664 5414 9716
rect 8110 9664 8116 9716
rect 8168 9704 8174 9716
rect 8665 9707 8723 9713
rect 8665 9704 8677 9707
rect 8168 9676 8677 9704
rect 8168 9664 8174 9676
rect 8665 9673 8677 9676
rect 8711 9673 8723 9707
rect 8665 9667 8723 9673
rect 9953 9707 10011 9713
rect 9953 9673 9965 9707
rect 9999 9704 10011 9707
rect 10226 9704 10232 9716
rect 9999 9676 10232 9704
rect 9999 9673 10011 9676
rect 9953 9667 10011 9673
rect 3786 9568 3792 9580
rect 3747 9540 3792 9568
rect 3786 9528 3792 9540
rect 3844 9528 3850 9580
rect 6730 9528 6736 9580
rect 6788 9568 6794 9580
rect 6825 9571 6883 9577
rect 6825 9568 6837 9571
rect 6788 9540 6837 9568
rect 6788 9528 6794 9540
rect 6825 9537 6837 9540
rect 6871 9537 6883 9571
rect 8680 9568 8708 9667
rect 10226 9664 10232 9676
rect 10284 9704 10290 9716
rect 10413 9707 10471 9713
rect 10413 9704 10425 9707
rect 10284 9676 10425 9704
rect 10284 9664 10290 9676
rect 10413 9673 10425 9676
rect 10459 9673 10471 9707
rect 10413 9667 10471 9673
rect 11517 9707 11575 9713
rect 11517 9673 11529 9707
rect 11563 9704 11575 9707
rect 12434 9704 12440 9716
rect 11563 9676 12440 9704
rect 11563 9673 11575 9676
rect 11517 9667 11575 9673
rect 9490 9568 9496 9580
rect 8680 9540 9352 9568
rect 9451 9540 9496 9568
rect 6825 9531 6883 9537
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9500 1455 9503
rect 1578 9500 1584 9512
rect 1443 9472 1584 9500
rect 1443 9469 1455 9472
rect 1397 9463 1455 9469
rect 1578 9460 1584 9472
rect 1636 9500 1642 9512
rect 3234 9500 3240 9512
rect 1636 9472 3240 9500
rect 1636 9460 1642 9472
rect 3234 9460 3240 9472
rect 3292 9460 3298 9512
rect 5721 9503 5779 9509
rect 5721 9469 5733 9503
rect 5767 9500 5779 9503
rect 8754 9500 8760 9512
rect 5767 9472 8760 9500
rect 5767 9469 5779 9472
rect 5721 9463 5779 9469
rect 8754 9460 8760 9472
rect 8812 9460 8818 9512
rect 9030 9500 9036 9512
rect 8991 9472 9036 9500
rect 9030 9460 9036 9472
rect 9088 9460 9094 9512
rect 9324 9509 9352 9540
rect 9490 9528 9496 9540
rect 9548 9528 9554 9580
rect 10428 9568 10456 9667
rect 12434 9664 12440 9676
rect 12492 9664 12498 9716
rect 14366 9704 14372 9716
rect 13096 9676 14372 9704
rect 11146 9596 11152 9648
rect 11204 9636 11210 9648
rect 11793 9639 11851 9645
rect 11793 9636 11805 9639
rect 11204 9608 11805 9636
rect 11204 9596 11210 9608
rect 11793 9605 11805 9608
rect 11839 9605 11851 9639
rect 11793 9599 11851 9605
rect 12253 9639 12311 9645
rect 12253 9605 12265 9639
rect 12299 9636 12311 9639
rect 12802 9636 12808 9648
rect 12299 9608 12808 9636
rect 12299 9605 12311 9608
rect 12253 9599 12311 9605
rect 12802 9596 12808 9608
rect 12860 9596 12866 9648
rect 10597 9571 10655 9577
rect 10428 9540 10548 9568
rect 9309 9503 9367 9509
rect 9309 9469 9321 9503
rect 9355 9469 9367 9503
rect 9309 9463 9367 9469
rect 1759 9435 1817 9441
rect 1759 9401 1771 9435
rect 1805 9401 1817 9435
rect 3605 9435 3663 9441
rect 3605 9432 3617 9435
rect 1759 9395 1817 9401
rect 2608 9404 3617 9432
rect 1774 9364 1802 9395
rect 1854 9364 1860 9376
rect 1774 9336 1860 9364
rect 1854 9324 1860 9336
rect 1912 9364 1918 9376
rect 2608 9373 2636 9404
rect 3605 9401 3617 9404
rect 3651 9432 3663 9435
rect 4151 9435 4209 9441
rect 4151 9432 4163 9435
rect 3651 9404 4163 9432
rect 3651 9401 3663 9404
rect 3605 9395 3663 9401
rect 4151 9401 4163 9404
rect 4197 9432 4209 9435
rect 4430 9432 4436 9444
rect 4197 9404 4436 9432
rect 4197 9401 4209 9404
rect 4151 9395 4209 9401
rect 4430 9392 4436 9404
rect 4488 9432 4494 9444
rect 10520 9432 10548 9540
rect 10597 9537 10609 9571
rect 10643 9568 10655 9571
rect 10778 9568 10784 9580
rect 10643 9540 10784 9568
rect 10643 9537 10655 9540
rect 10597 9531 10655 9537
rect 10778 9528 10784 9540
rect 10836 9528 10842 9580
rect 10962 9528 10968 9580
rect 11020 9568 11026 9580
rect 13096 9568 13124 9676
rect 14366 9664 14372 9676
rect 14424 9664 14430 9716
rect 14550 9704 14556 9716
rect 14511 9676 14556 9704
rect 14550 9664 14556 9676
rect 14608 9704 14614 9716
rect 14921 9707 14979 9713
rect 14921 9704 14933 9707
rect 14608 9676 14933 9704
rect 14608 9664 14614 9676
rect 14921 9673 14933 9676
rect 14967 9673 14979 9707
rect 14921 9667 14979 9673
rect 16025 9707 16083 9713
rect 16025 9673 16037 9707
rect 16071 9704 16083 9707
rect 16390 9704 16396 9716
rect 16071 9676 16396 9704
rect 16071 9673 16083 9676
rect 16025 9667 16083 9673
rect 13538 9596 13544 9648
rect 13596 9636 13602 9648
rect 13596 9608 13768 9636
rect 13596 9596 13602 9608
rect 11020 9540 13124 9568
rect 13449 9571 13507 9577
rect 11020 9528 11026 9540
rect 13449 9537 13461 9571
rect 13495 9568 13507 9571
rect 13630 9568 13636 9580
rect 13495 9540 13636 9568
rect 13495 9537 13507 9540
rect 13449 9531 13507 9537
rect 13630 9528 13636 9540
rect 13688 9528 13694 9580
rect 13740 9577 13768 9608
rect 13725 9571 13783 9577
rect 13725 9537 13737 9571
rect 13771 9537 13783 9571
rect 13725 9531 13783 9537
rect 11606 9460 11612 9512
rect 11664 9500 11670 9512
rect 12434 9500 12440 9512
rect 11664 9472 12440 9500
rect 11664 9460 11670 9472
rect 12434 9460 12440 9472
rect 12492 9460 12498 9512
rect 10959 9435 11017 9441
rect 10959 9432 10971 9435
rect 4488 9404 6684 9432
rect 10520 9404 10971 9432
rect 4488 9392 4494 9404
rect 2593 9367 2651 9373
rect 2593 9364 2605 9367
rect 1912 9336 2605 9364
rect 1912 9324 1918 9336
rect 2593 9333 2605 9336
rect 2639 9333 2651 9367
rect 2593 9327 2651 9333
rect 6273 9367 6331 9373
rect 6273 9333 6285 9367
rect 6319 9364 6331 9367
rect 6546 9364 6552 9376
rect 6319 9336 6552 9364
rect 6319 9333 6331 9336
rect 6273 9327 6331 9333
rect 6546 9324 6552 9336
rect 6604 9324 6610 9376
rect 6656 9373 6684 9404
rect 10959 9401 10971 9404
rect 11005 9432 11017 9435
rect 13541 9435 13599 9441
rect 11005 9404 11652 9432
rect 11005 9401 11017 9404
rect 10959 9395 11017 9401
rect 11624 9376 11652 9404
rect 13541 9401 13553 9435
rect 13587 9432 13599 9435
rect 13722 9432 13728 9444
rect 13587 9404 13728 9432
rect 13587 9401 13599 9404
rect 13541 9395 13599 9401
rect 6641 9367 6699 9373
rect 6641 9333 6653 9367
rect 6687 9364 6699 9367
rect 7193 9367 7251 9373
rect 7193 9364 7205 9367
rect 6687 9336 7205 9364
rect 6687 9333 6699 9336
rect 6641 9327 6699 9333
rect 7193 9333 7205 9336
rect 7239 9333 7251 9367
rect 7193 9327 7251 9333
rect 7650 9324 7656 9376
rect 7708 9364 7714 9376
rect 7745 9367 7803 9373
rect 7745 9364 7757 9367
rect 7708 9336 7757 9364
rect 7708 9324 7714 9336
rect 7745 9333 7757 9336
rect 7791 9364 7803 9367
rect 8021 9367 8079 9373
rect 8021 9364 8033 9367
rect 7791 9336 8033 9364
rect 7791 9333 7803 9336
rect 7745 9327 7803 9333
rect 8021 9333 8033 9336
rect 8067 9333 8079 9367
rect 8021 9327 8079 9333
rect 11606 9324 11612 9376
rect 11664 9364 11670 9376
rect 12805 9367 12863 9373
rect 12805 9364 12817 9367
rect 11664 9336 12817 9364
rect 11664 9324 11670 9336
rect 12805 9333 12817 9336
rect 12851 9364 12863 9367
rect 13170 9364 13176 9376
rect 12851 9336 13176 9364
rect 12851 9333 12863 9336
rect 12805 9327 12863 9333
rect 13170 9324 13176 9336
rect 13228 9324 13234 9376
rect 13265 9367 13323 9373
rect 13265 9333 13277 9367
rect 13311 9364 13323 9367
rect 13556 9364 13584 9395
rect 13722 9392 13728 9404
rect 13780 9392 13786 9444
rect 14936 9432 14964 9667
rect 16390 9664 16396 9676
rect 16448 9704 16454 9716
rect 16761 9707 16819 9713
rect 16761 9704 16773 9707
rect 16448 9676 16773 9704
rect 16448 9664 16454 9676
rect 16761 9673 16773 9676
rect 16807 9704 16819 9707
rect 17218 9704 17224 9716
rect 16807 9676 17224 9704
rect 16807 9673 16819 9676
rect 16761 9667 16819 9673
rect 17218 9664 17224 9676
rect 17276 9664 17282 9716
rect 18966 9664 18972 9716
rect 19024 9704 19030 9716
rect 19061 9707 19119 9713
rect 19061 9704 19073 9707
rect 19024 9676 19073 9704
rect 19024 9664 19030 9676
rect 19061 9673 19073 9676
rect 19107 9673 19119 9707
rect 19061 9667 19119 9673
rect 17037 9639 17095 9645
rect 17037 9605 17049 9639
rect 17083 9636 17095 9639
rect 21542 9636 21548 9648
rect 17083 9608 21548 9636
rect 17083 9605 17095 9608
rect 17037 9599 17095 9605
rect 21542 9596 21548 9608
rect 21600 9596 21606 9648
rect 15286 9528 15292 9580
rect 15344 9568 15350 9580
rect 16393 9571 16451 9577
rect 16393 9568 16405 9571
rect 15344 9540 16405 9568
rect 15344 9528 15350 9540
rect 16393 9537 16405 9540
rect 16439 9568 16451 9571
rect 17862 9568 17868 9580
rect 16439 9540 17868 9568
rect 16439 9537 16451 9540
rect 16393 9531 16451 9537
rect 17862 9528 17868 9540
rect 17920 9528 17926 9580
rect 18598 9528 18604 9580
rect 18656 9568 18662 9580
rect 18874 9568 18880 9580
rect 18656 9540 18880 9568
rect 18656 9528 18662 9540
rect 18874 9528 18880 9540
rect 18932 9568 18938 9580
rect 19429 9571 19487 9577
rect 19429 9568 19441 9571
rect 18932 9540 19441 9568
rect 18932 9528 18938 9540
rect 19429 9537 19441 9540
rect 19475 9537 19487 9571
rect 19429 9531 19487 9537
rect 15102 9500 15108 9512
rect 15063 9472 15108 9500
rect 15102 9460 15108 9472
rect 15160 9460 15166 9512
rect 16850 9500 16856 9512
rect 16811 9472 16856 9500
rect 16850 9460 16856 9472
rect 16908 9500 16914 9512
rect 17402 9500 17408 9512
rect 16908 9472 17408 9500
rect 16908 9460 16914 9472
rect 17402 9460 17408 9472
rect 17460 9460 17466 9512
rect 17770 9460 17776 9512
rect 17828 9500 17834 9512
rect 18046 9500 18052 9512
rect 17828 9472 18052 9500
rect 17828 9460 17834 9472
rect 18046 9460 18052 9472
rect 18104 9500 18110 9512
rect 18141 9503 18199 9509
rect 18141 9500 18153 9503
rect 18104 9472 18153 9500
rect 18104 9460 18110 9472
rect 18141 9469 18153 9472
rect 18187 9469 18199 9503
rect 18141 9463 18199 9469
rect 18506 9460 18512 9512
rect 18564 9500 18570 9512
rect 19150 9500 19156 9512
rect 18564 9472 19156 9500
rect 18564 9460 18570 9472
rect 19150 9460 19156 9472
rect 19208 9500 19214 9512
rect 19648 9503 19706 9509
rect 19648 9500 19660 9503
rect 19208 9472 19660 9500
rect 19208 9460 19214 9472
rect 19648 9469 19660 9472
rect 19694 9500 19706 9503
rect 20073 9503 20131 9509
rect 20073 9500 20085 9503
rect 19694 9472 20085 9500
rect 19694 9469 19706 9472
rect 19648 9463 19706 9469
rect 20073 9469 20085 9472
rect 20119 9469 20131 9503
rect 20073 9463 20131 9469
rect 15378 9432 15384 9444
rect 14936 9404 15384 9432
rect 15378 9392 15384 9404
rect 15436 9441 15442 9444
rect 15436 9435 15484 9441
rect 15436 9401 15438 9435
rect 15472 9401 15484 9435
rect 15436 9395 15484 9401
rect 15436 9392 15442 9395
rect 16942 9392 16948 9444
rect 17000 9432 17006 9444
rect 19751 9435 19809 9441
rect 19751 9432 19763 9435
rect 17000 9404 19763 9432
rect 17000 9392 17006 9404
rect 19751 9401 19763 9404
rect 19797 9401 19809 9435
rect 19751 9395 19809 9401
rect 17770 9364 17776 9376
rect 13311 9336 13584 9364
rect 17731 9336 17776 9364
rect 13311 9333 13323 9336
rect 13265 9327 13323 9333
rect 17770 9324 17776 9336
rect 17828 9324 17834 9376
rect 17862 9324 17868 9376
rect 17920 9364 17926 9376
rect 18325 9367 18383 9373
rect 18325 9364 18337 9367
rect 17920 9336 18337 9364
rect 17920 9324 17926 9336
rect 18325 9333 18337 9336
rect 18371 9333 18383 9367
rect 18325 9327 18383 9333
rect 1104 9274 20884 9296
rect 1104 9222 8315 9274
rect 8367 9222 8379 9274
rect 8431 9222 8443 9274
rect 8495 9222 8507 9274
rect 8559 9222 15648 9274
rect 15700 9222 15712 9274
rect 15764 9222 15776 9274
rect 15828 9222 15840 9274
rect 15892 9222 20884 9274
rect 1104 9200 20884 9222
rect 1578 9160 1584 9172
rect 1539 9132 1584 9160
rect 1578 9120 1584 9132
rect 1636 9120 1642 9172
rect 2314 9120 2320 9172
rect 2372 9160 2378 9172
rect 2869 9163 2927 9169
rect 2869 9160 2881 9163
rect 2372 9132 2881 9160
rect 2372 9120 2378 9132
rect 2869 9129 2881 9132
rect 2915 9129 2927 9163
rect 3234 9160 3240 9172
rect 3195 9132 3240 9160
rect 2869 9123 2927 9129
rect 3234 9120 3240 9132
rect 3292 9120 3298 9172
rect 3786 9160 3792 9172
rect 3747 9132 3792 9160
rect 3786 9120 3792 9132
rect 3844 9120 3850 9172
rect 4430 9160 4436 9172
rect 4391 9132 4436 9160
rect 4430 9120 4436 9132
rect 4488 9120 4494 9172
rect 7282 9160 7288 9172
rect 7243 9132 7288 9160
rect 7282 9120 7288 9132
rect 7340 9120 7346 9172
rect 7466 9120 7472 9172
rect 7524 9160 7530 9172
rect 8202 9160 8208 9172
rect 7524 9132 8208 9160
rect 7524 9120 7530 9132
rect 8202 9120 8208 9132
rect 8260 9120 8266 9172
rect 9950 9160 9956 9172
rect 9911 9132 9956 9160
rect 9950 9120 9956 9132
rect 10008 9120 10014 9172
rect 10318 9120 10324 9172
rect 10376 9120 10382 9172
rect 12342 9160 12348 9172
rect 12303 9132 12348 9160
rect 12342 9120 12348 9132
rect 12400 9160 12406 9172
rect 13541 9163 13599 9169
rect 12400 9132 12572 9160
rect 12400 9120 12406 9132
rect 5810 9092 5816 9104
rect 1780 9064 5816 9092
rect 1780 9036 1808 9064
rect 5810 9052 5816 9064
rect 5868 9052 5874 9104
rect 5902 9052 5908 9104
rect 5960 9092 5966 9104
rect 6365 9095 6423 9101
rect 6365 9092 6377 9095
rect 5960 9064 6377 9092
rect 5960 9052 5966 9064
rect 6365 9061 6377 9064
rect 6411 9092 6423 9095
rect 7650 9092 7656 9104
rect 6411 9064 7656 9092
rect 6411 9061 6423 9064
rect 6365 9055 6423 9061
rect 7650 9052 7656 9064
rect 7708 9052 7714 9104
rect 7834 9092 7840 9104
rect 7747 9064 7840 9092
rect 1762 9024 1768 9036
rect 1723 8996 1768 9024
rect 1762 8984 1768 8996
rect 1820 8984 1826 9036
rect 2041 9027 2099 9033
rect 2041 8993 2053 9027
rect 2087 9024 2099 9027
rect 2866 9024 2872 9036
rect 2087 8996 2872 9024
rect 2087 8993 2099 8996
rect 2041 8987 2099 8993
rect 2866 8984 2872 8996
rect 2924 8984 2930 9036
rect 3694 8984 3700 9036
rect 3752 9024 3758 9036
rect 5718 9024 5724 9036
rect 3752 8996 5724 9024
rect 3752 8984 3758 8996
rect 5718 8984 5724 8996
rect 5776 8984 5782 9036
rect 6914 8984 6920 9036
rect 6972 9024 6978 9036
rect 6972 8996 7017 9024
rect 6972 8984 6978 8996
rect 7466 8984 7472 9036
rect 7524 9024 7530 9036
rect 7760 9033 7788 9064
rect 7834 9052 7840 9064
rect 7892 9092 7898 9104
rect 9582 9092 9588 9104
rect 7892 9064 9588 9092
rect 7892 9052 7898 9064
rect 9582 9052 9588 9064
rect 9640 9052 9646 9104
rect 7745 9027 7803 9033
rect 7745 9024 7757 9027
rect 7524 8996 7757 9024
rect 7524 8984 7530 8996
rect 7745 8993 7757 8996
rect 7791 8993 7803 9027
rect 7745 8987 7803 8993
rect 8021 9027 8079 9033
rect 8021 8993 8033 9027
rect 8067 9024 8079 9027
rect 8110 9024 8116 9036
rect 8067 8996 8116 9024
rect 8067 8993 8079 8996
rect 8021 8987 8079 8993
rect 8110 8984 8116 8996
rect 8168 9024 8174 9036
rect 10336 9024 10364 9120
rect 11330 9092 11336 9104
rect 11291 9064 11336 9092
rect 11330 9052 11336 9064
rect 11388 9052 11394 9104
rect 12544 9101 12572 9132
rect 13541 9129 13553 9163
rect 13587 9160 13599 9163
rect 13630 9160 13636 9172
rect 13587 9132 13636 9160
rect 13587 9129 13599 9132
rect 13541 9123 13599 9129
rect 13630 9120 13636 9132
rect 13688 9120 13694 9172
rect 15102 9120 15108 9172
rect 15160 9160 15166 9172
rect 15565 9163 15623 9169
rect 15565 9160 15577 9163
rect 15160 9132 15577 9160
rect 15160 9120 15166 9132
rect 15565 9129 15577 9132
rect 15611 9160 15623 9163
rect 18690 9160 18696 9172
rect 15611 9132 18696 9160
rect 15611 9129 15623 9132
rect 15565 9123 15623 9129
rect 18690 9120 18696 9132
rect 18748 9120 18754 9172
rect 12529 9095 12587 9101
rect 12529 9061 12541 9095
rect 12575 9061 12587 9095
rect 12529 9055 12587 9061
rect 12618 9052 12624 9104
rect 12676 9092 12682 9104
rect 16390 9092 16396 9104
rect 12676 9064 12721 9092
rect 16351 9064 16396 9092
rect 12676 9052 12682 9064
rect 16390 9052 16396 9064
rect 16448 9052 16454 9104
rect 10597 9027 10655 9033
rect 10597 9024 10609 9027
rect 8168 8996 10364 9024
rect 10520 8996 10609 9024
rect 8168 8984 8174 8996
rect 4062 8956 4068 8968
rect 4023 8928 4068 8956
rect 4062 8916 4068 8928
rect 4120 8956 4126 8968
rect 6086 8956 6092 8968
rect 4120 8928 6092 8956
rect 4120 8916 4126 8928
rect 6086 8916 6092 8928
rect 6144 8916 6150 8968
rect 6270 8956 6276 8968
rect 6183 8928 6276 8956
rect 6270 8916 6276 8928
rect 6328 8956 6334 8968
rect 10410 8956 10416 8968
rect 6328 8928 10416 8956
rect 6328 8916 6334 8928
rect 10410 8916 10416 8928
rect 10468 8916 10474 8968
rect 7834 8888 7840 8900
rect 7747 8860 7840 8888
rect 7834 8848 7840 8860
rect 7892 8888 7898 8900
rect 8662 8888 8668 8900
rect 7892 8860 8668 8888
rect 7892 8848 7898 8860
rect 8662 8848 8668 8860
rect 8720 8848 8726 8900
rect 9858 8848 9864 8900
rect 9916 8888 9922 8900
rect 10520 8888 10548 8996
rect 10597 8993 10609 8996
rect 10643 8993 10655 9027
rect 10597 8987 10655 8993
rect 10962 8984 10968 9036
rect 11020 9024 11026 9036
rect 11057 9027 11115 9033
rect 11057 9024 11069 9027
rect 11020 8996 11069 9024
rect 11020 8984 11026 8996
rect 11057 8993 11069 8996
rect 11103 8993 11115 9027
rect 14090 9024 14096 9036
rect 14051 8996 14096 9024
rect 11057 8987 11115 8993
rect 14090 8984 14096 8996
rect 14148 8984 14154 9036
rect 17310 8984 17316 9036
rect 17368 9024 17374 9036
rect 17773 9027 17831 9033
rect 17773 9024 17785 9027
rect 17368 8996 17785 9024
rect 17368 8984 17374 8996
rect 17773 8993 17785 8996
rect 17819 8993 17831 9027
rect 17773 8987 17831 8993
rect 17920 9027 17978 9033
rect 17920 8993 17932 9027
rect 17966 9024 17978 9027
rect 18690 9024 18696 9036
rect 17966 8996 18696 9024
rect 17966 8993 17978 8996
rect 17920 8987 17978 8993
rect 18690 8984 18696 8996
rect 18748 8984 18754 9036
rect 18782 8984 18788 9036
rect 18840 9024 18846 9036
rect 19337 9027 19395 9033
rect 19337 9024 19349 9027
rect 18840 8996 19349 9024
rect 18840 8984 18846 8996
rect 19337 8993 19349 8996
rect 19383 8993 19395 9027
rect 19337 8987 19395 8993
rect 12526 8916 12532 8968
rect 12584 8956 12590 8968
rect 12805 8959 12863 8965
rect 12805 8956 12817 8959
rect 12584 8928 12817 8956
rect 12584 8916 12590 8928
rect 12805 8925 12817 8928
rect 12851 8956 12863 8959
rect 16298 8956 16304 8968
rect 12851 8928 13814 8956
rect 16259 8928 16304 8956
rect 12851 8925 12863 8928
rect 12805 8919 12863 8925
rect 9916 8860 10548 8888
rect 9916 8848 9922 8860
rect 10594 8848 10600 8900
rect 10652 8888 10658 8900
rect 11238 8888 11244 8900
rect 10652 8860 11244 8888
rect 10652 8848 10658 8860
rect 11238 8848 11244 8860
rect 11296 8848 11302 8900
rect 13786 8888 13814 8928
rect 16298 8916 16304 8928
rect 16356 8916 16362 8968
rect 16758 8956 16764 8968
rect 16719 8928 16764 8956
rect 16758 8916 16764 8928
rect 16816 8916 16822 8968
rect 17586 8956 17592 8968
rect 17547 8928 17592 8956
rect 17586 8916 17592 8928
rect 17644 8956 17650 8968
rect 18141 8959 18199 8965
rect 18141 8956 18153 8959
rect 17644 8928 18153 8956
rect 17644 8916 17650 8928
rect 18141 8925 18153 8928
rect 18187 8925 18199 8959
rect 18141 8919 18199 8925
rect 16776 8888 16804 8916
rect 13786 8860 16804 8888
rect 17313 8891 17371 8897
rect 17313 8857 17325 8891
rect 17359 8888 17371 8891
rect 18414 8888 18420 8900
rect 17359 8860 18420 8888
rect 17359 8857 17371 8860
rect 17313 8851 17371 8857
rect 18414 8848 18420 8860
rect 18472 8848 18478 8900
rect 1394 8780 1400 8832
rect 1452 8820 1458 8832
rect 2501 8823 2559 8829
rect 2501 8820 2513 8823
rect 1452 8792 2513 8820
rect 1452 8780 1458 8792
rect 2501 8789 2513 8792
rect 2547 8789 2559 8823
rect 2501 8783 2559 8789
rect 4522 8780 4528 8832
rect 4580 8820 4586 8832
rect 4985 8823 5043 8829
rect 4985 8820 4997 8823
rect 4580 8792 4997 8820
rect 4580 8780 4586 8792
rect 4985 8789 4997 8792
rect 5031 8789 5043 8823
rect 4985 8783 5043 8789
rect 5810 8780 5816 8832
rect 5868 8820 5874 8832
rect 8849 8823 8907 8829
rect 8849 8820 8861 8823
rect 5868 8792 8861 8820
rect 5868 8780 5874 8792
rect 8849 8789 8861 8792
rect 8895 8820 8907 8823
rect 9030 8820 9036 8832
rect 8895 8792 9036 8820
rect 8895 8789 8907 8792
rect 8849 8783 8907 8789
rect 9030 8780 9036 8792
rect 9088 8820 9094 8832
rect 10778 8820 10784 8832
rect 9088 8792 10784 8820
rect 9088 8780 9094 8792
rect 10778 8780 10784 8792
rect 10836 8780 10842 8832
rect 14277 8823 14335 8829
rect 14277 8789 14289 8823
rect 14323 8820 14335 8823
rect 15286 8820 15292 8832
rect 14323 8792 15292 8820
rect 14323 8789 14335 8792
rect 14277 8783 14335 8789
rect 15286 8780 15292 8792
rect 15344 8780 15350 8832
rect 18046 8820 18052 8832
rect 18007 8792 18052 8820
rect 18046 8780 18052 8792
rect 18104 8780 18110 8832
rect 18230 8820 18236 8832
rect 18191 8792 18236 8820
rect 18230 8780 18236 8792
rect 18288 8780 18294 8832
rect 18322 8780 18328 8832
rect 18380 8820 18386 8832
rect 18785 8823 18843 8829
rect 18785 8820 18797 8823
rect 18380 8792 18797 8820
rect 18380 8780 18386 8792
rect 18785 8789 18797 8792
rect 18831 8789 18843 8823
rect 18785 8783 18843 8789
rect 19150 8780 19156 8832
rect 19208 8820 19214 8832
rect 19521 8823 19579 8829
rect 19521 8820 19533 8823
rect 19208 8792 19533 8820
rect 19208 8780 19214 8792
rect 19521 8789 19533 8792
rect 19567 8789 19579 8823
rect 19521 8783 19579 8789
rect 1104 8730 20884 8752
rect 1104 8678 4648 8730
rect 4700 8678 4712 8730
rect 4764 8678 4776 8730
rect 4828 8678 4840 8730
rect 4892 8678 11982 8730
rect 12034 8678 12046 8730
rect 12098 8678 12110 8730
rect 12162 8678 12174 8730
rect 12226 8678 19315 8730
rect 19367 8678 19379 8730
rect 19431 8678 19443 8730
rect 19495 8678 19507 8730
rect 19559 8678 20884 8730
rect 1104 8656 20884 8678
rect 1673 8619 1731 8625
rect 1673 8585 1685 8619
rect 1719 8616 1731 8619
rect 1762 8616 1768 8628
rect 1719 8588 1768 8616
rect 1719 8585 1731 8588
rect 1673 8579 1731 8585
rect 1762 8576 1768 8588
rect 1820 8576 1826 8628
rect 2866 8616 2872 8628
rect 2827 8588 2872 8616
rect 2866 8576 2872 8588
rect 2924 8576 2930 8628
rect 3421 8619 3479 8625
rect 3421 8585 3433 8619
rect 3467 8616 3479 8619
rect 4062 8616 4068 8628
rect 3467 8588 4068 8616
rect 3467 8585 3479 8588
rect 3421 8579 3479 8585
rect 4062 8576 4068 8588
rect 4120 8576 4126 8628
rect 5902 8616 5908 8628
rect 5863 8588 5908 8616
rect 5902 8576 5908 8588
rect 5960 8576 5966 8628
rect 5994 8576 6000 8628
rect 6052 8616 6058 8628
rect 6457 8619 6515 8625
rect 6457 8616 6469 8619
rect 6052 8588 6469 8616
rect 6052 8576 6058 8588
rect 6457 8585 6469 8588
rect 6503 8616 6515 8619
rect 6549 8619 6607 8625
rect 6549 8616 6561 8619
rect 6503 8588 6561 8616
rect 6503 8585 6515 8588
rect 6457 8579 6515 8585
rect 6549 8585 6561 8588
rect 6595 8585 6607 8619
rect 6549 8579 6607 8585
rect 7558 8576 7564 8628
rect 7616 8616 7622 8628
rect 7834 8616 7840 8628
rect 7616 8588 7840 8616
rect 7616 8576 7622 8588
rect 7834 8576 7840 8588
rect 7892 8576 7898 8628
rect 8202 8616 8208 8628
rect 8163 8588 8208 8616
rect 8202 8576 8208 8588
rect 8260 8576 8266 8628
rect 8938 8576 8944 8628
rect 8996 8616 9002 8628
rect 9858 8616 9864 8628
rect 8996 8588 9864 8616
rect 8996 8576 9002 8588
rect 9858 8576 9864 8588
rect 9916 8616 9922 8628
rect 10045 8619 10103 8625
rect 10045 8616 10057 8619
rect 9916 8588 10057 8616
rect 9916 8576 9922 8588
rect 10045 8585 10057 8588
rect 10091 8585 10103 8619
rect 10045 8579 10103 8585
rect 11885 8619 11943 8625
rect 11885 8585 11897 8619
rect 11931 8616 11943 8619
rect 12710 8616 12716 8628
rect 11931 8588 12716 8616
rect 11931 8585 11943 8588
rect 11885 8579 11943 8585
rect 4982 8548 4988 8560
rect 4943 8520 4988 8548
rect 4982 8508 4988 8520
rect 5040 8508 5046 8560
rect 5537 8551 5595 8557
rect 5537 8517 5549 8551
rect 5583 8548 5595 8551
rect 6270 8548 6276 8560
rect 5583 8520 6276 8548
rect 5583 8517 5595 8520
rect 5537 8511 5595 8517
rect 6270 8508 6276 8520
rect 6328 8508 6334 8560
rect 6822 8508 6828 8560
rect 6880 8548 6886 8560
rect 6917 8551 6975 8557
rect 6917 8548 6929 8551
rect 6880 8520 6929 8548
rect 6880 8508 6886 8520
rect 6917 8517 6929 8520
rect 6963 8517 6975 8551
rect 6917 8511 6975 8517
rect 2406 8480 2412 8492
rect 2367 8452 2412 8480
rect 2406 8440 2412 8452
rect 2464 8440 2470 8492
rect 3789 8483 3847 8489
rect 3789 8449 3801 8483
rect 3835 8480 3847 8483
rect 4522 8480 4528 8492
rect 3835 8452 4528 8480
rect 3835 8449 3847 8452
rect 3789 8443 3847 8449
rect 4522 8440 4528 8452
rect 4580 8440 4586 8492
rect 6086 8440 6092 8492
rect 6144 8480 6150 8492
rect 8941 8483 8999 8489
rect 8941 8480 8953 8483
rect 6144 8452 8953 8480
rect 6144 8440 6150 8452
rect 8941 8449 8953 8452
rect 8987 8449 8999 8483
rect 8941 8443 8999 8449
rect 10597 8483 10655 8489
rect 10597 8449 10609 8483
rect 10643 8480 10655 8483
rect 11900 8480 11928 8579
rect 12710 8576 12716 8588
rect 12768 8576 12774 8628
rect 13909 8619 13967 8625
rect 13909 8585 13921 8619
rect 13955 8616 13967 8619
rect 14090 8616 14096 8628
rect 13955 8588 14096 8616
rect 13955 8585 13967 8588
rect 13909 8579 13967 8585
rect 14090 8576 14096 8588
rect 14148 8576 14154 8628
rect 15933 8619 15991 8625
rect 15933 8585 15945 8619
rect 15979 8616 15991 8619
rect 16390 8616 16396 8628
rect 15979 8588 16396 8616
rect 15979 8585 15991 8588
rect 15933 8579 15991 8585
rect 16390 8576 16396 8588
rect 16448 8576 16454 8628
rect 17865 8619 17923 8625
rect 17865 8585 17877 8619
rect 17911 8616 17923 8619
rect 18046 8616 18052 8628
rect 17911 8588 18052 8616
rect 17911 8585 17923 8588
rect 17865 8579 17923 8585
rect 18046 8576 18052 8588
rect 18104 8576 18110 8628
rect 18782 8576 18788 8628
rect 18840 8616 18846 8628
rect 19337 8619 19395 8625
rect 19337 8616 19349 8619
rect 18840 8588 19349 8616
rect 18840 8576 18846 8588
rect 19337 8585 19349 8588
rect 19383 8616 19395 8619
rect 19978 8616 19984 8628
rect 19383 8588 19984 8616
rect 19383 8585 19395 8588
rect 19337 8579 19395 8585
rect 19978 8576 19984 8588
rect 20036 8576 20042 8628
rect 12894 8548 12900 8560
rect 12544 8520 12900 8548
rect 12544 8489 12572 8520
rect 12894 8508 12900 8520
rect 12952 8548 12958 8560
rect 15565 8551 15623 8557
rect 12952 8520 14412 8548
rect 12952 8508 12958 8520
rect 10643 8452 11928 8480
rect 12529 8483 12587 8489
rect 10643 8449 10655 8452
rect 10597 8443 10655 8449
rect 12529 8449 12541 8483
rect 12575 8449 12587 8483
rect 12529 8443 12587 8449
rect 13173 8483 13231 8489
rect 13173 8449 13185 8483
rect 13219 8480 13231 8483
rect 13354 8480 13360 8492
rect 13219 8452 13360 8480
rect 13219 8449 13231 8452
rect 13173 8443 13231 8449
rect 13354 8440 13360 8452
rect 13412 8440 13418 8492
rect 14093 8483 14151 8489
rect 14093 8449 14105 8483
rect 14139 8480 14151 8483
rect 14274 8480 14280 8492
rect 14139 8452 14280 8480
rect 14139 8449 14151 8452
rect 14093 8443 14151 8449
rect 14274 8440 14280 8452
rect 14332 8440 14338 8492
rect 14384 8489 14412 8520
rect 15565 8517 15577 8551
rect 15611 8548 15623 8551
rect 16206 8548 16212 8560
rect 15611 8520 16212 8548
rect 15611 8517 15623 8520
rect 15565 8511 15623 8517
rect 16206 8508 16212 8520
rect 16264 8508 16270 8560
rect 16298 8508 16304 8560
rect 16356 8548 16362 8560
rect 16356 8520 19242 8548
rect 16356 8508 16362 8520
rect 14369 8483 14427 8489
rect 14369 8449 14381 8483
rect 14415 8480 14427 8483
rect 16761 8483 16819 8489
rect 16761 8480 16773 8483
rect 14415 8452 16773 8480
rect 14415 8449 14427 8452
rect 14369 8443 14427 8449
rect 16761 8449 16773 8452
rect 16807 8480 16819 8483
rect 17402 8480 17408 8492
rect 16807 8452 17408 8480
rect 16807 8449 16819 8452
rect 16761 8443 16819 8449
rect 17402 8440 17408 8452
rect 17460 8440 17466 8492
rect 18141 8483 18199 8489
rect 18141 8449 18153 8483
rect 18187 8480 18199 8483
rect 18414 8480 18420 8492
rect 18187 8452 18420 8480
rect 18187 8449 18199 8452
rect 18141 8443 18199 8449
rect 18414 8440 18420 8452
rect 18472 8440 18478 8492
rect 18598 8480 18604 8492
rect 18559 8452 18604 8480
rect 18598 8440 18604 8452
rect 18656 8440 18662 8492
rect 6457 8415 6515 8421
rect 6457 8381 6469 8415
rect 6503 8412 6515 8415
rect 6825 8415 6883 8421
rect 6825 8412 6837 8415
rect 6503 8384 6837 8412
rect 6503 8381 6515 8384
rect 6457 8375 6515 8381
rect 6825 8381 6837 8384
rect 6871 8381 6883 8415
rect 7098 8412 7104 8424
rect 7059 8384 7104 8412
rect 6825 8375 6883 8381
rect 7098 8372 7104 8384
rect 7156 8372 7162 8424
rect 7561 8415 7619 8421
rect 7561 8381 7573 8415
rect 7607 8412 7619 8415
rect 7742 8412 7748 8424
rect 7607 8384 7748 8412
rect 7607 8381 7619 8384
rect 7561 8375 7619 8381
rect 7742 8372 7748 8384
rect 7800 8372 7806 8424
rect 8662 8412 8668 8424
rect 8623 8384 8668 8412
rect 8662 8372 8668 8384
rect 8720 8372 8726 8424
rect 8849 8415 8907 8421
rect 8849 8381 8861 8415
rect 8895 8381 8907 8415
rect 8849 8375 8907 8381
rect 11517 8415 11575 8421
rect 11517 8381 11529 8415
rect 11563 8412 11575 8415
rect 12161 8415 12219 8421
rect 12161 8412 12173 8415
rect 11563 8384 12173 8412
rect 11563 8381 11575 8384
rect 11517 8375 11575 8381
rect 12161 8381 12173 8384
rect 12207 8381 12219 8415
rect 12161 8375 12219 8381
rect 1946 8344 1952 8356
rect 1907 8316 1952 8344
rect 1946 8304 1952 8316
rect 2004 8304 2010 8356
rect 2041 8347 2099 8353
rect 2041 8313 2053 8347
rect 2087 8344 2099 8347
rect 2314 8344 2320 8356
rect 2087 8316 2320 8344
rect 2087 8313 2099 8316
rect 2041 8307 2099 8313
rect 2314 8304 2320 8316
rect 2372 8304 2378 8356
rect 4430 8344 4436 8356
rect 4391 8316 4436 8344
rect 4430 8304 4436 8316
rect 4488 8304 4494 8356
rect 4522 8304 4528 8356
rect 4580 8344 4586 8356
rect 6273 8347 6331 8353
rect 4580 8316 4625 8344
rect 4580 8304 4586 8316
rect 6273 8313 6285 8347
rect 6319 8344 6331 8347
rect 7116 8344 7144 8372
rect 6319 8316 7144 8344
rect 6319 8313 6331 8316
rect 6273 8307 6331 8313
rect 8202 8304 8208 8356
rect 8260 8344 8266 8356
rect 8864 8344 8892 8375
rect 10686 8344 10692 8356
rect 8260 8316 8892 8344
rect 9294 8316 10692 8344
rect 8260 8304 8266 8316
rect 4062 8276 4068 8288
rect 4023 8248 4068 8276
rect 4062 8236 4068 8248
rect 4120 8236 4126 8288
rect 4154 8236 4160 8288
rect 4212 8276 4218 8288
rect 9294 8276 9322 8316
rect 10686 8304 10692 8316
rect 10744 8304 10750 8356
rect 10918 8347 10976 8353
rect 10918 8313 10930 8347
rect 10964 8313 10976 8347
rect 10918 8307 10976 8313
rect 4212 8248 9322 8276
rect 9493 8279 9551 8285
rect 4212 8236 4218 8248
rect 9493 8245 9505 8279
rect 9539 8276 9551 8279
rect 9582 8276 9588 8288
rect 9539 8248 9588 8276
rect 9539 8245 9551 8248
rect 9493 8239 9551 8245
rect 9582 8236 9588 8248
rect 9640 8236 9646 8288
rect 10505 8279 10563 8285
rect 10505 8245 10517 8279
rect 10551 8276 10563 8279
rect 10933 8276 10961 8307
rect 11606 8276 11612 8288
rect 10551 8248 11612 8276
rect 10551 8245 10563 8248
rect 10505 8239 10563 8245
rect 11606 8236 11612 8248
rect 11664 8236 11670 8288
rect 12176 8276 12204 8375
rect 14734 8372 14740 8424
rect 14792 8412 14798 8424
rect 16298 8412 16304 8424
rect 14792 8384 16304 8412
rect 14792 8372 14798 8384
rect 16298 8372 16304 8384
rect 16356 8372 16362 8424
rect 19214 8412 19242 8520
rect 19648 8415 19706 8421
rect 19648 8412 19660 8415
rect 19214 8384 19660 8412
rect 19648 8381 19660 8384
rect 19694 8412 19706 8415
rect 20073 8415 20131 8421
rect 20073 8412 20085 8415
rect 19694 8384 20085 8412
rect 19694 8381 19706 8384
rect 19648 8375 19706 8381
rect 20073 8381 20085 8384
rect 20119 8381 20131 8415
rect 20073 8375 20131 8381
rect 12621 8347 12679 8353
rect 12621 8313 12633 8347
rect 12667 8313 12679 8347
rect 14185 8347 14243 8353
rect 12621 8307 12679 8313
rect 13786 8316 13952 8344
rect 12636 8276 12664 8307
rect 13538 8276 13544 8288
rect 12176 8248 12664 8276
rect 13499 8248 13544 8276
rect 13538 8236 13544 8248
rect 13596 8276 13602 8288
rect 13786 8276 13814 8316
rect 13596 8248 13814 8276
rect 13924 8276 13952 8316
rect 14185 8313 14197 8347
rect 14231 8313 14243 8347
rect 14185 8307 14243 8313
rect 14200 8276 14228 8307
rect 16114 8304 16120 8356
rect 16172 8344 16178 8356
rect 16482 8344 16488 8356
rect 16172 8316 16488 8344
rect 16172 8304 16178 8316
rect 16482 8304 16488 8316
rect 16540 8304 16546 8356
rect 16577 8347 16635 8353
rect 16577 8313 16589 8347
rect 16623 8313 16635 8347
rect 16577 8307 16635 8313
rect 18233 8347 18291 8353
rect 18233 8313 18245 8347
rect 18279 8344 18291 8347
rect 18322 8344 18328 8356
rect 18279 8316 18328 8344
rect 18279 8313 18291 8316
rect 18233 8307 18291 8313
rect 16298 8276 16304 8288
rect 13924 8248 14228 8276
rect 16259 8248 16304 8276
rect 13596 8236 13602 8248
rect 16298 8236 16304 8248
rect 16356 8276 16362 8288
rect 16592 8276 16620 8307
rect 18322 8304 18328 8316
rect 18380 8304 18386 8356
rect 18414 8304 18420 8356
rect 18472 8344 18478 8356
rect 19751 8347 19809 8353
rect 19751 8344 19763 8347
rect 18472 8316 19763 8344
rect 18472 8304 18478 8316
rect 19751 8313 19763 8316
rect 19797 8313 19809 8347
rect 19751 8307 19809 8313
rect 16356 8248 16620 8276
rect 16356 8236 16362 8248
rect 17310 8236 17316 8288
rect 17368 8276 17374 8288
rect 17405 8279 17463 8285
rect 17405 8276 17417 8279
rect 17368 8248 17417 8276
rect 17368 8236 17374 8248
rect 17405 8245 17417 8248
rect 17451 8245 17463 8279
rect 17405 8239 17463 8245
rect 1104 8186 20884 8208
rect 1104 8134 8315 8186
rect 8367 8134 8379 8186
rect 8431 8134 8443 8186
rect 8495 8134 8507 8186
rect 8559 8134 15648 8186
rect 15700 8134 15712 8186
rect 15764 8134 15776 8186
rect 15828 8134 15840 8186
rect 15892 8134 20884 8186
rect 1104 8112 20884 8134
rect 3050 8072 3056 8084
rect 3011 8044 3056 8072
rect 3050 8032 3056 8044
rect 3108 8032 3114 8084
rect 3326 8072 3332 8084
rect 3287 8044 3332 8072
rect 3326 8032 3332 8044
rect 3384 8032 3390 8084
rect 4246 8072 4252 8084
rect 4207 8044 4252 8072
rect 4246 8032 4252 8044
rect 4304 8032 4310 8084
rect 4430 8032 4436 8084
rect 4488 8072 4494 8084
rect 5169 8075 5227 8081
rect 5169 8072 5181 8075
rect 4488 8044 5181 8072
rect 4488 8032 4494 8044
rect 5169 8041 5181 8044
rect 5215 8072 5227 8075
rect 6914 8072 6920 8084
rect 5215 8044 6920 8072
rect 5215 8041 5227 8044
rect 5169 8035 5227 8041
rect 6914 8032 6920 8044
rect 6972 8032 6978 8084
rect 7466 8072 7472 8084
rect 7392 8044 7472 8072
rect 1759 8007 1817 8013
rect 1759 7973 1771 8007
rect 1805 8004 1817 8007
rect 1854 8004 1860 8016
rect 1805 7976 1860 8004
rect 1805 7973 1817 7976
rect 1759 7967 1817 7973
rect 1854 7964 1860 7976
rect 1912 7964 1918 8016
rect 1946 7964 1952 8016
rect 2004 8004 2010 8016
rect 3697 8007 3755 8013
rect 3697 8004 3709 8007
rect 2004 7976 3709 8004
rect 2004 7964 2010 7976
rect 3697 7973 3709 7976
rect 3743 8004 3755 8007
rect 5258 8004 5264 8016
rect 3743 7976 5264 8004
rect 3743 7973 3755 7976
rect 3697 7967 3755 7973
rect 5258 7964 5264 7976
rect 5316 7964 5322 8016
rect 5994 8004 6000 8016
rect 5368 7976 6000 8004
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7936 1455 7939
rect 1578 7936 1584 7948
rect 1443 7908 1584 7936
rect 1443 7905 1455 7908
rect 1397 7899 1455 7905
rect 1578 7896 1584 7908
rect 1636 7896 1642 7948
rect 4065 7939 4123 7945
rect 4065 7905 4077 7939
rect 4111 7936 4123 7939
rect 4154 7936 4160 7948
rect 4111 7908 4160 7936
rect 4111 7905 4123 7908
rect 4065 7899 4123 7905
rect 4154 7896 4160 7908
rect 4212 7896 4218 7948
rect 5368 7945 5396 7976
rect 5994 7964 6000 7976
rect 6052 7964 6058 8016
rect 6549 8007 6607 8013
rect 6549 8004 6561 8007
rect 6104 7976 6561 8004
rect 5353 7939 5411 7945
rect 5353 7905 5365 7939
rect 5399 7905 5411 7939
rect 5353 7899 5411 7905
rect 5442 7896 5448 7948
rect 5500 7936 5506 7948
rect 5721 7939 5779 7945
rect 5721 7936 5733 7939
rect 5500 7908 5733 7936
rect 5500 7896 5506 7908
rect 5721 7905 5733 7908
rect 5767 7905 5779 7939
rect 5721 7899 5779 7905
rect 5810 7896 5816 7948
rect 5868 7936 5874 7948
rect 6104 7936 6132 7976
rect 6549 7973 6561 7976
rect 6595 8004 6607 8007
rect 7392 8004 7420 8044
rect 7466 8032 7472 8044
rect 7524 8032 7530 8084
rect 8110 8032 8116 8084
rect 8168 8072 8174 8084
rect 8389 8075 8447 8081
rect 8389 8072 8401 8075
rect 8168 8044 8401 8072
rect 8168 8032 8174 8044
rect 8389 8041 8401 8044
rect 8435 8041 8447 8075
rect 8389 8035 8447 8041
rect 8662 8032 8668 8084
rect 8720 8072 8726 8084
rect 8757 8075 8815 8081
rect 8757 8072 8769 8075
rect 8720 8044 8769 8072
rect 8720 8032 8726 8044
rect 8757 8041 8769 8044
rect 8803 8072 8815 8075
rect 9490 8072 9496 8084
rect 8803 8044 9496 8072
rect 8803 8041 8815 8044
rect 8757 8035 8815 8041
rect 9490 8032 9496 8044
rect 9548 8032 9554 8084
rect 10689 8075 10747 8081
rect 10689 8041 10701 8075
rect 10735 8072 10747 8075
rect 10962 8072 10968 8084
rect 10735 8044 10968 8072
rect 10735 8041 10747 8044
rect 10689 8035 10747 8041
rect 10962 8032 10968 8044
rect 11020 8032 11026 8084
rect 12529 8075 12587 8081
rect 12529 8041 12541 8075
rect 12575 8072 12587 8075
rect 12618 8072 12624 8084
rect 12575 8044 12624 8072
rect 12575 8041 12587 8044
rect 12529 8035 12587 8041
rect 12618 8032 12624 8044
rect 12676 8032 12682 8084
rect 12894 8072 12900 8084
rect 12855 8044 12900 8072
rect 12894 8032 12900 8044
rect 12952 8032 12958 8084
rect 14274 8032 14280 8084
rect 14332 8072 14338 8084
rect 14369 8075 14427 8081
rect 14369 8072 14381 8075
rect 14332 8044 14381 8072
rect 14332 8032 14338 8044
rect 14369 8041 14381 8044
rect 14415 8041 14427 8075
rect 16482 8072 16488 8084
rect 16443 8044 16488 8072
rect 14369 8035 14427 8041
rect 16482 8032 16488 8044
rect 16540 8032 16546 8084
rect 16574 8032 16580 8084
rect 16632 8072 16638 8084
rect 18693 8075 18751 8081
rect 18693 8072 18705 8075
rect 16632 8044 18705 8072
rect 16632 8032 16638 8044
rect 18693 8041 18705 8044
rect 18739 8041 18751 8075
rect 18693 8035 18751 8041
rect 6595 7976 7420 8004
rect 11327 8007 11385 8013
rect 6595 7973 6607 7976
rect 6549 7967 6607 7973
rect 11327 7973 11339 8007
rect 11373 8004 11385 8007
rect 11606 8004 11612 8016
rect 11373 7976 11612 8004
rect 11373 7973 11385 7976
rect 11327 7967 11385 7973
rect 11606 7964 11612 7976
rect 11664 7964 11670 8016
rect 13535 8007 13593 8013
rect 13535 7973 13547 8007
rect 13581 8004 13593 8007
rect 13998 8004 14004 8016
rect 13581 7976 14004 8004
rect 13581 7973 13593 7976
rect 13535 7967 13593 7973
rect 13998 7964 14004 7976
rect 14056 7964 14062 8016
rect 15378 7964 15384 8016
rect 15436 8004 15442 8016
rect 15610 8007 15668 8013
rect 15610 8004 15622 8007
rect 15436 7976 15622 8004
rect 15436 7964 15442 7976
rect 15610 7973 15622 7976
rect 15656 7973 15668 8007
rect 17126 8004 17132 8016
rect 17087 7976 17132 8004
rect 15610 7967 15668 7973
rect 17126 7964 17132 7976
rect 17184 7964 17190 8016
rect 17218 7964 17224 8016
rect 17276 8004 17282 8016
rect 18322 8004 18328 8016
rect 17276 7976 18328 8004
rect 17276 7964 17282 7976
rect 18322 7964 18328 7976
rect 18380 7964 18386 8016
rect 5868 7908 6132 7936
rect 6365 7939 6423 7945
rect 5868 7896 5874 7908
rect 6365 7905 6377 7939
rect 6411 7936 6423 7939
rect 6454 7936 6460 7948
rect 6411 7908 6460 7936
rect 6411 7905 6423 7908
rect 6365 7899 6423 7905
rect 6454 7896 6460 7908
rect 6512 7896 6518 7948
rect 7285 7939 7343 7945
rect 7285 7905 7297 7939
rect 7331 7936 7343 7939
rect 7377 7939 7435 7945
rect 7377 7936 7389 7939
rect 7331 7908 7389 7936
rect 7331 7905 7343 7908
rect 7285 7899 7343 7905
rect 7377 7905 7389 7908
rect 7423 7936 7435 7939
rect 7466 7936 7472 7948
rect 7423 7908 7472 7936
rect 7423 7905 7435 7908
rect 7377 7899 7435 7905
rect 7466 7896 7472 7908
rect 7524 7896 7530 7948
rect 9214 7936 9220 7948
rect 7668 7908 9220 7936
rect 4801 7871 4859 7877
rect 4801 7837 4813 7871
rect 4847 7868 4859 7871
rect 4982 7868 4988 7880
rect 4847 7840 4988 7868
rect 4847 7837 4859 7840
rect 4801 7831 4859 7837
rect 4982 7828 4988 7840
rect 5040 7868 5046 7880
rect 7668 7868 7696 7908
rect 9214 7896 9220 7908
rect 9272 7896 9278 7948
rect 10020 7939 10078 7945
rect 10020 7905 10032 7939
rect 10066 7936 10078 7939
rect 10226 7936 10232 7948
rect 10066 7908 10232 7936
rect 10066 7905 10078 7908
rect 10020 7899 10078 7905
rect 10226 7896 10232 7908
rect 10284 7896 10290 7948
rect 10965 7939 11023 7945
rect 10965 7905 10977 7939
rect 11011 7936 11023 7939
rect 11146 7936 11152 7948
rect 11011 7908 11152 7936
rect 11011 7905 11023 7908
rect 10965 7899 11023 7905
rect 11146 7896 11152 7908
rect 11204 7936 11210 7948
rect 12802 7936 12808 7948
rect 11204 7908 12808 7936
rect 11204 7896 11210 7908
rect 12802 7896 12808 7908
rect 12860 7896 12866 7948
rect 14918 7936 14924 7948
rect 12906 7908 14924 7936
rect 5040 7840 7696 7868
rect 7745 7871 7803 7877
rect 5040 7828 5046 7840
rect 7745 7837 7757 7871
rect 7791 7837 7803 7871
rect 7745 7831 7803 7837
rect 8113 7871 8171 7877
rect 8113 7837 8125 7871
rect 8159 7868 8171 7871
rect 9122 7868 9128 7880
rect 8159 7840 9128 7868
rect 8159 7837 8171 7840
rect 8113 7831 8171 7837
rect 7098 7760 7104 7812
rect 7156 7800 7162 7812
rect 7515 7803 7573 7809
rect 7515 7800 7527 7803
rect 7156 7772 7527 7800
rect 7156 7760 7162 7772
rect 7515 7769 7527 7772
rect 7561 7769 7573 7803
rect 7760 7800 7788 7831
rect 9122 7828 9128 7840
rect 9180 7828 9186 7880
rect 10778 7828 10784 7880
rect 10836 7868 10842 7880
rect 12906 7868 12934 7908
rect 14918 7896 14924 7908
rect 14976 7896 14982 7948
rect 15010 7896 15016 7948
rect 15068 7936 15074 7948
rect 15289 7939 15347 7945
rect 15289 7936 15301 7939
rect 15068 7908 15301 7936
rect 15068 7896 15074 7908
rect 15289 7905 15301 7908
rect 15335 7905 15347 7939
rect 15289 7899 15347 7905
rect 18138 7896 18144 7948
rect 18196 7936 18202 7948
rect 18601 7939 18659 7945
rect 18601 7936 18613 7939
rect 18196 7908 18613 7936
rect 18196 7896 18202 7908
rect 18601 7905 18613 7908
rect 18647 7905 18659 7939
rect 19058 7936 19064 7948
rect 19019 7908 19064 7936
rect 18601 7899 18659 7905
rect 19058 7896 19064 7908
rect 19116 7896 19122 7948
rect 13170 7868 13176 7880
rect 10836 7840 12934 7868
rect 13131 7840 13176 7868
rect 10836 7828 10842 7840
rect 13170 7828 13176 7840
rect 13228 7828 13234 7880
rect 17402 7868 17408 7880
rect 17363 7840 17408 7868
rect 17402 7828 17408 7840
rect 17460 7828 17466 7880
rect 17494 7828 17500 7880
rect 17552 7868 17558 7880
rect 18049 7871 18107 7877
rect 18049 7868 18061 7871
rect 17552 7840 18061 7868
rect 17552 7828 17558 7840
rect 18049 7837 18061 7840
rect 18095 7868 18107 7871
rect 18322 7868 18328 7880
rect 18095 7840 18328 7868
rect 18095 7837 18107 7840
rect 18049 7831 18107 7837
rect 18322 7828 18328 7840
rect 18380 7828 18386 7880
rect 8386 7800 8392 7812
rect 7760 7772 8392 7800
rect 7515 7763 7573 7769
rect 8386 7760 8392 7772
rect 8444 7800 8450 7812
rect 9030 7800 9036 7812
rect 8444 7772 9036 7800
rect 8444 7760 8450 7772
rect 9030 7760 9036 7772
rect 9088 7760 9094 7812
rect 11882 7800 11888 7812
rect 11843 7772 11888 7800
rect 11882 7760 11888 7772
rect 11940 7760 11946 7812
rect 16209 7803 16267 7809
rect 16209 7769 16221 7803
rect 16255 7800 16267 7803
rect 17218 7800 17224 7812
rect 16255 7772 17224 7800
rect 16255 7769 16267 7772
rect 16209 7763 16267 7769
rect 17218 7760 17224 7772
rect 17276 7760 17282 7812
rect 2314 7732 2320 7744
rect 2275 7704 2320 7732
rect 2314 7692 2320 7704
rect 2372 7732 2378 7744
rect 2593 7735 2651 7741
rect 2593 7732 2605 7735
rect 2372 7704 2605 7732
rect 2372 7692 2378 7704
rect 2593 7701 2605 7704
rect 2639 7701 2651 7735
rect 6822 7732 6828 7744
rect 6783 7704 6828 7732
rect 2593 7695 2651 7701
rect 6822 7692 6828 7704
rect 6880 7692 6886 7744
rect 7653 7735 7711 7741
rect 7653 7701 7665 7735
rect 7699 7732 7711 7735
rect 8110 7732 8116 7744
rect 7699 7704 8116 7732
rect 7699 7701 7711 7704
rect 7653 7695 7711 7701
rect 8110 7692 8116 7704
rect 8168 7692 8174 7744
rect 10091 7735 10149 7741
rect 10091 7701 10103 7735
rect 10137 7732 10149 7735
rect 10502 7732 10508 7744
rect 10137 7704 10508 7732
rect 10137 7701 10149 7704
rect 10091 7695 10149 7701
rect 10502 7692 10508 7704
rect 10560 7692 10566 7744
rect 13538 7692 13544 7744
rect 13596 7732 13602 7744
rect 14093 7735 14151 7741
rect 14093 7732 14105 7735
rect 13596 7704 14105 7732
rect 13596 7692 13602 7704
rect 14093 7701 14105 7704
rect 14139 7701 14151 7735
rect 14093 7695 14151 7701
rect 15194 7692 15200 7744
rect 15252 7732 15258 7744
rect 18509 7735 18567 7741
rect 18509 7732 18521 7735
rect 15252 7704 18521 7732
rect 15252 7692 15258 7704
rect 18509 7701 18521 7704
rect 18555 7732 18567 7735
rect 18690 7732 18696 7744
rect 18555 7704 18696 7732
rect 18555 7701 18567 7704
rect 18509 7695 18567 7701
rect 18690 7692 18696 7704
rect 18748 7692 18754 7744
rect 1104 7642 20884 7664
rect 1104 7590 4648 7642
rect 4700 7590 4712 7642
rect 4764 7590 4776 7642
rect 4828 7590 4840 7642
rect 4892 7590 11982 7642
rect 12034 7590 12046 7642
rect 12098 7590 12110 7642
rect 12162 7590 12174 7642
rect 12226 7590 19315 7642
rect 19367 7590 19379 7642
rect 19431 7590 19443 7642
rect 19495 7590 19507 7642
rect 19559 7590 20884 7642
rect 1104 7568 20884 7590
rect 3326 7528 3332 7540
rect 2056 7500 3332 7528
rect 1489 7395 1547 7401
rect 1489 7361 1501 7395
rect 1535 7392 1547 7395
rect 2056 7392 2084 7500
rect 3326 7488 3332 7500
rect 3384 7488 3390 7540
rect 4154 7488 4160 7540
rect 4212 7528 4218 7540
rect 5810 7528 5816 7540
rect 4212 7500 4257 7528
rect 5723 7500 5816 7528
rect 4212 7488 4218 7500
rect 5810 7488 5816 7500
rect 5868 7528 5874 7540
rect 5994 7528 6000 7540
rect 5868 7500 6000 7528
rect 5868 7488 5874 7500
rect 5994 7488 6000 7500
rect 6052 7488 6058 7540
rect 7282 7488 7288 7540
rect 7340 7528 7346 7540
rect 8018 7528 8024 7540
rect 7340 7500 8024 7528
rect 7340 7488 7346 7500
rect 8018 7488 8024 7500
rect 8076 7488 8082 7540
rect 8386 7528 8392 7540
rect 8347 7500 8392 7528
rect 8386 7488 8392 7500
rect 8444 7488 8450 7540
rect 10226 7528 10232 7540
rect 10187 7500 10232 7528
rect 10226 7488 10232 7500
rect 10284 7488 10290 7540
rect 13170 7488 13176 7540
rect 13228 7528 13234 7540
rect 15197 7531 15255 7537
rect 13228 7500 14320 7528
rect 13228 7488 13234 7500
rect 2130 7420 2136 7472
rect 2188 7460 2194 7472
rect 7193 7463 7251 7469
rect 2188 7432 5120 7460
rect 2188 7420 2194 7432
rect 1535 7364 2084 7392
rect 2961 7395 3019 7401
rect 1535 7361 1547 7364
rect 1489 7355 1547 7361
rect 2961 7361 2973 7395
rect 3007 7392 3019 7395
rect 3050 7392 3056 7404
rect 3007 7364 3056 7392
rect 3007 7361 3019 7364
rect 2961 7355 3019 7361
rect 3050 7352 3056 7364
rect 3108 7352 3114 7404
rect 4801 7395 4859 7401
rect 4801 7361 4813 7395
rect 4847 7392 4859 7395
rect 4982 7392 4988 7404
rect 4847 7364 4988 7392
rect 4847 7361 4859 7364
rect 4801 7355 4859 7361
rect 4982 7352 4988 7364
rect 5040 7352 5046 7404
rect 5092 7401 5120 7432
rect 7193 7429 7205 7463
rect 7239 7460 7251 7463
rect 7558 7460 7564 7472
rect 7239 7432 7564 7460
rect 7239 7429 7251 7432
rect 7193 7423 7251 7429
rect 7558 7420 7564 7432
rect 7616 7460 7622 7472
rect 7653 7463 7711 7469
rect 7653 7460 7665 7463
rect 7616 7432 7665 7460
rect 7616 7420 7622 7432
rect 7653 7429 7665 7432
rect 7699 7429 7711 7463
rect 8404 7460 8432 7488
rect 7653 7423 7711 7429
rect 7760 7432 8432 7460
rect 8849 7463 8907 7469
rect 5077 7395 5135 7401
rect 5077 7361 5089 7395
rect 5123 7361 5135 7395
rect 5077 7355 5135 7361
rect 5902 7352 5908 7404
rect 5960 7392 5966 7404
rect 7760 7401 7788 7432
rect 8849 7429 8861 7463
rect 8895 7460 8907 7463
rect 9214 7460 9220 7472
rect 8895 7432 9220 7460
rect 8895 7429 8907 7432
rect 8849 7423 8907 7429
rect 9214 7420 9220 7432
rect 9272 7460 9278 7472
rect 10870 7460 10876 7472
rect 9272 7432 10876 7460
rect 9272 7420 9278 7432
rect 10870 7420 10876 7432
rect 10928 7420 10934 7472
rect 11882 7420 11888 7472
rect 11940 7460 11946 7472
rect 12161 7463 12219 7469
rect 12161 7460 12173 7463
rect 11940 7432 12173 7460
rect 11940 7420 11946 7432
rect 12161 7429 12173 7432
rect 12207 7460 12219 7463
rect 12618 7460 12624 7472
rect 12207 7432 12624 7460
rect 12207 7429 12219 7432
rect 12161 7423 12219 7429
rect 12618 7420 12624 7432
rect 12676 7420 12682 7472
rect 13446 7420 13452 7472
rect 13504 7460 13510 7472
rect 14185 7463 14243 7469
rect 14185 7460 14197 7463
rect 13504 7432 14197 7460
rect 13504 7420 13510 7432
rect 14185 7429 14197 7432
rect 14231 7429 14243 7463
rect 14185 7423 14243 7429
rect 6641 7395 6699 7401
rect 6641 7392 6653 7395
rect 5960 7364 6653 7392
rect 5960 7352 5966 7364
rect 6641 7361 6653 7364
rect 6687 7392 6699 7395
rect 7745 7395 7803 7401
rect 7745 7392 7757 7395
rect 6687 7364 7757 7392
rect 6687 7361 6699 7364
rect 6641 7355 6699 7361
rect 7745 7361 7757 7364
rect 7791 7361 7803 7395
rect 7745 7355 7803 7361
rect 8113 7395 8171 7401
rect 8113 7361 8125 7395
rect 8159 7392 8171 7395
rect 10597 7395 10655 7401
rect 10597 7392 10609 7395
rect 8159 7364 10609 7392
rect 8159 7361 8171 7364
rect 8113 7355 8171 7361
rect 10597 7361 10609 7364
rect 10643 7392 10655 7395
rect 10643 7364 11284 7392
rect 10643 7361 10655 7364
rect 10597 7355 10655 7361
rect 3881 7327 3939 7333
rect 3881 7293 3893 7327
rect 3927 7324 3939 7327
rect 4246 7324 4252 7336
rect 3927 7296 4252 7324
rect 3927 7293 3939 7296
rect 3881 7287 3939 7293
rect 4246 7284 4252 7296
rect 4304 7324 4310 7336
rect 4525 7327 4583 7333
rect 4525 7324 4537 7327
rect 4304 7296 4537 7324
rect 4304 7284 4310 7296
rect 4525 7293 4537 7296
rect 4571 7293 4583 7327
rect 4525 7287 4583 7293
rect 1581 7259 1639 7265
rect 1581 7225 1593 7259
rect 1627 7256 1639 7259
rect 2130 7256 2136 7268
rect 1627 7228 1802 7256
rect 2091 7228 2136 7256
rect 1627 7225 1639 7228
rect 1581 7219 1639 7225
rect 1774 7188 1802 7228
rect 2130 7216 2136 7228
rect 2188 7216 2194 7268
rect 3282 7259 3340 7265
rect 3282 7256 3294 7259
rect 2792 7228 3294 7256
rect 2792 7200 2820 7228
rect 3282 7225 3294 7228
rect 3328 7256 3340 7259
rect 4062 7256 4068 7268
rect 3328 7228 4068 7256
rect 3328 7225 3340 7228
rect 3282 7219 3340 7225
rect 4062 7216 4068 7228
rect 4120 7216 4126 7268
rect 2314 7188 2320 7200
rect 1774 7160 2320 7188
rect 2314 7148 2320 7160
rect 2372 7188 2378 7200
rect 2409 7191 2467 7197
rect 2409 7188 2421 7191
rect 2372 7160 2421 7188
rect 2372 7148 2378 7160
rect 2409 7157 2421 7160
rect 2455 7157 2467 7191
rect 2774 7188 2780 7200
rect 2735 7160 2780 7188
rect 2409 7151 2467 7157
rect 2774 7148 2780 7160
rect 2832 7148 2838 7200
rect 4540 7188 4568 7287
rect 6914 7284 6920 7336
rect 6972 7324 6978 7336
rect 7098 7324 7104 7336
rect 6972 7296 7104 7324
rect 6972 7284 6978 7296
rect 7098 7284 7104 7296
rect 7156 7324 7162 7336
rect 7524 7327 7582 7333
rect 7524 7324 7536 7327
rect 7156 7296 7536 7324
rect 7156 7284 7162 7296
rect 7524 7293 7536 7296
rect 7570 7324 7582 7327
rect 7834 7324 7840 7336
rect 7570 7296 7840 7324
rect 7570 7293 7582 7296
rect 7524 7287 7582 7293
rect 7834 7284 7840 7296
rect 7892 7324 7898 7336
rect 8662 7324 8668 7336
rect 7892 7296 8668 7324
rect 7892 7284 7898 7296
rect 8662 7284 8668 7296
rect 8720 7284 8726 7336
rect 8941 7327 8999 7333
rect 8941 7293 8953 7327
rect 8987 7324 8999 7327
rect 9030 7324 9036 7336
rect 8987 7296 9036 7324
rect 8987 7293 8999 7296
rect 8941 7287 8999 7293
rect 9030 7284 9036 7296
rect 9088 7324 9094 7336
rect 9674 7324 9680 7336
rect 9088 7296 9680 7324
rect 9088 7284 9094 7296
rect 9674 7284 9680 7296
rect 9732 7284 9738 7336
rect 10778 7324 10784 7336
rect 10739 7296 10784 7324
rect 10778 7284 10784 7296
rect 10836 7284 10842 7336
rect 11256 7333 11284 7364
rect 11422 7352 11428 7404
rect 11480 7392 11486 7404
rect 13173 7395 13231 7401
rect 13173 7392 13185 7395
rect 11480 7364 13185 7392
rect 11480 7352 11486 7364
rect 13173 7361 13185 7364
rect 13219 7392 13231 7395
rect 13354 7392 13360 7404
rect 13219 7364 13360 7392
rect 13219 7361 13231 7364
rect 13173 7355 13231 7361
rect 13354 7352 13360 7364
rect 13412 7352 13418 7404
rect 13909 7395 13967 7401
rect 13909 7361 13921 7395
rect 13955 7392 13967 7395
rect 14292 7392 14320 7500
rect 15197 7497 15209 7531
rect 15243 7528 15255 7531
rect 15378 7528 15384 7540
rect 15243 7500 15384 7528
rect 15243 7497 15255 7500
rect 15197 7491 15255 7497
rect 15378 7488 15384 7500
rect 15436 7488 15442 7540
rect 15470 7488 15476 7540
rect 15528 7528 15534 7540
rect 17405 7531 17463 7537
rect 17405 7528 17417 7531
rect 15528 7500 17417 7528
rect 15528 7488 15534 7500
rect 17405 7497 17417 7500
rect 17451 7497 17463 7531
rect 17405 7491 17463 7497
rect 17865 7531 17923 7537
rect 17865 7497 17877 7531
rect 17911 7528 17923 7531
rect 18046 7528 18052 7540
rect 17911 7500 18052 7528
rect 17911 7497 17923 7500
rect 17865 7491 17923 7497
rect 14645 7463 14703 7469
rect 14645 7429 14657 7463
rect 14691 7460 14703 7463
rect 14734 7460 14740 7472
rect 14691 7432 14740 7460
rect 14691 7429 14703 7432
rect 14645 7423 14703 7429
rect 14734 7420 14740 7432
rect 14792 7420 14798 7472
rect 15010 7420 15016 7472
rect 15068 7460 15074 7472
rect 16485 7463 16543 7469
rect 16485 7460 16497 7463
rect 15068 7432 16497 7460
rect 15068 7420 15074 7432
rect 16485 7429 16497 7432
rect 16531 7429 16543 7463
rect 16485 7423 16543 7429
rect 17129 7463 17187 7469
rect 17129 7429 17141 7463
rect 17175 7460 17187 7463
rect 17218 7460 17224 7472
rect 17175 7432 17224 7460
rect 17175 7429 17187 7432
rect 17129 7423 17187 7429
rect 17218 7420 17224 7432
rect 17276 7420 17282 7472
rect 16574 7392 16580 7404
rect 13955 7364 16580 7392
rect 13955 7361 13967 7364
rect 13909 7355 13967 7361
rect 16574 7352 16580 7364
rect 16632 7352 16638 7404
rect 11241 7327 11299 7333
rect 11241 7293 11253 7327
rect 11287 7324 11299 7327
rect 11330 7324 11336 7336
rect 11287 7296 11336 7324
rect 11287 7293 11299 7296
rect 11241 7287 11299 7293
rect 11330 7284 11336 7296
rect 11388 7284 11394 7336
rect 14001 7327 14059 7333
rect 14001 7293 14013 7327
rect 14047 7324 14059 7327
rect 14734 7324 14740 7336
rect 14047 7296 14740 7324
rect 14047 7293 14059 7296
rect 14001 7287 14059 7293
rect 14734 7284 14740 7296
rect 14792 7284 14798 7336
rect 15102 7284 15108 7336
rect 15160 7324 15166 7336
rect 15289 7327 15347 7333
rect 15289 7324 15301 7327
rect 15160 7296 15301 7324
rect 15160 7284 15166 7296
rect 15289 7293 15301 7296
rect 15335 7324 15347 7327
rect 15930 7324 15936 7336
rect 15335 7296 15936 7324
rect 15335 7293 15347 7296
rect 15289 7287 15347 7293
rect 15930 7284 15936 7296
rect 15988 7284 15994 7336
rect 16209 7327 16267 7333
rect 16209 7293 16221 7327
rect 16255 7324 16267 7327
rect 16298 7324 16304 7336
rect 16255 7296 16304 7324
rect 16255 7293 16267 7296
rect 16209 7287 16267 7293
rect 16298 7284 16304 7296
rect 16356 7324 16362 7336
rect 16850 7324 16856 7336
rect 16356 7296 16856 7324
rect 16356 7284 16362 7296
rect 16850 7284 16856 7296
rect 16908 7284 16914 7336
rect 17420 7324 17448 7491
rect 18046 7488 18052 7500
rect 18104 7488 18110 7540
rect 19058 7528 19064 7540
rect 19019 7500 19064 7528
rect 19058 7488 19064 7500
rect 19116 7488 19122 7540
rect 18064 7460 18092 7488
rect 18141 7463 18199 7469
rect 18141 7460 18153 7463
rect 18064 7432 18153 7460
rect 18141 7429 18153 7432
rect 18187 7429 18199 7463
rect 18141 7423 18199 7429
rect 17494 7352 17500 7404
rect 17552 7392 17558 7404
rect 19751 7395 19809 7401
rect 19751 7392 19763 7395
rect 17552 7364 19763 7392
rect 17552 7352 17558 7364
rect 19751 7361 19763 7364
rect 19797 7361 19809 7395
rect 19751 7355 19809 7361
rect 18049 7327 18107 7333
rect 18049 7324 18061 7327
rect 17420 7296 18061 7324
rect 18049 7293 18061 7296
rect 18095 7293 18107 7327
rect 18322 7324 18328 7336
rect 18283 7296 18328 7324
rect 18049 7287 18107 7293
rect 18322 7284 18328 7296
rect 18380 7284 18386 7336
rect 19610 7324 19616 7336
rect 19574 7296 19616 7324
rect 19610 7284 19616 7296
rect 19668 7333 19674 7336
rect 19668 7327 19722 7333
rect 19668 7293 19676 7327
rect 19710 7324 19722 7327
rect 19710 7296 20208 7324
rect 19710 7293 19722 7296
rect 19668 7287 19722 7293
rect 19668 7284 19674 7287
rect 4893 7259 4951 7265
rect 4893 7225 4905 7259
rect 4939 7225 4951 7259
rect 4893 7219 4951 7225
rect 7377 7259 7435 7265
rect 7377 7225 7389 7259
rect 7423 7225 7435 7259
rect 11514 7256 11520 7268
rect 11475 7228 11520 7256
rect 7377 7219 7435 7225
rect 4908 7188 4936 7219
rect 4540 7160 4936 7188
rect 6181 7191 6239 7197
rect 6181 7157 6193 7191
rect 6227 7188 6239 7191
rect 6454 7188 6460 7200
rect 6227 7160 6460 7188
rect 6227 7157 6239 7160
rect 6181 7151 6239 7157
rect 6454 7148 6460 7160
rect 6512 7148 6518 7200
rect 7392 7188 7420 7219
rect 11514 7216 11520 7228
rect 11572 7216 11578 7268
rect 12526 7256 12532 7268
rect 12487 7228 12532 7256
rect 12526 7216 12532 7228
rect 12584 7216 12590 7268
rect 12618 7216 12624 7268
rect 12676 7256 12682 7268
rect 12676 7228 12721 7256
rect 12676 7216 12682 7228
rect 15378 7216 15384 7268
rect 15436 7256 15442 7268
rect 15610 7259 15668 7265
rect 15610 7256 15622 7259
rect 15436 7228 15622 7256
rect 15436 7216 15442 7228
rect 15610 7225 15622 7228
rect 15656 7225 15668 7259
rect 18782 7256 18788 7268
rect 18743 7228 18788 7256
rect 15610 7219 15668 7225
rect 18782 7216 18788 7228
rect 18840 7216 18846 7268
rect 20180 7200 20208 7296
rect 7466 7188 7472 7200
rect 7392 7160 7472 7188
rect 7466 7148 7472 7160
rect 7524 7148 7530 7200
rect 9214 7148 9220 7200
rect 9272 7188 9278 7200
rect 9309 7191 9367 7197
rect 9309 7188 9321 7191
rect 9272 7160 9321 7188
rect 9272 7148 9278 7160
rect 9309 7157 9321 7160
rect 9355 7157 9367 7191
rect 9858 7188 9864 7200
rect 9819 7160 9864 7188
rect 9309 7151 9367 7157
rect 9858 7148 9864 7160
rect 9916 7148 9922 7200
rect 10870 7148 10876 7200
rect 10928 7188 10934 7200
rect 11606 7188 11612 7200
rect 10928 7160 11612 7188
rect 10928 7148 10934 7160
rect 11606 7148 11612 7160
rect 11664 7188 11670 7200
rect 11885 7191 11943 7197
rect 11885 7188 11897 7191
rect 11664 7160 11897 7188
rect 11664 7148 11670 7160
rect 11885 7157 11897 7160
rect 11931 7188 11943 7191
rect 13541 7191 13599 7197
rect 13541 7188 13553 7191
rect 11931 7160 13553 7188
rect 11931 7157 11943 7160
rect 11885 7151 11943 7157
rect 13541 7157 13553 7160
rect 13587 7188 13599 7191
rect 13998 7188 14004 7200
rect 13587 7160 14004 7188
rect 13587 7157 13599 7160
rect 13541 7151 13599 7157
rect 13998 7148 14004 7160
rect 14056 7148 14062 7200
rect 14182 7148 14188 7200
rect 14240 7188 14246 7200
rect 18506 7188 18512 7200
rect 14240 7160 18512 7188
rect 14240 7148 14246 7160
rect 18506 7148 18512 7160
rect 18564 7148 18570 7200
rect 19058 7148 19064 7200
rect 19116 7188 19122 7200
rect 19429 7191 19487 7197
rect 19429 7188 19441 7191
rect 19116 7160 19441 7188
rect 19116 7148 19122 7160
rect 19429 7157 19441 7160
rect 19475 7157 19487 7191
rect 20162 7188 20168 7200
rect 20123 7160 20168 7188
rect 19429 7151 19487 7157
rect 20162 7148 20168 7160
rect 20220 7148 20226 7200
rect 1104 7098 20884 7120
rect 1104 7046 8315 7098
rect 8367 7046 8379 7098
rect 8431 7046 8443 7098
rect 8495 7046 8507 7098
rect 8559 7046 15648 7098
rect 15700 7046 15712 7098
rect 15764 7046 15776 7098
rect 15828 7046 15840 7098
rect 15892 7046 20884 7098
rect 1104 7024 20884 7046
rect 1394 6984 1400 6996
rect 1355 6956 1400 6984
rect 1394 6944 1400 6956
rect 1452 6944 1458 6996
rect 1578 6944 1584 6996
rect 1636 6984 1642 6996
rect 2225 6987 2283 6993
rect 2225 6984 2237 6987
rect 1636 6956 2237 6984
rect 1636 6944 1642 6956
rect 2225 6953 2237 6956
rect 2271 6953 2283 6987
rect 6362 6984 6368 6996
rect 2225 6947 2283 6953
rect 3988 6956 6368 6984
rect 2682 6848 2688 6860
rect 2643 6820 2688 6848
rect 2682 6808 2688 6820
rect 2740 6808 2746 6860
rect 2866 6848 2872 6860
rect 2827 6820 2872 6848
rect 2866 6808 2872 6820
rect 2924 6808 2930 6860
rect 3142 6780 3148 6792
rect 3103 6752 3148 6780
rect 3142 6740 3148 6752
rect 3200 6740 3206 6792
rect 3881 6783 3939 6789
rect 3881 6749 3893 6783
rect 3927 6780 3939 6783
rect 3988 6780 4016 6956
rect 6362 6944 6368 6956
rect 6420 6944 6426 6996
rect 6914 6984 6920 6996
rect 6875 6956 6920 6984
rect 6914 6944 6920 6956
rect 6972 6944 6978 6996
rect 7285 6987 7343 6993
rect 7285 6953 7297 6987
rect 7331 6984 7343 6987
rect 7466 6984 7472 6996
rect 7331 6956 7472 6984
rect 7331 6953 7343 6956
rect 7285 6947 7343 6953
rect 4246 6916 4252 6928
rect 4207 6888 4252 6916
rect 4246 6876 4252 6888
rect 4304 6876 4310 6928
rect 5994 6876 6000 6928
rect 6052 6916 6058 6928
rect 7300 6916 7328 6947
rect 7466 6944 7472 6956
rect 7524 6944 7530 6996
rect 9030 6984 9036 6996
rect 8991 6956 9036 6984
rect 9030 6944 9036 6956
rect 9088 6944 9094 6996
rect 9306 6984 9312 6996
rect 9267 6956 9312 6984
rect 9306 6944 9312 6956
rect 9364 6944 9370 6996
rect 10778 6984 10784 6996
rect 10739 6956 10784 6984
rect 10778 6944 10784 6956
rect 10836 6944 10842 6996
rect 11146 6984 11152 6996
rect 11107 6956 11152 6984
rect 11146 6944 11152 6956
rect 11204 6944 11210 6996
rect 11514 6944 11520 6996
rect 11572 6984 11578 6996
rect 14090 6984 14096 6996
rect 11572 6956 14096 6984
rect 11572 6944 11578 6956
rect 14090 6944 14096 6956
rect 14148 6984 14154 6996
rect 14369 6987 14427 6993
rect 14369 6984 14381 6987
rect 14148 6956 14381 6984
rect 14148 6944 14154 6956
rect 14369 6953 14381 6956
rect 14415 6953 14427 6987
rect 15102 6984 15108 6996
rect 15063 6956 15108 6984
rect 14369 6947 14427 6953
rect 15102 6944 15108 6956
rect 15160 6944 15166 6996
rect 15378 6944 15384 6996
rect 15436 6984 15442 6996
rect 15841 6987 15899 6993
rect 15841 6984 15853 6987
rect 15436 6956 15853 6984
rect 15436 6944 15442 6956
rect 15841 6953 15853 6956
rect 15887 6953 15899 6987
rect 15841 6947 15899 6953
rect 15948 6956 16988 6984
rect 8938 6916 8944 6928
rect 6052 6888 7328 6916
rect 7852 6888 8944 6916
rect 6052 6876 6058 6888
rect 5629 6851 5687 6857
rect 5629 6817 5641 6851
rect 5675 6848 5687 6851
rect 5718 6848 5724 6860
rect 5675 6820 5724 6848
rect 5675 6817 5687 6820
rect 5629 6811 5687 6817
rect 5718 6808 5724 6820
rect 5776 6808 5782 6860
rect 5902 6848 5908 6860
rect 5863 6820 5908 6848
rect 5902 6808 5908 6820
rect 5960 6848 5966 6860
rect 6270 6848 6276 6860
rect 5960 6820 6276 6848
rect 5960 6808 5966 6820
rect 6270 6808 6276 6820
rect 6328 6808 6334 6860
rect 7190 6808 7196 6860
rect 7248 6848 7254 6860
rect 7377 6851 7435 6857
rect 7377 6848 7389 6851
rect 7248 6820 7389 6848
rect 7248 6808 7254 6820
rect 7377 6817 7389 6820
rect 7423 6817 7435 6851
rect 7377 6811 7435 6817
rect 7466 6808 7472 6860
rect 7524 6848 7530 6860
rect 7852 6857 7880 6888
rect 8938 6876 8944 6888
rect 8996 6876 9002 6928
rect 9858 6916 9864 6928
rect 9819 6888 9864 6916
rect 9858 6876 9864 6888
rect 9916 6876 9922 6928
rect 10413 6919 10471 6925
rect 10413 6885 10425 6919
rect 10459 6916 10471 6919
rect 11422 6916 11428 6928
rect 10459 6888 11428 6916
rect 10459 6885 10471 6888
rect 10413 6879 10471 6885
rect 11422 6876 11428 6888
rect 11480 6876 11486 6928
rect 11790 6916 11796 6928
rect 11751 6888 11796 6916
rect 11790 6876 11796 6888
rect 11848 6876 11854 6928
rect 12986 6916 12992 6928
rect 12947 6888 12992 6916
rect 12986 6876 12992 6888
rect 13044 6876 13050 6928
rect 13538 6916 13544 6928
rect 13499 6888 13544 6916
rect 13538 6876 13544 6888
rect 13596 6876 13602 6928
rect 15948 6916 15976 6956
rect 14108 6888 15976 6916
rect 16669 6919 16727 6925
rect 7837 6851 7895 6857
rect 7837 6848 7849 6851
rect 7524 6820 7849 6848
rect 7524 6808 7530 6820
rect 7837 6817 7849 6820
rect 7883 6817 7895 6851
rect 7837 6811 7895 6817
rect 8110 6808 8116 6860
rect 8168 6848 8174 6860
rect 8478 6848 8484 6860
rect 8168 6820 8484 6848
rect 8168 6808 8174 6820
rect 8478 6808 8484 6820
rect 8536 6808 8542 6860
rect 14108 6857 14136 6888
rect 16669 6885 16681 6919
rect 16715 6916 16727 6919
rect 16850 6916 16856 6928
rect 16715 6888 16856 6916
rect 16715 6885 16727 6888
rect 16669 6879 16727 6885
rect 16850 6876 16856 6888
rect 16908 6876 16914 6928
rect 16960 6916 16988 6956
rect 17126 6944 17132 6996
rect 17184 6984 17190 6996
rect 17497 6987 17555 6993
rect 17497 6984 17509 6987
rect 17184 6956 17509 6984
rect 17184 6944 17190 6956
rect 17497 6953 17509 6956
rect 17543 6953 17555 6987
rect 18138 6984 18144 6996
rect 18099 6956 18144 6984
rect 17497 6947 17555 6953
rect 18138 6944 18144 6956
rect 18196 6944 18202 6996
rect 19794 6944 19800 6996
rect 19852 6984 19858 6996
rect 21634 6984 21640 6996
rect 19852 6956 21640 6984
rect 19852 6944 19858 6956
rect 21634 6944 21640 6956
rect 21692 6944 21698 6996
rect 17221 6919 17279 6925
rect 17221 6916 17233 6919
rect 16960 6888 17233 6916
rect 17221 6885 17233 6888
rect 17267 6916 17279 6919
rect 18598 6916 18604 6928
rect 17267 6888 18604 6916
rect 17267 6885 17279 6888
rect 17221 6879 17279 6885
rect 18598 6876 18604 6888
rect 18656 6876 18662 6928
rect 14093 6851 14151 6857
rect 14093 6817 14105 6851
rect 14139 6817 14151 6851
rect 14093 6811 14151 6817
rect 15289 6851 15347 6857
rect 15289 6817 15301 6851
rect 15335 6848 15347 6851
rect 15378 6848 15384 6860
rect 15335 6820 15384 6848
rect 15335 6817 15347 6820
rect 15289 6811 15347 6817
rect 4157 6783 4215 6789
rect 4157 6780 4169 6783
rect 3927 6752 4169 6780
rect 3927 6749 3939 6752
rect 3881 6743 3939 6749
rect 4157 6749 4169 6752
rect 4203 6749 4215 6783
rect 6089 6783 6147 6789
rect 6089 6780 6101 6783
rect 4157 6743 4215 6749
rect 4264 6752 6101 6780
rect 2866 6672 2872 6724
rect 2924 6712 2930 6724
rect 4264 6712 4292 6752
rect 6089 6749 6101 6752
rect 6135 6749 6147 6783
rect 7926 6780 7932 6792
rect 7887 6752 7932 6780
rect 6089 6743 6147 6749
rect 7926 6740 7932 6752
rect 7984 6740 7990 6792
rect 8754 6740 8760 6792
rect 8812 6780 8818 6792
rect 9766 6780 9772 6792
rect 8812 6752 9772 6780
rect 8812 6740 8818 6752
rect 9766 6740 9772 6752
rect 9824 6740 9830 6792
rect 11698 6780 11704 6792
rect 11659 6752 11704 6780
rect 11698 6740 11704 6752
rect 11756 6740 11762 6792
rect 12345 6783 12403 6789
rect 12345 6749 12357 6783
rect 12391 6780 12403 6783
rect 12802 6780 12808 6792
rect 12391 6752 12808 6780
rect 12391 6749 12403 6752
rect 12345 6743 12403 6749
rect 12802 6740 12808 6752
rect 12860 6740 12866 6792
rect 13078 6740 13084 6792
rect 13136 6780 13142 6792
rect 13449 6783 13507 6789
rect 13449 6780 13461 6783
rect 13136 6752 13461 6780
rect 13136 6740 13142 6752
rect 13449 6749 13461 6752
rect 13495 6749 13507 6783
rect 13449 6743 13507 6749
rect 2924 6684 4292 6712
rect 2924 6672 2930 6684
rect 4338 6672 4344 6724
rect 4396 6712 4402 6724
rect 4709 6715 4767 6721
rect 4709 6712 4721 6715
rect 4396 6684 4721 6712
rect 4396 6672 4402 6684
rect 4709 6681 4721 6684
rect 4755 6681 4767 6715
rect 5721 6715 5779 6721
rect 5721 6712 5733 6715
rect 4709 6675 4767 6681
rect 4816 6684 5733 6712
rect 1854 6644 1860 6656
rect 1815 6616 1860 6644
rect 1854 6604 1860 6616
rect 1912 6644 1918 6656
rect 2774 6644 2780 6656
rect 1912 6616 2780 6644
rect 1912 6604 1918 6616
rect 2774 6604 2780 6616
rect 2832 6604 2838 6656
rect 4430 6604 4436 6656
rect 4488 6644 4494 6656
rect 4816 6644 4844 6684
rect 5721 6681 5733 6684
rect 5767 6681 5779 6715
rect 5721 6675 5779 6681
rect 5350 6644 5356 6656
rect 4488 6616 4844 6644
rect 5311 6616 5356 6644
rect 4488 6604 4494 6616
rect 5350 6604 5356 6616
rect 5408 6604 5414 6656
rect 5736 6644 5764 6675
rect 6546 6672 6552 6724
rect 6604 6712 6610 6724
rect 10042 6712 10048 6724
rect 6604 6684 10048 6712
rect 6604 6672 6610 6684
rect 10042 6672 10048 6684
rect 10100 6712 10106 6724
rect 11606 6712 11612 6724
rect 10100 6684 11612 6712
rect 10100 6672 10106 6684
rect 11606 6672 11612 6684
rect 11664 6672 11670 6724
rect 12526 6672 12532 6724
rect 12584 6712 12590 6724
rect 12713 6715 12771 6721
rect 12713 6712 12725 6715
rect 12584 6684 12725 6712
rect 12584 6672 12590 6684
rect 12713 6681 12725 6684
rect 12759 6712 12771 6715
rect 14108 6712 14136 6811
rect 15378 6808 15384 6820
rect 15436 6808 15442 6860
rect 18230 6848 18236 6860
rect 18191 6820 18236 6848
rect 18230 6808 18236 6820
rect 18288 6808 18294 6860
rect 18506 6848 18512 6860
rect 18467 6820 18512 6848
rect 18506 6808 18512 6820
rect 18564 6808 18570 6860
rect 19648 6851 19706 6857
rect 19648 6817 19660 6851
rect 19694 6817 19706 6851
rect 19648 6811 19706 6817
rect 16577 6783 16635 6789
rect 16577 6749 16589 6783
rect 16623 6780 16635 6783
rect 16666 6780 16672 6792
rect 16623 6752 16672 6780
rect 16623 6749 16635 6752
rect 16577 6743 16635 6749
rect 16666 6740 16672 6752
rect 16724 6740 16730 6792
rect 17678 6740 17684 6792
rect 17736 6780 17742 6792
rect 19663 6780 19691 6811
rect 20438 6780 20444 6792
rect 17736 6752 20444 6780
rect 17736 6740 17742 6752
rect 20438 6740 20444 6752
rect 20496 6740 20502 6792
rect 12759 6684 14136 6712
rect 12759 6681 12771 6684
rect 12713 6675 12771 6681
rect 14642 6672 14648 6724
rect 14700 6712 14706 6724
rect 15473 6715 15531 6721
rect 15473 6712 15485 6715
rect 14700 6684 15485 6712
rect 14700 6672 14706 6684
rect 15473 6681 15485 6684
rect 15519 6681 15531 6715
rect 15473 6675 15531 6681
rect 5902 6644 5908 6656
rect 5736 6616 5908 6644
rect 5902 6604 5908 6616
rect 5960 6644 5966 6656
rect 8110 6644 8116 6656
rect 5960 6616 8116 6644
rect 5960 6604 5966 6616
rect 8110 6604 8116 6616
rect 8168 6604 8174 6656
rect 15930 6604 15936 6656
rect 15988 6644 15994 6656
rect 16209 6647 16267 6653
rect 16209 6644 16221 6647
rect 15988 6616 16221 6644
rect 15988 6604 15994 6616
rect 16209 6613 16221 6616
rect 16255 6613 16267 6647
rect 16209 6607 16267 6613
rect 16298 6604 16304 6656
rect 16356 6644 16362 6656
rect 19751 6647 19809 6653
rect 19751 6644 19763 6647
rect 16356 6616 19763 6644
rect 16356 6604 16362 6616
rect 19751 6613 19763 6616
rect 19797 6613 19809 6647
rect 19751 6607 19809 6613
rect 1104 6554 20884 6576
rect 1104 6502 4648 6554
rect 4700 6502 4712 6554
rect 4764 6502 4776 6554
rect 4828 6502 4840 6554
rect 4892 6502 11982 6554
rect 12034 6502 12046 6554
rect 12098 6502 12110 6554
rect 12162 6502 12174 6554
rect 12226 6502 19315 6554
rect 19367 6502 19379 6554
rect 19431 6502 19443 6554
rect 19495 6502 19507 6554
rect 19559 6502 20884 6554
rect 1104 6480 20884 6502
rect 842 6400 848 6452
rect 900 6440 906 6452
rect 900 6412 2544 6440
rect 900 6400 906 6412
rect 2406 6372 2412 6384
rect 2367 6344 2412 6372
rect 2406 6332 2412 6344
rect 2464 6332 2470 6384
rect 2516 6372 2544 6412
rect 2866 6400 2872 6452
rect 2924 6440 2930 6452
rect 3145 6443 3203 6449
rect 3145 6440 3157 6443
rect 2924 6412 3157 6440
rect 2924 6400 2930 6412
rect 3145 6409 3157 6412
rect 3191 6440 3203 6443
rect 3234 6440 3240 6452
rect 3191 6412 3240 6440
rect 3191 6409 3203 6412
rect 3145 6403 3203 6409
rect 3234 6400 3240 6412
rect 3292 6400 3298 6452
rect 3973 6443 4031 6449
rect 3973 6409 3985 6443
rect 4019 6440 4031 6443
rect 4246 6440 4252 6452
rect 4019 6412 4252 6440
rect 4019 6409 4031 6412
rect 3973 6403 4031 6409
rect 4246 6400 4252 6412
rect 4304 6400 4310 6452
rect 5261 6443 5319 6449
rect 5261 6409 5273 6443
rect 5307 6440 5319 6443
rect 5718 6440 5724 6452
rect 5307 6412 5724 6440
rect 5307 6409 5319 6412
rect 5261 6403 5319 6409
rect 5718 6400 5724 6412
rect 5776 6400 5782 6452
rect 5859 6443 5917 6449
rect 5859 6409 5871 6443
rect 5905 6440 5917 6443
rect 11514 6440 11520 6452
rect 5905 6412 11520 6440
rect 5905 6409 5917 6412
rect 5859 6403 5917 6409
rect 11514 6400 11520 6412
rect 11572 6400 11578 6452
rect 11606 6400 11612 6452
rect 11664 6440 11670 6452
rect 13538 6440 13544 6452
rect 11664 6412 13124 6440
rect 13499 6412 13544 6440
rect 11664 6400 11670 6412
rect 6454 6372 6460 6384
rect 2516 6344 6460 6372
rect 6454 6332 6460 6344
rect 6512 6332 6518 6384
rect 6546 6332 6552 6384
rect 6604 6372 6610 6384
rect 7469 6375 7527 6381
rect 7469 6372 7481 6375
rect 6604 6344 7481 6372
rect 6604 6332 6610 6344
rect 7469 6341 7481 6344
rect 7515 6372 7527 6375
rect 9217 6375 9275 6381
rect 9217 6372 9229 6375
rect 7515 6344 9229 6372
rect 7515 6341 7527 6344
rect 7469 6335 7527 6341
rect 9217 6341 9229 6344
rect 9263 6341 9275 6375
rect 9766 6372 9772 6384
rect 9727 6344 9772 6372
rect 9217 6335 9275 6341
rect 9766 6332 9772 6344
rect 9824 6332 9830 6384
rect 12986 6372 12992 6384
rect 12544 6344 12992 6372
rect 1857 6307 1915 6313
rect 1857 6273 1869 6307
rect 1903 6304 1915 6307
rect 3050 6304 3056 6316
rect 1903 6276 3056 6304
rect 1903 6273 1915 6276
rect 1857 6267 1915 6273
rect 3050 6264 3056 6276
rect 3108 6264 3114 6316
rect 3418 6264 3424 6316
rect 3476 6304 3482 6316
rect 4157 6307 4215 6313
rect 4157 6304 4169 6307
rect 3476 6276 4169 6304
rect 3476 6264 3482 6276
rect 4157 6273 4169 6276
rect 4203 6304 4215 6307
rect 4338 6304 4344 6316
rect 4203 6276 4344 6304
rect 4203 6273 4215 6276
rect 4157 6267 4215 6273
rect 4338 6264 4344 6276
rect 4396 6264 4402 6316
rect 4801 6307 4859 6313
rect 4801 6273 4813 6307
rect 4847 6304 4859 6307
rect 4982 6304 4988 6316
rect 4847 6276 4988 6304
rect 4847 6273 4859 6276
rect 4801 6267 4859 6273
rect 4982 6264 4988 6276
rect 5040 6304 5046 6316
rect 5442 6304 5448 6316
rect 5040 6276 5448 6304
rect 5040 6264 5046 6276
rect 5442 6264 5448 6276
rect 5500 6264 5506 6316
rect 5534 6264 5540 6316
rect 5592 6304 5598 6316
rect 6917 6307 6975 6313
rect 6917 6304 6929 6307
rect 5592 6276 6929 6304
rect 5592 6264 5598 6276
rect 6917 6273 6929 6276
rect 6963 6304 6975 6307
rect 7650 6304 7656 6316
rect 6963 6276 7656 6304
rect 6963 6273 6975 6276
rect 6917 6267 6975 6273
rect 7650 6264 7656 6276
rect 7708 6264 7714 6316
rect 7834 6304 7840 6316
rect 7795 6276 7840 6304
rect 7834 6264 7840 6276
rect 7892 6264 7898 6316
rect 8665 6307 8723 6313
rect 8665 6273 8677 6307
rect 8711 6304 8723 6307
rect 9306 6304 9312 6316
rect 8711 6276 9312 6304
rect 8711 6273 8723 6276
rect 8665 6267 8723 6273
rect 9306 6264 9312 6276
rect 9364 6264 9370 6316
rect 12544 6313 12572 6344
rect 12986 6332 12992 6344
rect 13044 6332 13050 6384
rect 13096 6372 13124 6412
rect 13538 6400 13544 6412
rect 13596 6400 13602 6452
rect 15378 6440 15384 6452
rect 13786 6412 15384 6440
rect 13786 6372 13814 6412
rect 15378 6400 15384 6412
rect 15436 6440 15442 6452
rect 16850 6440 16856 6452
rect 15436 6412 16620 6440
rect 16811 6412 16856 6440
rect 15436 6400 15442 6412
rect 13096 6344 13814 6372
rect 16022 6332 16028 6384
rect 16080 6372 16086 6384
rect 16485 6375 16543 6381
rect 16485 6372 16497 6375
rect 16080 6344 16497 6372
rect 16080 6332 16086 6344
rect 16485 6341 16497 6344
rect 16531 6341 16543 6375
rect 16592 6372 16620 6412
rect 16850 6400 16856 6412
rect 16908 6400 16914 6452
rect 17497 6443 17555 6449
rect 17497 6409 17509 6443
rect 17543 6440 17555 6443
rect 18230 6440 18236 6452
rect 17543 6412 18236 6440
rect 17543 6409 17555 6412
rect 17497 6403 17555 6409
rect 18230 6400 18236 6412
rect 18288 6440 18294 6452
rect 19058 6440 19064 6452
rect 18288 6412 19064 6440
rect 18288 6400 18294 6412
rect 19058 6400 19064 6412
rect 19116 6400 19122 6452
rect 20438 6440 20444 6452
rect 20399 6412 20444 6440
rect 20438 6400 20444 6412
rect 20496 6400 20502 6452
rect 17586 6372 17592 6384
rect 16592 6344 17592 6372
rect 16485 6335 16543 6341
rect 17586 6332 17592 6344
rect 17644 6332 17650 6384
rect 12529 6307 12587 6313
rect 12529 6273 12541 6307
rect 12575 6273 12587 6307
rect 12894 6304 12900 6316
rect 12855 6276 12900 6304
rect 12529 6267 12587 6273
rect 12894 6264 12900 6276
rect 12952 6264 12958 6316
rect 14090 6304 14096 6316
rect 14051 6276 14096 6304
rect 14090 6264 14096 6276
rect 14148 6264 14154 6316
rect 15010 6264 15016 6316
rect 15068 6304 15074 6316
rect 19751 6307 19809 6313
rect 19751 6304 19763 6307
rect 15068 6276 19763 6304
rect 15068 6264 15074 6276
rect 19751 6273 19763 6276
rect 19797 6273 19809 6307
rect 19751 6267 19809 6273
rect 2682 6196 2688 6248
rect 2740 6236 2746 6248
rect 2869 6239 2927 6245
rect 2869 6236 2881 6239
rect 2740 6208 2881 6236
rect 2740 6196 2746 6208
rect 2869 6205 2881 6208
rect 2915 6236 2927 6239
rect 3970 6236 3976 6248
rect 2915 6208 3976 6236
rect 2915 6205 2927 6208
rect 2869 6199 2927 6205
rect 3970 6196 3976 6208
rect 4028 6196 4034 6248
rect 5626 6196 5632 6248
rect 5684 6236 5690 6248
rect 5756 6239 5814 6245
rect 5756 6236 5768 6239
rect 5684 6208 5768 6236
rect 5684 6196 5690 6208
rect 5756 6205 5768 6208
rect 5802 6236 5814 6239
rect 6549 6239 6607 6245
rect 6549 6236 6561 6239
rect 5802 6208 6561 6236
rect 5802 6205 5814 6208
rect 5756 6199 5814 6205
rect 6549 6205 6561 6208
rect 6595 6205 6607 6239
rect 10318 6236 10324 6248
rect 10279 6208 10324 6236
rect 6549 6199 6607 6205
rect 10318 6196 10324 6208
rect 10376 6196 10382 6248
rect 18230 6236 18236 6248
rect 18191 6208 18236 6236
rect 18230 6196 18236 6208
rect 18288 6196 18294 6248
rect 18509 6239 18567 6245
rect 18509 6205 18521 6239
rect 18555 6205 18567 6239
rect 18509 6199 18567 6205
rect 19664 6239 19722 6245
rect 19664 6205 19676 6239
rect 19710 6236 19722 6239
rect 19978 6236 19984 6248
rect 19710 6208 19984 6236
rect 19710 6205 19722 6208
rect 19664 6199 19722 6205
rect 1949 6171 2007 6177
rect 1949 6137 1961 6171
rect 1995 6137 2007 6171
rect 1949 6131 2007 6137
rect 3605 6171 3663 6177
rect 3605 6137 3617 6171
rect 3651 6168 3663 6171
rect 4246 6168 4252 6180
rect 3651 6140 4252 6168
rect 3651 6137 3663 6140
rect 3605 6131 3663 6137
rect 1673 6103 1731 6109
rect 1673 6069 1685 6103
rect 1719 6100 1731 6103
rect 1964 6100 1992 6131
rect 4246 6128 4252 6140
rect 4304 6128 4310 6180
rect 5442 6128 5448 6180
rect 5500 6168 5506 6180
rect 6270 6168 6276 6180
rect 5500 6140 6276 6168
rect 5500 6128 5506 6140
rect 6270 6128 6276 6140
rect 6328 6128 6334 6180
rect 7006 6128 7012 6180
rect 7064 6168 7070 6180
rect 7064 6140 7109 6168
rect 7064 6128 7070 6140
rect 7190 6128 7196 6180
rect 7248 6168 7254 6180
rect 8205 6171 8263 6177
rect 8205 6168 8217 6171
rect 7248 6140 8217 6168
rect 7248 6128 7254 6140
rect 8205 6137 8217 6140
rect 8251 6137 8263 6171
rect 8205 6131 8263 6137
rect 2314 6100 2320 6112
rect 1719 6072 2320 6100
rect 1719 6069 1731 6072
rect 1673 6063 1731 6069
rect 2314 6060 2320 6072
rect 2372 6060 2378 6112
rect 5629 6103 5687 6109
rect 5629 6069 5641 6103
rect 5675 6100 5687 6103
rect 5902 6100 5908 6112
rect 5675 6072 5908 6100
rect 5675 6069 5687 6072
rect 5629 6063 5687 6069
rect 5902 6060 5908 6072
rect 5960 6060 5966 6112
rect 8220 6100 8248 6131
rect 8754 6128 8760 6180
rect 8812 6168 8818 6180
rect 10229 6171 10287 6177
rect 8812 6140 8857 6168
rect 8812 6128 8818 6140
rect 10229 6137 10241 6171
rect 10275 6168 10287 6171
rect 10683 6171 10741 6177
rect 10683 6168 10695 6171
rect 10275 6140 10695 6168
rect 10275 6137 10287 6140
rect 10229 6131 10287 6137
rect 10683 6137 10695 6140
rect 10729 6168 10741 6171
rect 10870 6168 10876 6180
rect 10729 6140 10876 6168
rect 10729 6137 10741 6140
rect 10683 6131 10741 6137
rect 10870 6128 10876 6140
rect 10928 6128 10934 6180
rect 12621 6171 12679 6177
rect 12621 6137 12633 6171
rect 12667 6137 12679 6171
rect 12621 6131 12679 6137
rect 14001 6171 14059 6177
rect 14001 6137 14013 6171
rect 14047 6168 14059 6171
rect 14090 6168 14096 6180
rect 14047 6140 14096 6168
rect 14047 6137 14059 6140
rect 14001 6131 14059 6137
rect 9582 6100 9588 6112
rect 8220 6072 9588 6100
rect 9582 6060 9588 6072
rect 9640 6060 9646 6112
rect 11238 6100 11244 6112
rect 11199 6072 11244 6100
rect 11238 6060 11244 6072
rect 11296 6060 11302 6112
rect 11606 6100 11612 6112
rect 11567 6072 11612 6100
rect 11606 6060 11612 6072
rect 11664 6100 11670 6112
rect 11790 6100 11796 6112
rect 11664 6072 11796 6100
rect 11664 6060 11670 6072
rect 11790 6060 11796 6072
rect 11848 6100 11854 6112
rect 12161 6103 12219 6109
rect 12161 6100 12173 6103
rect 11848 6072 12173 6100
rect 11848 6060 11854 6072
rect 12161 6069 12173 6072
rect 12207 6100 12219 6103
rect 12636 6100 12664 6131
rect 14090 6128 14096 6140
rect 14148 6168 14154 6180
rect 14414 6171 14472 6177
rect 14414 6168 14426 6171
rect 14148 6140 14426 6168
rect 14148 6128 14154 6140
rect 14414 6137 14426 6140
rect 14460 6137 14472 6171
rect 14414 6131 14472 6137
rect 14918 6128 14924 6180
rect 14976 6168 14982 6180
rect 15657 6171 15715 6177
rect 15657 6168 15669 6171
rect 14976 6140 15669 6168
rect 14976 6128 14982 6140
rect 15657 6137 15669 6140
rect 15703 6137 15715 6171
rect 15930 6168 15936 6180
rect 15891 6140 15936 6168
rect 15657 6131 15715 6137
rect 12207 6072 12664 6100
rect 15013 6103 15071 6109
rect 12207 6069 12219 6072
rect 12161 6063 12219 6069
rect 15013 6069 15025 6103
rect 15059 6100 15071 6103
rect 15194 6100 15200 6112
rect 15059 6072 15200 6100
rect 15059 6069 15071 6072
rect 15013 6063 15071 6069
rect 15194 6060 15200 6072
rect 15252 6060 15258 6112
rect 15672 6100 15700 6131
rect 15930 6128 15936 6140
rect 15988 6128 15994 6180
rect 16025 6171 16083 6177
rect 16025 6137 16037 6171
rect 16071 6137 16083 6171
rect 16025 6131 16083 6137
rect 16040 6100 16068 6131
rect 17310 6128 17316 6180
rect 17368 6168 17374 6180
rect 17773 6171 17831 6177
rect 17773 6168 17785 6171
rect 17368 6140 17785 6168
rect 17368 6128 17374 6140
rect 17773 6137 17785 6140
rect 17819 6168 17831 6171
rect 18524 6168 18552 6199
rect 19978 6196 19984 6208
rect 20036 6236 20042 6248
rect 20073 6239 20131 6245
rect 20073 6236 20085 6239
rect 20036 6208 20085 6236
rect 20036 6196 20042 6208
rect 20073 6205 20085 6208
rect 20119 6205 20131 6239
rect 20073 6199 20131 6205
rect 17819 6140 18552 6168
rect 17819 6137 17831 6140
rect 17773 6131 17831 6137
rect 15672 6072 16068 6100
rect 17862 6060 17868 6112
rect 17920 6100 17926 6112
rect 18141 6103 18199 6109
rect 18141 6100 18153 6103
rect 17920 6072 18153 6100
rect 17920 6060 17926 6072
rect 18141 6069 18153 6072
rect 18187 6069 18199 6103
rect 18141 6063 18199 6069
rect 1104 6010 20884 6032
rect 1104 5958 8315 6010
rect 8367 5958 8379 6010
rect 8431 5958 8443 6010
rect 8495 5958 8507 6010
rect 8559 5958 15648 6010
rect 15700 5958 15712 6010
rect 15764 5958 15776 6010
rect 15828 5958 15840 6010
rect 15892 5958 20884 6010
rect 1104 5936 20884 5958
rect 2314 5896 2320 5908
rect 2275 5868 2320 5896
rect 2314 5856 2320 5868
rect 2372 5856 2378 5908
rect 2406 5856 2412 5908
rect 2464 5896 2470 5908
rect 3418 5896 3424 5908
rect 2464 5868 3424 5896
rect 2464 5856 2470 5868
rect 3418 5856 3424 5868
rect 3476 5856 3482 5908
rect 4246 5856 4252 5908
rect 4304 5896 4310 5908
rect 4985 5899 5043 5905
rect 4985 5896 4997 5899
rect 4304 5868 4997 5896
rect 4304 5856 4310 5868
rect 4985 5865 4997 5868
rect 5031 5865 5043 5899
rect 5534 5896 5540 5908
rect 5495 5868 5540 5896
rect 4985 5859 5043 5865
rect 5534 5856 5540 5868
rect 5592 5856 5598 5908
rect 7466 5896 7472 5908
rect 7427 5868 7472 5896
rect 7466 5856 7472 5868
rect 7524 5856 7530 5908
rect 9858 5896 9864 5908
rect 9819 5868 9864 5896
rect 9858 5856 9864 5868
rect 9916 5856 9922 5908
rect 11333 5899 11391 5905
rect 11333 5865 11345 5899
rect 11379 5896 11391 5899
rect 11606 5896 11612 5908
rect 11379 5868 11612 5896
rect 11379 5865 11391 5868
rect 11333 5859 11391 5865
rect 11606 5856 11612 5868
rect 11664 5856 11670 5908
rect 11698 5856 11704 5908
rect 11756 5896 11762 5908
rect 15010 5896 15016 5908
rect 11756 5868 15016 5896
rect 11756 5856 11762 5868
rect 15010 5856 15016 5868
rect 15068 5856 15074 5908
rect 18509 5899 18567 5905
rect 18509 5896 18521 5899
rect 15120 5868 18521 5896
rect 1759 5831 1817 5837
rect 1759 5797 1771 5831
rect 1805 5828 1817 5831
rect 1854 5828 1860 5840
rect 1805 5800 1860 5828
rect 1805 5797 1817 5800
rect 1759 5791 1817 5797
rect 1854 5788 1860 5800
rect 1912 5788 1918 5840
rect 2498 5788 2504 5840
rect 2556 5828 2562 5840
rect 2593 5831 2651 5837
rect 2593 5828 2605 5831
rect 2556 5800 2605 5828
rect 2556 5788 2562 5800
rect 2593 5797 2605 5800
rect 2639 5797 2651 5831
rect 2593 5791 2651 5797
rect 3694 5788 3700 5840
rect 3752 5828 3758 5840
rect 4427 5831 4485 5837
rect 4427 5828 4439 5831
rect 3752 5800 4439 5828
rect 3752 5788 3758 5800
rect 4427 5797 4439 5800
rect 4473 5828 4485 5831
rect 6359 5831 6417 5837
rect 6359 5828 6371 5831
rect 4473 5800 6371 5828
rect 4473 5797 4485 5800
rect 4427 5791 4485 5797
rect 6359 5797 6371 5800
rect 6405 5828 6417 5831
rect 6638 5828 6644 5840
rect 6405 5800 6644 5828
rect 6405 5797 6417 5800
rect 6359 5791 6417 5797
rect 6638 5788 6644 5800
rect 6696 5828 6702 5840
rect 8199 5831 8257 5837
rect 8199 5828 8211 5831
rect 6696 5800 8211 5828
rect 6696 5788 6702 5800
rect 8199 5797 8211 5800
rect 8245 5828 8257 5831
rect 9214 5828 9220 5840
rect 8245 5800 9220 5828
rect 8245 5797 8257 5800
rect 8199 5791 8257 5797
rect 9214 5788 9220 5800
rect 9272 5788 9278 5840
rect 10775 5831 10833 5837
rect 10775 5797 10787 5831
rect 10821 5828 10833 5831
rect 10870 5828 10876 5840
rect 10821 5800 10876 5828
rect 10821 5797 10833 5800
rect 10775 5791 10833 5797
rect 10870 5788 10876 5800
rect 10928 5788 10934 5840
rect 11238 5788 11244 5840
rect 11296 5828 11302 5840
rect 12342 5828 12348 5840
rect 11296 5800 12348 5828
rect 11296 5788 11302 5800
rect 12342 5788 12348 5800
rect 12400 5788 12406 5840
rect 13078 5788 13084 5840
rect 13136 5828 13142 5840
rect 13357 5831 13415 5837
rect 13357 5828 13369 5831
rect 13136 5800 13369 5828
rect 13136 5788 13142 5800
rect 13357 5797 13369 5800
rect 13403 5797 13415 5831
rect 13357 5791 13415 5797
rect 3050 5760 3056 5772
rect 3011 5732 3056 5760
rect 3050 5720 3056 5732
rect 3108 5720 3114 5772
rect 3142 5720 3148 5772
rect 3200 5760 3206 5772
rect 4062 5760 4068 5772
rect 3200 5732 4068 5760
rect 3200 5720 3206 5732
rect 4062 5720 4068 5732
rect 4120 5720 4126 5772
rect 7837 5763 7895 5769
rect 7837 5729 7849 5763
rect 7883 5760 7895 5763
rect 7926 5760 7932 5772
rect 7883 5732 7932 5760
rect 7883 5729 7895 5732
rect 7837 5723 7895 5729
rect 7926 5720 7932 5732
rect 7984 5720 7990 5772
rect 14093 5763 14151 5769
rect 14093 5729 14105 5763
rect 14139 5760 14151 5763
rect 14182 5760 14188 5772
rect 14139 5732 14188 5760
rect 14139 5729 14151 5732
rect 14093 5723 14151 5729
rect 14182 5720 14188 5732
rect 14240 5720 14246 5772
rect 1394 5692 1400 5704
rect 1355 5664 1400 5692
rect 1394 5652 1400 5664
rect 1452 5652 1458 5704
rect 5626 5652 5632 5704
rect 5684 5692 5690 5704
rect 5997 5695 6055 5701
rect 5997 5692 6009 5695
rect 5684 5664 6009 5692
rect 5684 5652 5690 5664
rect 5997 5661 6009 5664
rect 6043 5661 6055 5695
rect 10410 5692 10416 5704
rect 10371 5664 10416 5692
rect 5997 5655 6055 5661
rect 10410 5652 10416 5664
rect 10468 5652 10474 5704
rect 11514 5652 11520 5704
rect 11572 5692 11578 5704
rect 12253 5695 12311 5701
rect 12253 5692 12265 5695
rect 11572 5664 12265 5692
rect 11572 5652 11578 5664
rect 12253 5661 12265 5664
rect 12299 5692 12311 5695
rect 12710 5692 12716 5704
rect 12299 5664 12716 5692
rect 12299 5661 12311 5664
rect 12253 5655 12311 5661
rect 12710 5652 12716 5664
rect 12768 5652 12774 5704
rect 12894 5692 12900 5704
rect 12855 5664 12900 5692
rect 12894 5652 12900 5664
rect 12952 5652 12958 5704
rect 3970 5584 3976 5636
rect 4028 5624 4034 5636
rect 10042 5624 10048 5636
rect 4028 5596 10048 5624
rect 4028 5584 4034 5596
rect 10042 5584 10048 5596
rect 10100 5584 10106 5636
rect 10318 5624 10324 5636
rect 10231 5596 10324 5624
rect 10318 5584 10324 5596
rect 10376 5624 10382 5636
rect 15120 5624 15148 5868
rect 18509 5865 18521 5868
rect 18555 5865 18567 5899
rect 18509 5859 18567 5865
rect 15194 5788 15200 5840
rect 15252 5828 15258 5840
rect 15473 5831 15531 5837
rect 15473 5828 15485 5831
rect 15252 5800 15485 5828
rect 15252 5788 15258 5800
rect 15473 5797 15485 5800
rect 15519 5797 15531 5831
rect 15473 5791 15531 5797
rect 16577 5831 16635 5837
rect 16577 5797 16589 5831
rect 16623 5828 16635 5831
rect 16666 5828 16672 5840
rect 16623 5800 16672 5828
rect 16623 5797 16635 5800
rect 16577 5791 16635 5797
rect 16666 5788 16672 5800
rect 16724 5788 16730 5840
rect 17034 5828 17040 5840
rect 16995 5800 17040 5828
rect 17034 5788 17040 5800
rect 17092 5788 17098 5840
rect 18598 5760 18604 5772
rect 18559 5732 18604 5760
rect 18598 5720 18604 5732
rect 18656 5720 18662 5772
rect 18877 5763 18935 5769
rect 18877 5729 18889 5763
rect 18923 5729 18935 5763
rect 18877 5723 18935 5729
rect 15381 5695 15439 5701
rect 15381 5661 15393 5695
rect 15427 5661 15439 5695
rect 16022 5692 16028 5704
rect 15983 5664 16028 5692
rect 15381 5655 15439 5661
rect 10376 5596 15148 5624
rect 15396 5624 15424 5655
rect 16022 5652 16028 5664
rect 16080 5652 16086 5704
rect 16942 5692 16948 5704
rect 16903 5664 16948 5692
rect 16942 5652 16948 5664
rect 17000 5652 17006 5704
rect 17218 5692 17224 5704
rect 17179 5664 17224 5692
rect 17218 5652 17224 5664
rect 17276 5652 17282 5704
rect 18506 5692 18512 5704
rect 18064 5664 18512 5692
rect 16298 5624 16304 5636
rect 15396 5596 16304 5624
rect 10376 5584 10382 5596
rect 3786 5556 3792 5568
rect 3747 5528 3792 5556
rect 3786 5516 3792 5528
rect 3844 5516 3850 5568
rect 5905 5559 5963 5565
rect 5905 5525 5917 5559
rect 5951 5556 5963 5559
rect 6917 5559 6975 5565
rect 6917 5556 6929 5559
rect 5951 5528 6929 5556
rect 5951 5525 5963 5528
rect 5905 5519 5963 5525
rect 6917 5525 6929 5528
rect 6963 5556 6975 5559
rect 7006 5556 7012 5568
rect 6963 5528 7012 5556
rect 6963 5525 6975 5528
rect 6917 5519 6975 5525
rect 7006 5516 7012 5528
rect 7064 5516 7070 5568
rect 8754 5556 8760 5568
rect 8715 5528 8760 5556
rect 8754 5516 8760 5528
rect 8812 5556 8818 5568
rect 9033 5559 9091 5565
rect 9033 5556 9045 5559
rect 8812 5528 9045 5556
rect 8812 5516 8818 5528
rect 9033 5525 9045 5528
rect 9079 5525 9091 5559
rect 14274 5556 14280 5568
rect 14235 5528 14280 5556
rect 9033 5519 9091 5525
rect 14274 5516 14280 5528
rect 14332 5516 14338 5568
rect 15105 5559 15163 5565
rect 15105 5525 15117 5559
rect 15151 5556 15163 5559
rect 15396 5556 15424 5596
rect 16298 5584 16304 5596
rect 16356 5584 16362 5636
rect 15151 5528 15424 5556
rect 15151 5525 15163 5528
rect 15105 5519 15163 5525
rect 15838 5516 15844 5568
rect 15896 5556 15902 5568
rect 17494 5556 17500 5568
rect 15896 5528 17500 5556
rect 15896 5516 15902 5528
rect 17494 5516 17500 5528
rect 17552 5516 17558 5568
rect 17678 5516 17684 5568
rect 17736 5556 17742 5568
rect 18064 5565 18092 5664
rect 18506 5652 18512 5664
rect 18564 5692 18570 5704
rect 18892 5692 18920 5723
rect 19058 5692 19064 5704
rect 18564 5664 19064 5692
rect 18564 5652 18570 5664
rect 19058 5652 19064 5664
rect 19116 5652 19122 5704
rect 18049 5559 18107 5565
rect 18049 5556 18061 5559
rect 17736 5528 18061 5556
rect 17736 5516 17742 5528
rect 18049 5525 18061 5528
rect 18095 5525 18107 5559
rect 18049 5519 18107 5525
rect 1104 5466 20884 5488
rect 1104 5414 4648 5466
rect 4700 5414 4712 5466
rect 4764 5414 4776 5466
rect 4828 5414 4840 5466
rect 4892 5414 11982 5466
rect 12034 5414 12046 5466
rect 12098 5414 12110 5466
rect 12162 5414 12174 5466
rect 12226 5414 19315 5466
rect 19367 5414 19379 5466
rect 19431 5414 19443 5466
rect 19495 5414 19507 5466
rect 19559 5414 20884 5466
rect 1104 5392 20884 5414
rect 1394 5312 1400 5364
rect 1452 5352 1458 5364
rect 2866 5352 2872 5364
rect 1452 5324 2872 5352
rect 1452 5312 1458 5324
rect 2866 5312 2872 5324
rect 2924 5352 2930 5364
rect 3053 5355 3111 5361
rect 3053 5352 3065 5355
rect 2924 5324 3065 5352
rect 2924 5312 2930 5324
rect 3053 5321 3065 5324
rect 3099 5321 3111 5355
rect 3053 5315 3111 5321
rect 4062 5312 4068 5364
rect 4120 5352 4126 5364
rect 4985 5355 5043 5361
rect 4985 5352 4997 5355
rect 4120 5324 4997 5352
rect 4120 5312 4126 5324
rect 4985 5321 4997 5324
rect 5031 5321 5043 5355
rect 6638 5352 6644 5364
rect 6599 5324 6644 5352
rect 4985 5315 5043 5321
rect 6638 5312 6644 5324
rect 6696 5352 6702 5364
rect 7837 5355 7895 5361
rect 7837 5352 7849 5355
rect 6696 5324 7849 5352
rect 6696 5312 6702 5324
rect 7837 5321 7849 5324
rect 7883 5321 7895 5355
rect 7837 5315 7895 5321
rect 9769 5355 9827 5361
rect 9769 5321 9781 5355
rect 9815 5352 9827 5355
rect 10410 5352 10416 5364
rect 9815 5324 10416 5352
rect 9815 5321 9827 5324
rect 9769 5315 9827 5321
rect 10410 5312 10416 5324
rect 10468 5312 10474 5364
rect 10502 5312 10508 5364
rect 10560 5352 10566 5364
rect 11793 5355 11851 5361
rect 11793 5352 11805 5355
rect 10560 5324 11805 5352
rect 10560 5312 10566 5324
rect 11793 5321 11805 5324
rect 11839 5352 11851 5355
rect 12069 5355 12127 5361
rect 12069 5352 12081 5355
rect 11839 5324 12081 5352
rect 11839 5321 11851 5324
rect 11793 5315 11851 5321
rect 12069 5321 12081 5324
rect 12115 5321 12127 5355
rect 12069 5315 12127 5321
rect 12253 5355 12311 5361
rect 12253 5321 12265 5355
rect 12299 5352 12311 5355
rect 12342 5352 12348 5364
rect 12299 5324 12348 5352
rect 12299 5321 12311 5324
rect 12253 5315 12311 5321
rect 12342 5312 12348 5324
rect 12400 5312 12406 5364
rect 13909 5355 13967 5361
rect 13909 5321 13921 5355
rect 13955 5352 13967 5355
rect 14182 5352 14188 5364
rect 13955 5324 14188 5352
rect 13955 5321 13967 5324
rect 13909 5315 13967 5321
rect 14182 5312 14188 5324
rect 14240 5312 14246 5364
rect 14918 5352 14924 5364
rect 14879 5324 14924 5352
rect 14918 5312 14924 5324
rect 14976 5312 14982 5364
rect 15194 5312 15200 5364
rect 15252 5352 15258 5364
rect 15289 5355 15347 5361
rect 15289 5352 15301 5355
rect 15252 5324 15301 5352
rect 15252 5312 15258 5324
rect 15289 5321 15301 5324
rect 15335 5321 15347 5355
rect 15289 5315 15347 5321
rect 15930 5312 15936 5364
rect 15988 5352 15994 5364
rect 19058 5352 19064 5364
rect 15988 5324 17816 5352
rect 19019 5324 19064 5352
rect 15988 5312 15994 5324
rect 2130 5244 2136 5296
rect 2188 5284 2194 5296
rect 2317 5287 2375 5293
rect 2317 5284 2329 5287
rect 2188 5256 2329 5284
rect 2188 5244 2194 5256
rect 2317 5253 2329 5256
rect 2363 5253 2375 5287
rect 2317 5247 2375 5253
rect 2774 5244 2780 5296
rect 2832 5284 2838 5296
rect 3605 5287 3663 5293
rect 3605 5284 3617 5287
rect 2832 5256 3617 5284
rect 2832 5244 2838 5256
rect 3605 5253 3617 5256
rect 3651 5284 3663 5287
rect 3694 5284 3700 5296
rect 3651 5256 3700 5284
rect 3651 5253 3663 5256
rect 3605 5247 3663 5253
rect 3694 5244 3700 5256
rect 3752 5244 3758 5296
rect 10042 5284 10048 5296
rect 10003 5256 10048 5284
rect 10042 5244 10048 5256
rect 10100 5244 10106 5296
rect 14936 5284 14964 5312
rect 16853 5287 16911 5293
rect 16853 5284 16865 5287
rect 14936 5256 16865 5284
rect 16853 5253 16865 5256
rect 16899 5284 16911 5287
rect 17034 5284 17040 5296
rect 16899 5256 17040 5284
rect 16899 5253 16911 5256
rect 16853 5247 16911 5253
rect 17034 5244 17040 5256
rect 17092 5244 17098 5296
rect 17788 5284 17816 5324
rect 19058 5312 19064 5324
rect 19116 5312 19122 5364
rect 19751 5287 19809 5293
rect 19751 5284 19763 5287
rect 17788 5256 19763 5284
rect 19751 5253 19763 5256
rect 19797 5253 19809 5287
rect 19751 5247 19809 5253
rect 1765 5219 1823 5225
rect 1765 5185 1777 5219
rect 1811 5216 1823 5219
rect 2498 5216 2504 5228
rect 1811 5188 2504 5216
rect 1811 5185 1823 5188
rect 1765 5179 1823 5185
rect 2498 5176 2504 5188
rect 2556 5176 2562 5228
rect 5258 5176 5264 5228
rect 5316 5216 5322 5228
rect 7193 5219 7251 5225
rect 7193 5216 7205 5219
rect 5316 5188 7205 5216
rect 5316 5176 5322 5188
rect 7193 5185 7205 5188
rect 7239 5216 7251 5219
rect 8662 5216 8668 5228
rect 7239 5188 8668 5216
rect 7239 5185 7251 5188
rect 7193 5179 7251 5185
rect 8662 5176 8668 5188
rect 8720 5216 8726 5228
rect 8849 5219 8907 5225
rect 8849 5216 8861 5219
rect 8720 5188 8861 5216
rect 8720 5176 8726 5188
rect 8849 5185 8861 5188
rect 8895 5185 8907 5219
rect 8849 5179 8907 5185
rect 3142 5108 3148 5160
rect 3200 5148 3206 5160
rect 3786 5148 3792 5160
rect 3200 5120 3792 5148
rect 3200 5108 3206 5120
rect 3786 5108 3792 5120
rect 3844 5108 3850 5160
rect 5788 5151 5846 5157
rect 5788 5117 5800 5151
rect 5834 5148 5846 5151
rect 10060 5148 10088 5244
rect 10505 5219 10563 5225
rect 10505 5185 10517 5219
rect 10551 5216 10563 5219
rect 10870 5216 10876 5228
rect 10551 5188 10876 5216
rect 10551 5185 10563 5188
rect 10505 5179 10563 5185
rect 10870 5176 10876 5188
rect 10928 5176 10934 5228
rect 11514 5176 11520 5228
rect 11572 5216 11578 5228
rect 12802 5216 12808 5228
rect 11572 5188 12808 5216
rect 11572 5176 11578 5188
rect 12802 5176 12808 5188
rect 12860 5216 12866 5228
rect 13354 5216 13360 5228
rect 12860 5188 13360 5216
rect 12860 5176 12866 5188
rect 13354 5176 13360 5188
rect 13412 5176 13418 5228
rect 13541 5219 13599 5225
rect 13541 5185 13553 5219
rect 13587 5216 13599 5219
rect 14001 5219 14059 5225
rect 14001 5216 14013 5219
rect 13587 5188 14013 5216
rect 13587 5185 13599 5188
rect 13541 5179 13599 5185
rect 14001 5185 14013 5188
rect 14047 5216 14059 5219
rect 17862 5216 17868 5228
rect 14047 5188 17868 5216
rect 14047 5185 14059 5188
rect 14001 5179 14059 5185
rect 17862 5176 17868 5188
rect 17920 5176 17926 5228
rect 10778 5148 10784 5160
rect 5834 5120 6316 5148
rect 10060 5120 10784 5148
rect 5834 5117 5846 5120
rect 5788 5111 5846 5117
rect 1857 5083 1915 5089
rect 1857 5049 1869 5083
rect 1903 5080 1915 5083
rect 2222 5080 2228 5092
rect 1903 5052 2228 5080
rect 1903 5049 1915 5052
rect 1857 5043 1915 5049
rect 2222 5040 2228 5052
rect 2280 5040 2286 5092
rect 3694 5040 3700 5092
rect 3752 5080 3758 5092
rect 4110 5083 4168 5089
rect 4110 5080 4122 5083
rect 3752 5052 4122 5080
rect 3752 5040 3758 5052
rect 4110 5049 4122 5052
rect 4156 5049 4168 5083
rect 4110 5043 4168 5049
rect 2240 5012 2268 5040
rect 6288 5024 6316 5120
rect 10778 5108 10784 5120
rect 10836 5108 10842 5160
rect 11330 5148 11336 5160
rect 11291 5120 11336 5148
rect 11330 5108 11336 5120
rect 11388 5108 11394 5160
rect 16482 5108 16488 5160
rect 16540 5148 16546 5160
rect 17218 5148 17224 5160
rect 16540 5120 17224 5148
rect 16540 5108 16546 5120
rect 17218 5108 17224 5120
rect 17276 5108 17282 5160
rect 17770 5108 17776 5160
rect 17828 5148 17834 5160
rect 18141 5151 18199 5157
rect 18141 5148 18153 5151
rect 17828 5120 18153 5148
rect 17828 5108 17834 5120
rect 18141 5117 18153 5120
rect 18187 5117 18199 5151
rect 18141 5111 18199 5117
rect 19680 5151 19738 5157
rect 19680 5117 19692 5151
rect 19726 5148 19738 5151
rect 20070 5148 20076 5160
rect 19726 5120 20076 5148
rect 19726 5117 19738 5120
rect 19680 5111 19738 5117
rect 20070 5108 20076 5120
rect 20128 5108 20134 5160
rect 6914 5080 6920 5092
rect 6875 5052 6920 5080
rect 6914 5040 6920 5052
rect 6972 5040 6978 5092
rect 7006 5040 7012 5092
rect 7064 5080 7070 5092
rect 7064 5052 7109 5080
rect 7064 5040 7070 5052
rect 8110 5040 8116 5092
rect 8168 5080 8174 5092
rect 8573 5083 8631 5089
rect 8573 5080 8585 5083
rect 8168 5052 8585 5080
rect 8168 5040 8174 5052
rect 8573 5049 8585 5052
rect 8619 5049 8631 5083
rect 8573 5043 8631 5049
rect 8665 5083 8723 5089
rect 8665 5049 8677 5083
rect 8711 5080 8723 5083
rect 8754 5080 8760 5092
rect 8711 5052 8760 5080
rect 8711 5049 8723 5052
rect 8665 5043 8723 5049
rect 2685 5015 2743 5021
rect 2685 5012 2697 5015
rect 2240 4984 2697 5012
rect 2685 4981 2697 4984
rect 2731 4981 2743 5015
rect 4706 5012 4712 5024
rect 4667 4984 4712 5012
rect 2685 4975 2743 4981
rect 4706 4972 4712 4984
rect 4764 4972 4770 5024
rect 5626 5012 5632 5024
rect 5587 4984 5632 5012
rect 5626 4972 5632 4984
rect 5684 4972 5690 5024
rect 5859 5015 5917 5021
rect 5859 4981 5871 5015
rect 5905 5012 5917 5015
rect 6086 5012 6092 5024
rect 5905 4984 6092 5012
rect 5905 4981 5917 4984
rect 5859 4975 5917 4981
rect 6086 4972 6092 4984
rect 6144 4972 6150 5024
rect 6270 5012 6276 5024
rect 6231 4984 6276 5012
rect 6270 4972 6276 4984
rect 6328 4972 6334 5024
rect 8389 5015 8447 5021
rect 8389 4981 8401 5015
rect 8435 5012 8447 5015
rect 8680 5012 8708 5043
rect 8754 5040 8760 5052
rect 8812 5040 8818 5092
rect 11422 5040 11428 5092
rect 11480 5080 11486 5092
rect 11517 5083 11575 5089
rect 11517 5080 11529 5083
rect 11480 5052 11529 5080
rect 11480 5040 11486 5052
rect 11517 5049 11529 5052
rect 11563 5049 11575 5083
rect 11517 5043 11575 5049
rect 12069 5083 12127 5089
rect 12069 5049 12081 5083
rect 12115 5080 12127 5083
rect 12529 5083 12587 5089
rect 12529 5080 12541 5083
rect 12115 5052 12541 5080
rect 12115 5049 12127 5052
rect 12069 5043 12127 5049
rect 12529 5049 12541 5052
rect 12575 5049 12587 5083
rect 12529 5043 12587 5049
rect 12621 5083 12679 5089
rect 12621 5049 12633 5083
rect 12667 5049 12679 5083
rect 12621 5043 12679 5049
rect 8435 4984 8708 5012
rect 8435 4981 8447 4984
rect 8389 4975 8447 4981
rect 12342 4972 12348 5024
rect 12400 5012 12406 5024
rect 12636 5012 12664 5043
rect 14090 5040 14096 5092
rect 14148 5080 14154 5092
rect 14322 5083 14380 5089
rect 14322 5080 14334 5083
rect 14148 5052 14334 5080
rect 14148 5040 14154 5052
rect 14322 5049 14334 5052
rect 14368 5049 14380 5083
rect 14322 5043 14380 5049
rect 15102 5040 15108 5092
rect 15160 5080 15166 5092
rect 15838 5080 15844 5092
rect 15160 5052 15844 5080
rect 15160 5040 15166 5052
rect 15838 5040 15844 5052
rect 15896 5040 15902 5092
rect 15933 5083 15991 5089
rect 15933 5049 15945 5083
rect 15979 5049 15991 5083
rect 18046 5080 18052 5092
rect 18007 5052 18052 5080
rect 15933 5043 15991 5049
rect 12400 4984 12664 5012
rect 12400 4972 12406 4984
rect 15194 4972 15200 5024
rect 15252 5012 15258 5024
rect 15948 5012 15976 5043
rect 18046 5040 18052 5052
rect 18104 5040 18110 5092
rect 16298 5012 16304 5024
rect 15252 4984 16304 5012
rect 15252 4972 15258 4984
rect 16298 4972 16304 4984
rect 16356 4972 16362 5024
rect 16942 4972 16948 5024
rect 17000 5012 17006 5024
rect 17221 5015 17279 5021
rect 17221 5012 17233 5015
rect 17000 4984 17233 5012
rect 17000 4972 17006 4984
rect 17221 4981 17233 4984
rect 17267 4981 17279 5015
rect 17770 5012 17776 5024
rect 17731 4984 17776 5012
rect 17221 4975 17279 4981
rect 17770 4972 17776 4984
rect 17828 4972 17834 5024
rect 19521 5015 19579 5021
rect 19521 4981 19533 5015
rect 19567 5012 19579 5015
rect 19702 5012 19708 5024
rect 19567 4984 19708 5012
rect 19567 4981 19579 4984
rect 19521 4975 19579 4981
rect 19702 4972 19708 4984
rect 19760 4972 19766 5024
rect 1104 4922 20884 4944
rect 1104 4870 8315 4922
rect 8367 4870 8379 4922
rect 8431 4870 8443 4922
rect 8495 4870 8507 4922
rect 8559 4870 15648 4922
rect 15700 4870 15712 4922
rect 15764 4870 15776 4922
rect 15828 4870 15840 4922
rect 15892 4870 20884 4922
rect 1104 4848 20884 4870
rect 2130 4768 2136 4820
rect 2188 4808 2194 4820
rect 3421 4811 3479 4817
rect 3421 4808 3433 4811
rect 2188 4780 3433 4808
rect 2188 4768 2194 4780
rect 3421 4777 3433 4780
rect 3467 4808 3479 4811
rect 3467 4780 4292 4808
rect 3467 4777 3479 4780
rect 3421 4771 3479 4777
rect 1397 4743 1455 4749
rect 1397 4709 1409 4743
rect 1443 4740 1455 4743
rect 1443 4712 3280 4740
rect 1443 4709 1455 4712
rect 1397 4703 1455 4709
rect 2682 4672 2688 4684
rect 2643 4644 2688 4672
rect 2682 4632 2688 4644
rect 2740 4632 2746 4684
rect 2869 4675 2927 4681
rect 2869 4641 2881 4675
rect 2915 4641 2927 4675
rect 3142 4672 3148 4684
rect 3103 4644 3148 4672
rect 2869 4635 2927 4641
rect 1762 4496 1768 4548
rect 1820 4536 1826 4548
rect 2317 4539 2375 4545
rect 2317 4536 2329 4539
rect 1820 4508 2329 4536
rect 1820 4496 1826 4508
rect 2317 4505 2329 4508
rect 2363 4536 2375 4539
rect 2774 4536 2780 4548
rect 2363 4508 2780 4536
rect 2363 4505 2375 4508
rect 2317 4499 2375 4505
rect 2774 4496 2780 4508
rect 2832 4536 2838 4548
rect 2884 4536 2912 4635
rect 3142 4632 3148 4644
rect 3200 4632 3206 4684
rect 3252 4604 3280 4712
rect 3694 4700 3700 4752
rect 3752 4740 3758 4752
rect 4264 4749 4292 4780
rect 7006 4768 7012 4820
rect 7064 4808 7070 4820
rect 7469 4811 7527 4817
rect 7469 4808 7481 4811
rect 7064 4780 7481 4808
rect 7064 4768 7070 4780
rect 7469 4777 7481 4780
rect 7515 4777 7527 4811
rect 7926 4808 7932 4820
rect 7887 4780 7932 4808
rect 7469 4771 7527 4777
rect 7926 4768 7932 4780
rect 7984 4768 7990 4820
rect 8110 4768 8116 4820
rect 8168 4808 8174 4820
rect 9125 4811 9183 4817
rect 9125 4808 9137 4811
rect 8168 4780 9137 4808
rect 8168 4768 8174 4780
rect 9125 4777 9137 4780
rect 9171 4808 9183 4811
rect 10134 4808 10140 4820
rect 9171 4780 10140 4808
rect 9171 4777 9183 4780
rect 9125 4771 9183 4777
rect 10134 4768 10140 4780
rect 10192 4768 10198 4820
rect 10965 4811 11023 4817
rect 10965 4777 10977 4811
rect 11011 4808 11023 4811
rect 11238 4808 11244 4820
rect 11011 4780 11244 4808
rect 11011 4777 11023 4780
rect 10965 4771 11023 4777
rect 3789 4743 3847 4749
rect 3789 4740 3801 4743
rect 3752 4712 3801 4740
rect 3752 4700 3758 4712
rect 3789 4709 3801 4712
rect 3835 4709 3847 4743
rect 3789 4703 3847 4709
rect 4249 4743 4307 4749
rect 4249 4709 4261 4743
rect 4295 4709 4307 4743
rect 4249 4703 4307 4709
rect 4341 4743 4399 4749
rect 4341 4709 4353 4743
rect 4387 4740 4399 4743
rect 4522 4740 4528 4752
rect 4387 4712 4528 4740
rect 4387 4709 4399 4712
rect 4341 4703 4399 4709
rect 4522 4700 4528 4712
rect 4580 4740 4586 4752
rect 4706 4740 4712 4752
rect 4580 4712 4712 4740
rect 4580 4700 4586 4712
rect 4706 4700 4712 4712
rect 4764 4700 4770 4752
rect 4893 4743 4951 4749
rect 4893 4709 4905 4743
rect 4939 4740 4951 4743
rect 4982 4740 4988 4752
rect 4939 4712 4988 4740
rect 4939 4709 4951 4712
rect 4893 4703 4951 4709
rect 4982 4700 4988 4712
rect 5040 4700 5046 4752
rect 6638 4740 6644 4752
rect 6599 4712 6644 4740
rect 6638 4700 6644 4712
rect 6696 4700 6702 4752
rect 7193 4743 7251 4749
rect 7193 4709 7205 4743
rect 7239 4740 7251 4743
rect 7282 4740 7288 4752
rect 7239 4712 7288 4740
rect 7239 4709 7251 4712
rect 7193 4703 7251 4709
rect 7282 4700 7288 4712
rect 7340 4700 7346 4752
rect 8202 4740 8208 4752
rect 8163 4712 8208 4740
rect 8202 4700 8208 4712
rect 8260 4700 8266 4752
rect 8754 4632 8760 4684
rect 8812 4672 8818 4684
rect 9490 4672 9496 4684
rect 8812 4644 9496 4672
rect 8812 4632 8818 4644
rect 9490 4632 9496 4644
rect 9548 4672 9554 4684
rect 9858 4672 9864 4684
rect 9548 4644 9864 4672
rect 9548 4632 9554 4644
rect 9858 4632 9864 4644
rect 9916 4632 9922 4684
rect 9950 4632 9956 4684
rect 10008 4672 10014 4684
rect 10413 4675 10471 4681
rect 10413 4672 10425 4675
rect 10008 4644 10425 4672
rect 10008 4632 10014 4644
rect 10413 4641 10425 4644
rect 10459 4672 10471 4675
rect 10980 4672 11008 4771
rect 11238 4768 11244 4780
rect 11296 4808 11302 4820
rect 11296 4780 12296 4808
rect 11296 4768 11302 4780
rect 11333 4743 11391 4749
rect 11333 4709 11345 4743
rect 11379 4740 11391 4743
rect 11514 4740 11520 4752
rect 11379 4712 11520 4740
rect 11379 4709 11391 4712
rect 11333 4703 11391 4709
rect 11514 4700 11520 4712
rect 11572 4700 11578 4752
rect 11609 4743 11667 4749
rect 11609 4709 11621 4743
rect 11655 4740 11667 4743
rect 11698 4740 11704 4752
rect 11655 4712 11704 4740
rect 11655 4709 11667 4712
rect 11609 4703 11667 4709
rect 11698 4700 11704 4712
rect 11756 4700 11762 4752
rect 12268 4740 12296 4780
rect 12342 4768 12348 4820
rect 12400 4808 12406 4820
rect 12437 4811 12495 4817
rect 12437 4808 12449 4811
rect 12400 4780 12449 4808
rect 12400 4768 12406 4780
rect 12437 4777 12449 4780
rect 12483 4777 12495 4811
rect 12437 4771 12495 4777
rect 12710 4768 12716 4820
rect 12768 4808 12774 4820
rect 12805 4811 12863 4817
rect 12805 4808 12817 4811
rect 12768 4780 12817 4808
rect 12768 4768 12774 4780
rect 12805 4777 12817 4780
rect 12851 4777 12863 4811
rect 15102 4808 15108 4820
rect 12805 4771 12863 4777
rect 12906 4780 13814 4808
rect 15063 4780 15108 4808
rect 12906 4740 12934 4780
rect 12268 4712 12934 4740
rect 13173 4743 13231 4749
rect 13173 4709 13185 4743
rect 13219 4740 13231 4743
rect 13262 4740 13268 4752
rect 13219 4712 13268 4740
rect 13219 4709 13231 4712
rect 13173 4703 13231 4709
rect 13262 4700 13268 4712
rect 13320 4700 13326 4752
rect 13786 4740 13814 4780
rect 15102 4768 15108 4780
rect 15160 4768 15166 4820
rect 16298 4808 16304 4820
rect 15304 4780 16160 4808
rect 16259 4780 16304 4808
rect 15304 4740 15332 4780
rect 15470 4740 15476 4752
rect 13786 4712 15332 4740
rect 15431 4712 15476 4740
rect 15470 4700 15476 4712
rect 15528 4700 15534 4752
rect 16132 4740 16160 4780
rect 16298 4768 16304 4780
rect 16356 4768 16362 4820
rect 16942 4808 16948 4820
rect 16903 4780 16948 4808
rect 16942 4768 16948 4780
rect 17000 4768 17006 4820
rect 18690 4808 18696 4820
rect 18651 4780 18696 4808
rect 18690 4768 18696 4780
rect 18748 4768 18754 4820
rect 18141 4743 18199 4749
rect 16132 4712 17356 4740
rect 17328 4684 17356 4712
rect 18141 4709 18153 4743
rect 18187 4740 18199 4743
rect 18874 4740 18880 4752
rect 18187 4712 18880 4740
rect 18187 4709 18199 4712
rect 18141 4703 18199 4709
rect 10459 4644 11008 4672
rect 10459 4641 10471 4644
rect 10413 4635 10471 4641
rect 16298 4632 16304 4684
rect 16356 4672 16362 4684
rect 17129 4675 17187 4681
rect 17129 4672 17141 4675
rect 16356 4644 17141 4672
rect 16356 4632 16362 4644
rect 17129 4641 17141 4644
rect 17175 4641 17187 4675
rect 17310 4672 17316 4684
rect 17223 4644 17316 4672
rect 17129 4635 17187 4641
rect 5534 4604 5540 4616
rect 3252 4576 5540 4604
rect 5534 4564 5540 4576
rect 5592 4564 5598 4616
rect 5997 4607 6055 4613
rect 5997 4573 6009 4607
rect 6043 4604 6055 4607
rect 6546 4604 6552 4616
rect 6043 4576 6552 4604
rect 6043 4573 6055 4576
rect 5997 4567 6055 4573
rect 6546 4564 6552 4576
rect 6604 4604 6610 4616
rect 7466 4604 7472 4616
rect 6604 4576 7472 4604
rect 6604 4564 6610 4576
rect 7466 4564 7472 4576
rect 7524 4564 7530 4616
rect 8113 4607 8171 4613
rect 8113 4573 8125 4607
rect 8159 4573 8171 4607
rect 10594 4604 10600 4616
rect 10555 4576 10600 4604
rect 8113 4567 8171 4573
rect 3234 4536 3240 4548
rect 2832 4508 3240 4536
rect 2832 4496 2838 4508
rect 3234 4496 3240 4508
rect 3292 4496 3298 4548
rect 6365 4539 6423 4545
rect 6365 4505 6377 4539
rect 6411 4536 6423 4539
rect 6914 4536 6920 4548
rect 6411 4508 6920 4536
rect 6411 4505 6423 4508
rect 6365 4499 6423 4505
rect 6914 4496 6920 4508
rect 6972 4536 6978 4548
rect 7374 4536 7380 4548
rect 6972 4508 7380 4536
rect 6972 4496 6978 4508
rect 7374 4496 7380 4508
rect 7432 4496 7438 4548
rect 8128 4480 8156 4567
rect 10594 4564 10600 4576
rect 10652 4564 10658 4616
rect 12161 4607 12219 4613
rect 12161 4573 12173 4607
rect 12207 4604 12219 4607
rect 12342 4604 12348 4616
rect 12207 4576 12348 4604
rect 12207 4573 12219 4576
rect 12161 4567 12219 4573
rect 12342 4564 12348 4576
rect 12400 4564 12406 4616
rect 13078 4604 13084 4616
rect 13039 4576 13084 4604
rect 13078 4564 13084 4576
rect 13136 4564 13142 4616
rect 13354 4604 13360 4616
rect 13315 4576 13360 4604
rect 13354 4564 13360 4576
rect 13412 4564 13418 4616
rect 14737 4607 14795 4613
rect 14737 4573 14749 4607
rect 14783 4604 14795 4607
rect 15381 4607 15439 4613
rect 15381 4604 15393 4607
rect 14783 4576 15393 4604
rect 14783 4573 14795 4576
rect 14737 4567 14795 4573
rect 15381 4573 15393 4576
rect 15427 4604 15439 4607
rect 16390 4604 16396 4616
rect 15427 4576 16396 4604
rect 15427 4573 15439 4576
rect 15381 4567 15439 4573
rect 16390 4564 16396 4576
rect 16448 4564 16454 4616
rect 17144 4604 17172 4635
rect 17310 4632 17316 4644
rect 17368 4632 17374 4684
rect 18156 4616 18184 4703
rect 18874 4700 18880 4712
rect 18932 4700 18938 4752
rect 18506 4672 18512 4684
rect 18467 4644 18512 4672
rect 18506 4632 18512 4644
rect 18564 4632 18570 4684
rect 18138 4604 18144 4616
rect 17144 4576 18144 4604
rect 18138 4564 18144 4576
rect 18196 4564 18202 4616
rect 8662 4536 8668 4548
rect 8623 4508 8668 4536
rect 8662 4496 8668 4508
rect 8720 4496 8726 4548
rect 15930 4536 15936 4548
rect 15891 4508 15936 4536
rect 15930 4496 15936 4508
rect 15988 4496 15994 4548
rect 1854 4468 1860 4480
rect 1815 4440 1860 4468
rect 1854 4428 1860 4440
rect 1912 4428 1918 4480
rect 8110 4428 8116 4480
rect 8168 4468 8174 4480
rect 11054 4468 11060 4480
rect 8168 4440 11060 4468
rect 8168 4428 8174 4440
rect 11054 4428 11060 4440
rect 11112 4428 11118 4480
rect 14090 4468 14096 4480
rect 14051 4440 14096 4468
rect 14090 4428 14096 4440
rect 14148 4428 14154 4480
rect 16482 4428 16488 4480
rect 16540 4468 16546 4480
rect 16669 4471 16727 4477
rect 16669 4468 16681 4471
rect 16540 4440 16681 4468
rect 16540 4428 16546 4440
rect 16669 4437 16681 4440
rect 16715 4437 16727 4471
rect 16669 4431 16727 4437
rect 18598 4428 18604 4480
rect 18656 4468 18662 4480
rect 19702 4468 19708 4480
rect 18656 4440 19708 4468
rect 18656 4428 18662 4440
rect 19702 4428 19708 4440
rect 19760 4428 19766 4480
rect 1104 4378 20884 4400
rect 1104 4326 4648 4378
rect 4700 4326 4712 4378
rect 4764 4326 4776 4378
rect 4828 4326 4840 4378
rect 4892 4326 11982 4378
rect 12034 4326 12046 4378
rect 12098 4326 12110 4378
rect 12162 4326 12174 4378
rect 12226 4326 19315 4378
rect 19367 4326 19379 4378
rect 19431 4326 19443 4378
rect 19495 4326 19507 4378
rect 19559 4326 20884 4378
rect 1104 4304 20884 4326
rect 1762 4264 1768 4276
rect 1723 4236 1768 4264
rect 1762 4224 1768 4236
rect 1820 4224 1826 4276
rect 2133 4267 2191 4273
rect 2133 4233 2145 4267
rect 2179 4264 2191 4267
rect 2406 4264 2412 4276
rect 2179 4236 2412 4264
rect 2179 4233 2191 4236
rect 2133 4227 2191 4233
rect 2148 4196 2176 4227
rect 2406 4224 2412 4236
rect 2464 4224 2470 4276
rect 2682 4224 2688 4276
rect 2740 4264 2746 4276
rect 3237 4267 3295 4273
rect 3237 4264 3249 4267
rect 2740 4236 3249 4264
rect 2740 4224 2746 4236
rect 3237 4233 3249 4236
rect 3283 4264 3295 4267
rect 3283 4236 4154 4264
rect 3283 4233 3295 4236
rect 3237 4227 3295 4233
rect 2056 4168 2176 4196
rect 4126 4196 4154 4236
rect 4522 4224 4528 4276
rect 4580 4264 4586 4276
rect 4801 4267 4859 4273
rect 4801 4264 4813 4267
rect 4580 4236 4813 4264
rect 4580 4224 4586 4236
rect 4801 4233 4813 4236
rect 4847 4233 4859 4267
rect 4801 4227 4859 4233
rect 8113 4267 8171 4273
rect 8113 4233 8125 4267
rect 8159 4264 8171 4267
rect 8202 4264 8208 4276
rect 8159 4236 8208 4264
rect 8159 4233 8171 4236
rect 8113 4227 8171 4233
rect 8202 4224 8208 4236
rect 8260 4264 8266 4276
rect 9493 4267 9551 4273
rect 9493 4264 9505 4267
rect 8260 4236 9505 4264
rect 8260 4224 8266 4236
rect 9493 4233 9505 4236
rect 9539 4233 9551 4267
rect 9950 4264 9956 4276
rect 9911 4236 9956 4264
rect 9493 4227 9551 4233
rect 9950 4224 9956 4236
rect 10008 4224 10014 4276
rect 13909 4267 13967 4273
rect 13909 4264 13921 4267
rect 13786 4236 13921 4264
rect 8754 4196 8760 4208
rect 4126 4168 8760 4196
rect 2056 4128 2084 4168
rect 8754 4156 8760 4168
rect 8812 4156 8818 4208
rect 10318 4156 10324 4208
rect 10376 4196 10382 4208
rect 10376 4168 13032 4196
rect 10376 4156 10382 4168
rect 3510 4128 3516 4140
rect 2056 4100 3516 4128
rect 2516 4069 2544 4100
rect 3510 4088 3516 4100
rect 3568 4088 3574 4140
rect 4525 4131 4583 4137
rect 4525 4097 4537 4131
rect 4571 4128 4583 4131
rect 4982 4128 4988 4140
rect 4571 4100 4988 4128
rect 4571 4097 4583 4100
rect 4525 4091 4583 4097
rect 4982 4088 4988 4100
rect 5040 4088 5046 4140
rect 5261 4131 5319 4137
rect 5261 4097 5273 4131
rect 5307 4128 5319 4131
rect 5350 4128 5356 4140
rect 5307 4100 5356 4128
rect 5307 4097 5319 4100
rect 5261 4091 5319 4097
rect 5350 4088 5356 4100
rect 5408 4128 5414 4140
rect 5902 4128 5908 4140
rect 5408 4100 5580 4128
rect 5863 4100 5908 4128
rect 5408 4088 5414 4100
rect 2501 4063 2559 4069
rect 2501 4029 2513 4063
rect 2547 4029 2559 4063
rect 2774 4060 2780 4072
rect 2735 4032 2780 4060
rect 2501 4023 2559 4029
rect 2774 4020 2780 4032
rect 2832 4020 2838 4072
rect 5552 4069 5580 4100
rect 5902 4088 5908 4100
rect 5960 4088 5966 4140
rect 11790 4088 11796 4140
rect 11848 4128 11854 4140
rect 12805 4131 12863 4137
rect 12805 4128 12817 4131
rect 11848 4100 12817 4128
rect 11848 4088 11854 4100
rect 12805 4097 12817 4100
rect 12851 4128 12863 4131
rect 12894 4128 12900 4140
rect 12851 4100 12900 4128
rect 12851 4097 12863 4100
rect 12805 4091 12863 4097
rect 12894 4088 12900 4100
rect 12952 4088 12958 4140
rect 13004 4128 13032 4168
rect 13078 4156 13084 4208
rect 13136 4196 13142 4208
rect 13786 4196 13814 4236
rect 13909 4233 13921 4236
rect 13955 4264 13967 4267
rect 13955 4236 14641 4264
rect 13955 4233 13967 4236
rect 13909 4227 13967 4233
rect 13136 4168 13814 4196
rect 14613 4196 14641 4236
rect 15102 4224 15108 4276
rect 15160 4264 15166 4276
rect 18414 4264 18420 4276
rect 15160 4236 18420 4264
rect 15160 4224 15166 4236
rect 18414 4224 18420 4236
rect 18472 4224 18478 4276
rect 18506 4224 18512 4276
rect 18564 4264 18570 4276
rect 19061 4267 19119 4273
rect 19061 4264 19073 4267
rect 18564 4236 19073 4264
rect 18564 4224 18570 4236
rect 19061 4233 19073 4236
rect 19107 4233 19119 4267
rect 19061 4227 19119 4233
rect 14613 4168 19196 4196
rect 13136 4156 13142 4168
rect 16209 4131 16267 4137
rect 16209 4128 16221 4131
rect 13004 4100 16221 4128
rect 16209 4097 16221 4100
rect 16255 4128 16267 4131
rect 16298 4128 16304 4140
rect 16255 4100 16304 4128
rect 16255 4097 16267 4100
rect 16209 4091 16267 4097
rect 16298 4088 16304 4100
rect 16356 4088 16362 4140
rect 16482 4128 16488 4140
rect 16395 4100 16488 4128
rect 16482 4088 16488 4100
rect 16540 4128 16546 4140
rect 16758 4128 16764 4140
rect 16540 4100 16764 4128
rect 16540 4088 16546 4100
rect 16758 4088 16764 4100
rect 16816 4088 16822 4140
rect 19168 4128 19196 4168
rect 19751 4131 19809 4137
rect 19751 4128 19763 4131
rect 19168 4100 19763 4128
rect 19751 4097 19763 4100
rect 19797 4097 19809 4131
rect 19751 4091 19809 4097
rect 5537 4063 5595 4069
rect 5537 4029 5549 4063
rect 5583 4029 5595 4063
rect 5537 4023 5595 4029
rect 6825 4063 6883 4069
rect 6825 4029 6837 4063
rect 6871 4060 6883 4063
rect 7558 4060 7564 4072
rect 6871 4032 7564 4060
rect 6871 4029 6883 4032
rect 6825 4023 6883 4029
rect 7558 4020 7564 4032
rect 7616 4020 7622 4072
rect 8573 4063 8631 4069
rect 8573 4029 8585 4063
rect 8619 4060 8631 4063
rect 9030 4060 9036 4072
rect 8619 4032 9036 4060
rect 8619 4029 8631 4032
rect 8573 4023 8631 4029
rect 9030 4020 9036 4032
rect 9088 4020 9094 4072
rect 10505 4063 10563 4069
rect 10505 4029 10517 4063
rect 10551 4060 10563 4063
rect 11146 4060 11152 4072
rect 10551 4032 11152 4060
rect 10551 4029 10563 4032
rect 10505 4023 10563 4029
rect 11146 4020 11152 4032
rect 11204 4020 11210 4072
rect 11425 4063 11483 4069
rect 11425 4029 11437 4063
rect 11471 4060 11483 4063
rect 12161 4063 12219 4069
rect 12161 4060 12173 4063
rect 11471 4032 12173 4060
rect 11471 4029 11483 4032
rect 11425 4023 11483 4029
rect 12161 4029 12173 4032
rect 12207 4029 12219 4063
rect 12161 4023 12219 4029
rect 14645 4063 14703 4069
rect 14645 4029 14657 4063
rect 14691 4060 14703 4063
rect 14734 4060 14740 4072
rect 14691 4032 14740 4060
rect 14691 4029 14703 4032
rect 14645 4023 14703 4029
rect 2961 3995 3019 4001
rect 2961 3961 2973 3995
rect 3007 3992 3019 3995
rect 3418 3992 3424 4004
rect 3007 3964 3424 3992
rect 3007 3961 3019 3964
rect 2961 3955 3019 3961
rect 3418 3952 3424 3964
rect 3476 3952 3482 4004
rect 3881 3995 3939 4001
rect 3881 3992 3893 3995
rect 3620 3964 3893 3992
rect 3620 3936 3648 3964
rect 3881 3961 3893 3964
rect 3927 3961 3939 3995
rect 3881 3955 3939 3961
rect 3973 3995 4031 4001
rect 3973 3961 3985 3995
rect 4019 3992 4031 3995
rect 4154 3992 4160 4004
rect 4019 3964 4160 3992
rect 4019 3961 4031 3964
rect 3973 3955 4031 3961
rect 4154 3952 4160 3964
rect 4212 3952 4218 4004
rect 5353 3995 5411 4001
rect 5353 3961 5365 3995
rect 5399 3992 5411 3995
rect 5810 3992 5816 4004
rect 5399 3964 5816 3992
rect 5399 3961 5411 3964
rect 5353 3955 5411 3961
rect 5810 3952 5816 3964
rect 5868 3992 5874 4004
rect 6181 3995 6239 4001
rect 6181 3992 6193 3995
rect 5868 3964 6193 3992
rect 5868 3952 5874 3964
rect 6181 3961 6193 3964
rect 6227 3961 6239 3995
rect 7146 3995 7204 4001
rect 7146 3992 7158 3995
rect 6181 3955 6239 3961
rect 6564 3964 7158 3992
rect 6564 3936 6592 3964
rect 7146 3961 7158 3964
rect 7192 3992 7204 3995
rect 7834 3992 7840 4004
rect 7192 3964 7840 3992
rect 7192 3961 7204 3964
rect 7146 3955 7204 3961
rect 7834 3952 7840 3964
rect 7892 3992 7898 4004
rect 8389 3995 8447 4001
rect 8389 3992 8401 3995
rect 7892 3964 8401 3992
rect 7892 3952 7898 3964
rect 8389 3961 8401 3964
rect 8435 3992 8447 3995
rect 8894 3995 8952 4001
rect 8894 3992 8906 3995
rect 8435 3964 8906 3992
rect 8435 3961 8447 3964
rect 8389 3955 8447 3961
rect 8894 3961 8906 3964
rect 8940 3992 8952 3995
rect 10321 3995 10379 4001
rect 10321 3992 10333 3995
rect 8940 3964 10333 3992
rect 8940 3961 8952 3964
rect 8894 3955 8952 3961
rect 10321 3961 10333 3964
rect 10367 3992 10379 3995
rect 10826 3995 10884 4001
rect 10826 3992 10838 3995
rect 10367 3964 10838 3992
rect 10367 3961 10379 3964
rect 10321 3955 10379 3961
rect 10826 3961 10838 3964
rect 10872 3961 10884 3995
rect 10826 3955 10884 3961
rect 3602 3924 3608 3936
rect 3563 3896 3608 3924
rect 3602 3884 3608 3896
rect 3660 3884 3666 3936
rect 6546 3924 6552 3936
rect 6507 3896 6552 3924
rect 6546 3884 6552 3896
rect 6604 3884 6610 3936
rect 6638 3884 6644 3936
rect 6696 3924 6702 3936
rect 7745 3927 7803 3933
rect 7745 3924 7757 3927
rect 6696 3896 7757 3924
rect 6696 3884 6702 3896
rect 7745 3893 7757 3896
rect 7791 3893 7803 3927
rect 11698 3924 11704 3936
rect 11659 3896 11704 3924
rect 7745 3887 7803 3893
rect 11698 3884 11704 3896
rect 11756 3884 11762 3936
rect 12176 3924 12204 4023
rect 14734 4020 14740 4032
rect 14792 4020 14798 4072
rect 15565 4063 15623 4069
rect 15565 4029 15577 4063
rect 15611 4060 15623 4063
rect 18138 4060 18144 4072
rect 15611 4032 16344 4060
rect 18099 4032 18144 4060
rect 15611 4029 15623 4032
rect 15565 4023 15623 4029
rect 12342 3952 12348 4004
rect 12400 3992 12406 4004
rect 12529 3995 12587 4001
rect 12529 3992 12541 3995
rect 12400 3964 12541 3992
rect 12400 3952 12406 3964
rect 12529 3961 12541 3964
rect 12575 3961 12587 3995
rect 12529 3955 12587 3961
rect 12621 3995 12679 4001
rect 12621 3961 12633 3995
rect 12667 3961 12679 3995
rect 12621 3955 12679 3961
rect 12636 3924 12664 3955
rect 14182 3952 14188 4004
rect 14240 3992 14246 4004
rect 15470 3992 15476 4004
rect 14240 3964 15476 3992
rect 14240 3952 14246 3964
rect 15470 3952 15476 3964
rect 15528 3992 15534 4004
rect 15841 3995 15899 4001
rect 15841 3992 15853 3995
rect 15528 3964 15853 3992
rect 15528 3952 15534 3964
rect 15841 3961 15853 3964
rect 15887 3961 15899 3995
rect 15841 3955 15899 3961
rect 13262 3924 13268 3936
rect 12176 3896 13268 3924
rect 13262 3884 13268 3896
rect 13320 3924 13326 3936
rect 13449 3927 13507 3933
rect 13449 3924 13461 3927
rect 13320 3896 13461 3924
rect 13320 3884 13326 3896
rect 13449 3893 13461 3896
rect 13495 3893 13507 3927
rect 13449 3887 13507 3893
rect 14090 3884 14096 3936
rect 14148 3924 14154 3936
rect 14553 3927 14611 3933
rect 14553 3924 14565 3927
rect 14148 3896 14565 3924
rect 14148 3884 14154 3896
rect 14553 3893 14565 3896
rect 14599 3924 14611 3927
rect 15013 3927 15071 3933
rect 15013 3924 15025 3927
rect 14599 3896 15025 3924
rect 14599 3893 14611 3896
rect 14553 3887 14611 3893
rect 15013 3893 15025 3896
rect 15059 3893 15071 3927
rect 15013 3887 15071 3893
rect 15378 3884 15384 3936
rect 15436 3924 15442 3936
rect 16022 3924 16028 3936
rect 15436 3896 16028 3924
rect 15436 3884 15442 3896
rect 16022 3884 16028 3896
rect 16080 3884 16086 3936
rect 16316 3924 16344 4032
rect 18138 4020 18144 4032
rect 18196 4020 18202 4072
rect 18509 4063 18567 4069
rect 18509 4029 18521 4063
rect 18555 4029 18567 4063
rect 18509 4023 18567 4029
rect 16574 3952 16580 4004
rect 16632 3992 16638 4004
rect 17126 3992 17132 4004
rect 16632 3964 16677 3992
rect 17087 3964 17132 3992
rect 16632 3952 16638 3964
rect 17126 3952 17132 3964
rect 17184 3952 17190 4004
rect 18524 3992 18552 4023
rect 18598 4020 18604 4072
rect 18656 4060 18662 4072
rect 19648 4063 19706 4069
rect 19648 4060 19660 4063
rect 18656 4032 19660 4060
rect 18656 4020 18662 4032
rect 19648 4029 19660 4032
rect 19694 4060 19706 4063
rect 20073 4063 20131 4069
rect 20073 4060 20085 4063
rect 19694 4032 20085 4060
rect 19694 4029 19706 4032
rect 19648 4023 19706 4029
rect 20073 4029 20085 4032
rect 20119 4029 20131 4063
rect 20073 4023 20131 4029
rect 17788 3964 18552 3992
rect 16592 3924 16620 3952
rect 16316 3896 16620 3924
rect 17310 3884 17316 3936
rect 17368 3924 17374 3936
rect 17405 3927 17463 3933
rect 17405 3924 17417 3927
rect 17368 3896 17417 3924
rect 17368 3884 17374 3896
rect 17405 3893 17417 3896
rect 17451 3893 17463 3927
rect 17405 3887 17463 3893
rect 17678 3884 17684 3936
rect 17736 3924 17742 3936
rect 17788 3933 17816 3964
rect 17773 3927 17831 3933
rect 17773 3924 17785 3927
rect 17736 3896 17785 3924
rect 17736 3884 17742 3896
rect 17773 3893 17785 3896
rect 17819 3893 17831 3927
rect 18138 3924 18144 3936
rect 18099 3896 18144 3924
rect 17773 3887 17831 3893
rect 18138 3884 18144 3896
rect 18196 3884 18202 3936
rect 1104 3834 20884 3856
rect 1104 3782 8315 3834
rect 8367 3782 8379 3834
rect 8431 3782 8443 3834
rect 8495 3782 8507 3834
rect 8559 3782 15648 3834
rect 15700 3782 15712 3834
rect 15764 3782 15776 3834
rect 15828 3782 15840 3834
rect 15892 3782 20884 3834
rect 1104 3760 20884 3782
rect 1397 3723 1455 3729
rect 1397 3689 1409 3723
rect 1443 3720 1455 3723
rect 3602 3720 3608 3732
rect 1443 3692 3608 3720
rect 1443 3689 1455 3692
rect 1397 3683 1455 3689
rect 3602 3680 3608 3692
rect 3660 3680 3666 3732
rect 5258 3720 5264 3732
rect 5219 3692 5264 3720
rect 5258 3680 5264 3692
rect 5316 3680 5322 3732
rect 6638 3680 6644 3732
rect 6696 3720 6702 3732
rect 7101 3723 7159 3729
rect 7101 3720 7113 3723
rect 6696 3692 7113 3720
rect 6696 3680 6702 3692
rect 7101 3689 7113 3692
rect 7147 3689 7159 3723
rect 7101 3683 7159 3689
rect 7929 3723 7987 3729
rect 7929 3689 7941 3723
rect 7975 3720 7987 3723
rect 8110 3720 8116 3732
rect 7975 3692 8116 3720
rect 7975 3689 7987 3692
rect 7929 3683 7987 3689
rect 8110 3680 8116 3692
rect 8168 3680 8174 3732
rect 9030 3720 9036 3732
rect 8991 3692 9036 3720
rect 9030 3680 9036 3692
rect 9088 3720 9094 3732
rect 9769 3723 9827 3729
rect 9769 3720 9781 3723
rect 9088 3692 9781 3720
rect 9088 3680 9094 3692
rect 9769 3689 9781 3692
rect 9815 3689 9827 3723
rect 9769 3683 9827 3689
rect 10594 3680 10600 3732
rect 10652 3720 10658 3732
rect 13081 3723 13139 3729
rect 13081 3720 13093 3723
rect 10652 3692 13093 3720
rect 10652 3680 10658 3692
rect 13081 3689 13093 3692
rect 13127 3720 13139 3723
rect 14182 3720 14188 3732
rect 13127 3692 13308 3720
rect 14143 3692 14188 3720
rect 13127 3689 13139 3692
rect 13081 3683 13139 3689
rect 2038 3612 2044 3664
rect 2096 3652 2102 3664
rect 2317 3655 2375 3661
rect 2317 3652 2329 3655
rect 2096 3624 2329 3652
rect 2096 3612 2102 3624
rect 2317 3621 2329 3624
rect 2363 3652 2375 3655
rect 2774 3652 2780 3664
rect 2363 3624 2780 3652
rect 2363 3621 2375 3624
rect 2317 3615 2375 3621
rect 2774 3612 2780 3624
rect 2832 3612 2838 3664
rect 3418 3652 3424 3664
rect 3379 3624 3424 3652
rect 3418 3612 3424 3624
rect 3476 3612 3482 3664
rect 3786 3612 3792 3664
rect 3844 3652 3850 3664
rect 4386 3655 4444 3661
rect 4386 3652 4398 3655
rect 3844 3624 4398 3652
rect 3844 3612 3850 3624
rect 4386 3621 4398 3624
rect 4432 3652 4444 3655
rect 4522 3652 4528 3664
rect 4432 3624 4528 3652
rect 4432 3621 4444 3624
rect 4386 3615 4444 3621
rect 4522 3612 4528 3624
rect 4580 3652 4586 3664
rect 6226 3655 6284 3661
rect 6226 3652 6238 3655
rect 4580 3624 6238 3652
rect 4580 3612 4586 3624
rect 6226 3621 6238 3624
rect 6272 3652 6284 3655
rect 6546 3652 6552 3664
rect 6272 3624 6552 3652
rect 6272 3621 6284 3624
rect 6226 3615 6284 3621
rect 6546 3612 6552 3624
rect 6604 3612 6610 3664
rect 8202 3652 8208 3664
rect 8163 3624 8208 3652
rect 8202 3612 8208 3624
rect 8260 3612 8266 3664
rect 9398 3652 9404 3664
rect 9359 3624 9404 3652
rect 9398 3612 9404 3624
rect 9456 3612 9462 3664
rect 11606 3652 11612 3664
rect 11567 3624 11612 3652
rect 11606 3612 11612 3624
rect 11664 3612 11670 3664
rect 12161 3655 12219 3661
rect 12161 3621 12173 3655
rect 12207 3652 12219 3655
rect 12250 3652 12256 3664
rect 12207 3624 12256 3652
rect 12207 3621 12219 3624
rect 12161 3615 12219 3621
rect 2682 3584 2688 3596
rect 2643 3556 2688 3584
rect 2682 3544 2688 3556
rect 2740 3544 2746 3596
rect 2958 3584 2964 3596
rect 2919 3556 2964 3584
rect 2958 3544 2964 3556
rect 3016 3544 3022 3596
rect 3145 3519 3203 3525
rect 3145 3485 3157 3519
rect 3191 3516 3203 3519
rect 3326 3516 3332 3528
rect 3191 3488 3332 3516
rect 3191 3485 3203 3488
rect 3145 3479 3203 3485
rect 3326 3476 3332 3488
rect 3384 3476 3390 3528
rect 3436 3516 3464 3612
rect 3881 3587 3939 3593
rect 3881 3553 3893 3587
rect 3927 3584 3939 3587
rect 4154 3584 4160 3596
rect 3927 3556 4160 3584
rect 3927 3553 3939 3556
rect 3881 3547 3939 3553
rect 4154 3544 4160 3556
rect 4212 3584 4218 3596
rect 4985 3587 5043 3593
rect 4985 3584 4997 3587
rect 4212 3556 4997 3584
rect 4212 3544 4218 3556
rect 4985 3553 4997 3556
rect 5031 3553 5043 3587
rect 4985 3547 5043 3553
rect 9582 3544 9588 3596
rect 9640 3584 9646 3596
rect 9950 3584 9956 3596
rect 9640 3556 9956 3584
rect 9640 3544 9646 3556
rect 9950 3544 9956 3556
rect 10008 3544 10014 3596
rect 10042 3544 10048 3596
rect 10100 3584 10106 3596
rect 10137 3587 10195 3593
rect 10137 3584 10149 3587
rect 10100 3556 10149 3584
rect 10100 3544 10106 3556
rect 10137 3553 10149 3556
rect 10183 3584 10195 3587
rect 10318 3584 10324 3596
rect 10183 3556 10324 3584
rect 10183 3553 10195 3556
rect 10137 3547 10195 3553
rect 10318 3544 10324 3556
rect 10376 3544 10382 3596
rect 4065 3519 4123 3525
rect 4065 3516 4077 3519
rect 3436 3488 4077 3516
rect 4065 3485 4077 3488
rect 4111 3485 4123 3519
rect 4065 3479 4123 3485
rect 5905 3519 5963 3525
rect 5905 3485 5917 3519
rect 5951 3516 5963 3519
rect 6362 3516 6368 3528
rect 5951 3488 6368 3516
rect 5951 3485 5963 3488
rect 5905 3479 5963 3485
rect 6362 3476 6368 3488
rect 6420 3476 6426 3528
rect 7466 3476 7472 3528
rect 7524 3476 7530 3528
rect 8110 3516 8116 3528
rect 8071 3488 8116 3516
rect 8110 3476 8116 3488
rect 8168 3476 8174 3528
rect 8389 3519 8447 3525
rect 8389 3516 8401 3519
rect 8220 3488 8401 3516
rect 1762 3408 1768 3460
rect 1820 3448 1826 3460
rect 1949 3451 2007 3457
rect 1949 3448 1961 3451
rect 1820 3420 1961 3448
rect 1820 3408 1826 3420
rect 1949 3417 1961 3420
rect 1995 3448 2007 3451
rect 5166 3448 5172 3460
rect 1995 3420 5172 3448
rect 1995 3417 2007 3420
rect 1949 3411 2007 3417
rect 5166 3408 5172 3420
rect 5224 3408 5230 3460
rect 5350 3408 5356 3460
rect 5408 3448 5414 3460
rect 6825 3451 6883 3457
rect 6825 3448 6837 3451
rect 5408 3420 6837 3448
rect 5408 3408 5414 3420
rect 6825 3417 6837 3420
rect 6871 3417 6883 3451
rect 7484 3448 7512 3476
rect 8220 3448 8248 3488
rect 8389 3485 8401 3488
rect 8435 3485 8447 3519
rect 11146 3516 11152 3528
rect 11107 3488 11152 3516
rect 8389 3479 8447 3485
rect 11146 3476 11152 3488
rect 11204 3476 11210 3528
rect 11517 3519 11575 3525
rect 11517 3485 11529 3519
rect 11563 3516 11575 3519
rect 11790 3516 11796 3528
rect 11563 3488 11796 3516
rect 11563 3485 11575 3488
rect 11517 3479 11575 3485
rect 11790 3476 11796 3488
rect 11848 3476 11854 3528
rect 7484 3420 8248 3448
rect 6825 3411 6883 3417
rect 9582 3408 9588 3460
rect 9640 3448 9646 3460
rect 12176 3448 12204 3615
rect 12250 3612 12256 3624
rect 12308 3612 12314 3664
rect 12342 3612 12348 3664
rect 12400 3652 12406 3664
rect 12437 3655 12495 3661
rect 12437 3652 12449 3655
rect 12400 3624 12449 3652
rect 12400 3612 12406 3624
rect 12437 3621 12449 3624
rect 12483 3621 12495 3655
rect 12437 3615 12495 3621
rect 13280 3593 13308 3692
rect 14182 3680 14188 3692
rect 14240 3680 14246 3732
rect 15102 3720 15108 3732
rect 15063 3692 15108 3720
rect 15102 3680 15108 3692
rect 15160 3680 15166 3732
rect 16485 3723 16543 3729
rect 15212 3692 15700 3720
rect 13627 3655 13685 3661
rect 13627 3621 13639 3655
rect 13673 3652 13685 3655
rect 13814 3652 13820 3664
rect 13673 3624 13820 3652
rect 13673 3621 13685 3624
rect 13627 3615 13685 3621
rect 13814 3612 13820 3624
rect 13872 3612 13878 3664
rect 14645 3655 14703 3661
rect 14645 3621 14657 3655
rect 14691 3652 14703 3655
rect 14734 3652 14740 3664
rect 14691 3624 14740 3652
rect 14691 3621 14703 3624
rect 14645 3615 14703 3621
rect 14734 3612 14740 3624
rect 14792 3652 14798 3664
rect 15212 3652 15240 3692
rect 15470 3652 15476 3664
rect 14792 3624 15240 3652
rect 15431 3624 15476 3652
rect 14792 3612 14798 3624
rect 15470 3612 15476 3624
rect 15528 3612 15534 3664
rect 15672 3652 15700 3692
rect 16485 3689 16497 3723
rect 16531 3720 16543 3723
rect 16574 3720 16580 3732
rect 16531 3692 16580 3720
rect 16531 3689 16543 3692
rect 16485 3683 16543 3689
rect 16574 3680 16580 3692
rect 16632 3680 16638 3732
rect 18506 3720 18512 3732
rect 18467 3692 18512 3720
rect 18506 3680 18512 3692
rect 18564 3680 18570 3732
rect 16942 3652 16948 3664
rect 15672 3624 16948 3652
rect 16942 3612 16948 3624
rect 17000 3612 17006 3664
rect 13265 3587 13323 3593
rect 13265 3553 13277 3587
rect 13311 3553 13323 3587
rect 13265 3547 13323 3553
rect 17129 3587 17187 3593
rect 17129 3553 17141 3587
rect 17175 3584 17187 3587
rect 17218 3584 17224 3596
rect 17175 3556 17224 3584
rect 17175 3553 17187 3556
rect 17129 3547 17187 3553
rect 17218 3544 17224 3556
rect 17276 3544 17282 3596
rect 17310 3544 17316 3596
rect 17368 3584 17374 3596
rect 17368 3556 17413 3584
rect 17368 3544 17374 3556
rect 17770 3544 17776 3596
rect 17828 3584 17834 3596
rect 18417 3587 18475 3593
rect 18417 3584 18429 3587
rect 17828 3556 18429 3584
rect 17828 3544 17834 3556
rect 18417 3553 18429 3556
rect 18463 3584 18475 3587
rect 18782 3584 18788 3596
rect 18463 3556 18788 3584
rect 18463 3553 18475 3556
rect 18417 3547 18475 3553
rect 18782 3544 18788 3556
rect 18840 3544 18846 3596
rect 18966 3584 18972 3596
rect 18927 3556 18972 3584
rect 18966 3544 18972 3556
rect 19024 3544 19030 3596
rect 15378 3516 15384 3528
rect 15339 3488 15384 3516
rect 15378 3476 15384 3488
rect 15436 3476 15442 3528
rect 17405 3519 17463 3525
rect 17405 3516 17417 3519
rect 15488 3488 17417 3516
rect 9640 3420 12204 3448
rect 9640 3408 9646 3420
rect 13354 3408 13360 3460
rect 13412 3448 13418 3460
rect 15488 3448 15516 3488
rect 17405 3485 17417 3488
rect 17451 3485 17463 3519
rect 17405 3479 17463 3485
rect 15930 3448 15936 3460
rect 13412 3420 15516 3448
rect 15891 3420 15936 3448
rect 13412 3408 13418 3420
rect 15930 3408 15936 3420
rect 15988 3408 15994 3460
rect 16040 3420 18184 3448
rect 5813 3383 5871 3389
rect 5813 3349 5825 3383
rect 5859 3380 5871 3383
rect 7098 3380 7104 3392
rect 5859 3352 7104 3380
rect 5859 3349 5871 3352
rect 5813 3343 5871 3349
rect 7098 3340 7104 3352
rect 7156 3340 7162 3392
rect 7558 3380 7564 3392
rect 7519 3352 7564 3380
rect 7558 3340 7564 3352
rect 7616 3340 7622 3392
rect 8110 3340 8116 3392
rect 8168 3380 8174 3392
rect 9398 3380 9404 3392
rect 8168 3352 9404 3380
rect 8168 3340 8174 3352
rect 9398 3340 9404 3352
rect 9456 3340 9462 3392
rect 9858 3340 9864 3392
rect 9916 3380 9922 3392
rect 10781 3383 10839 3389
rect 10781 3380 10793 3383
rect 9916 3352 10793 3380
rect 9916 3340 9922 3352
rect 10781 3349 10793 3352
rect 10827 3380 10839 3383
rect 16040 3380 16068 3420
rect 18156 3392 18184 3420
rect 10827 3352 16068 3380
rect 10827 3349 10839 3352
rect 10781 3343 10839 3349
rect 16482 3340 16488 3392
rect 16540 3380 16546 3392
rect 17678 3380 17684 3392
rect 16540 3352 17684 3380
rect 16540 3340 16546 3352
rect 17678 3340 17684 3352
rect 17736 3340 17742 3392
rect 18138 3380 18144 3392
rect 18099 3352 18144 3380
rect 18138 3340 18144 3352
rect 18196 3340 18202 3392
rect 1104 3290 20884 3312
rect 1104 3238 4648 3290
rect 4700 3238 4712 3290
rect 4764 3238 4776 3290
rect 4828 3238 4840 3290
rect 4892 3238 11982 3290
rect 12034 3238 12046 3290
rect 12098 3238 12110 3290
rect 12162 3238 12174 3290
rect 12226 3238 19315 3290
rect 19367 3238 19379 3290
rect 19431 3238 19443 3290
rect 19495 3238 19507 3290
rect 19559 3238 20884 3290
rect 1104 3216 20884 3238
rect 2682 3136 2688 3188
rect 2740 3176 2746 3188
rect 2869 3179 2927 3185
rect 2869 3176 2881 3179
rect 2740 3148 2881 3176
rect 2740 3136 2746 3148
rect 2869 3145 2881 3148
rect 2915 3145 2927 3179
rect 2869 3139 2927 3145
rect 8113 3179 8171 3185
rect 8113 3145 8125 3179
rect 8159 3176 8171 3179
rect 8202 3176 8208 3188
rect 8159 3148 8208 3176
rect 8159 3145 8171 3148
rect 8113 3139 8171 3145
rect 8202 3136 8208 3148
rect 8260 3136 8266 3188
rect 8757 3179 8815 3185
rect 8757 3145 8769 3179
rect 8803 3176 8815 3179
rect 8846 3176 8852 3188
rect 8803 3148 8852 3176
rect 8803 3145 8815 3148
rect 8757 3139 8815 3145
rect 8846 3136 8852 3148
rect 8904 3136 8910 3188
rect 11425 3179 11483 3185
rect 11425 3145 11437 3179
rect 11471 3176 11483 3179
rect 11698 3176 11704 3188
rect 11471 3148 11704 3176
rect 11471 3145 11483 3148
rect 11425 3139 11483 3145
rect 11698 3136 11704 3148
rect 11756 3136 11762 3188
rect 13078 3176 13084 3188
rect 13039 3148 13084 3176
rect 13078 3136 13084 3148
rect 13136 3136 13142 3188
rect 14829 3179 14887 3185
rect 14829 3145 14841 3179
rect 14875 3176 14887 3179
rect 15197 3179 15255 3185
rect 15197 3176 15209 3179
rect 14875 3148 15209 3176
rect 14875 3145 14887 3148
rect 14829 3139 14887 3145
rect 15197 3145 15209 3148
rect 15243 3176 15255 3179
rect 15470 3176 15476 3188
rect 15243 3148 15476 3176
rect 15243 3145 15255 3148
rect 15197 3139 15255 3145
rect 15470 3136 15476 3148
rect 15528 3136 15534 3188
rect 15565 3179 15623 3185
rect 15565 3145 15577 3179
rect 15611 3176 15623 3179
rect 15838 3176 15844 3188
rect 15611 3148 15844 3176
rect 15611 3145 15623 3148
rect 15565 3139 15623 3145
rect 15838 3136 15844 3148
rect 15896 3176 15902 3188
rect 16574 3176 16580 3188
rect 15896 3148 16580 3176
rect 15896 3136 15902 3148
rect 16574 3136 16580 3148
rect 16632 3136 16638 3188
rect 17218 3176 17224 3188
rect 17179 3148 17224 3176
rect 17218 3136 17224 3148
rect 17276 3136 17282 3188
rect 18966 3136 18972 3188
rect 19024 3176 19030 3188
rect 19429 3179 19487 3185
rect 19429 3176 19441 3179
rect 19024 3148 19441 3176
rect 19024 3136 19030 3148
rect 19429 3145 19441 3148
rect 19475 3176 19487 3179
rect 19702 3176 19708 3188
rect 19475 3148 19708 3176
rect 19475 3145 19487 3148
rect 19429 3139 19487 3145
rect 19702 3136 19708 3148
rect 19760 3136 19766 3188
rect 4522 3068 4528 3120
rect 4580 3108 4586 3120
rect 4617 3111 4675 3117
rect 4617 3108 4629 3111
rect 4580 3080 4629 3108
rect 4580 3068 4586 3080
rect 4617 3077 4629 3080
rect 4663 3077 4675 3111
rect 6549 3111 6607 3117
rect 6549 3108 6561 3111
rect 4617 3071 4675 3077
rect 5092 3080 6561 3108
rect 1394 3000 1400 3052
rect 1452 3040 1458 3052
rect 5092 3040 5120 3080
rect 6549 3077 6561 3080
rect 6595 3077 6607 3111
rect 6549 3071 6607 3077
rect 5258 3040 5264 3052
rect 1452 3012 5120 3040
rect 5219 3012 5264 3040
rect 1452 3000 1458 3012
rect 5258 3000 5264 3012
rect 5316 3000 5322 3052
rect 6564 3040 6592 3071
rect 6917 3043 6975 3049
rect 6917 3040 6929 3043
rect 6564 3012 6929 3040
rect 6917 3009 6929 3012
rect 6963 3009 6975 3043
rect 6917 3003 6975 3009
rect 7098 3000 7104 3052
rect 7156 3040 7162 3052
rect 8864 3040 8892 3136
rect 9030 3068 9036 3120
rect 9088 3108 9094 3120
rect 9088 3080 10548 3108
rect 9088 3068 9094 3080
rect 8941 3043 8999 3049
rect 8941 3040 8953 3043
rect 7156 3012 8064 3040
rect 8864 3012 8953 3040
rect 7156 3000 7162 3012
rect 1762 2972 1768 2984
rect 1723 2944 1768 2972
rect 1762 2932 1768 2944
rect 1820 2932 1826 2984
rect 2038 2972 2044 2984
rect 1999 2944 2044 2972
rect 2038 2932 2044 2944
rect 2096 2932 2102 2984
rect 2225 2975 2283 2981
rect 2225 2941 2237 2975
rect 2271 2972 2283 2975
rect 2866 2972 2872 2984
rect 2271 2944 2872 2972
rect 2271 2941 2283 2944
rect 2225 2935 2283 2941
rect 2866 2932 2872 2944
rect 2924 2932 2930 2984
rect 3602 2972 3608 2984
rect 3563 2944 3608 2972
rect 3602 2932 3608 2944
rect 3660 2932 3666 2984
rect 4203 2975 4261 2981
rect 4203 2941 4215 2975
rect 4249 2972 4261 2975
rect 4982 2972 4988 2984
rect 4249 2944 4988 2972
rect 4249 2941 4261 2944
rect 4203 2935 4261 2941
rect 2593 2839 2651 2845
rect 2593 2805 2605 2839
rect 2639 2836 2651 2839
rect 2958 2836 2964 2848
rect 2639 2808 2964 2836
rect 2639 2805 2651 2808
rect 2593 2799 2651 2805
rect 2958 2796 2964 2808
rect 3016 2836 3022 2848
rect 3513 2839 3571 2845
rect 3513 2836 3525 2839
rect 3016 2808 3525 2836
rect 3016 2796 3022 2808
rect 3513 2805 3525 2808
rect 3559 2836 3571 2839
rect 4218 2836 4246 2935
rect 4982 2932 4988 2944
rect 5040 2932 5046 2984
rect 4338 2904 4344 2916
rect 4299 2876 4344 2904
rect 4338 2864 4344 2876
rect 4396 2864 4402 2916
rect 5077 2907 5135 2913
rect 5077 2873 5089 2907
rect 5123 2904 5135 2907
rect 5350 2904 5356 2916
rect 5123 2876 5356 2904
rect 5123 2873 5135 2876
rect 5077 2867 5135 2873
rect 5350 2864 5356 2876
rect 5408 2864 5414 2916
rect 5905 2907 5963 2913
rect 5905 2873 5917 2907
rect 5951 2904 5963 2907
rect 5951 2876 6960 2904
rect 5951 2873 5963 2876
rect 5905 2867 5963 2873
rect 3559 2808 4246 2836
rect 3559 2805 3571 2808
rect 3513 2799 3571 2805
rect 4522 2796 4528 2848
rect 4580 2836 4586 2848
rect 5258 2836 5264 2848
rect 4580 2808 5264 2836
rect 4580 2796 4586 2808
rect 5258 2796 5264 2808
rect 5316 2836 5322 2848
rect 6181 2839 6239 2845
rect 6181 2836 6193 2839
rect 5316 2808 6193 2836
rect 5316 2796 5322 2808
rect 6181 2805 6193 2808
rect 6227 2805 6239 2839
rect 6932 2836 6960 2876
rect 7006 2864 7012 2916
rect 7064 2904 7070 2916
rect 7561 2907 7619 2913
rect 7064 2876 7109 2904
rect 7064 2864 7070 2876
rect 7561 2873 7573 2907
rect 7607 2873 7619 2907
rect 7561 2867 7619 2873
rect 7282 2836 7288 2848
rect 6932 2808 7288 2836
rect 6181 2799 6239 2805
rect 7282 2796 7288 2808
rect 7340 2836 7346 2848
rect 7576 2836 7604 2867
rect 7340 2808 7604 2836
rect 8036 2836 8064 3012
rect 8941 3009 8953 3012
rect 8987 3009 8999 3043
rect 9950 3040 9956 3052
rect 9911 3012 9956 3040
rect 8941 3003 8999 3009
rect 9950 3000 9956 3012
rect 10008 3000 10014 3052
rect 10520 3049 10548 3080
rect 10870 3068 10876 3120
rect 10928 3108 10934 3120
rect 12621 3111 12679 3117
rect 12621 3108 12633 3111
rect 10928 3080 12633 3108
rect 10928 3068 10934 3080
rect 12621 3077 12633 3080
rect 12667 3077 12679 3111
rect 12621 3071 12679 3077
rect 16945 3111 17003 3117
rect 16945 3077 16957 3111
rect 16991 3108 17003 3111
rect 17310 3108 17316 3120
rect 16991 3080 17316 3108
rect 16991 3077 17003 3080
rect 16945 3071 17003 3077
rect 17310 3068 17316 3080
rect 17368 3068 17374 3120
rect 10505 3043 10563 3049
rect 10505 3009 10517 3043
rect 10551 3040 10563 3043
rect 11701 3043 11759 3049
rect 11701 3040 11713 3043
rect 10551 3012 11713 3040
rect 10551 3009 10563 3012
rect 10505 3003 10563 3009
rect 11701 3009 11713 3012
rect 11747 3009 11759 3043
rect 11701 3003 11759 3009
rect 12176 3012 13814 3040
rect 11422 2932 11428 2984
rect 11480 2972 11486 2984
rect 12176 2972 12204 3012
rect 12434 2972 12440 2984
rect 11480 2944 12204 2972
rect 12347 2944 12440 2972
rect 11480 2932 11486 2944
rect 12434 2932 12440 2944
rect 12492 2972 12498 2984
rect 13078 2972 13084 2984
rect 12492 2944 13084 2972
rect 12492 2932 12498 2944
rect 13078 2932 13084 2944
rect 13136 2932 13142 2984
rect 13786 2972 13814 3012
rect 15102 3000 15108 3052
rect 15160 3040 15166 3052
rect 15749 3043 15807 3049
rect 15749 3040 15761 3043
rect 15160 3012 15761 3040
rect 15160 3000 15166 3012
rect 15749 3009 15761 3012
rect 15795 3009 15807 3043
rect 16390 3040 16396 3052
rect 16351 3012 16396 3040
rect 15749 3003 15807 3009
rect 16390 3000 16396 3012
rect 16448 3000 16454 3052
rect 16758 3000 16764 3052
rect 16816 3040 16822 3052
rect 19751 3043 19809 3049
rect 19751 3040 19763 3043
rect 16816 3012 19763 3040
rect 16816 3000 16822 3012
rect 19751 3009 19763 3012
rect 19797 3009 19809 3043
rect 19751 3003 19809 3009
rect 13906 2972 13912 2984
rect 13786 2944 13912 2972
rect 13906 2932 13912 2944
rect 13964 2932 13970 2984
rect 17770 2932 17776 2984
rect 17828 2972 17834 2984
rect 18049 2975 18107 2981
rect 18049 2972 18061 2975
rect 17828 2944 18061 2972
rect 17828 2932 17834 2944
rect 18049 2941 18061 2944
rect 18095 2941 18107 2975
rect 18049 2935 18107 2941
rect 9030 2864 9036 2916
rect 9088 2904 9094 2916
rect 9582 2904 9588 2916
rect 9088 2876 9133 2904
rect 9495 2876 9588 2904
rect 9088 2864 9094 2876
rect 9582 2864 9588 2876
rect 9640 2864 9646 2916
rect 10826 2907 10884 2913
rect 10826 2904 10838 2907
rect 10336 2876 10838 2904
rect 9600 2836 9628 2864
rect 10336 2848 10364 2876
rect 10826 2873 10838 2876
rect 10872 2873 10884 2907
rect 13725 2907 13783 2913
rect 13725 2904 13737 2907
rect 10826 2867 10884 2873
rect 13372 2876 13737 2904
rect 10318 2836 10324 2848
rect 8036 2808 9628 2836
rect 10279 2808 10324 2836
rect 7340 2796 7346 2808
rect 10318 2796 10324 2808
rect 10376 2796 10382 2848
rect 12066 2836 12072 2848
rect 12027 2808 12072 2836
rect 12066 2796 12072 2808
rect 12124 2796 12130 2848
rect 13262 2796 13268 2848
rect 13320 2836 13326 2848
rect 13372 2845 13400 2876
rect 13725 2873 13737 2876
rect 13771 2873 13783 2907
rect 13725 2867 13783 2873
rect 13814 2864 13820 2916
rect 13872 2904 13878 2916
rect 14230 2907 14288 2913
rect 14230 2904 14242 2907
rect 13872 2876 14242 2904
rect 13872 2864 13878 2876
rect 14230 2873 14242 2876
rect 14276 2873 14288 2907
rect 15838 2904 15844 2916
rect 15799 2876 15844 2904
rect 14230 2867 14288 2873
rect 15838 2864 15844 2876
rect 15896 2864 15902 2916
rect 18064 2904 18092 2935
rect 18138 2932 18144 2984
rect 18196 2972 18202 2984
rect 18509 2975 18567 2981
rect 18509 2972 18521 2975
rect 18196 2944 18521 2972
rect 18196 2932 18202 2944
rect 18509 2941 18521 2944
rect 18555 2941 18567 2975
rect 18509 2935 18567 2941
rect 19664 2975 19722 2981
rect 19664 2941 19676 2975
rect 19710 2972 19722 2975
rect 20070 2972 20076 2984
rect 19710 2944 20076 2972
rect 19710 2941 19722 2944
rect 19664 2935 19722 2941
rect 19812 2916 19840 2944
rect 20070 2932 20076 2944
rect 20128 2932 20134 2984
rect 19061 2907 19119 2913
rect 19061 2904 19073 2907
rect 18064 2876 19073 2904
rect 19061 2873 19073 2876
rect 19107 2873 19119 2907
rect 19061 2867 19119 2873
rect 19794 2864 19800 2916
rect 19852 2864 19858 2916
rect 13357 2839 13415 2845
rect 13357 2836 13369 2839
rect 13320 2808 13369 2836
rect 13320 2796 13326 2808
rect 13357 2805 13369 2808
rect 13403 2805 13415 2839
rect 17770 2836 17776 2848
rect 17731 2808 17776 2836
rect 13357 2799 13415 2805
rect 17770 2796 17776 2808
rect 17828 2796 17834 2848
rect 18138 2836 18144 2848
rect 18099 2808 18144 2836
rect 18138 2796 18144 2808
rect 18196 2796 18202 2848
rect 1104 2746 20884 2768
rect 1104 2694 8315 2746
rect 8367 2694 8379 2746
rect 8431 2694 8443 2746
rect 8495 2694 8507 2746
rect 8559 2694 15648 2746
rect 15700 2694 15712 2746
rect 15764 2694 15776 2746
rect 15828 2694 15840 2746
rect 15892 2694 20884 2746
rect 1104 2672 20884 2694
rect 1394 2632 1400 2644
rect 1355 2604 1400 2632
rect 1394 2592 1400 2604
rect 1452 2592 1458 2644
rect 3602 2632 3608 2644
rect 3563 2604 3608 2632
rect 3602 2592 3608 2604
rect 3660 2592 3666 2644
rect 4338 2592 4344 2644
rect 4396 2632 4402 2644
rect 5997 2635 6055 2641
rect 4396 2604 5580 2632
rect 4396 2592 4402 2604
rect 2317 2567 2375 2573
rect 2317 2533 2329 2567
rect 2363 2564 2375 2567
rect 3142 2564 3148 2576
rect 2363 2536 3004 2564
rect 3103 2536 3148 2564
rect 2363 2533 2375 2536
rect 2317 2527 2375 2533
rect 2976 2508 3004 2536
rect 3142 2524 3148 2536
rect 3200 2524 3206 2576
rect 4617 2567 4675 2573
rect 4617 2533 4629 2567
rect 4663 2564 4675 2567
rect 4663 2536 5120 2564
rect 4663 2533 4675 2536
rect 4617 2527 4675 2533
rect 1949 2499 2007 2505
rect 1949 2465 1961 2499
rect 1995 2496 2007 2499
rect 2498 2496 2504 2508
rect 1995 2468 2504 2496
rect 1995 2465 2007 2468
rect 1949 2459 2007 2465
rect 2498 2456 2504 2468
rect 2556 2456 2562 2508
rect 2958 2496 2964 2508
rect 2919 2468 2964 2496
rect 2958 2456 2964 2468
rect 3016 2456 3022 2508
rect 4132 2499 4190 2505
rect 4132 2465 4144 2499
rect 4178 2496 4190 2499
rect 4890 2496 4896 2508
rect 4178 2468 4896 2496
rect 4178 2465 4190 2468
rect 4132 2459 4190 2465
rect 4890 2456 4896 2468
rect 4948 2456 4954 2508
rect 5092 2505 5120 2536
rect 5258 2524 5264 2576
rect 5316 2564 5322 2576
rect 5398 2567 5456 2573
rect 5398 2564 5410 2567
rect 5316 2536 5410 2564
rect 5316 2524 5322 2536
rect 5398 2533 5410 2536
rect 5444 2533 5456 2567
rect 5552 2564 5580 2604
rect 5997 2601 6009 2635
rect 6043 2632 6055 2635
rect 7006 2632 7012 2644
rect 6043 2604 7012 2632
rect 6043 2601 6055 2604
rect 5997 2595 6055 2601
rect 7006 2592 7012 2604
rect 7064 2632 7070 2644
rect 7377 2635 7435 2641
rect 7377 2632 7389 2635
rect 7064 2604 7389 2632
rect 7064 2592 7070 2604
rect 7377 2601 7389 2604
rect 7423 2601 7435 2635
rect 7834 2632 7840 2644
rect 7795 2604 7840 2632
rect 7377 2595 7435 2601
rect 7834 2592 7840 2604
rect 7892 2632 7898 2644
rect 8849 2635 8907 2641
rect 7892 2604 8293 2632
rect 7892 2592 7898 2604
rect 6730 2564 6736 2576
rect 5552 2536 6736 2564
rect 5398 2527 5456 2533
rect 6730 2524 6736 2536
rect 6788 2524 6794 2576
rect 7190 2524 7196 2576
rect 7248 2564 7254 2576
rect 8265 2573 8293 2604
rect 8849 2601 8861 2635
rect 8895 2632 8907 2635
rect 9030 2632 9036 2644
rect 8895 2604 9036 2632
rect 8895 2601 8907 2604
rect 8849 2595 8907 2601
rect 9030 2592 9036 2604
rect 9088 2632 9094 2644
rect 9125 2635 9183 2641
rect 9125 2632 9137 2635
rect 9088 2604 9137 2632
rect 9088 2592 9094 2604
rect 9125 2601 9137 2604
rect 9171 2601 9183 2635
rect 10042 2632 10048 2644
rect 10003 2604 10048 2632
rect 9125 2595 9183 2601
rect 10042 2592 10048 2604
rect 10100 2592 10106 2644
rect 11425 2635 11483 2641
rect 11425 2601 11437 2635
rect 11471 2632 11483 2635
rect 11606 2632 11612 2644
rect 11471 2604 11612 2632
rect 11471 2601 11483 2604
rect 11425 2595 11483 2601
rect 11606 2592 11612 2604
rect 11664 2632 11670 2644
rect 12066 2632 12072 2644
rect 11664 2604 12072 2632
rect 11664 2592 11670 2604
rect 12066 2592 12072 2604
rect 12124 2592 12130 2644
rect 14277 2635 14335 2641
rect 14277 2601 14289 2635
rect 14323 2632 14335 2635
rect 16945 2635 17003 2641
rect 14323 2604 15700 2632
rect 14323 2601 14335 2604
rect 14277 2595 14335 2601
rect 8250 2567 8308 2573
rect 7248 2536 8156 2564
rect 7248 2524 7254 2536
rect 5077 2499 5135 2505
rect 5077 2465 5089 2499
rect 5123 2496 5135 2499
rect 6178 2496 6184 2508
rect 5123 2468 6184 2496
rect 5123 2465 5135 2468
rect 5077 2459 5135 2465
rect 6178 2456 6184 2468
rect 6236 2456 6242 2508
rect 6984 2499 7042 2505
rect 6984 2465 6996 2499
rect 7030 2496 7042 2499
rect 7098 2496 7104 2508
rect 7030 2468 7104 2496
rect 7030 2465 7042 2468
rect 6984 2459 7042 2465
rect 7098 2456 7104 2468
rect 7156 2456 7162 2508
rect 8128 2496 8156 2536
rect 8250 2533 8262 2567
rect 8296 2564 8308 2567
rect 10318 2564 10324 2576
rect 8296 2536 10324 2564
rect 8296 2533 8308 2536
rect 8250 2527 8308 2533
rect 10318 2524 10324 2536
rect 10376 2564 10382 2576
rect 10826 2567 10884 2573
rect 10826 2564 10838 2567
rect 10376 2536 10838 2564
rect 10376 2524 10382 2536
rect 10826 2533 10838 2536
rect 10872 2564 10884 2567
rect 13173 2567 13231 2573
rect 13173 2564 13185 2567
rect 10872 2536 13185 2564
rect 10872 2533 10884 2536
rect 10826 2527 10884 2533
rect 13173 2533 13185 2536
rect 13219 2564 13231 2567
rect 13262 2564 13268 2576
rect 13219 2536 13268 2564
rect 13219 2533 13231 2536
rect 13173 2527 13231 2533
rect 13262 2524 13268 2536
rect 13320 2564 13326 2576
rect 13678 2567 13736 2573
rect 13678 2564 13690 2567
rect 13320 2536 13690 2564
rect 13320 2524 13326 2536
rect 13678 2533 13690 2536
rect 13724 2564 13736 2567
rect 13814 2564 13820 2576
rect 13724 2536 13820 2564
rect 13724 2533 13736 2536
rect 13678 2527 13736 2533
rect 13814 2524 13820 2536
rect 13872 2524 13878 2576
rect 13906 2524 13912 2576
rect 13964 2564 13970 2576
rect 14553 2567 14611 2573
rect 14553 2564 14565 2567
rect 13964 2536 14565 2564
rect 13964 2524 13970 2536
rect 14553 2533 14565 2536
rect 14599 2533 14611 2567
rect 15562 2564 15568 2576
rect 14553 2527 14611 2533
rect 14660 2536 15568 2564
rect 10505 2499 10563 2505
rect 10505 2496 10517 2499
rect 8128 2468 10517 2496
rect 10505 2465 10517 2468
rect 10551 2496 10563 2499
rect 11701 2499 11759 2505
rect 11701 2496 11713 2499
rect 10551 2468 11713 2496
rect 10551 2465 10563 2468
rect 10505 2459 10563 2465
rect 11701 2465 11713 2468
rect 11747 2465 11759 2499
rect 11701 2459 11759 2465
rect 11790 2456 11796 2508
rect 11848 2496 11854 2508
rect 12069 2499 12127 2505
rect 12069 2496 12081 2499
rect 11848 2468 12081 2496
rect 11848 2456 11854 2468
rect 12069 2465 12081 2468
rect 12115 2465 12127 2499
rect 12069 2459 12127 2465
rect 12897 2499 12955 2505
rect 12897 2465 12909 2499
rect 12943 2496 12955 2499
rect 13354 2496 13360 2508
rect 12943 2468 13360 2496
rect 12943 2465 12955 2468
rect 12897 2459 12955 2465
rect 13354 2456 13360 2468
rect 13412 2456 13418 2508
rect 14660 2496 14688 2536
rect 15562 2524 15568 2536
rect 15620 2524 15626 2576
rect 15672 2573 15700 2604
rect 16945 2601 16957 2635
rect 16991 2632 17003 2635
rect 17126 2632 17132 2644
rect 16991 2604 17132 2632
rect 16991 2601 17003 2604
rect 16945 2595 17003 2601
rect 17126 2592 17132 2604
rect 17184 2592 17190 2644
rect 17770 2592 17776 2644
rect 17828 2632 17834 2644
rect 18049 2635 18107 2641
rect 18049 2632 18061 2635
rect 17828 2604 18061 2632
rect 17828 2592 17834 2604
rect 18049 2601 18061 2604
rect 18095 2601 18107 2635
rect 18414 2632 18420 2644
rect 18375 2604 18420 2632
rect 18049 2595 18107 2601
rect 15657 2567 15715 2573
rect 15657 2533 15669 2567
rect 15703 2564 15715 2567
rect 16485 2567 16543 2573
rect 16485 2564 16497 2567
rect 15703 2536 16497 2564
rect 15703 2533 15715 2536
rect 15657 2527 15715 2533
rect 16485 2533 16497 2536
rect 16531 2533 16543 2567
rect 16485 2527 16543 2533
rect 14429 2468 14688 2496
rect 6822 2388 6828 2440
rect 6880 2428 6886 2440
rect 7929 2431 7987 2437
rect 7929 2428 7941 2431
rect 6880 2400 7941 2428
rect 6880 2388 6886 2400
rect 7929 2397 7941 2400
rect 7975 2428 7987 2431
rect 9493 2431 9551 2437
rect 9493 2428 9505 2431
rect 7975 2400 9505 2428
rect 7975 2397 7987 2400
rect 7929 2391 7987 2397
rect 9493 2397 9505 2400
rect 9539 2397 9551 2431
rect 14429 2428 14457 2468
rect 17034 2456 17040 2508
rect 17092 2496 17098 2508
rect 17129 2499 17187 2505
rect 17129 2496 17141 2499
rect 17092 2468 17141 2496
rect 17092 2456 17098 2468
rect 17129 2465 17141 2468
rect 17175 2496 17187 2499
rect 17681 2499 17739 2505
rect 17681 2496 17693 2499
rect 17175 2468 17693 2496
rect 17175 2465 17187 2468
rect 17129 2459 17187 2465
rect 17681 2465 17693 2468
rect 17727 2465 17739 2499
rect 18064 2496 18092 2595
rect 18414 2592 18420 2604
rect 18472 2592 18478 2644
rect 18782 2524 18788 2576
rect 18840 2564 18846 2576
rect 19337 2567 19395 2573
rect 19337 2564 19349 2567
rect 18840 2536 19349 2564
rect 18840 2524 18846 2536
rect 18892 2505 18920 2536
rect 19337 2533 19349 2536
rect 19383 2533 19395 2567
rect 19337 2527 19395 2533
rect 18325 2499 18383 2505
rect 18325 2496 18337 2499
rect 18064 2468 18337 2496
rect 17681 2459 17739 2465
rect 18325 2465 18337 2468
rect 18371 2465 18383 2499
rect 18325 2459 18383 2465
rect 18877 2499 18935 2505
rect 18877 2465 18889 2499
rect 18923 2465 18935 2499
rect 18877 2459 18935 2465
rect 15565 2431 15623 2437
rect 15565 2428 15577 2431
rect 9493 2391 9551 2397
rect 9646 2400 14457 2428
rect 15304 2400 15577 2428
rect 4203 2363 4261 2369
rect 4203 2329 4215 2363
rect 4249 2360 4261 2363
rect 6086 2360 6092 2372
rect 4249 2332 6092 2360
rect 4249 2329 4261 2332
rect 4203 2323 4261 2329
rect 6086 2320 6092 2332
rect 6144 2320 6150 2372
rect 6733 2363 6791 2369
rect 6733 2360 6745 2363
rect 6196 2332 6745 2360
rect 4522 2252 4528 2304
rect 4580 2292 4586 2304
rect 4893 2295 4951 2301
rect 4893 2292 4905 2295
rect 4580 2264 4905 2292
rect 4580 2252 4586 2264
rect 4893 2261 4905 2264
rect 4939 2261 4951 2295
rect 4893 2255 4951 2261
rect 4982 2252 4988 2304
rect 5040 2292 5046 2304
rect 6196 2292 6224 2332
rect 6733 2329 6745 2332
rect 6779 2360 6791 2363
rect 9646 2360 9674 2400
rect 6779 2332 9674 2360
rect 6779 2329 6791 2332
rect 6733 2323 6791 2329
rect 6362 2292 6368 2304
rect 5040 2264 6224 2292
rect 6323 2264 6368 2292
rect 5040 2252 5046 2264
rect 6362 2252 6368 2264
rect 6420 2252 6426 2304
rect 7055 2295 7113 2301
rect 7055 2261 7067 2295
rect 7101 2292 7113 2295
rect 7282 2292 7288 2304
rect 7101 2264 7288 2292
rect 7101 2261 7113 2264
rect 7055 2255 7113 2261
rect 7282 2252 7288 2264
rect 7340 2252 7346 2304
rect 15194 2292 15200 2304
rect 15155 2264 15200 2292
rect 15194 2252 15200 2264
rect 15252 2292 15258 2304
rect 15304 2292 15332 2400
rect 15565 2397 15577 2400
rect 15611 2397 15623 2431
rect 15565 2391 15623 2397
rect 15654 2388 15660 2440
rect 15712 2428 15718 2440
rect 15841 2431 15899 2437
rect 15841 2428 15853 2431
rect 15712 2400 15853 2428
rect 15712 2388 15718 2400
rect 15841 2397 15853 2400
rect 15887 2428 15899 2431
rect 15930 2428 15936 2440
rect 15887 2400 15936 2428
rect 15887 2397 15899 2400
rect 15841 2391 15899 2397
rect 15930 2388 15936 2400
rect 15988 2388 15994 2440
rect 17696 2428 17724 2459
rect 20070 2428 20076 2440
rect 17696 2400 20076 2428
rect 20070 2388 20076 2400
rect 20128 2388 20134 2440
rect 17313 2363 17371 2369
rect 17313 2329 17325 2363
rect 17359 2360 17371 2363
rect 21450 2360 21456 2372
rect 17359 2332 21456 2360
rect 17359 2329 17371 2332
rect 17313 2323 17371 2329
rect 21450 2320 21456 2332
rect 21508 2320 21514 2372
rect 15252 2264 15332 2292
rect 15252 2252 15258 2264
rect 1104 2202 20884 2224
rect 1104 2150 4648 2202
rect 4700 2150 4712 2202
rect 4764 2150 4776 2202
rect 4828 2150 4840 2202
rect 4892 2150 11982 2202
rect 12034 2150 12046 2202
rect 12098 2150 12110 2202
rect 12162 2150 12174 2202
rect 12226 2150 19315 2202
rect 19367 2150 19379 2202
rect 19431 2150 19443 2202
rect 19495 2150 19507 2202
rect 19559 2150 20884 2202
rect 1104 2128 20884 2150
rect 9766 76 9772 128
rect 9824 116 9830 128
rect 10502 116 10508 128
rect 9824 88 10508 116
rect 9824 76 9830 88
rect 10502 76 10508 88
rect 10560 76 10566 128
<< via1 >>
rect 4648 19558 4700 19610
rect 4712 19558 4764 19610
rect 4776 19558 4828 19610
rect 4840 19558 4892 19610
rect 11982 19558 12034 19610
rect 12046 19558 12098 19610
rect 12110 19558 12162 19610
rect 12174 19558 12226 19610
rect 19315 19558 19367 19610
rect 19379 19558 19431 19610
rect 19443 19558 19495 19610
rect 19507 19558 19559 19610
rect 4252 19456 4304 19508
rect 6736 19388 6788 19440
rect 4160 19363 4212 19372
rect 4160 19329 4169 19363
rect 4169 19329 4203 19363
rect 4203 19329 4212 19363
rect 4160 19320 4212 19329
rect 5448 19320 5500 19372
rect 7012 19320 7064 19372
rect 2136 19295 2188 19304
rect 2136 19261 2145 19295
rect 2145 19261 2179 19295
rect 2179 19261 2188 19295
rect 2136 19252 2188 19261
rect 4068 19295 4120 19304
rect 4068 19261 4077 19295
rect 4077 19261 4111 19295
rect 4111 19261 4120 19295
rect 4068 19252 4120 19261
rect 4344 19295 4396 19304
rect 2320 19184 2372 19236
rect 4344 19261 4353 19295
rect 4353 19261 4387 19295
rect 4387 19261 4396 19295
rect 4344 19252 4396 19261
rect 4988 19252 5040 19304
rect 5540 19252 5592 19304
rect 6460 19252 6512 19304
rect 7288 19252 7340 19304
rect 10324 19252 10376 19304
rect 2596 19116 2648 19168
rect 2872 19116 2924 19168
rect 3424 19159 3476 19168
rect 3424 19125 3433 19159
rect 3433 19125 3467 19159
rect 3467 19125 3476 19159
rect 3424 19116 3476 19125
rect 4068 19116 4120 19168
rect 6184 19184 6236 19236
rect 5172 19116 5224 19168
rect 6460 19116 6512 19168
rect 7104 19184 7156 19236
rect 11704 19252 11756 19304
rect 13268 19252 13320 19304
rect 11244 19227 11296 19236
rect 11244 19193 11253 19227
rect 11253 19193 11287 19227
rect 11287 19193 11296 19227
rect 11244 19184 11296 19193
rect 8944 19116 8996 19168
rect 9496 19116 9548 19168
rect 8315 19014 8367 19066
rect 8379 19014 8431 19066
rect 8443 19014 8495 19066
rect 8507 19014 8559 19066
rect 15648 19014 15700 19066
rect 15712 19014 15764 19066
rect 15776 19014 15828 19066
rect 15840 19014 15892 19066
rect 5816 18912 5868 18964
rect 11244 18912 11296 18964
rect 19064 18912 19116 18964
rect 5356 18844 5408 18896
rect 2320 18776 2372 18828
rect 4344 18819 4396 18828
rect 1400 18751 1452 18760
rect 1400 18717 1409 18751
rect 1409 18717 1443 18751
rect 1443 18717 1452 18751
rect 1400 18708 1452 18717
rect 3148 18751 3200 18760
rect 3148 18717 3157 18751
rect 3157 18717 3191 18751
rect 3191 18717 3200 18751
rect 3148 18708 3200 18717
rect 4344 18785 4353 18819
rect 4353 18785 4387 18819
rect 4387 18785 4396 18819
rect 4344 18776 4396 18785
rect 5632 18819 5684 18828
rect 5632 18785 5641 18819
rect 5641 18785 5675 18819
rect 5675 18785 5684 18819
rect 5632 18776 5684 18785
rect 6644 18776 6696 18828
rect 7472 18819 7524 18828
rect 7472 18785 7481 18819
rect 7481 18785 7515 18819
rect 7515 18785 7524 18819
rect 7472 18776 7524 18785
rect 11152 18776 11204 18828
rect 11520 18776 11572 18828
rect 12808 18776 12860 18828
rect 13728 18819 13780 18828
rect 13728 18785 13737 18819
rect 13737 18785 13771 18819
rect 13771 18785 13780 18819
rect 13728 18776 13780 18785
rect 5080 18708 5132 18760
rect 5448 18708 5500 18760
rect 6000 18708 6052 18760
rect 6276 18751 6328 18760
rect 6276 18717 6285 18751
rect 6285 18717 6319 18751
rect 6319 18717 6328 18751
rect 6276 18708 6328 18717
rect 6828 18708 6880 18760
rect 9404 18708 9456 18760
rect 4252 18640 4304 18692
rect 7380 18640 7432 18692
rect 10600 18640 10652 18692
rect 1860 18615 1912 18624
rect 1860 18581 1869 18615
rect 1869 18581 1903 18615
rect 1903 18581 1912 18615
rect 1860 18572 1912 18581
rect 7196 18572 7248 18624
rect 8208 18615 8260 18624
rect 8208 18581 8217 18615
rect 8217 18581 8251 18615
rect 8251 18581 8260 18615
rect 8208 18572 8260 18581
rect 9128 18572 9180 18624
rect 12624 18572 12676 18624
rect 4648 18470 4700 18522
rect 4712 18470 4764 18522
rect 4776 18470 4828 18522
rect 4840 18470 4892 18522
rect 11982 18470 12034 18522
rect 12046 18470 12098 18522
rect 12110 18470 12162 18522
rect 12174 18470 12226 18522
rect 19315 18470 19367 18522
rect 19379 18470 19431 18522
rect 19443 18470 19495 18522
rect 19507 18470 19559 18522
rect 1584 18411 1636 18420
rect 1584 18377 1593 18411
rect 1593 18377 1627 18411
rect 1627 18377 1636 18411
rect 1584 18368 1636 18377
rect 3148 18368 3200 18420
rect 5356 18411 5408 18420
rect 5356 18377 5365 18411
rect 5365 18377 5399 18411
rect 5399 18377 5408 18411
rect 5356 18368 5408 18377
rect 5632 18411 5684 18420
rect 5632 18377 5641 18411
rect 5641 18377 5675 18411
rect 5675 18377 5684 18411
rect 5632 18368 5684 18377
rect 6000 18411 6052 18420
rect 6000 18377 6009 18411
rect 6009 18377 6043 18411
rect 6043 18377 6052 18411
rect 6000 18368 6052 18377
rect 6644 18411 6696 18420
rect 6644 18377 6653 18411
rect 6653 18377 6687 18411
rect 6687 18377 6696 18411
rect 6644 18368 6696 18377
rect 7380 18411 7432 18420
rect 7380 18377 7389 18411
rect 7389 18377 7423 18411
rect 7423 18377 7432 18411
rect 7380 18368 7432 18377
rect 7472 18368 7524 18420
rect 19708 18368 19760 18420
rect 2044 18300 2096 18352
rect 2688 18300 2740 18352
rect 4712 18343 4764 18352
rect 4712 18309 4721 18343
rect 4721 18309 4755 18343
rect 4755 18309 4764 18343
rect 4712 18300 4764 18309
rect 7564 18300 7616 18352
rect 112 18232 164 18284
rect 11152 18232 11204 18284
rect 13084 18232 13136 18284
rect 1492 18164 1544 18216
rect 2872 18207 2924 18216
rect 2872 18173 2881 18207
rect 2881 18173 2915 18207
rect 2915 18173 2924 18207
rect 2872 18164 2924 18173
rect 3608 18164 3660 18216
rect 4068 18164 4120 18216
rect 4712 18164 4764 18216
rect 4252 18096 4304 18148
rect 5632 18164 5684 18216
rect 7932 18207 7984 18216
rect 7932 18173 7941 18207
rect 7941 18173 7975 18207
rect 7975 18173 7984 18207
rect 7932 18164 7984 18173
rect 8208 18207 8260 18216
rect 8208 18173 8217 18207
rect 8217 18173 8251 18207
rect 8251 18173 8260 18207
rect 8208 18164 8260 18173
rect 10508 18164 10560 18216
rect 10692 18164 10744 18216
rect 13728 18232 13780 18284
rect 2320 18028 2372 18080
rect 9680 18096 9732 18148
rect 6920 18071 6972 18080
rect 6920 18037 6929 18071
rect 6929 18037 6963 18071
rect 6963 18037 6972 18071
rect 6920 18028 6972 18037
rect 9864 18028 9916 18080
rect 12808 18096 12860 18148
rect 13728 18096 13780 18148
rect 14556 18207 14608 18216
rect 14556 18173 14574 18207
rect 14574 18173 14608 18207
rect 14556 18164 14608 18173
rect 14740 18164 14792 18216
rect 18420 18164 18472 18216
rect 14372 18096 14424 18148
rect 10876 18028 10928 18080
rect 11520 18028 11572 18080
rect 12440 18028 12492 18080
rect 12716 18028 12768 18080
rect 14188 18028 14240 18080
rect 16764 18028 16816 18080
rect 8315 17926 8367 17978
rect 8379 17926 8431 17978
rect 8443 17926 8495 17978
rect 8507 17926 8559 17978
rect 15648 17926 15700 17978
rect 15712 17926 15764 17978
rect 15776 17926 15828 17978
rect 15840 17926 15892 17978
rect 4344 17824 4396 17876
rect 6000 17824 6052 17876
rect 12532 17824 12584 17876
rect 1308 17756 1360 17808
rect 1860 17688 1912 17740
rect 2412 17731 2464 17740
rect 2412 17697 2421 17731
rect 2421 17697 2455 17731
rect 2455 17697 2464 17731
rect 2412 17688 2464 17697
rect 4252 17756 4304 17808
rect 10416 17756 10468 17808
rect 2320 17620 2372 17672
rect 3976 17688 4028 17740
rect 4988 17688 5040 17740
rect 5632 17731 5684 17740
rect 5632 17697 5641 17731
rect 5641 17697 5675 17731
rect 5675 17697 5684 17731
rect 5632 17688 5684 17697
rect 5908 17731 5960 17740
rect 5908 17697 5917 17731
rect 5917 17697 5951 17731
rect 5951 17697 5960 17731
rect 5908 17688 5960 17697
rect 7656 17688 7708 17740
rect 8208 17688 8260 17740
rect 9312 17688 9364 17740
rect 10140 17731 10192 17740
rect 10140 17697 10149 17731
rect 10149 17697 10183 17731
rect 10183 17697 10192 17731
rect 10140 17688 10192 17697
rect 11520 17688 11572 17740
rect 12992 17688 13044 17740
rect 14096 17688 14148 17740
rect 15476 17688 15528 17740
rect 17224 17688 17276 17740
rect 4436 17620 4488 17672
rect 6736 17620 6788 17672
rect 10048 17620 10100 17672
rect 1492 17552 1544 17604
rect 4068 17552 4120 17604
rect 7104 17552 7156 17604
rect 7564 17552 7616 17604
rect 9036 17552 9088 17604
rect 3884 17484 3936 17536
rect 7196 17527 7248 17536
rect 7196 17493 7205 17527
rect 7205 17493 7239 17527
rect 7239 17493 7248 17527
rect 7196 17484 7248 17493
rect 10692 17484 10744 17536
rect 11060 17484 11112 17536
rect 13820 17484 13872 17536
rect 14188 17484 14240 17536
rect 16120 17484 16172 17536
rect 4648 17382 4700 17434
rect 4712 17382 4764 17434
rect 4776 17382 4828 17434
rect 4840 17382 4892 17434
rect 11982 17382 12034 17434
rect 12046 17382 12098 17434
rect 12110 17382 12162 17434
rect 12174 17382 12226 17434
rect 19315 17382 19367 17434
rect 19379 17382 19431 17434
rect 19443 17382 19495 17434
rect 19507 17382 19559 17434
rect 1584 17323 1636 17332
rect 1584 17289 1593 17323
rect 1593 17289 1627 17323
rect 1627 17289 1636 17323
rect 1584 17280 1636 17289
rect 6368 17280 6420 17332
rect 12716 17280 12768 17332
rect 3976 17144 4028 17196
rect 2780 17119 2832 17128
rect 2780 17085 2789 17119
rect 2789 17085 2823 17119
rect 2823 17085 2832 17119
rect 2780 17076 2832 17085
rect 5632 17212 5684 17264
rect 6828 17212 6880 17264
rect 5080 17187 5132 17196
rect 5080 17153 5089 17187
rect 5089 17153 5123 17187
rect 5123 17153 5132 17187
rect 5080 17144 5132 17153
rect 3240 17051 3292 17060
rect 3240 17017 3249 17051
rect 3249 17017 3283 17051
rect 3283 17017 3292 17051
rect 3240 17008 3292 17017
rect 5264 17076 5316 17128
rect 5724 17076 5776 17128
rect 6828 17076 6880 17128
rect 7196 17076 7248 17128
rect 9772 17144 9824 17196
rect 10692 17212 10744 17264
rect 10232 17144 10284 17196
rect 5908 17008 5960 17060
rect 7656 17008 7708 17060
rect 8208 17051 8260 17060
rect 8208 17017 8217 17051
rect 8217 17017 8251 17051
rect 8251 17017 8260 17051
rect 8208 17008 8260 17017
rect 8852 17008 8904 17060
rect 2320 16983 2372 16992
rect 2320 16949 2329 16983
rect 2329 16949 2363 16983
rect 2363 16949 2372 16983
rect 2320 16940 2372 16949
rect 3332 16940 3384 16992
rect 3976 16940 4028 16992
rect 6092 16940 6144 16992
rect 7380 16983 7432 16992
rect 7380 16949 7389 16983
rect 7389 16949 7423 16983
rect 7423 16949 7432 16983
rect 7380 16940 7432 16949
rect 8760 16983 8812 16992
rect 8760 16949 8769 16983
rect 8769 16949 8803 16983
rect 8803 16949 8812 16983
rect 10140 17076 10192 17128
rect 11336 17144 11388 17196
rect 12992 17144 13044 17196
rect 13912 17280 13964 17332
rect 14096 17280 14148 17332
rect 17224 17323 17276 17332
rect 17224 17289 17233 17323
rect 17233 17289 17267 17323
rect 17267 17289 17276 17323
rect 17224 17280 17276 17289
rect 18788 17280 18840 17332
rect 15476 17212 15528 17264
rect 13636 17144 13688 17196
rect 10416 17051 10468 17060
rect 10416 17017 10425 17051
rect 10425 17017 10459 17051
rect 10459 17017 10468 17051
rect 12256 17076 12308 17128
rect 10416 17008 10468 17017
rect 9220 16983 9272 16992
rect 8760 16940 8812 16949
rect 9220 16949 9229 16983
rect 9229 16949 9263 16983
rect 9263 16949 9272 16983
rect 9220 16940 9272 16949
rect 10784 16983 10836 16992
rect 10784 16949 10793 16983
rect 10793 16949 10827 16983
rect 10827 16949 10836 16983
rect 10784 16940 10836 16949
rect 11520 16983 11572 16992
rect 11520 16949 11529 16983
rect 11529 16949 11563 16983
rect 11563 16949 11572 16983
rect 11520 16940 11572 16949
rect 12348 16940 12400 16992
rect 12532 16983 12584 16992
rect 12532 16949 12541 16983
rect 12541 16949 12575 16983
rect 12575 16949 12584 16983
rect 12532 16940 12584 16949
rect 12808 16940 12860 16992
rect 14096 17008 14148 17060
rect 14004 16940 14056 16992
rect 16028 17008 16080 17060
rect 18328 17008 18380 17060
rect 15384 16940 15436 16992
rect 8315 16838 8367 16890
rect 8379 16838 8431 16890
rect 8443 16838 8495 16890
rect 8507 16838 8559 16890
rect 15648 16838 15700 16890
rect 15712 16838 15764 16890
rect 15776 16838 15828 16890
rect 15840 16838 15892 16890
rect 1860 16736 1912 16788
rect 2228 16711 2280 16720
rect 2228 16677 2237 16711
rect 2237 16677 2271 16711
rect 2271 16677 2280 16711
rect 2228 16668 2280 16677
rect 6552 16736 6604 16788
rect 7564 16736 7616 16788
rect 9312 16736 9364 16788
rect 9588 16736 9640 16788
rect 10232 16736 10284 16788
rect 6920 16668 6972 16720
rect 7748 16668 7800 16720
rect 16212 16736 16264 16788
rect 12256 16668 12308 16720
rect 4988 16643 5040 16652
rect 4988 16609 4997 16643
rect 4997 16609 5031 16643
rect 5031 16609 5040 16643
rect 4988 16600 5040 16609
rect 5264 16643 5316 16652
rect 5264 16609 5273 16643
rect 5273 16609 5307 16643
rect 5307 16609 5316 16643
rect 5264 16600 5316 16609
rect 5632 16600 5684 16652
rect 8024 16600 8076 16652
rect 8116 16600 8168 16652
rect 9956 16600 10008 16652
rect 10140 16643 10192 16652
rect 10140 16609 10149 16643
rect 10149 16609 10183 16643
rect 10183 16609 10192 16643
rect 10140 16600 10192 16609
rect 11428 16600 11480 16652
rect 12716 16643 12768 16652
rect 12716 16609 12725 16643
rect 12725 16609 12759 16643
rect 12759 16609 12768 16643
rect 12716 16600 12768 16609
rect 13176 16643 13228 16652
rect 13176 16609 13185 16643
rect 13185 16609 13219 16643
rect 13219 16609 13228 16643
rect 13176 16600 13228 16609
rect 13360 16668 13412 16720
rect 3056 16532 3108 16584
rect 5448 16575 5500 16584
rect 5448 16541 5457 16575
rect 5457 16541 5491 16575
rect 5491 16541 5500 16575
rect 5448 16532 5500 16541
rect 6828 16575 6880 16584
rect 6828 16541 6837 16575
rect 6837 16541 6871 16575
rect 6871 16541 6880 16575
rect 6828 16532 6880 16541
rect 10232 16575 10284 16584
rect 10232 16541 10241 16575
rect 10241 16541 10275 16575
rect 10275 16541 10284 16575
rect 10232 16532 10284 16541
rect 13544 16532 13596 16584
rect 15476 16600 15528 16652
rect 16304 16643 16356 16652
rect 16304 16609 16313 16643
rect 16313 16609 16347 16643
rect 16347 16609 16356 16643
rect 16304 16600 16356 16609
rect 17316 16643 17368 16652
rect 17316 16609 17325 16643
rect 17325 16609 17359 16643
rect 17359 16609 17368 16643
rect 17316 16600 17368 16609
rect 18512 16600 18564 16652
rect 18236 16532 18288 16584
rect 2780 16464 2832 16516
rect 3148 16464 3200 16516
rect 6092 16464 6144 16516
rect 16028 16464 16080 16516
rect 2412 16396 2464 16448
rect 3608 16396 3660 16448
rect 9772 16396 9824 16448
rect 14280 16439 14332 16448
rect 14280 16405 14289 16439
rect 14289 16405 14323 16439
rect 14323 16405 14332 16439
rect 14280 16396 14332 16405
rect 15108 16396 15160 16448
rect 15936 16396 15988 16448
rect 17132 16396 17184 16448
rect 4648 16294 4700 16346
rect 4712 16294 4764 16346
rect 4776 16294 4828 16346
rect 4840 16294 4892 16346
rect 11982 16294 12034 16346
rect 12046 16294 12098 16346
rect 12110 16294 12162 16346
rect 12174 16294 12226 16346
rect 19315 16294 19367 16346
rect 19379 16294 19431 16346
rect 19443 16294 19495 16346
rect 19507 16294 19559 16346
rect 5264 16192 5316 16244
rect 6920 16192 6972 16244
rect 9956 16192 10008 16244
rect 12716 16192 12768 16244
rect 13912 16192 13964 16244
rect 16304 16235 16356 16244
rect 16304 16201 16313 16235
rect 16313 16201 16347 16235
rect 16347 16201 16356 16235
rect 16304 16192 16356 16201
rect 1400 15920 1452 15972
rect 9680 16124 9732 16176
rect 13636 16124 13688 16176
rect 14096 16167 14148 16176
rect 14096 16133 14105 16167
rect 14105 16133 14139 16167
rect 14139 16133 14148 16167
rect 17408 16192 17460 16244
rect 17960 16192 18012 16244
rect 14096 16124 14148 16133
rect 1860 16056 1912 16108
rect 2228 16056 2280 16108
rect 6828 16099 6880 16108
rect 6828 16065 6837 16099
rect 6837 16065 6871 16099
rect 6871 16065 6880 16099
rect 6828 16056 6880 16065
rect 4436 16031 4488 16040
rect 4436 15997 4445 16031
rect 4445 15997 4479 16031
rect 4479 15997 4488 16031
rect 4436 15988 4488 15997
rect 5264 15988 5316 16040
rect 8208 15988 8260 16040
rect 14648 16056 14700 16108
rect 6460 15920 6512 15972
rect 7104 15852 7156 15904
rect 7748 15895 7800 15904
rect 7748 15861 7757 15895
rect 7757 15861 7791 15895
rect 7791 15861 7800 15895
rect 7748 15852 7800 15861
rect 8116 15852 8168 15904
rect 8760 15920 8812 15972
rect 9312 15963 9364 15972
rect 9312 15929 9321 15963
rect 9321 15929 9355 15963
rect 9355 15929 9364 15963
rect 9312 15920 9364 15929
rect 9956 15920 10008 15972
rect 10324 15963 10376 15972
rect 10324 15929 10333 15963
rect 10333 15929 10367 15963
rect 10367 15929 10376 15963
rect 10324 15920 10376 15929
rect 10508 15920 10560 15972
rect 12164 15920 12216 15972
rect 13176 15988 13228 16040
rect 14280 16031 14332 16040
rect 14280 15997 14289 16031
rect 14289 15997 14323 16031
rect 14323 15997 14332 16031
rect 14280 15988 14332 15997
rect 17040 16124 17092 16176
rect 15476 16056 15528 16108
rect 16304 16056 16356 16108
rect 16580 16056 16632 16108
rect 16028 15988 16080 16040
rect 17960 16031 18012 16040
rect 13452 15920 13504 15972
rect 14924 15920 14976 15972
rect 16212 15920 16264 15972
rect 17960 15997 17969 16031
rect 17969 15997 18003 16031
rect 18003 15997 18012 16031
rect 17960 15988 18012 15997
rect 19156 16031 19208 16040
rect 19156 15997 19174 16031
rect 19174 15997 19208 16031
rect 19156 15988 19208 15997
rect 18972 15920 19024 15972
rect 12348 15852 12400 15904
rect 16396 15852 16448 15904
rect 17316 15852 17368 15904
rect 18512 15895 18564 15904
rect 18512 15861 18521 15895
rect 18521 15861 18555 15895
rect 18555 15861 18564 15895
rect 18512 15852 18564 15861
rect 8315 15750 8367 15802
rect 8379 15750 8431 15802
rect 8443 15750 8495 15802
rect 8507 15750 8559 15802
rect 15648 15750 15700 15802
rect 15712 15750 15764 15802
rect 15776 15750 15828 15802
rect 15840 15750 15892 15802
rect 1676 15648 1728 15700
rect 2228 15648 2280 15700
rect 4252 15691 4304 15700
rect 4252 15657 4261 15691
rect 4261 15657 4295 15691
rect 4295 15657 4304 15691
rect 4252 15648 4304 15657
rect 4988 15648 5040 15700
rect 5264 15691 5316 15700
rect 5264 15657 5273 15691
rect 5273 15657 5307 15691
rect 5307 15657 5316 15691
rect 5264 15648 5316 15657
rect 7748 15648 7800 15700
rect 8208 15648 8260 15700
rect 10324 15648 10376 15700
rect 2596 15623 2648 15632
rect 2596 15589 2605 15623
rect 2605 15589 2639 15623
rect 2639 15589 2648 15623
rect 2596 15580 2648 15589
rect 7104 15580 7156 15632
rect 7472 15623 7524 15632
rect 7472 15589 7481 15623
rect 7481 15589 7515 15623
rect 7515 15589 7524 15623
rect 7472 15580 7524 15589
rect 8024 15623 8076 15632
rect 8024 15589 8033 15623
rect 8033 15589 8067 15623
rect 8067 15589 8076 15623
rect 8024 15580 8076 15589
rect 9772 15580 9824 15632
rect 3976 15512 4028 15564
rect 5448 15512 5500 15564
rect 9312 15512 9364 15564
rect 2872 15444 2924 15496
rect 3424 15444 3476 15496
rect 7564 15444 7616 15496
rect 8024 15444 8076 15496
rect 11428 15648 11480 15700
rect 12716 15648 12768 15700
rect 18052 15648 18104 15700
rect 19616 15648 19668 15700
rect 11612 15623 11664 15632
rect 11612 15589 11621 15623
rect 11621 15589 11655 15623
rect 11655 15589 11664 15623
rect 11612 15580 11664 15589
rect 13268 15580 13320 15632
rect 15476 15623 15528 15632
rect 13452 15555 13504 15564
rect 13452 15521 13461 15555
rect 13461 15521 13495 15555
rect 13495 15521 13504 15555
rect 13452 15512 13504 15521
rect 15476 15589 15485 15623
rect 15485 15589 15519 15623
rect 15519 15589 15528 15623
rect 15476 15580 15528 15589
rect 16028 15623 16080 15632
rect 16028 15589 16037 15623
rect 16037 15589 16071 15623
rect 16071 15589 16080 15623
rect 16028 15580 16080 15589
rect 17316 15512 17368 15564
rect 17776 15512 17828 15564
rect 18604 15512 18656 15564
rect 11796 15444 11848 15496
rect 12164 15487 12216 15496
rect 12164 15453 12173 15487
rect 12173 15453 12207 15487
rect 12207 15453 12216 15487
rect 12164 15444 12216 15453
rect 12992 15444 13044 15496
rect 15384 15487 15436 15496
rect 15384 15453 15393 15487
rect 15393 15453 15427 15487
rect 15427 15453 15436 15487
rect 15384 15444 15436 15453
rect 3792 15376 3844 15428
rect 5264 15376 5316 15428
rect 6092 15376 6144 15428
rect 12624 15376 12676 15428
rect 13636 15376 13688 15428
rect 2964 15351 3016 15360
rect 2964 15317 2973 15351
rect 2973 15317 3007 15351
rect 3007 15317 3016 15351
rect 2964 15308 3016 15317
rect 6460 15351 6512 15360
rect 6460 15317 6469 15351
rect 6469 15317 6503 15351
rect 6503 15317 6512 15351
rect 6460 15308 6512 15317
rect 9956 15308 10008 15360
rect 12348 15308 12400 15360
rect 16488 15308 16540 15360
rect 4648 15206 4700 15258
rect 4712 15206 4764 15258
rect 4776 15206 4828 15258
rect 4840 15206 4892 15258
rect 11982 15206 12034 15258
rect 12046 15206 12098 15258
rect 12110 15206 12162 15258
rect 12174 15206 12226 15258
rect 19315 15206 19367 15258
rect 19379 15206 19431 15258
rect 19443 15206 19495 15258
rect 19507 15206 19559 15258
rect 5908 15104 5960 15156
rect 6460 15104 6512 15156
rect 7472 15104 7524 15156
rect 9312 15104 9364 15156
rect 9772 15147 9824 15156
rect 9772 15113 9781 15147
rect 9781 15113 9815 15147
rect 9815 15113 9824 15147
rect 9772 15104 9824 15113
rect 11612 15104 11664 15156
rect 15384 15104 15436 15156
rect 15476 15104 15528 15156
rect 17316 15147 17368 15156
rect 17316 15113 17325 15147
rect 17325 15113 17359 15147
rect 17359 15113 17368 15147
rect 17316 15104 17368 15113
rect 17776 15147 17828 15156
rect 17776 15113 17785 15147
rect 17785 15113 17819 15147
rect 17819 15113 17828 15147
rect 17776 15104 17828 15113
rect 3056 15079 3108 15088
rect 3056 15045 3065 15079
rect 3065 15045 3099 15079
rect 3099 15045 3108 15079
rect 3056 15036 3108 15045
rect 3424 15079 3476 15088
rect 3424 15045 3433 15079
rect 3433 15045 3467 15079
rect 3467 15045 3476 15079
rect 3424 15036 3476 15045
rect 2964 14968 3016 15020
rect 3516 14900 3568 14952
rect 11152 15036 11204 15088
rect 12624 15036 12676 15088
rect 8024 14968 8076 15020
rect 10232 14968 10284 15020
rect 10416 14968 10468 15020
rect 11244 14968 11296 15020
rect 7564 14900 7616 14952
rect 2596 14875 2648 14884
rect 2596 14841 2605 14875
rect 2605 14841 2639 14875
rect 2639 14841 2648 14875
rect 2596 14832 2648 14841
rect 1676 14764 1728 14816
rect 3700 14764 3752 14816
rect 3976 14764 4028 14816
rect 5264 14875 5316 14884
rect 5264 14841 5273 14875
rect 5273 14841 5307 14875
rect 5307 14841 5316 14875
rect 5264 14832 5316 14841
rect 5632 14832 5684 14884
rect 7104 14832 7156 14884
rect 7196 14832 7248 14884
rect 7012 14764 7064 14816
rect 8024 14832 8076 14884
rect 11704 14900 11756 14952
rect 13544 15011 13596 15020
rect 13544 14977 13553 15011
rect 13553 14977 13587 15011
rect 13587 14977 13596 15011
rect 13544 14968 13596 14977
rect 15476 14968 15528 15020
rect 16028 15011 16080 15020
rect 16028 14977 16037 15011
rect 16037 14977 16071 15011
rect 16071 14977 16080 15011
rect 16028 14968 16080 14977
rect 17316 14968 17368 15020
rect 18696 14968 18748 15020
rect 15200 14900 15252 14952
rect 16764 14943 16816 14952
rect 16764 14909 16773 14943
rect 16773 14909 16807 14943
rect 16807 14909 16816 14943
rect 16764 14900 16816 14909
rect 8208 14764 8260 14816
rect 9496 14764 9548 14816
rect 9772 14764 9824 14816
rect 10140 14764 10192 14816
rect 11796 14807 11848 14816
rect 11796 14773 11805 14807
rect 11805 14773 11839 14807
rect 11839 14773 11848 14807
rect 11796 14764 11848 14773
rect 11888 14764 11940 14816
rect 12900 14764 12952 14816
rect 13268 14764 13320 14816
rect 18420 14900 18472 14952
rect 16856 14764 16908 14816
rect 17592 14764 17644 14816
rect 17684 14764 17736 14816
rect 18604 14764 18656 14816
rect 8315 14662 8367 14714
rect 8379 14662 8431 14714
rect 8443 14662 8495 14714
rect 8507 14662 8559 14714
rect 15648 14662 15700 14714
rect 15712 14662 15764 14714
rect 15776 14662 15828 14714
rect 15840 14662 15892 14714
rect 1676 14603 1728 14612
rect 1676 14569 1685 14603
rect 1685 14569 1719 14603
rect 1719 14569 1728 14603
rect 1676 14560 1728 14569
rect 2964 14560 3016 14612
rect 4436 14560 4488 14612
rect 5264 14560 5316 14612
rect 5448 14560 5500 14612
rect 7012 14603 7064 14612
rect 7012 14569 7021 14603
rect 7021 14569 7055 14603
rect 7055 14569 7064 14603
rect 7012 14560 7064 14569
rect 8208 14560 8260 14612
rect 9956 14603 10008 14612
rect 9956 14569 9965 14603
rect 9965 14569 9999 14603
rect 9999 14569 10008 14603
rect 9956 14560 10008 14569
rect 10232 14560 10284 14612
rect 13544 14560 13596 14612
rect 15292 14560 15344 14612
rect 2136 14492 2188 14544
rect 3056 14492 3108 14544
rect 3332 14492 3384 14544
rect 3608 14492 3660 14544
rect 7104 14492 7156 14544
rect 8300 14492 8352 14544
rect 9496 14492 9548 14544
rect 11152 14535 11204 14544
rect 11152 14501 11161 14535
rect 11161 14501 11195 14535
rect 11195 14501 11204 14535
rect 11152 14492 11204 14501
rect 12716 14535 12768 14544
rect 12716 14501 12725 14535
rect 12725 14501 12759 14535
rect 12759 14501 12768 14535
rect 12716 14492 12768 14501
rect 12900 14492 12952 14544
rect 15384 14492 15436 14544
rect 16028 14535 16080 14544
rect 16028 14501 16037 14535
rect 16037 14501 16071 14535
rect 16071 14501 16080 14535
rect 16028 14492 16080 14501
rect 16672 14560 16724 14612
rect 5264 14424 5316 14476
rect 5632 14467 5684 14476
rect 5632 14433 5641 14467
rect 5641 14433 5675 14467
rect 5675 14433 5684 14467
rect 5632 14424 5684 14433
rect 5908 14424 5960 14476
rect 6644 14424 6696 14476
rect 7380 14424 7432 14476
rect 8208 14424 8260 14476
rect 13268 14424 13320 14476
rect 13728 14424 13780 14476
rect 14096 14467 14148 14476
rect 14096 14433 14140 14467
rect 14140 14433 14148 14467
rect 14096 14424 14148 14433
rect 17224 14424 17276 14476
rect 17408 14467 17460 14476
rect 17408 14433 17417 14467
rect 17417 14433 17451 14467
rect 17451 14433 17460 14467
rect 17408 14424 17460 14433
rect 18420 14467 18472 14476
rect 18420 14433 18429 14467
rect 18429 14433 18463 14467
rect 18463 14433 18472 14467
rect 18420 14424 18472 14433
rect 19064 14424 19116 14476
rect 19892 14424 19944 14476
rect 1676 14356 1728 14408
rect 4528 14356 4580 14408
rect 7472 14356 7524 14408
rect 9680 14356 9732 14408
rect 10048 14356 10100 14408
rect 10692 14356 10744 14408
rect 11060 14399 11112 14408
rect 11060 14365 11069 14399
rect 11069 14365 11103 14399
rect 11103 14365 11112 14399
rect 11060 14356 11112 14365
rect 11704 14399 11756 14408
rect 11704 14365 11713 14399
rect 11713 14365 11747 14399
rect 11747 14365 11756 14399
rect 11704 14356 11756 14365
rect 12992 14399 13044 14408
rect 12992 14365 13001 14399
rect 13001 14365 13035 14399
rect 13035 14365 13044 14399
rect 12992 14356 13044 14365
rect 13452 14356 13504 14408
rect 6920 14288 6972 14340
rect 7196 14288 7248 14340
rect 3056 14263 3108 14272
rect 3056 14229 3065 14263
rect 3065 14229 3099 14263
rect 3099 14229 3108 14263
rect 3056 14220 3108 14229
rect 5724 14220 5776 14272
rect 7472 14263 7524 14272
rect 7472 14229 7481 14263
rect 7481 14229 7515 14263
rect 7515 14229 7524 14263
rect 7472 14220 7524 14229
rect 10968 14220 11020 14272
rect 15016 14356 15068 14408
rect 16764 14356 16816 14408
rect 17776 14356 17828 14408
rect 15476 14220 15528 14272
rect 4648 14118 4700 14170
rect 4712 14118 4764 14170
rect 4776 14118 4828 14170
rect 4840 14118 4892 14170
rect 11982 14118 12034 14170
rect 12046 14118 12098 14170
rect 12110 14118 12162 14170
rect 12174 14118 12226 14170
rect 19315 14118 19367 14170
rect 19379 14118 19431 14170
rect 19443 14118 19495 14170
rect 19507 14118 19559 14170
rect 2136 14016 2188 14068
rect 2596 13948 2648 14000
rect 3056 13880 3108 13932
rect 3700 13948 3752 14000
rect 5264 14016 5316 14068
rect 5356 14016 5408 14068
rect 6092 14016 6144 14068
rect 6644 14059 6696 14068
rect 6644 14025 6653 14059
rect 6653 14025 6687 14059
rect 6687 14025 6696 14059
rect 6644 14016 6696 14025
rect 7472 14016 7524 14068
rect 9220 14059 9272 14068
rect 9220 14025 9229 14059
rect 9229 14025 9263 14059
rect 9263 14025 9272 14059
rect 9220 14016 9272 14025
rect 9496 14016 9548 14068
rect 9864 14016 9916 14068
rect 11060 14016 11112 14068
rect 11428 14016 11480 14068
rect 12716 14016 12768 14068
rect 14096 14059 14148 14068
rect 14096 14025 14105 14059
rect 14105 14025 14139 14059
rect 14139 14025 14148 14059
rect 14096 14016 14148 14025
rect 15200 14016 15252 14068
rect 2596 13855 2648 13864
rect 2596 13821 2605 13855
rect 2605 13821 2639 13855
rect 2639 13821 2648 13855
rect 2596 13812 2648 13821
rect 6276 13880 6328 13932
rect 3700 13812 3752 13864
rect 1768 13719 1820 13728
rect 1768 13685 1777 13719
rect 1777 13685 1811 13719
rect 1811 13685 1820 13719
rect 1768 13676 1820 13685
rect 3424 13676 3476 13728
rect 3608 13676 3660 13728
rect 5632 13812 5684 13864
rect 6644 13880 6696 13932
rect 7748 13948 7800 14000
rect 7932 13948 7984 14000
rect 8208 13991 8260 14000
rect 8208 13957 8217 13991
rect 8217 13957 8251 13991
rect 8251 13957 8260 13991
rect 8208 13948 8260 13957
rect 10140 13948 10192 14000
rect 8300 13812 8352 13864
rect 4344 13787 4396 13796
rect 4344 13753 4353 13787
rect 4353 13753 4387 13787
rect 4387 13753 4396 13787
rect 4344 13744 4396 13753
rect 7012 13787 7064 13796
rect 7012 13753 7021 13787
rect 7021 13753 7055 13787
rect 7055 13753 7064 13787
rect 7012 13744 7064 13753
rect 7196 13744 7248 13796
rect 7564 13787 7616 13796
rect 7564 13753 7573 13787
rect 7573 13753 7607 13787
rect 7607 13753 7616 13787
rect 7564 13744 7616 13753
rect 8208 13744 8260 13796
rect 9036 13744 9088 13796
rect 9864 13744 9916 13796
rect 11336 13744 11388 13796
rect 11980 13744 12032 13796
rect 15384 13948 15436 14000
rect 12532 13923 12584 13932
rect 12532 13889 12541 13923
rect 12541 13889 12575 13923
rect 12575 13889 12584 13923
rect 12532 13880 12584 13889
rect 16948 13948 17000 14000
rect 17408 13948 17460 14000
rect 16396 13880 16448 13932
rect 18604 14016 18656 14068
rect 19892 14059 19944 14068
rect 19892 14025 19901 14059
rect 19901 14025 19935 14059
rect 19935 14025 19944 14059
rect 19892 14016 19944 14025
rect 18420 13948 18472 14000
rect 18328 13880 18380 13932
rect 12900 13744 12952 13796
rect 14096 13744 14148 13796
rect 9680 13676 9732 13728
rect 11152 13676 11204 13728
rect 11612 13676 11664 13728
rect 15384 13676 15436 13728
rect 16764 13787 16816 13796
rect 16764 13753 16773 13787
rect 16773 13753 16807 13787
rect 16807 13753 16816 13787
rect 16764 13744 16816 13753
rect 16672 13676 16724 13728
rect 17040 13676 17092 13728
rect 17224 13676 17276 13728
rect 17500 13676 17552 13728
rect 18604 13676 18656 13728
rect 8315 13574 8367 13626
rect 8379 13574 8431 13626
rect 8443 13574 8495 13626
rect 8507 13574 8559 13626
rect 15648 13574 15700 13626
rect 15712 13574 15764 13626
rect 15776 13574 15828 13626
rect 15840 13574 15892 13626
rect 1676 13472 1728 13524
rect 2320 13515 2372 13524
rect 2320 13481 2329 13515
rect 2329 13481 2363 13515
rect 2363 13481 2372 13515
rect 2320 13472 2372 13481
rect 3516 13472 3568 13524
rect 3700 13515 3752 13524
rect 3700 13481 3709 13515
rect 3709 13481 3743 13515
rect 3743 13481 3752 13515
rect 3700 13472 3752 13481
rect 4528 13404 4580 13456
rect 1308 13336 1360 13388
rect 1768 13336 1820 13388
rect 2596 13379 2648 13388
rect 2596 13345 2605 13379
rect 2605 13345 2639 13379
rect 2639 13345 2648 13379
rect 2596 13336 2648 13345
rect 3792 13336 3844 13388
rect 4068 13336 4120 13388
rect 8208 13472 8260 13524
rect 10968 13515 11020 13524
rect 10968 13481 10977 13515
rect 10977 13481 11011 13515
rect 11011 13481 11020 13515
rect 10968 13472 11020 13481
rect 11152 13472 11204 13524
rect 11520 13472 11572 13524
rect 12532 13515 12584 13524
rect 12532 13481 12541 13515
rect 12541 13481 12575 13515
rect 12575 13481 12584 13515
rect 12532 13472 12584 13481
rect 13912 13472 13964 13524
rect 14372 13472 14424 13524
rect 16948 13515 17000 13524
rect 16948 13481 16957 13515
rect 16957 13481 16991 13515
rect 16991 13481 17000 13515
rect 16948 13472 17000 13481
rect 5264 13404 5316 13456
rect 6276 13404 6328 13456
rect 9864 13404 9916 13456
rect 11612 13447 11664 13456
rect 11612 13413 11621 13447
rect 11621 13413 11655 13447
rect 11655 13413 11664 13447
rect 11612 13404 11664 13413
rect 7932 13336 7984 13388
rect 9680 13379 9732 13388
rect 9680 13345 9689 13379
rect 9689 13345 9723 13379
rect 9723 13345 9732 13379
rect 9680 13336 9732 13345
rect 13728 13404 13780 13456
rect 14096 13404 14148 13456
rect 15384 13404 15436 13456
rect 13452 13379 13504 13388
rect 13452 13345 13461 13379
rect 13461 13345 13495 13379
rect 13495 13345 13504 13379
rect 13452 13336 13504 13345
rect 13912 13336 13964 13388
rect 17224 13404 17276 13456
rect 17040 13336 17092 13388
rect 18788 13472 18840 13524
rect 20168 13472 20220 13524
rect 5080 13311 5132 13320
rect 5080 13277 5089 13311
rect 5089 13277 5123 13311
rect 5123 13277 5132 13311
rect 5080 13268 5132 13277
rect 5540 13268 5592 13320
rect 11520 13311 11572 13320
rect 11520 13277 11529 13311
rect 11529 13277 11563 13311
rect 11563 13277 11572 13311
rect 11520 13268 11572 13277
rect 11888 13268 11940 13320
rect 13544 13311 13596 13320
rect 13544 13277 13553 13311
rect 13553 13277 13587 13311
rect 13587 13277 13596 13311
rect 13544 13268 13596 13277
rect 15200 13268 15252 13320
rect 15476 13268 15528 13320
rect 18236 13336 18288 13388
rect 18880 13379 18932 13388
rect 18880 13345 18889 13379
rect 18889 13345 18923 13379
rect 18923 13345 18932 13379
rect 18880 13336 18932 13345
rect 7472 13243 7524 13252
rect 7472 13209 7481 13243
rect 7481 13209 7515 13243
rect 7515 13209 7524 13243
rect 7472 13200 7524 13209
rect 11428 13200 11480 13252
rect 2596 13132 2648 13184
rect 2964 13132 3016 13184
rect 6092 13132 6144 13184
rect 10416 13132 10468 13184
rect 11796 13132 11848 13184
rect 12900 13200 12952 13252
rect 16396 13243 16448 13252
rect 16396 13209 16405 13243
rect 16405 13209 16439 13243
rect 16439 13209 16448 13243
rect 16396 13200 16448 13209
rect 18604 13200 18656 13252
rect 12808 13132 12860 13184
rect 15016 13132 15068 13184
rect 16764 13132 16816 13184
rect 4648 13030 4700 13082
rect 4712 13030 4764 13082
rect 4776 13030 4828 13082
rect 4840 13030 4892 13082
rect 11982 13030 12034 13082
rect 12046 13030 12098 13082
rect 12110 13030 12162 13082
rect 12174 13030 12226 13082
rect 19315 13030 19367 13082
rect 19379 13030 19431 13082
rect 19443 13030 19495 13082
rect 19507 13030 19559 13082
rect 2688 12928 2740 12980
rect 3792 12971 3844 12980
rect 3792 12937 3801 12971
rect 3801 12937 3835 12971
rect 3835 12937 3844 12971
rect 3792 12928 3844 12937
rect 5264 12928 5316 12980
rect 5724 12928 5776 12980
rect 6276 12971 6328 12980
rect 6276 12937 6285 12971
rect 6285 12937 6319 12971
rect 6319 12937 6328 12971
rect 6276 12928 6328 12937
rect 9680 12928 9732 12980
rect 11612 12971 11664 12980
rect 11612 12937 11621 12971
rect 11621 12937 11655 12971
rect 11655 12937 11664 12971
rect 11612 12928 11664 12937
rect 2780 12903 2832 12912
rect 2780 12869 2789 12903
rect 2789 12869 2823 12903
rect 2823 12869 2832 12903
rect 2780 12860 2832 12869
rect 7472 12903 7524 12912
rect 7472 12869 7481 12903
rect 7481 12869 7515 12903
rect 7515 12869 7524 12903
rect 7472 12860 7524 12869
rect 9588 12860 9640 12912
rect 9864 12860 9916 12912
rect 12348 12928 12400 12980
rect 13452 12971 13504 12980
rect 13452 12937 13461 12971
rect 13461 12937 13495 12971
rect 13495 12937 13504 12971
rect 13452 12928 13504 12937
rect 13728 12928 13780 12980
rect 15384 12971 15436 12980
rect 15384 12937 15393 12971
rect 15393 12937 15427 12971
rect 15427 12937 15436 12971
rect 15384 12928 15436 12937
rect 17408 12928 17460 12980
rect 6092 12792 6144 12844
rect 6920 12835 6972 12844
rect 6920 12801 6929 12835
rect 6929 12801 6963 12835
rect 6963 12801 6972 12835
rect 6920 12792 6972 12801
rect 112 12724 164 12776
rect 2320 12724 2372 12776
rect 2688 12767 2740 12776
rect 2688 12733 2697 12767
rect 2697 12733 2731 12767
rect 2731 12733 2740 12767
rect 2688 12724 2740 12733
rect 2964 12767 3016 12776
rect 2964 12733 2973 12767
rect 2973 12733 3007 12767
rect 3007 12733 3016 12767
rect 2964 12724 3016 12733
rect 7748 12724 7800 12776
rect 8208 12724 8260 12776
rect 11796 12860 11848 12912
rect 17500 12860 17552 12912
rect 10968 12792 11020 12844
rect 12808 12835 12860 12844
rect 12808 12801 12817 12835
rect 12817 12801 12851 12835
rect 12851 12801 12860 12835
rect 12808 12792 12860 12801
rect 13912 12835 13964 12844
rect 13912 12801 13921 12835
rect 13921 12801 13955 12835
rect 13955 12801 13964 12835
rect 13912 12792 13964 12801
rect 14372 12835 14424 12844
rect 14372 12801 14381 12835
rect 14381 12801 14415 12835
rect 14415 12801 14424 12835
rect 14372 12792 14424 12801
rect 15016 12835 15068 12844
rect 15016 12801 15025 12835
rect 15025 12801 15059 12835
rect 15059 12801 15068 12835
rect 15016 12792 15068 12801
rect 16396 12792 16448 12844
rect 16764 12792 16816 12844
rect 18236 12860 18288 12912
rect 2412 12656 2464 12708
rect 3148 12656 3200 12708
rect 3516 12656 3568 12708
rect 3792 12656 3844 12708
rect 5080 12656 5132 12708
rect 5908 12699 5960 12708
rect 20 12588 72 12640
rect 1952 12588 2004 12640
rect 4068 12631 4120 12640
rect 4068 12597 4077 12631
rect 4077 12597 4111 12631
rect 4111 12597 4120 12631
rect 4068 12588 4120 12597
rect 4252 12588 4304 12640
rect 5264 12588 5316 12640
rect 5908 12665 5917 12699
rect 5917 12665 5951 12699
rect 5951 12665 5960 12699
rect 5908 12656 5960 12665
rect 7012 12699 7064 12708
rect 7012 12665 7021 12699
rect 7021 12665 7055 12699
rect 7055 12665 7064 12699
rect 7012 12656 7064 12665
rect 6276 12588 6328 12640
rect 9588 12724 9640 12776
rect 11612 12724 11664 12776
rect 11888 12724 11940 12776
rect 18052 12767 18104 12776
rect 18052 12733 18061 12767
rect 18061 12733 18095 12767
rect 18095 12733 18104 12767
rect 18052 12724 18104 12733
rect 18972 12792 19024 12844
rect 18880 12724 18932 12776
rect 8668 12588 8720 12640
rect 9680 12631 9732 12640
rect 9680 12597 9689 12631
rect 9689 12597 9723 12631
rect 9723 12597 9732 12631
rect 9680 12588 9732 12597
rect 10508 12631 10560 12640
rect 10508 12597 10517 12631
rect 10517 12597 10551 12631
rect 10551 12597 10560 12631
rect 11704 12656 11756 12708
rect 12072 12656 12124 12708
rect 12532 12699 12584 12708
rect 12532 12665 12541 12699
rect 12541 12665 12575 12699
rect 12575 12665 12584 12699
rect 12532 12656 12584 12665
rect 14464 12699 14516 12708
rect 10508 12588 10560 12597
rect 11888 12588 11940 12640
rect 14464 12665 14473 12699
rect 14473 12665 14507 12699
rect 14507 12665 14516 12699
rect 14464 12656 14516 12665
rect 16028 12699 16080 12708
rect 16028 12665 16037 12699
rect 16037 12665 16071 12699
rect 16071 12665 16080 12699
rect 16028 12656 16080 12665
rect 18420 12656 18472 12708
rect 17040 12588 17092 12640
rect 17316 12631 17368 12640
rect 17316 12597 17325 12631
rect 17325 12597 17359 12631
rect 17359 12597 17368 12631
rect 17316 12588 17368 12597
rect 18144 12631 18196 12640
rect 18144 12597 18153 12631
rect 18153 12597 18187 12631
rect 18187 12597 18196 12631
rect 18144 12588 18196 12597
rect 20076 12631 20128 12640
rect 20076 12597 20085 12631
rect 20085 12597 20119 12631
rect 20119 12597 20128 12631
rect 20076 12588 20128 12597
rect 8315 12486 8367 12538
rect 8379 12486 8431 12538
rect 8443 12486 8495 12538
rect 8507 12486 8559 12538
rect 15648 12486 15700 12538
rect 15712 12486 15764 12538
rect 15776 12486 15828 12538
rect 15840 12486 15892 12538
rect 2780 12384 2832 12436
rect 3332 12384 3384 12436
rect 5264 12427 5316 12436
rect 5264 12393 5273 12427
rect 5273 12393 5307 12427
rect 5307 12393 5316 12427
rect 5264 12384 5316 12393
rect 5540 12427 5592 12436
rect 5540 12393 5549 12427
rect 5549 12393 5583 12427
rect 5583 12393 5592 12427
rect 5540 12384 5592 12393
rect 6920 12384 6972 12436
rect 7472 12384 7524 12436
rect 8208 12384 8260 12436
rect 11520 12427 11572 12436
rect 2872 12359 2924 12368
rect 2872 12325 2881 12359
rect 2881 12325 2915 12359
rect 2915 12325 2924 12359
rect 2872 12316 2924 12325
rect 1676 12291 1728 12300
rect 1676 12257 1685 12291
rect 1685 12257 1719 12291
rect 1719 12257 1728 12291
rect 1676 12248 1728 12257
rect 2136 12291 2188 12300
rect 2136 12257 2145 12291
rect 2145 12257 2179 12291
rect 2179 12257 2188 12291
rect 2136 12248 2188 12257
rect 2412 12291 2464 12300
rect 2412 12257 2421 12291
rect 2421 12257 2455 12291
rect 2455 12257 2464 12291
rect 2412 12248 2464 12257
rect 5724 12316 5776 12368
rect 6276 12316 6328 12368
rect 3516 12248 3568 12300
rect 4436 12291 4488 12300
rect 4436 12257 4445 12291
rect 4445 12257 4479 12291
rect 4479 12257 4488 12291
rect 4436 12248 4488 12257
rect 5080 12248 5132 12300
rect 7012 12316 7064 12368
rect 7840 12316 7892 12368
rect 7932 12316 7984 12368
rect 5724 12223 5776 12232
rect 5724 12189 5733 12223
rect 5733 12189 5767 12223
rect 5767 12189 5776 12223
rect 5724 12180 5776 12189
rect 8208 12180 8260 12232
rect 9680 12316 9732 12368
rect 11520 12393 11529 12427
rect 11529 12393 11563 12427
rect 11563 12393 11572 12427
rect 11520 12384 11572 12393
rect 13544 12384 13596 12436
rect 14464 12384 14516 12436
rect 15200 12384 15252 12436
rect 15292 12384 15344 12436
rect 11888 12359 11940 12368
rect 11888 12325 11897 12359
rect 11897 12325 11931 12359
rect 11931 12325 11940 12359
rect 11888 12316 11940 12325
rect 14096 12316 14148 12368
rect 16488 12384 16540 12436
rect 16580 12384 16632 12436
rect 18052 12427 18104 12436
rect 18052 12393 18061 12427
rect 18061 12393 18095 12427
rect 18095 12393 18104 12427
rect 18052 12384 18104 12393
rect 18512 12427 18564 12436
rect 18512 12393 18521 12427
rect 18521 12393 18555 12427
rect 18555 12393 18564 12427
rect 18512 12384 18564 12393
rect 16028 12316 16080 12368
rect 9956 12291 10008 12300
rect 9956 12257 9965 12291
rect 9965 12257 9999 12291
rect 9999 12257 10008 12291
rect 9956 12248 10008 12257
rect 17040 12291 17092 12300
rect 17040 12257 17049 12291
rect 17049 12257 17083 12291
rect 17083 12257 17092 12291
rect 17040 12248 17092 12257
rect 17500 12248 17552 12300
rect 18696 12248 18748 12300
rect 18880 12291 18932 12300
rect 18880 12257 18889 12291
rect 18889 12257 18923 12291
rect 18923 12257 18932 12291
rect 18880 12248 18932 12257
rect 11612 12180 11664 12232
rect 11796 12223 11848 12232
rect 11796 12189 11805 12223
rect 11805 12189 11839 12223
rect 11839 12189 11848 12223
rect 11796 12180 11848 12189
rect 12072 12223 12124 12232
rect 12072 12189 12081 12223
rect 12081 12189 12115 12223
rect 12115 12189 12124 12223
rect 12072 12180 12124 12189
rect 14556 12180 14608 12232
rect 15476 12180 15528 12232
rect 5908 12112 5960 12164
rect 12532 12112 12584 12164
rect 7012 12087 7064 12096
rect 7012 12053 7021 12087
rect 7021 12053 7055 12087
rect 7055 12053 7064 12087
rect 7012 12044 7064 12053
rect 7564 12044 7616 12096
rect 9220 12044 9272 12096
rect 12624 12044 12676 12096
rect 16028 12112 16080 12164
rect 14924 12044 14976 12096
rect 4648 11942 4700 11994
rect 4712 11942 4764 11994
rect 4776 11942 4828 11994
rect 4840 11942 4892 11994
rect 11982 11942 12034 11994
rect 12046 11942 12098 11994
rect 12110 11942 12162 11994
rect 12174 11942 12226 11994
rect 19315 11942 19367 11994
rect 19379 11942 19431 11994
rect 19443 11942 19495 11994
rect 19507 11942 19559 11994
rect 112 11840 164 11892
rect 4436 11840 4488 11892
rect 6276 11840 6328 11892
rect 7840 11883 7892 11892
rect 6092 11815 6144 11824
rect 6092 11781 6101 11815
rect 6101 11781 6135 11815
rect 6135 11781 6144 11815
rect 6092 11772 6144 11781
rect 7840 11849 7849 11883
rect 7849 11849 7883 11883
rect 7883 11849 7892 11883
rect 7840 11840 7892 11849
rect 8208 11883 8260 11892
rect 8208 11849 8217 11883
rect 8217 11849 8251 11883
rect 8251 11849 8260 11883
rect 8208 11840 8260 11849
rect 9956 11840 10008 11892
rect 11336 11840 11388 11892
rect 12348 11840 12400 11892
rect 14096 11840 14148 11892
rect 14464 11840 14516 11892
rect 16028 11883 16080 11892
rect 9680 11772 9732 11824
rect 3056 11704 3108 11756
rect 3424 11704 3476 11756
rect 4804 11704 4856 11756
rect 1676 11679 1728 11688
rect 1676 11645 1685 11679
rect 1685 11645 1719 11679
rect 1719 11645 1728 11679
rect 2136 11679 2188 11688
rect 1676 11636 1728 11645
rect 2136 11645 2145 11679
rect 2145 11645 2179 11679
rect 2179 11645 2188 11679
rect 2136 11636 2188 11645
rect 2412 11679 2464 11688
rect 2412 11645 2421 11679
rect 2421 11645 2455 11679
rect 2455 11645 2464 11679
rect 2412 11636 2464 11645
rect 2688 11679 2740 11688
rect 2688 11645 2697 11679
rect 2697 11645 2731 11679
rect 2731 11645 2740 11679
rect 2688 11636 2740 11645
rect 3332 11636 3384 11688
rect 3884 11636 3936 11688
rect 5632 11636 5684 11688
rect 6552 11704 6604 11756
rect 7104 11704 7156 11756
rect 3424 11568 3476 11620
rect 4068 11611 4120 11620
rect 4068 11577 4077 11611
rect 4077 11577 4111 11611
rect 4111 11577 4120 11611
rect 4068 11568 4120 11577
rect 4252 11568 4304 11620
rect 3700 11500 3752 11552
rect 5080 11543 5132 11552
rect 5080 11509 5089 11543
rect 5089 11509 5123 11543
rect 5123 11509 5132 11543
rect 5080 11500 5132 11509
rect 7012 11611 7064 11620
rect 7012 11577 7021 11611
rect 7021 11577 7055 11611
rect 7055 11577 7064 11611
rect 7012 11568 7064 11577
rect 6920 11500 6972 11552
rect 9496 11636 9548 11688
rect 10968 11636 11020 11688
rect 11152 11636 11204 11688
rect 11888 11772 11940 11824
rect 13544 11704 13596 11756
rect 13084 11636 13136 11688
rect 13452 11636 13504 11688
rect 14188 11636 14240 11688
rect 9680 11568 9732 11620
rect 9956 11568 10008 11620
rect 10140 11568 10192 11620
rect 13360 11568 13412 11620
rect 14096 11568 14148 11620
rect 16028 11849 16037 11883
rect 16037 11849 16071 11883
rect 16071 11849 16080 11883
rect 16028 11840 16080 11849
rect 16304 11840 16356 11892
rect 21640 11840 21692 11892
rect 14924 11772 14976 11824
rect 15108 11747 15160 11756
rect 15108 11713 15117 11747
rect 15117 11713 15151 11747
rect 15151 11713 15160 11747
rect 15108 11704 15160 11713
rect 15476 11747 15528 11756
rect 15476 11713 15485 11747
rect 15485 11713 15519 11747
rect 15519 11713 15528 11747
rect 15476 11704 15528 11713
rect 17408 11704 17460 11756
rect 17500 11679 17552 11688
rect 9036 11500 9088 11552
rect 10508 11543 10560 11552
rect 10508 11509 10517 11543
rect 10517 11509 10551 11543
rect 10551 11509 10560 11543
rect 10508 11500 10560 11509
rect 14556 11543 14608 11552
rect 14556 11509 14565 11543
rect 14565 11509 14599 11543
rect 14599 11509 14608 11543
rect 14556 11500 14608 11509
rect 14648 11500 14700 11552
rect 17040 11568 17092 11620
rect 16856 11500 16908 11552
rect 17500 11645 17509 11679
rect 17509 11645 17543 11679
rect 17543 11645 17552 11679
rect 17500 11636 17552 11645
rect 17960 11636 18012 11688
rect 17592 11568 17644 11620
rect 17224 11500 17276 11552
rect 17500 11500 17552 11552
rect 18880 11636 18932 11688
rect 19064 11679 19116 11688
rect 19064 11645 19073 11679
rect 19073 11645 19107 11679
rect 19107 11645 19116 11679
rect 19064 11636 19116 11645
rect 20076 11679 20128 11688
rect 20076 11645 20085 11679
rect 20085 11645 20119 11679
rect 20119 11645 20128 11679
rect 20076 11636 20128 11645
rect 8315 11398 8367 11450
rect 8379 11398 8431 11450
rect 8443 11398 8495 11450
rect 8507 11398 8559 11450
rect 15648 11398 15700 11450
rect 15712 11398 15764 11450
rect 15776 11398 15828 11450
rect 15840 11398 15892 11450
rect 2688 11296 2740 11348
rect 3424 11339 3476 11348
rect 3424 11305 3433 11339
rect 3433 11305 3467 11339
rect 3467 11305 3476 11339
rect 3424 11296 3476 11305
rect 3884 11339 3936 11348
rect 3884 11305 3893 11339
rect 3893 11305 3927 11339
rect 3927 11305 3936 11339
rect 3884 11296 3936 11305
rect 4068 11296 4120 11348
rect 5356 11296 5408 11348
rect 5724 11339 5776 11348
rect 5724 11305 5733 11339
rect 5733 11305 5767 11339
rect 5767 11305 5776 11339
rect 5724 11296 5776 11305
rect 6092 11296 6144 11348
rect 6276 11339 6328 11348
rect 6276 11305 6285 11339
rect 6285 11305 6319 11339
rect 6319 11305 6328 11339
rect 6276 11296 6328 11305
rect 7012 11296 7064 11348
rect 7104 11339 7156 11348
rect 7104 11305 7113 11339
rect 7113 11305 7147 11339
rect 7147 11305 7156 11339
rect 7104 11296 7156 11305
rect 8116 11296 8168 11348
rect 3516 11228 3568 11280
rect 4252 11271 4304 11280
rect 4252 11237 4261 11271
rect 4261 11237 4295 11271
rect 4295 11237 4304 11271
rect 4252 11228 4304 11237
rect 7196 11228 7248 11280
rect 10876 11296 10928 11348
rect 11796 11296 11848 11348
rect 10508 11228 10560 11280
rect 12348 11228 12400 11280
rect 14004 11296 14056 11348
rect 15108 11339 15160 11348
rect 15108 11305 15117 11339
rect 15117 11305 15151 11339
rect 15151 11305 15160 11339
rect 15108 11296 15160 11305
rect 15292 11296 15344 11348
rect 16028 11296 16080 11348
rect 18696 11339 18748 11348
rect 18696 11305 18705 11339
rect 18705 11305 18739 11339
rect 18739 11305 18748 11339
rect 18696 11296 18748 11305
rect 19708 11296 19760 11348
rect 13268 11271 13320 11280
rect 13268 11237 13277 11271
rect 13277 11237 13311 11271
rect 13311 11237 13320 11271
rect 16304 11271 16356 11280
rect 13268 11228 13320 11237
rect 16304 11237 16313 11271
rect 16313 11237 16347 11271
rect 16347 11237 16356 11271
rect 16304 11228 16356 11237
rect 17224 11228 17276 11280
rect 18604 11228 18656 11280
rect 2872 11203 2924 11212
rect 2872 11169 2881 11203
rect 2881 11169 2915 11203
rect 2915 11169 2924 11203
rect 2872 11160 2924 11169
rect 4804 11160 4856 11212
rect 7472 11160 7524 11212
rect 8208 11203 8260 11212
rect 8208 11169 8217 11203
rect 8217 11169 8251 11203
rect 8251 11169 8260 11203
rect 8208 11160 8260 11169
rect 8852 11160 8904 11212
rect 17868 11203 17920 11212
rect 17868 11169 17877 11203
rect 17877 11169 17911 11203
rect 17911 11169 17920 11203
rect 17868 11160 17920 11169
rect 17960 11160 18012 11212
rect 18236 11203 18288 11212
rect 18236 11169 18245 11203
rect 18245 11169 18279 11203
rect 18279 11169 18288 11203
rect 18236 11160 18288 11169
rect 19616 11160 19668 11212
rect 3056 11135 3108 11144
rect 3056 11101 3065 11135
rect 3065 11101 3099 11135
rect 3099 11101 3108 11135
rect 3056 11092 3108 11101
rect 4068 11024 4120 11076
rect 112 10956 164 11008
rect 3700 10956 3752 11008
rect 4344 11092 4396 11144
rect 6276 11092 6328 11144
rect 6644 11092 6696 11144
rect 10692 11092 10744 11144
rect 11336 11135 11388 11144
rect 11336 11101 11345 11135
rect 11345 11101 11379 11135
rect 11379 11101 11388 11135
rect 11336 11092 11388 11101
rect 13636 11135 13688 11144
rect 13636 11101 13645 11135
rect 13645 11101 13679 11135
rect 13679 11101 13688 11135
rect 13636 11092 13688 11101
rect 16488 11092 16540 11144
rect 4528 11024 4580 11076
rect 8668 11024 8720 11076
rect 10416 11067 10468 11076
rect 10416 11033 10425 11067
rect 10425 11033 10459 11067
rect 10459 11033 10468 11067
rect 10416 11024 10468 11033
rect 12624 11024 12676 11076
rect 13268 11024 13320 11076
rect 16764 11067 16816 11076
rect 16764 11033 16773 11067
rect 16773 11033 16807 11067
rect 16807 11033 16816 11067
rect 16764 11024 16816 11033
rect 17684 11024 17736 11076
rect 5816 10956 5868 11008
rect 7656 10956 7708 11008
rect 7840 10956 7892 11008
rect 9496 10999 9548 11008
rect 9496 10965 9505 10999
rect 9505 10965 9539 10999
rect 9539 10965 9548 10999
rect 9496 10956 9548 10965
rect 12716 10956 12768 11008
rect 18144 10956 18196 11008
rect 4648 10854 4700 10906
rect 4712 10854 4764 10906
rect 4776 10854 4828 10906
rect 4840 10854 4892 10906
rect 11982 10854 12034 10906
rect 12046 10854 12098 10906
rect 12110 10854 12162 10906
rect 12174 10854 12226 10906
rect 19315 10854 19367 10906
rect 19379 10854 19431 10906
rect 19443 10854 19495 10906
rect 19507 10854 19559 10906
rect 4252 10752 4304 10804
rect 6092 10752 6144 10804
rect 6276 10795 6328 10804
rect 6276 10761 6285 10795
rect 6285 10761 6319 10795
rect 6319 10761 6328 10795
rect 6276 10752 6328 10761
rect 7012 10752 7064 10804
rect 7472 10752 7524 10804
rect 7748 10752 7800 10804
rect 10508 10795 10560 10804
rect 10508 10761 10517 10795
rect 10517 10761 10551 10795
rect 10551 10761 10560 10795
rect 10508 10752 10560 10761
rect 10692 10752 10744 10804
rect 12348 10752 12400 10804
rect 13268 10752 13320 10804
rect 13728 10752 13780 10804
rect 16304 10752 16356 10804
rect 20168 10795 20220 10804
rect 20168 10761 20177 10795
rect 20177 10761 20211 10795
rect 20211 10761 20220 10795
rect 20168 10752 20220 10761
rect 3608 10684 3660 10736
rect 3240 10616 3292 10668
rect 2596 10480 2648 10532
rect 9404 10684 9456 10736
rect 4988 10591 5040 10600
rect 4988 10557 4997 10591
rect 4997 10557 5031 10591
rect 5031 10557 5040 10591
rect 4988 10548 5040 10557
rect 7472 10616 7524 10668
rect 7564 10616 7616 10668
rect 3792 10480 3844 10532
rect 1584 10455 1636 10464
rect 1584 10421 1593 10455
rect 1593 10421 1627 10455
rect 1627 10421 1636 10455
rect 1584 10412 1636 10421
rect 7196 10480 7248 10532
rect 9588 10523 9640 10532
rect 7012 10412 7064 10464
rect 9588 10489 9597 10523
rect 9597 10489 9631 10523
rect 9631 10489 9640 10523
rect 9588 10480 9640 10489
rect 13544 10684 13596 10736
rect 14372 10684 14424 10736
rect 18236 10684 18288 10736
rect 18512 10684 18564 10736
rect 12992 10616 13044 10668
rect 10692 10548 10744 10600
rect 10968 10548 11020 10600
rect 14096 10616 14148 10668
rect 14556 10659 14608 10668
rect 14556 10625 14565 10659
rect 14565 10625 14599 10659
rect 14599 10625 14608 10659
rect 14556 10616 14608 10625
rect 12532 10523 12584 10532
rect 8668 10412 8720 10464
rect 8760 10412 8812 10464
rect 12532 10489 12541 10523
rect 12541 10489 12575 10523
rect 12575 10489 12584 10523
rect 12532 10480 12584 10489
rect 11336 10412 11388 10464
rect 12440 10412 12492 10464
rect 13728 10480 13780 10532
rect 17316 10548 17368 10600
rect 18236 10591 18288 10600
rect 18236 10557 18245 10591
rect 18245 10557 18279 10591
rect 18279 10557 18288 10591
rect 18236 10548 18288 10557
rect 18512 10591 18564 10600
rect 18512 10557 18521 10591
rect 18521 10557 18555 10591
rect 18555 10557 18564 10591
rect 18512 10548 18564 10557
rect 20168 10548 20220 10600
rect 16304 10523 16356 10532
rect 16304 10489 16313 10523
rect 16313 10489 16347 10523
rect 16347 10489 16356 10523
rect 16304 10480 16356 10489
rect 13820 10412 13872 10464
rect 17316 10412 17368 10464
rect 17868 10412 17920 10464
rect 19616 10412 19668 10464
rect 8315 10310 8367 10362
rect 8379 10310 8431 10362
rect 8443 10310 8495 10362
rect 8507 10310 8559 10362
rect 15648 10310 15700 10362
rect 15712 10310 15764 10362
rect 15776 10310 15828 10362
rect 15840 10310 15892 10362
rect 2136 10208 2188 10260
rect 3240 10208 3292 10260
rect 4252 10251 4304 10260
rect 4252 10217 4261 10251
rect 4261 10217 4295 10251
rect 4295 10217 4304 10251
rect 4252 10208 4304 10217
rect 5816 10208 5868 10260
rect 6644 10208 6696 10260
rect 6736 10208 6788 10260
rect 9956 10208 10008 10260
rect 10232 10208 10284 10260
rect 10784 10208 10836 10260
rect 12532 10208 12584 10260
rect 2320 10140 2372 10192
rect 4528 10140 4580 10192
rect 5448 10140 5500 10192
rect 7656 10140 7708 10192
rect 11152 10140 11204 10192
rect 2596 10072 2648 10124
rect 6552 10072 6604 10124
rect 9588 10072 9640 10124
rect 1400 10004 1452 10056
rect 4620 10004 4672 10056
rect 5356 10004 5408 10056
rect 6828 10004 6880 10056
rect 7288 10047 7340 10056
rect 7288 10013 7297 10047
rect 7297 10013 7331 10047
rect 7331 10013 7340 10047
rect 7288 10004 7340 10013
rect 7564 10047 7616 10056
rect 7564 10013 7573 10047
rect 7573 10013 7607 10047
rect 7607 10013 7616 10047
rect 7564 10004 7616 10013
rect 9956 10004 10008 10056
rect 13268 10140 13320 10192
rect 14556 10140 14608 10192
rect 16304 10208 16356 10260
rect 16488 10251 16540 10260
rect 16488 10217 16497 10251
rect 16497 10217 16531 10251
rect 16531 10217 16540 10251
rect 16488 10208 16540 10217
rect 16856 10251 16908 10260
rect 16856 10217 16865 10251
rect 16865 10217 16899 10251
rect 16899 10217 16908 10251
rect 16856 10208 16908 10217
rect 17960 10208 18012 10260
rect 18696 10251 18748 10260
rect 18696 10217 18705 10251
rect 18705 10217 18739 10251
rect 18739 10217 18748 10251
rect 18696 10208 18748 10217
rect 16580 10140 16632 10192
rect 17224 10183 17276 10192
rect 17224 10149 17233 10183
rect 17233 10149 17267 10183
rect 17267 10149 17276 10183
rect 17224 10140 17276 10149
rect 18512 10140 18564 10192
rect 18972 10140 19024 10192
rect 12808 10047 12860 10056
rect 12808 10013 12817 10047
rect 12817 10013 12851 10047
rect 12851 10013 12860 10047
rect 16028 10072 16080 10124
rect 18604 10115 18656 10124
rect 18604 10081 18613 10115
rect 18613 10081 18647 10115
rect 18647 10081 18656 10115
rect 18604 10072 18656 10081
rect 15292 10047 15344 10056
rect 12808 10004 12860 10013
rect 15292 10013 15301 10047
rect 15301 10013 15335 10047
rect 15335 10013 15344 10047
rect 15292 10004 15344 10013
rect 17316 10004 17368 10056
rect 4988 9936 5040 9988
rect 3516 9868 3568 9920
rect 4068 9868 4120 9920
rect 8760 9936 8812 9988
rect 9404 9936 9456 9988
rect 13452 9936 13504 9988
rect 13636 9936 13688 9988
rect 13820 9936 13872 9988
rect 16488 9936 16540 9988
rect 18328 9936 18380 9988
rect 8208 9911 8260 9920
rect 8208 9877 8217 9911
rect 8217 9877 8251 9911
rect 8251 9877 8260 9911
rect 8208 9868 8260 9877
rect 11796 9868 11848 9920
rect 12440 9911 12492 9920
rect 12440 9877 12449 9911
rect 12449 9877 12483 9911
rect 12483 9877 12492 9911
rect 12440 9868 12492 9877
rect 13728 9911 13780 9920
rect 13728 9877 13737 9911
rect 13737 9877 13771 9911
rect 13771 9877 13780 9911
rect 13728 9868 13780 9877
rect 14096 9911 14148 9920
rect 14096 9877 14105 9911
rect 14105 9877 14139 9911
rect 14139 9877 14148 9911
rect 14096 9868 14148 9877
rect 18236 9868 18288 9920
rect 19708 9868 19760 9920
rect 4648 9766 4700 9818
rect 4712 9766 4764 9818
rect 4776 9766 4828 9818
rect 4840 9766 4892 9818
rect 11982 9766 12034 9818
rect 12046 9766 12098 9818
rect 12110 9766 12162 9818
rect 12174 9766 12226 9818
rect 19315 9766 19367 9818
rect 19379 9766 19431 9818
rect 19443 9766 19495 9818
rect 19507 9766 19559 9818
rect 2320 9707 2372 9716
rect 2320 9673 2329 9707
rect 2329 9673 2363 9707
rect 2363 9673 2372 9707
rect 2320 9664 2372 9673
rect 2872 9664 2924 9716
rect 4528 9664 4580 9716
rect 5356 9707 5408 9716
rect 5356 9673 5365 9707
rect 5365 9673 5399 9707
rect 5399 9673 5408 9707
rect 5356 9664 5408 9673
rect 8116 9664 8168 9716
rect 3792 9571 3844 9580
rect 3792 9537 3801 9571
rect 3801 9537 3835 9571
rect 3835 9537 3844 9571
rect 3792 9528 3844 9537
rect 6736 9528 6788 9580
rect 10232 9664 10284 9716
rect 9496 9571 9548 9580
rect 1584 9460 1636 9512
rect 3240 9460 3292 9512
rect 8760 9460 8812 9512
rect 9036 9503 9088 9512
rect 9036 9469 9045 9503
rect 9045 9469 9079 9503
rect 9079 9469 9088 9503
rect 9036 9460 9088 9469
rect 9496 9537 9505 9571
rect 9505 9537 9539 9571
rect 9539 9537 9548 9571
rect 9496 9528 9548 9537
rect 12440 9664 12492 9716
rect 11152 9596 11204 9648
rect 12808 9596 12860 9648
rect 1860 9324 1912 9376
rect 4436 9392 4488 9444
rect 10784 9528 10836 9580
rect 10968 9528 11020 9580
rect 14372 9664 14424 9716
rect 14556 9707 14608 9716
rect 14556 9673 14565 9707
rect 14565 9673 14599 9707
rect 14599 9673 14608 9707
rect 14556 9664 14608 9673
rect 13544 9596 13596 9648
rect 13636 9528 13688 9580
rect 11612 9460 11664 9512
rect 12440 9460 12492 9512
rect 6552 9324 6604 9376
rect 7656 9324 7708 9376
rect 11612 9324 11664 9376
rect 13176 9324 13228 9376
rect 13728 9392 13780 9444
rect 16396 9664 16448 9716
rect 17224 9664 17276 9716
rect 18972 9664 19024 9716
rect 21548 9596 21600 9648
rect 15292 9528 15344 9580
rect 17868 9528 17920 9580
rect 18604 9528 18656 9580
rect 18880 9528 18932 9580
rect 15108 9503 15160 9512
rect 15108 9469 15117 9503
rect 15117 9469 15151 9503
rect 15151 9469 15160 9503
rect 15108 9460 15160 9469
rect 16856 9503 16908 9512
rect 16856 9469 16865 9503
rect 16865 9469 16899 9503
rect 16899 9469 16908 9503
rect 17408 9503 17460 9512
rect 16856 9460 16908 9469
rect 17408 9469 17417 9503
rect 17417 9469 17451 9503
rect 17451 9469 17460 9503
rect 17408 9460 17460 9469
rect 17776 9460 17828 9512
rect 18052 9460 18104 9512
rect 18512 9460 18564 9512
rect 19156 9460 19208 9512
rect 15384 9392 15436 9444
rect 16948 9392 17000 9444
rect 17776 9367 17828 9376
rect 17776 9333 17785 9367
rect 17785 9333 17819 9367
rect 17819 9333 17828 9367
rect 17776 9324 17828 9333
rect 17868 9324 17920 9376
rect 8315 9222 8367 9274
rect 8379 9222 8431 9274
rect 8443 9222 8495 9274
rect 8507 9222 8559 9274
rect 15648 9222 15700 9274
rect 15712 9222 15764 9274
rect 15776 9222 15828 9274
rect 15840 9222 15892 9274
rect 1584 9163 1636 9172
rect 1584 9129 1593 9163
rect 1593 9129 1627 9163
rect 1627 9129 1636 9163
rect 1584 9120 1636 9129
rect 2320 9120 2372 9172
rect 3240 9163 3292 9172
rect 3240 9129 3249 9163
rect 3249 9129 3283 9163
rect 3283 9129 3292 9163
rect 3240 9120 3292 9129
rect 3792 9163 3844 9172
rect 3792 9129 3801 9163
rect 3801 9129 3835 9163
rect 3835 9129 3844 9163
rect 3792 9120 3844 9129
rect 4436 9163 4488 9172
rect 4436 9129 4445 9163
rect 4445 9129 4479 9163
rect 4479 9129 4488 9163
rect 4436 9120 4488 9129
rect 7288 9163 7340 9172
rect 7288 9129 7297 9163
rect 7297 9129 7331 9163
rect 7331 9129 7340 9163
rect 7288 9120 7340 9129
rect 7472 9120 7524 9172
rect 8208 9163 8260 9172
rect 8208 9129 8217 9163
rect 8217 9129 8251 9163
rect 8251 9129 8260 9163
rect 8208 9120 8260 9129
rect 9956 9163 10008 9172
rect 9956 9129 9965 9163
rect 9965 9129 9999 9163
rect 9999 9129 10008 9163
rect 9956 9120 10008 9129
rect 10324 9120 10376 9172
rect 12348 9163 12400 9172
rect 12348 9129 12357 9163
rect 12357 9129 12391 9163
rect 12391 9129 12400 9163
rect 12348 9120 12400 9129
rect 5816 9052 5868 9104
rect 5908 9052 5960 9104
rect 7656 9052 7708 9104
rect 1768 9027 1820 9036
rect 1768 8993 1777 9027
rect 1777 8993 1811 9027
rect 1811 8993 1820 9027
rect 1768 8984 1820 8993
rect 2872 8984 2924 9036
rect 3700 8984 3752 9036
rect 5724 8984 5776 9036
rect 6920 9027 6972 9036
rect 6920 8993 6929 9027
rect 6929 8993 6963 9027
rect 6963 8993 6972 9027
rect 6920 8984 6972 8993
rect 7472 8984 7524 9036
rect 7840 9052 7892 9104
rect 9588 9052 9640 9104
rect 8116 8984 8168 9036
rect 11336 9095 11388 9104
rect 11336 9061 11345 9095
rect 11345 9061 11379 9095
rect 11379 9061 11388 9095
rect 11336 9052 11388 9061
rect 13636 9120 13688 9172
rect 15108 9120 15160 9172
rect 18696 9120 18748 9172
rect 12624 9095 12676 9104
rect 12624 9061 12633 9095
rect 12633 9061 12667 9095
rect 12667 9061 12676 9095
rect 16396 9095 16448 9104
rect 12624 9052 12676 9061
rect 16396 9061 16405 9095
rect 16405 9061 16439 9095
rect 16439 9061 16448 9095
rect 16396 9052 16448 9061
rect 4068 8959 4120 8968
rect 4068 8925 4077 8959
rect 4077 8925 4111 8959
rect 4111 8925 4120 8959
rect 4068 8916 4120 8925
rect 6092 8916 6144 8968
rect 6276 8959 6328 8968
rect 6276 8925 6285 8959
rect 6285 8925 6319 8959
rect 6319 8925 6328 8959
rect 6276 8916 6328 8925
rect 10416 8916 10468 8968
rect 7840 8891 7892 8900
rect 7840 8857 7849 8891
rect 7849 8857 7883 8891
rect 7883 8857 7892 8891
rect 7840 8848 7892 8857
rect 8668 8848 8720 8900
rect 9864 8848 9916 8900
rect 10968 8984 11020 9036
rect 14096 9027 14148 9036
rect 14096 8993 14105 9027
rect 14105 8993 14139 9027
rect 14139 8993 14148 9027
rect 14096 8984 14148 8993
rect 17316 8984 17368 9036
rect 18696 8984 18748 9036
rect 18788 8984 18840 9036
rect 12532 8916 12584 8968
rect 16304 8959 16356 8968
rect 10600 8848 10652 8900
rect 11244 8848 11296 8900
rect 16304 8925 16313 8959
rect 16313 8925 16347 8959
rect 16347 8925 16356 8959
rect 16304 8916 16356 8925
rect 16764 8959 16816 8968
rect 16764 8925 16773 8959
rect 16773 8925 16807 8959
rect 16807 8925 16816 8959
rect 16764 8916 16816 8925
rect 17592 8959 17644 8968
rect 17592 8925 17601 8959
rect 17601 8925 17635 8959
rect 17635 8925 17644 8959
rect 17592 8916 17644 8925
rect 18420 8848 18472 8900
rect 1400 8780 1452 8832
rect 4528 8780 4580 8832
rect 5816 8780 5868 8832
rect 9036 8780 9088 8832
rect 10784 8780 10836 8832
rect 15292 8780 15344 8832
rect 18052 8823 18104 8832
rect 18052 8789 18061 8823
rect 18061 8789 18095 8823
rect 18095 8789 18104 8823
rect 18052 8780 18104 8789
rect 18236 8823 18288 8832
rect 18236 8789 18245 8823
rect 18245 8789 18279 8823
rect 18279 8789 18288 8823
rect 18236 8780 18288 8789
rect 18328 8780 18380 8832
rect 19156 8780 19208 8832
rect 4648 8678 4700 8730
rect 4712 8678 4764 8730
rect 4776 8678 4828 8730
rect 4840 8678 4892 8730
rect 11982 8678 12034 8730
rect 12046 8678 12098 8730
rect 12110 8678 12162 8730
rect 12174 8678 12226 8730
rect 19315 8678 19367 8730
rect 19379 8678 19431 8730
rect 19443 8678 19495 8730
rect 19507 8678 19559 8730
rect 1768 8576 1820 8628
rect 2872 8619 2924 8628
rect 2872 8585 2881 8619
rect 2881 8585 2915 8619
rect 2915 8585 2924 8619
rect 2872 8576 2924 8585
rect 4068 8576 4120 8628
rect 5908 8619 5960 8628
rect 5908 8585 5917 8619
rect 5917 8585 5951 8619
rect 5951 8585 5960 8619
rect 5908 8576 5960 8585
rect 6000 8576 6052 8628
rect 7564 8576 7616 8628
rect 7840 8619 7892 8628
rect 7840 8585 7849 8619
rect 7849 8585 7883 8619
rect 7883 8585 7892 8619
rect 7840 8576 7892 8585
rect 8208 8619 8260 8628
rect 8208 8585 8217 8619
rect 8217 8585 8251 8619
rect 8251 8585 8260 8619
rect 8208 8576 8260 8585
rect 8944 8576 8996 8628
rect 9864 8576 9916 8628
rect 4988 8551 5040 8560
rect 4988 8517 4997 8551
rect 4997 8517 5031 8551
rect 5031 8517 5040 8551
rect 4988 8508 5040 8517
rect 6276 8508 6328 8560
rect 6828 8508 6880 8560
rect 2412 8483 2464 8492
rect 2412 8449 2421 8483
rect 2421 8449 2455 8483
rect 2455 8449 2464 8483
rect 2412 8440 2464 8449
rect 4528 8440 4580 8492
rect 6092 8440 6144 8492
rect 12716 8576 12768 8628
rect 14096 8576 14148 8628
rect 16396 8576 16448 8628
rect 18052 8576 18104 8628
rect 18788 8576 18840 8628
rect 19984 8576 20036 8628
rect 12900 8508 12952 8560
rect 13360 8440 13412 8492
rect 14280 8440 14332 8492
rect 16212 8508 16264 8560
rect 16304 8508 16356 8560
rect 17408 8440 17460 8492
rect 18420 8440 18472 8492
rect 18604 8483 18656 8492
rect 18604 8449 18613 8483
rect 18613 8449 18647 8483
rect 18647 8449 18656 8483
rect 18604 8440 18656 8449
rect 7104 8415 7156 8424
rect 7104 8381 7113 8415
rect 7113 8381 7147 8415
rect 7147 8381 7156 8415
rect 7104 8372 7156 8381
rect 7748 8372 7800 8424
rect 8668 8415 8720 8424
rect 8668 8381 8677 8415
rect 8677 8381 8711 8415
rect 8711 8381 8720 8415
rect 8668 8372 8720 8381
rect 1952 8347 2004 8356
rect 1952 8313 1961 8347
rect 1961 8313 1995 8347
rect 1995 8313 2004 8347
rect 1952 8304 2004 8313
rect 2320 8304 2372 8356
rect 4436 8347 4488 8356
rect 4436 8313 4445 8347
rect 4445 8313 4479 8347
rect 4479 8313 4488 8347
rect 4436 8304 4488 8313
rect 4528 8347 4580 8356
rect 4528 8313 4537 8347
rect 4537 8313 4571 8347
rect 4571 8313 4580 8347
rect 4528 8304 4580 8313
rect 8208 8304 8260 8356
rect 4068 8279 4120 8288
rect 4068 8245 4077 8279
rect 4077 8245 4111 8279
rect 4111 8245 4120 8279
rect 4068 8236 4120 8245
rect 4160 8236 4212 8288
rect 10692 8304 10744 8356
rect 9588 8236 9640 8288
rect 11612 8236 11664 8288
rect 14740 8372 14792 8424
rect 16304 8372 16356 8424
rect 13544 8279 13596 8288
rect 13544 8245 13553 8279
rect 13553 8245 13587 8279
rect 13587 8245 13596 8279
rect 16120 8304 16172 8356
rect 16488 8347 16540 8356
rect 16488 8313 16497 8347
rect 16497 8313 16531 8347
rect 16531 8313 16540 8347
rect 16488 8304 16540 8313
rect 16304 8279 16356 8288
rect 13544 8236 13596 8245
rect 16304 8245 16313 8279
rect 16313 8245 16347 8279
rect 16347 8245 16356 8279
rect 18328 8304 18380 8356
rect 18420 8304 18472 8356
rect 16304 8236 16356 8245
rect 17316 8236 17368 8288
rect 8315 8134 8367 8186
rect 8379 8134 8431 8186
rect 8443 8134 8495 8186
rect 8507 8134 8559 8186
rect 15648 8134 15700 8186
rect 15712 8134 15764 8186
rect 15776 8134 15828 8186
rect 15840 8134 15892 8186
rect 3056 8075 3108 8084
rect 3056 8041 3065 8075
rect 3065 8041 3099 8075
rect 3099 8041 3108 8075
rect 3056 8032 3108 8041
rect 3332 8075 3384 8084
rect 3332 8041 3341 8075
rect 3341 8041 3375 8075
rect 3375 8041 3384 8075
rect 3332 8032 3384 8041
rect 4252 8075 4304 8084
rect 4252 8041 4261 8075
rect 4261 8041 4295 8075
rect 4295 8041 4304 8075
rect 4252 8032 4304 8041
rect 4436 8032 4488 8084
rect 6920 8032 6972 8084
rect 1860 7964 1912 8016
rect 1952 7964 2004 8016
rect 5264 7964 5316 8016
rect 1584 7896 1636 7948
rect 4160 7896 4212 7948
rect 6000 7964 6052 8016
rect 5448 7896 5500 7948
rect 5816 7896 5868 7948
rect 7472 8032 7524 8084
rect 8116 8032 8168 8084
rect 8668 8032 8720 8084
rect 9496 8032 9548 8084
rect 10968 8032 11020 8084
rect 12624 8032 12676 8084
rect 12900 8075 12952 8084
rect 12900 8041 12909 8075
rect 12909 8041 12943 8075
rect 12943 8041 12952 8075
rect 12900 8032 12952 8041
rect 14280 8032 14332 8084
rect 16488 8075 16540 8084
rect 16488 8041 16497 8075
rect 16497 8041 16531 8075
rect 16531 8041 16540 8075
rect 16488 8032 16540 8041
rect 16580 8032 16632 8084
rect 11612 7964 11664 8016
rect 14004 7964 14056 8016
rect 15384 7964 15436 8016
rect 17132 8007 17184 8016
rect 17132 7973 17141 8007
rect 17141 7973 17175 8007
rect 17175 7973 17184 8007
rect 17132 7964 17184 7973
rect 17224 8007 17276 8016
rect 17224 7973 17233 8007
rect 17233 7973 17267 8007
rect 17267 7973 17276 8007
rect 17224 7964 17276 7973
rect 18328 7964 18380 8016
rect 6460 7896 6512 7948
rect 7472 7896 7524 7948
rect 4988 7828 5040 7880
rect 9220 7896 9272 7948
rect 10232 7896 10284 7948
rect 11152 7896 11204 7948
rect 12808 7896 12860 7948
rect 7104 7760 7156 7812
rect 9128 7828 9180 7880
rect 10784 7828 10836 7880
rect 14924 7896 14976 7948
rect 15016 7896 15068 7948
rect 18144 7896 18196 7948
rect 19064 7939 19116 7948
rect 19064 7905 19073 7939
rect 19073 7905 19107 7939
rect 19107 7905 19116 7939
rect 19064 7896 19116 7905
rect 13176 7871 13228 7880
rect 13176 7837 13185 7871
rect 13185 7837 13219 7871
rect 13219 7837 13228 7871
rect 13176 7828 13228 7837
rect 17408 7871 17460 7880
rect 17408 7837 17417 7871
rect 17417 7837 17451 7871
rect 17451 7837 17460 7871
rect 17408 7828 17460 7837
rect 17500 7828 17552 7880
rect 18328 7828 18380 7880
rect 8392 7760 8444 7812
rect 9036 7760 9088 7812
rect 11888 7803 11940 7812
rect 11888 7769 11897 7803
rect 11897 7769 11931 7803
rect 11931 7769 11940 7803
rect 11888 7760 11940 7769
rect 17224 7760 17276 7812
rect 2320 7735 2372 7744
rect 2320 7701 2329 7735
rect 2329 7701 2363 7735
rect 2363 7701 2372 7735
rect 2320 7692 2372 7701
rect 6828 7735 6880 7744
rect 6828 7701 6837 7735
rect 6837 7701 6871 7735
rect 6871 7701 6880 7735
rect 6828 7692 6880 7701
rect 8116 7692 8168 7744
rect 10508 7692 10560 7744
rect 13544 7692 13596 7744
rect 15200 7692 15252 7744
rect 18696 7692 18748 7744
rect 4648 7590 4700 7642
rect 4712 7590 4764 7642
rect 4776 7590 4828 7642
rect 4840 7590 4892 7642
rect 11982 7590 12034 7642
rect 12046 7590 12098 7642
rect 12110 7590 12162 7642
rect 12174 7590 12226 7642
rect 19315 7590 19367 7642
rect 19379 7590 19431 7642
rect 19443 7590 19495 7642
rect 19507 7590 19559 7642
rect 3332 7488 3384 7540
rect 4160 7531 4212 7540
rect 4160 7497 4169 7531
rect 4169 7497 4203 7531
rect 4203 7497 4212 7531
rect 5816 7531 5868 7540
rect 4160 7488 4212 7497
rect 5816 7497 5825 7531
rect 5825 7497 5859 7531
rect 5859 7497 5868 7531
rect 5816 7488 5868 7497
rect 6000 7488 6052 7540
rect 7288 7488 7340 7540
rect 8024 7488 8076 7540
rect 8392 7531 8444 7540
rect 8392 7497 8401 7531
rect 8401 7497 8435 7531
rect 8435 7497 8444 7531
rect 8392 7488 8444 7497
rect 10232 7531 10284 7540
rect 10232 7497 10241 7531
rect 10241 7497 10275 7531
rect 10275 7497 10284 7531
rect 10232 7488 10284 7497
rect 13176 7488 13228 7540
rect 2136 7420 2188 7472
rect 3056 7352 3108 7404
rect 4988 7352 5040 7404
rect 7564 7420 7616 7472
rect 5908 7352 5960 7404
rect 9220 7420 9272 7472
rect 10876 7420 10928 7472
rect 11888 7420 11940 7472
rect 12624 7420 12676 7472
rect 13452 7420 13504 7472
rect 4252 7284 4304 7336
rect 2136 7259 2188 7268
rect 2136 7225 2145 7259
rect 2145 7225 2179 7259
rect 2179 7225 2188 7259
rect 2136 7216 2188 7225
rect 4068 7216 4120 7268
rect 2320 7148 2372 7200
rect 2780 7191 2832 7200
rect 2780 7157 2789 7191
rect 2789 7157 2823 7191
rect 2823 7157 2832 7191
rect 2780 7148 2832 7157
rect 6920 7284 6972 7336
rect 7104 7284 7156 7336
rect 7840 7284 7892 7336
rect 8668 7284 8720 7336
rect 9036 7284 9088 7336
rect 9680 7284 9732 7336
rect 10784 7327 10836 7336
rect 10784 7293 10793 7327
rect 10793 7293 10827 7327
rect 10827 7293 10836 7327
rect 10784 7284 10836 7293
rect 11428 7352 11480 7404
rect 13360 7352 13412 7404
rect 15384 7488 15436 7540
rect 15476 7488 15528 7540
rect 14740 7420 14792 7472
rect 15016 7420 15068 7472
rect 17224 7420 17276 7472
rect 16580 7352 16632 7404
rect 11336 7284 11388 7336
rect 14740 7284 14792 7336
rect 15108 7284 15160 7336
rect 15936 7284 15988 7336
rect 16304 7284 16356 7336
rect 16856 7284 16908 7336
rect 18052 7488 18104 7540
rect 19064 7531 19116 7540
rect 19064 7497 19073 7531
rect 19073 7497 19107 7531
rect 19107 7497 19116 7531
rect 19064 7488 19116 7497
rect 17500 7352 17552 7404
rect 18328 7327 18380 7336
rect 18328 7293 18337 7327
rect 18337 7293 18371 7327
rect 18371 7293 18380 7327
rect 18328 7284 18380 7293
rect 19616 7284 19668 7336
rect 11520 7259 11572 7268
rect 6460 7148 6512 7200
rect 11520 7225 11529 7259
rect 11529 7225 11563 7259
rect 11563 7225 11572 7259
rect 11520 7216 11572 7225
rect 12532 7259 12584 7268
rect 12532 7225 12541 7259
rect 12541 7225 12575 7259
rect 12575 7225 12584 7259
rect 12532 7216 12584 7225
rect 12624 7259 12676 7268
rect 12624 7225 12633 7259
rect 12633 7225 12667 7259
rect 12667 7225 12676 7259
rect 12624 7216 12676 7225
rect 15384 7216 15436 7268
rect 18788 7259 18840 7268
rect 18788 7225 18797 7259
rect 18797 7225 18831 7259
rect 18831 7225 18840 7259
rect 18788 7216 18840 7225
rect 7472 7148 7524 7200
rect 9220 7148 9272 7200
rect 9864 7191 9916 7200
rect 9864 7157 9873 7191
rect 9873 7157 9907 7191
rect 9907 7157 9916 7191
rect 9864 7148 9916 7157
rect 10876 7148 10928 7200
rect 11612 7148 11664 7200
rect 14004 7148 14056 7200
rect 14188 7148 14240 7200
rect 18512 7148 18564 7200
rect 19064 7148 19116 7200
rect 20168 7191 20220 7200
rect 20168 7157 20177 7191
rect 20177 7157 20211 7191
rect 20211 7157 20220 7191
rect 20168 7148 20220 7157
rect 8315 7046 8367 7098
rect 8379 7046 8431 7098
rect 8443 7046 8495 7098
rect 8507 7046 8559 7098
rect 15648 7046 15700 7098
rect 15712 7046 15764 7098
rect 15776 7046 15828 7098
rect 15840 7046 15892 7098
rect 1400 6987 1452 6996
rect 1400 6953 1409 6987
rect 1409 6953 1443 6987
rect 1443 6953 1452 6987
rect 1400 6944 1452 6953
rect 1584 6944 1636 6996
rect 2688 6851 2740 6860
rect 2688 6817 2697 6851
rect 2697 6817 2731 6851
rect 2731 6817 2740 6851
rect 2688 6808 2740 6817
rect 2872 6851 2924 6860
rect 2872 6817 2881 6851
rect 2881 6817 2915 6851
rect 2915 6817 2924 6851
rect 2872 6808 2924 6817
rect 3148 6783 3200 6792
rect 3148 6749 3157 6783
rect 3157 6749 3191 6783
rect 3191 6749 3200 6783
rect 3148 6740 3200 6749
rect 6368 6944 6420 6996
rect 6920 6987 6972 6996
rect 6920 6953 6929 6987
rect 6929 6953 6963 6987
rect 6963 6953 6972 6987
rect 6920 6944 6972 6953
rect 4252 6919 4304 6928
rect 4252 6885 4261 6919
rect 4261 6885 4295 6919
rect 4295 6885 4304 6919
rect 4252 6876 4304 6885
rect 6000 6876 6052 6928
rect 7472 6944 7524 6996
rect 9036 6987 9088 6996
rect 9036 6953 9045 6987
rect 9045 6953 9079 6987
rect 9079 6953 9088 6987
rect 9036 6944 9088 6953
rect 9312 6987 9364 6996
rect 9312 6953 9321 6987
rect 9321 6953 9355 6987
rect 9355 6953 9364 6987
rect 9312 6944 9364 6953
rect 10784 6987 10836 6996
rect 10784 6953 10793 6987
rect 10793 6953 10827 6987
rect 10827 6953 10836 6987
rect 10784 6944 10836 6953
rect 11152 6987 11204 6996
rect 11152 6953 11161 6987
rect 11161 6953 11195 6987
rect 11195 6953 11204 6987
rect 11152 6944 11204 6953
rect 11520 6944 11572 6996
rect 14096 6944 14148 6996
rect 15108 6987 15160 6996
rect 15108 6953 15117 6987
rect 15117 6953 15151 6987
rect 15151 6953 15160 6987
rect 15108 6944 15160 6953
rect 15384 6944 15436 6996
rect 5724 6808 5776 6860
rect 5908 6851 5960 6860
rect 5908 6817 5917 6851
rect 5917 6817 5951 6851
rect 5951 6817 5960 6851
rect 5908 6808 5960 6817
rect 6276 6808 6328 6860
rect 7196 6808 7248 6860
rect 7472 6808 7524 6860
rect 8944 6876 8996 6928
rect 9864 6919 9916 6928
rect 9864 6885 9873 6919
rect 9873 6885 9907 6919
rect 9907 6885 9916 6919
rect 9864 6876 9916 6885
rect 11428 6876 11480 6928
rect 11796 6919 11848 6928
rect 11796 6885 11805 6919
rect 11805 6885 11839 6919
rect 11839 6885 11848 6919
rect 11796 6876 11848 6885
rect 12992 6919 13044 6928
rect 12992 6885 13001 6919
rect 13001 6885 13035 6919
rect 13035 6885 13044 6919
rect 12992 6876 13044 6885
rect 13544 6919 13596 6928
rect 13544 6885 13553 6919
rect 13553 6885 13587 6919
rect 13587 6885 13596 6919
rect 13544 6876 13596 6885
rect 8116 6808 8168 6860
rect 8484 6851 8536 6860
rect 8484 6817 8493 6851
rect 8493 6817 8527 6851
rect 8527 6817 8536 6851
rect 8484 6808 8536 6817
rect 16856 6876 16908 6928
rect 17132 6944 17184 6996
rect 18144 6987 18196 6996
rect 18144 6953 18153 6987
rect 18153 6953 18187 6987
rect 18187 6953 18196 6987
rect 18144 6944 18196 6953
rect 19800 6944 19852 6996
rect 21640 6944 21692 6996
rect 18604 6876 18656 6928
rect 2872 6672 2924 6724
rect 7932 6783 7984 6792
rect 7932 6749 7941 6783
rect 7941 6749 7975 6783
rect 7975 6749 7984 6783
rect 7932 6740 7984 6749
rect 8760 6740 8812 6792
rect 9772 6783 9824 6792
rect 9772 6749 9781 6783
rect 9781 6749 9815 6783
rect 9815 6749 9824 6783
rect 9772 6740 9824 6749
rect 11704 6783 11756 6792
rect 11704 6749 11713 6783
rect 11713 6749 11747 6783
rect 11747 6749 11756 6783
rect 11704 6740 11756 6749
rect 12808 6740 12860 6792
rect 13084 6740 13136 6792
rect 4344 6672 4396 6724
rect 1860 6647 1912 6656
rect 1860 6613 1869 6647
rect 1869 6613 1903 6647
rect 1903 6613 1912 6647
rect 1860 6604 1912 6613
rect 2780 6604 2832 6656
rect 4436 6604 4488 6656
rect 5356 6647 5408 6656
rect 5356 6613 5365 6647
rect 5365 6613 5399 6647
rect 5399 6613 5408 6647
rect 5356 6604 5408 6613
rect 6552 6672 6604 6724
rect 10048 6672 10100 6724
rect 11612 6672 11664 6724
rect 12532 6672 12584 6724
rect 15384 6808 15436 6860
rect 18236 6851 18288 6860
rect 18236 6817 18245 6851
rect 18245 6817 18279 6851
rect 18279 6817 18288 6851
rect 18236 6808 18288 6817
rect 18512 6851 18564 6860
rect 18512 6817 18521 6851
rect 18521 6817 18555 6851
rect 18555 6817 18564 6851
rect 18512 6808 18564 6817
rect 16672 6740 16724 6792
rect 17684 6740 17736 6792
rect 20444 6740 20496 6792
rect 14648 6672 14700 6724
rect 5908 6604 5960 6656
rect 8116 6604 8168 6656
rect 15936 6604 15988 6656
rect 16304 6604 16356 6656
rect 4648 6502 4700 6554
rect 4712 6502 4764 6554
rect 4776 6502 4828 6554
rect 4840 6502 4892 6554
rect 11982 6502 12034 6554
rect 12046 6502 12098 6554
rect 12110 6502 12162 6554
rect 12174 6502 12226 6554
rect 19315 6502 19367 6554
rect 19379 6502 19431 6554
rect 19443 6502 19495 6554
rect 19507 6502 19559 6554
rect 848 6400 900 6452
rect 2412 6375 2464 6384
rect 2412 6341 2421 6375
rect 2421 6341 2455 6375
rect 2455 6341 2464 6375
rect 2412 6332 2464 6341
rect 2872 6400 2924 6452
rect 3240 6400 3292 6452
rect 4252 6400 4304 6452
rect 5724 6400 5776 6452
rect 11520 6400 11572 6452
rect 11612 6400 11664 6452
rect 13544 6443 13596 6452
rect 6460 6332 6512 6384
rect 6552 6332 6604 6384
rect 9772 6375 9824 6384
rect 9772 6341 9781 6375
rect 9781 6341 9815 6375
rect 9815 6341 9824 6375
rect 9772 6332 9824 6341
rect 3056 6264 3108 6316
rect 3424 6264 3476 6316
rect 4344 6264 4396 6316
rect 4988 6264 5040 6316
rect 5448 6264 5500 6316
rect 5540 6264 5592 6316
rect 7656 6264 7708 6316
rect 7840 6307 7892 6316
rect 7840 6273 7849 6307
rect 7849 6273 7883 6307
rect 7883 6273 7892 6307
rect 7840 6264 7892 6273
rect 9312 6264 9364 6316
rect 12992 6332 13044 6384
rect 13544 6409 13553 6443
rect 13553 6409 13587 6443
rect 13587 6409 13596 6443
rect 13544 6400 13596 6409
rect 15384 6443 15436 6452
rect 15384 6409 15393 6443
rect 15393 6409 15427 6443
rect 15427 6409 15436 6443
rect 16856 6443 16908 6452
rect 15384 6400 15436 6409
rect 16028 6332 16080 6384
rect 16856 6409 16865 6443
rect 16865 6409 16899 6443
rect 16899 6409 16908 6443
rect 16856 6400 16908 6409
rect 18236 6400 18288 6452
rect 19064 6443 19116 6452
rect 19064 6409 19073 6443
rect 19073 6409 19107 6443
rect 19107 6409 19116 6443
rect 19064 6400 19116 6409
rect 20444 6443 20496 6452
rect 20444 6409 20453 6443
rect 20453 6409 20487 6443
rect 20487 6409 20496 6443
rect 20444 6400 20496 6409
rect 17592 6332 17644 6384
rect 12900 6307 12952 6316
rect 12900 6273 12909 6307
rect 12909 6273 12943 6307
rect 12943 6273 12952 6307
rect 12900 6264 12952 6273
rect 14096 6307 14148 6316
rect 14096 6273 14105 6307
rect 14105 6273 14139 6307
rect 14139 6273 14148 6307
rect 14096 6264 14148 6273
rect 15016 6264 15068 6316
rect 2688 6196 2740 6248
rect 3976 6196 4028 6248
rect 5632 6196 5684 6248
rect 10324 6239 10376 6248
rect 10324 6205 10333 6239
rect 10333 6205 10367 6239
rect 10367 6205 10376 6239
rect 10324 6196 10376 6205
rect 18236 6239 18288 6248
rect 18236 6205 18245 6239
rect 18245 6205 18279 6239
rect 18279 6205 18288 6239
rect 18236 6196 18288 6205
rect 4252 6171 4304 6180
rect 4252 6137 4261 6171
rect 4261 6137 4295 6171
rect 4295 6137 4304 6171
rect 4252 6128 4304 6137
rect 5448 6128 5500 6180
rect 6276 6171 6328 6180
rect 6276 6137 6285 6171
rect 6285 6137 6319 6171
rect 6319 6137 6328 6171
rect 6276 6128 6328 6137
rect 7012 6171 7064 6180
rect 7012 6137 7021 6171
rect 7021 6137 7055 6171
rect 7055 6137 7064 6171
rect 7012 6128 7064 6137
rect 7196 6128 7248 6180
rect 2320 6060 2372 6112
rect 5908 6060 5960 6112
rect 8760 6171 8812 6180
rect 8760 6137 8769 6171
rect 8769 6137 8803 6171
rect 8803 6137 8812 6171
rect 8760 6128 8812 6137
rect 10876 6128 10928 6180
rect 9588 6060 9640 6112
rect 11244 6103 11296 6112
rect 11244 6069 11253 6103
rect 11253 6069 11287 6103
rect 11287 6069 11296 6103
rect 11244 6060 11296 6069
rect 11612 6103 11664 6112
rect 11612 6069 11621 6103
rect 11621 6069 11655 6103
rect 11655 6069 11664 6103
rect 11612 6060 11664 6069
rect 11796 6060 11848 6112
rect 14096 6128 14148 6180
rect 14924 6128 14976 6180
rect 15936 6171 15988 6180
rect 15200 6060 15252 6112
rect 15936 6137 15945 6171
rect 15945 6137 15979 6171
rect 15979 6137 15988 6171
rect 15936 6128 15988 6137
rect 17316 6128 17368 6180
rect 19984 6196 20036 6248
rect 17868 6060 17920 6112
rect 8315 5958 8367 6010
rect 8379 5958 8431 6010
rect 8443 5958 8495 6010
rect 8507 5958 8559 6010
rect 15648 5958 15700 6010
rect 15712 5958 15764 6010
rect 15776 5958 15828 6010
rect 15840 5958 15892 6010
rect 2320 5899 2372 5908
rect 2320 5865 2329 5899
rect 2329 5865 2363 5899
rect 2363 5865 2372 5899
rect 2320 5856 2372 5865
rect 2412 5856 2464 5908
rect 3424 5899 3476 5908
rect 3424 5865 3433 5899
rect 3433 5865 3467 5899
rect 3467 5865 3476 5899
rect 3424 5856 3476 5865
rect 4252 5856 4304 5908
rect 5540 5899 5592 5908
rect 5540 5865 5549 5899
rect 5549 5865 5583 5899
rect 5583 5865 5592 5899
rect 5540 5856 5592 5865
rect 7472 5899 7524 5908
rect 7472 5865 7481 5899
rect 7481 5865 7515 5899
rect 7515 5865 7524 5899
rect 7472 5856 7524 5865
rect 9864 5899 9916 5908
rect 9864 5865 9873 5899
rect 9873 5865 9907 5899
rect 9907 5865 9916 5899
rect 9864 5856 9916 5865
rect 11612 5856 11664 5908
rect 11704 5899 11756 5908
rect 11704 5865 11713 5899
rect 11713 5865 11747 5899
rect 11747 5865 11756 5899
rect 11704 5856 11756 5865
rect 15016 5856 15068 5908
rect 1860 5788 1912 5840
rect 2504 5788 2556 5840
rect 3700 5788 3752 5840
rect 6644 5788 6696 5840
rect 9220 5788 9272 5840
rect 10876 5788 10928 5840
rect 11244 5788 11296 5840
rect 12348 5831 12400 5840
rect 12348 5797 12357 5831
rect 12357 5797 12391 5831
rect 12391 5797 12400 5831
rect 12348 5788 12400 5797
rect 13084 5788 13136 5840
rect 3056 5763 3108 5772
rect 3056 5729 3065 5763
rect 3065 5729 3099 5763
rect 3099 5729 3108 5763
rect 3056 5720 3108 5729
rect 3148 5720 3200 5772
rect 4068 5763 4120 5772
rect 4068 5729 4077 5763
rect 4077 5729 4111 5763
rect 4111 5729 4120 5763
rect 4068 5720 4120 5729
rect 7932 5720 7984 5772
rect 14188 5720 14240 5772
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 5632 5652 5684 5704
rect 10416 5695 10468 5704
rect 10416 5661 10425 5695
rect 10425 5661 10459 5695
rect 10459 5661 10468 5695
rect 10416 5652 10468 5661
rect 11520 5652 11572 5704
rect 12716 5652 12768 5704
rect 12900 5695 12952 5704
rect 12900 5661 12909 5695
rect 12909 5661 12943 5695
rect 12943 5661 12952 5695
rect 12900 5652 12952 5661
rect 3976 5584 4028 5636
rect 10048 5584 10100 5636
rect 10324 5627 10376 5636
rect 10324 5593 10333 5627
rect 10333 5593 10367 5627
rect 10367 5593 10376 5627
rect 15200 5788 15252 5840
rect 16672 5788 16724 5840
rect 17040 5831 17092 5840
rect 17040 5797 17049 5831
rect 17049 5797 17083 5831
rect 17083 5797 17092 5831
rect 17040 5788 17092 5797
rect 18604 5763 18656 5772
rect 18604 5729 18613 5763
rect 18613 5729 18647 5763
rect 18647 5729 18656 5763
rect 18604 5720 18656 5729
rect 16028 5695 16080 5704
rect 16028 5661 16037 5695
rect 16037 5661 16071 5695
rect 16071 5661 16080 5695
rect 16028 5652 16080 5661
rect 16948 5695 17000 5704
rect 16948 5661 16957 5695
rect 16957 5661 16991 5695
rect 16991 5661 17000 5695
rect 16948 5652 17000 5661
rect 17224 5695 17276 5704
rect 17224 5661 17233 5695
rect 17233 5661 17267 5695
rect 17267 5661 17276 5695
rect 17224 5652 17276 5661
rect 10324 5584 10376 5593
rect 3792 5559 3844 5568
rect 3792 5525 3801 5559
rect 3801 5525 3835 5559
rect 3835 5525 3844 5559
rect 3792 5516 3844 5525
rect 7012 5516 7064 5568
rect 8760 5559 8812 5568
rect 8760 5525 8769 5559
rect 8769 5525 8803 5559
rect 8803 5525 8812 5559
rect 8760 5516 8812 5525
rect 14280 5559 14332 5568
rect 14280 5525 14289 5559
rect 14289 5525 14323 5559
rect 14323 5525 14332 5559
rect 14280 5516 14332 5525
rect 16304 5584 16356 5636
rect 15844 5516 15896 5568
rect 17500 5516 17552 5568
rect 17684 5516 17736 5568
rect 18512 5652 18564 5704
rect 19064 5652 19116 5704
rect 4648 5414 4700 5466
rect 4712 5414 4764 5466
rect 4776 5414 4828 5466
rect 4840 5414 4892 5466
rect 11982 5414 12034 5466
rect 12046 5414 12098 5466
rect 12110 5414 12162 5466
rect 12174 5414 12226 5466
rect 19315 5414 19367 5466
rect 19379 5414 19431 5466
rect 19443 5414 19495 5466
rect 19507 5414 19559 5466
rect 1400 5312 1452 5364
rect 2872 5312 2924 5364
rect 4068 5312 4120 5364
rect 6644 5355 6696 5364
rect 6644 5321 6653 5355
rect 6653 5321 6687 5355
rect 6687 5321 6696 5355
rect 6644 5312 6696 5321
rect 10416 5312 10468 5364
rect 10508 5312 10560 5364
rect 12348 5312 12400 5364
rect 14188 5312 14240 5364
rect 14924 5355 14976 5364
rect 14924 5321 14933 5355
rect 14933 5321 14967 5355
rect 14967 5321 14976 5355
rect 14924 5312 14976 5321
rect 15200 5312 15252 5364
rect 15936 5312 15988 5364
rect 19064 5355 19116 5364
rect 2136 5244 2188 5296
rect 2780 5244 2832 5296
rect 3700 5244 3752 5296
rect 10048 5287 10100 5296
rect 10048 5253 10057 5287
rect 10057 5253 10091 5287
rect 10091 5253 10100 5287
rect 10048 5244 10100 5253
rect 17040 5244 17092 5296
rect 19064 5321 19073 5355
rect 19073 5321 19107 5355
rect 19107 5321 19116 5355
rect 19064 5312 19116 5321
rect 2504 5176 2556 5228
rect 5264 5176 5316 5228
rect 8668 5176 8720 5228
rect 3148 5108 3200 5160
rect 3792 5151 3844 5160
rect 3792 5117 3801 5151
rect 3801 5117 3835 5151
rect 3835 5117 3844 5151
rect 3792 5108 3844 5117
rect 10876 5176 10928 5228
rect 11520 5176 11572 5228
rect 12808 5219 12860 5228
rect 12808 5185 12817 5219
rect 12817 5185 12851 5219
rect 12851 5185 12860 5219
rect 12808 5176 12860 5185
rect 13360 5176 13412 5228
rect 17868 5176 17920 5228
rect 10784 5151 10836 5160
rect 2228 5040 2280 5092
rect 3700 5040 3752 5092
rect 10784 5117 10793 5151
rect 10793 5117 10827 5151
rect 10827 5117 10836 5151
rect 10784 5108 10836 5117
rect 11336 5151 11388 5160
rect 11336 5117 11345 5151
rect 11345 5117 11379 5151
rect 11379 5117 11388 5151
rect 11336 5108 11388 5117
rect 16488 5151 16540 5160
rect 16488 5117 16497 5151
rect 16497 5117 16531 5151
rect 16531 5117 16540 5151
rect 16488 5108 16540 5117
rect 17224 5108 17276 5160
rect 17776 5108 17828 5160
rect 20076 5151 20128 5160
rect 20076 5117 20085 5151
rect 20085 5117 20119 5151
rect 20119 5117 20128 5151
rect 20076 5108 20128 5117
rect 6920 5083 6972 5092
rect 6920 5049 6929 5083
rect 6929 5049 6963 5083
rect 6963 5049 6972 5083
rect 6920 5040 6972 5049
rect 7012 5083 7064 5092
rect 7012 5049 7021 5083
rect 7021 5049 7055 5083
rect 7055 5049 7064 5083
rect 7012 5040 7064 5049
rect 8116 5040 8168 5092
rect 4712 5015 4764 5024
rect 4712 4981 4721 5015
rect 4721 4981 4755 5015
rect 4755 4981 4764 5015
rect 4712 4972 4764 4981
rect 5632 5015 5684 5024
rect 5632 4981 5641 5015
rect 5641 4981 5675 5015
rect 5675 4981 5684 5015
rect 5632 4972 5684 4981
rect 6092 4972 6144 5024
rect 6276 5015 6328 5024
rect 6276 4981 6285 5015
rect 6285 4981 6319 5015
rect 6319 4981 6328 5015
rect 6276 4972 6328 4981
rect 8760 5040 8812 5092
rect 11428 5040 11480 5092
rect 12348 4972 12400 5024
rect 14096 5040 14148 5092
rect 15108 5040 15160 5092
rect 15844 5083 15896 5092
rect 15844 5049 15853 5083
rect 15853 5049 15887 5083
rect 15887 5049 15896 5083
rect 15844 5040 15896 5049
rect 18052 5083 18104 5092
rect 15200 4972 15252 5024
rect 18052 5049 18061 5083
rect 18061 5049 18095 5083
rect 18095 5049 18104 5083
rect 18052 5040 18104 5049
rect 16304 4972 16356 5024
rect 16948 4972 17000 5024
rect 17776 5015 17828 5024
rect 17776 4981 17785 5015
rect 17785 4981 17819 5015
rect 17819 4981 17828 5015
rect 17776 4972 17828 4981
rect 19708 4972 19760 5024
rect 8315 4870 8367 4922
rect 8379 4870 8431 4922
rect 8443 4870 8495 4922
rect 8507 4870 8559 4922
rect 15648 4870 15700 4922
rect 15712 4870 15764 4922
rect 15776 4870 15828 4922
rect 15840 4870 15892 4922
rect 2136 4768 2188 4820
rect 2688 4675 2740 4684
rect 2688 4641 2697 4675
rect 2697 4641 2731 4675
rect 2731 4641 2740 4675
rect 2688 4632 2740 4641
rect 3148 4675 3200 4684
rect 1768 4496 1820 4548
rect 2780 4496 2832 4548
rect 3148 4641 3157 4675
rect 3157 4641 3191 4675
rect 3191 4641 3200 4675
rect 3148 4632 3200 4641
rect 3700 4700 3752 4752
rect 7012 4768 7064 4820
rect 7932 4811 7984 4820
rect 7932 4777 7941 4811
rect 7941 4777 7975 4811
rect 7975 4777 7984 4811
rect 7932 4768 7984 4777
rect 8116 4768 8168 4820
rect 10140 4768 10192 4820
rect 4528 4700 4580 4752
rect 4712 4700 4764 4752
rect 4988 4700 5040 4752
rect 6644 4743 6696 4752
rect 6644 4709 6653 4743
rect 6653 4709 6687 4743
rect 6687 4709 6696 4743
rect 6644 4700 6696 4709
rect 7288 4700 7340 4752
rect 8208 4743 8260 4752
rect 8208 4709 8217 4743
rect 8217 4709 8251 4743
rect 8251 4709 8260 4743
rect 8208 4700 8260 4709
rect 8760 4632 8812 4684
rect 9496 4632 9548 4684
rect 9864 4675 9916 4684
rect 9864 4641 9873 4675
rect 9873 4641 9907 4675
rect 9907 4641 9916 4675
rect 9864 4632 9916 4641
rect 9956 4632 10008 4684
rect 11244 4768 11296 4820
rect 11520 4743 11572 4752
rect 11520 4709 11529 4743
rect 11529 4709 11563 4743
rect 11563 4709 11572 4743
rect 11520 4700 11572 4709
rect 11704 4700 11756 4752
rect 12348 4768 12400 4820
rect 12716 4768 12768 4820
rect 15108 4811 15160 4820
rect 13268 4700 13320 4752
rect 15108 4777 15117 4811
rect 15117 4777 15151 4811
rect 15151 4777 15160 4811
rect 15108 4768 15160 4777
rect 16304 4811 16356 4820
rect 15476 4743 15528 4752
rect 15476 4709 15485 4743
rect 15485 4709 15519 4743
rect 15519 4709 15528 4743
rect 15476 4700 15528 4709
rect 16304 4777 16313 4811
rect 16313 4777 16347 4811
rect 16347 4777 16356 4811
rect 16304 4768 16356 4777
rect 16948 4811 17000 4820
rect 16948 4777 16957 4811
rect 16957 4777 16991 4811
rect 16991 4777 17000 4811
rect 16948 4768 17000 4777
rect 18696 4811 18748 4820
rect 18696 4777 18705 4811
rect 18705 4777 18739 4811
rect 18739 4777 18748 4811
rect 18696 4768 18748 4777
rect 16304 4632 16356 4684
rect 17316 4675 17368 4684
rect 5540 4564 5592 4616
rect 6552 4607 6604 4616
rect 6552 4573 6561 4607
rect 6561 4573 6595 4607
rect 6595 4573 6604 4607
rect 6552 4564 6604 4573
rect 7472 4564 7524 4616
rect 10600 4607 10652 4616
rect 3240 4496 3292 4548
rect 6920 4496 6972 4548
rect 7380 4496 7432 4548
rect 10600 4573 10609 4607
rect 10609 4573 10643 4607
rect 10643 4573 10652 4607
rect 10600 4564 10652 4573
rect 12348 4564 12400 4616
rect 13084 4607 13136 4616
rect 13084 4573 13093 4607
rect 13093 4573 13127 4607
rect 13127 4573 13136 4607
rect 13084 4564 13136 4573
rect 13360 4607 13412 4616
rect 13360 4573 13369 4607
rect 13369 4573 13403 4607
rect 13403 4573 13412 4607
rect 13360 4564 13412 4573
rect 16396 4564 16448 4616
rect 17316 4641 17325 4675
rect 17325 4641 17359 4675
rect 17359 4641 17368 4675
rect 17316 4632 17368 4641
rect 18880 4700 18932 4752
rect 18512 4675 18564 4684
rect 18512 4641 18521 4675
rect 18521 4641 18555 4675
rect 18555 4641 18564 4675
rect 18512 4632 18564 4641
rect 18144 4564 18196 4616
rect 8668 4539 8720 4548
rect 8668 4505 8677 4539
rect 8677 4505 8711 4539
rect 8711 4505 8720 4539
rect 8668 4496 8720 4505
rect 15936 4539 15988 4548
rect 15936 4505 15945 4539
rect 15945 4505 15979 4539
rect 15979 4505 15988 4539
rect 15936 4496 15988 4505
rect 1860 4471 1912 4480
rect 1860 4437 1869 4471
rect 1869 4437 1903 4471
rect 1903 4437 1912 4471
rect 1860 4428 1912 4437
rect 8116 4428 8168 4480
rect 11060 4428 11112 4480
rect 14096 4471 14148 4480
rect 14096 4437 14105 4471
rect 14105 4437 14139 4471
rect 14139 4437 14148 4471
rect 14096 4428 14148 4437
rect 16488 4428 16540 4480
rect 18604 4428 18656 4480
rect 19708 4428 19760 4480
rect 4648 4326 4700 4378
rect 4712 4326 4764 4378
rect 4776 4326 4828 4378
rect 4840 4326 4892 4378
rect 11982 4326 12034 4378
rect 12046 4326 12098 4378
rect 12110 4326 12162 4378
rect 12174 4326 12226 4378
rect 19315 4326 19367 4378
rect 19379 4326 19431 4378
rect 19443 4326 19495 4378
rect 19507 4326 19559 4378
rect 1768 4267 1820 4276
rect 1768 4233 1777 4267
rect 1777 4233 1811 4267
rect 1811 4233 1820 4267
rect 1768 4224 1820 4233
rect 2412 4224 2464 4276
rect 2688 4224 2740 4276
rect 4528 4224 4580 4276
rect 8208 4224 8260 4276
rect 9956 4267 10008 4276
rect 9956 4233 9965 4267
rect 9965 4233 9999 4267
rect 9999 4233 10008 4267
rect 9956 4224 10008 4233
rect 8760 4156 8812 4208
rect 10324 4156 10376 4208
rect 3516 4088 3568 4140
rect 4988 4088 5040 4140
rect 5356 4088 5408 4140
rect 5908 4131 5960 4140
rect 2780 4063 2832 4072
rect 2780 4029 2789 4063
rect 2789 4029 2823 4063
rect 2823 4029 2832 4063
rect 2780 4020 2832 4029
rect 5908 4097 5917 4131
rect 5917 4097 5951 4131
rect 5951 4097 5960 4131
rect 5908 4088 5960 4097
rect 11796 4088 11848 4140
rect 12900 4088 12952 4140
rect 13084 4156 13136 4208
rect 15108 4224 15160 4276
rect 18420 4224 18472 4276
rect 18512 4224 18564 4276
rect 16304 4088 16356 4140
rect 16488 4131 16540 4140
rect 16488 4097 16497 4131
rect 16497 4097 16531 4131
rect 16531 4097 16540 4131
rect 16488 4088 16540 4097
rect 16764 4088 16816 4140
rect 7564 4020 7616 4072
rect 9036 4020 9088 4072
rect 11152 4020 11204 4072
rect 3424 3952 3476 4004
rect 4160 3952 4212 4004
rect 5816 3952 5868 4004
rect 7840 3952 7892 4004
rect 3608 3927 3660 3936
rect 3608 3893 3617 3927
rect 3617 3893 3651 3927
rect 3651 3893 3660 3927
rect 3608 3884 3660 3893
rect 6552 3927 6604 3936
rect 6552 3893 6561 3927
rect 6561 3893 6595 3927
rect 6595 3893 6604 3927
rect 6552 3884 6604 3893
rect 6644 3884 6696 3936
rect 11704 3927 11756 3936
rect 11704 3893 11713 3927
rect 11713 3893 11747 3927
rect 11747 3893 11756 3927
rect 11704 3884 11756 3893
rect 14740 4020 14792 4072
rect 18144 4063 18196 4072
rect 12348 3952 12400 4004
rect 14188 3952 14240 4004
rect 15476 3952 15528 4004
rect 13268 3884 13320 3936
rect 14096 3884 14148 3936
rect 15384 3884 15436 3936
rect 16028 3884 16080 3936
rect 18144 4029 18153 4063
rect 18153 4029 18187 4063
rect 18187 4029 18196 4063
rect 18144 4020 18196 4029
rect 16580 3995 16632 4004
rect 16580 3961 16589 3995
rect 16589 3961 16623 3995
rect 16623 3961 16632 3995
rect 17132 3995 17184 4004
rect 16580 3952 16632 3961
rect 17132 3961 17141 3995
rect 17141 3961 17175 3995
rect 17175 3961 17184 3995
rect 17132 3952 17184 3961
rect 18604 4020 18656 4072
rect 17316 3884 17368 3936
rect 17684 3884 17736 3936
rect 18144 3927 18196 3936
rect 18144 3893 18153 3927
rect 18153 3893 18187 3927
rect 18187 3893 18196 3927
rect 18144 3884 18196 3893
rect 8315 3782 8367 3834
rect 8379 3782 8431 3834
rect 8443 3782 8495 3834
rect 8507 3782 8559 3834
rect 15648 3782 15700 3834
rect 15712 3782 15764 3834
rect 15776 3782 15828 3834
rect 15840 3782 15892 3834
rect 3608 3680 3660 3732
rect 5264 3723 5316 3732
rect 5264 3689 5273 3723
rect 5273 3689 5307 3723
rect 5307 3689 5316 3723
rect 5264 3680 5316 3689
rect 6644 3680 6696 3732
rect 8116 3680 8168 3732
rect 9036 3723 9088 3732
rect 9036 3689 9045 3723
rect 9045 3689 9079 3723
rect 9079 3689 9088 3723
rect 9036 3680 9088 3689
rect 10600 3680 10652 3732
rect 14188 3723 14240 3732
rect 2044 3612 2096 3664
rect 2780 3612 2832 3664
rect 3424 3655 3476 3664
rect 3424 3621 3433 3655
rect 3433 3621 3467 3655
rect 3467 3621 3476 3655
rect 3424 3612 3476 3621
rect 3792 3612 3844 3664
rect 4528 3612 4580 3664
rect 6552 3612 6604 3664
rect 8208 3655 8260 3664
rect 8208 3621 8217 3655
rect 8217 3621 8251 3655
rect 8251 3621 8260 3655
rect 8208 3612 8260 3621
rect 9404 3655 9456 3664
rect 9404 3621 9413 3655
rect 9413 3621 9447 3655
rect 9447 3621 9456 3655
rect 9404 3612 9456 3621
rect 11612 3655 11664 3664
rect 11612 3621 11621 3655
rect 11621 3621 11655 3655
rect 11655 3621 11664 3655
rect 11612 3612 11664 3621
rect 2688 3587 2740 3596
rect 2688 3553 2697 3587
rect 2697 3553 2731 3587
rect 2731 3553 2740 3587
rect 2688 3544 2740 3553
rect 2964 3587 3016 3596
rect 2964 3553 2973 3587
rect 2973 3553 3007 3587
rect 3007 3553 3016 3587
rect 2964 3544 3016 3553
rect 3332 3476 3384 3528
rect 4160 3544 4212 3596
rect 9588 3544 9640 3596
rect 9956 3587 10008 3596
rect 9956 3553 9965 3587
rect 9965 3553 9999 3587
rect 9999 3553 10008 3587
rect 9956 3544 10008 3553
rect 10048 3544 10100 3596
rect 10324 3544 10376 3596
rect 6368 3476 6420 3528
rect 7472 3476 7524 3528
rect 8116 3519 8168 3528
rect 8116 3485 8125 3519
rect 8125 3485 8159 3519
rect 8159 3485 8168 3519
rect 8116 3476 8168 3485
rect 1768 3408 1820 3460
rect 5172 3408 5224 3460
rect 5356 3408 5408 3460
rect 11152 3519 11204 3528
rect 11152 3485 11161 3519
rect 11161 3485 11195 3519
rect 11195 3485 11204 3519
rect 11152 3476 11204 3485
rect 11796 3476 11848 3528
rect 9588 3408 9640 3460
rect 12256 3612 12308 3664
rect 12348 3612 12400 3664
rect 14188 3689 14197 3723
rect 14197 3689 14231 3723
rect 14231 3689 14240 3723
rect 14188 3680 14240 3689
rect 15108 3723 15160 3732
rect 15108 3689 15117 3723
rect 15117 3689 15151 3723
rect 15151 3689 15160 3723
rect 15108 3680 15160 3689
rect 13820 3612 13872 3664
rect 14740 3612 14792 3664
rect 15476 3655 15528 3664
rect 15476 3621 15485 3655
rect 15485 3621 15519 3655
rect 15519 3621 15528 3655
rect 15476 3612 15528 3621
rect 16580 3680 16632 3732
rect 18512 3723 18564 3732
rect 18512 3689 18521 3723
rect 18521 3689 18555 3723
rect 18555 3689 18564 3723
rect 18512 3680 18564 3689
rect 16948 3612 17000 3664
rect 17224 3544 17276 3596
rect 17316 3587 17368 3596
rect 17316 3553 17325 3587
rect 17325 3553 17359 3587
rect 17359 3553 17368 3587
rect 17316 3544 17368 3553
rect 17776 3544 17828 3596
rect 18788 3544 18840 3596
rect 18972 3587 19024 3596
rect 18972 3553 18981 3587
rect 18981 3553 19015 3587
rect 19015 3553 19024 3587
rect 18972 3544 19024 3553
rect 15384 3519 15436 3528
rect 15384 3485 15393 3519
rect 15393 3485 15427 3519
rect 15427 3485 15436 3519
rect 15384 3476 15436 3485
rect 13360 3408 13412 3460
rect 15936 3451 15988 3460
rect 15936 3417 15945 3451
rect 15945 3417 15979 3451
rect 15979 3417 15988 3451
rect 15936 3408 15988 3417
rect 7104 3340 7156 3392
rect 7564 3383 7616 3392
rect 7564 3349 7573 3383
rect 7573 3349 7607 3383
rect 7607 3349 7616 3383
rect 7564 3340 7616 3349
rect 8116 3340 8168 3392
rect 9404 3340 9456 3392
rect 9864 3340 9916 3392
rect 16488 3340 16540 3392
rect 17684 3340 17736 3392
rect 18144 3383 18196 3392
rect 18144 3349 18153 3383
rect 18153 3349 18187 3383
rect 18187 3349 18196 3383
rect 18144 3340 18196 3349
rect 4648 3238 4700 3290
rect 4712 3238 4764 3290
rect 4776 3238 4828 3290
rect 4840 3238 4892 3290
rect 11982 3238 12034 3290
rect 12046 3238 12098 3290
rect 12110 3238 12162 3290
rect 12174 3238 12226 3290
rect 19315 3238 19367 3290
rect 19379 3238 19431 3290
rect 19443 3238 19495 3290
rect 19507 3238 19559 3290
rect 2688 3136 2740 3188
rect 8208 3136 8260 3188
rect 8852 3136 8904 3188
rect 11704 3136 11756 3188
rect 13084 3179 13136 3188
rect 13084 3145 13093 3179
rect 13093 3145 13127 3179
rect 13127 3145 13136 3179
rect 13084 3136 13136 3145
rect 15476 3136 15528 3188
rect 15844 3136 15896 3188
rect 16580 3136 16632 3188
rect 17224 3179 17276 3188
rect 17224 3145 17233 3179
rect 17233 3145 17267 3179
rect 17267 3145 17276 3179
rect 17224 3136 17276 3145
rect 18972 3136 19024 3188
rect 19708 3136 19760 3188
rect 4528 3068 4580 3120
rect 1400 3000 1452 3052
rect 5264 3043 5316 3052
rect 5264 3009 5273 3043
rect 5273 3009 5307 3043
rect 5307 3009 5316 3043
rect 5264 3000 5316 3009
rect 7104 3000 7156 3052
rect 9036 3068 9088 3120
rect 1768 2975 1820 2984
rect 1768 2941 1777 2975
rect 1777 2941 1811 2975
rect 1811 2941 1820 2975
rect 1768 2932 1820 2941
rect 2044 2975 2096 2984
rect 2044 2941 2053 2975
rect 2053 2941 2087 2975
rect 2087 2941 2096 2975
rect 2044 2932 2096 2941
rect 2872 2932 2924 2984
rect 3608 2975 3660 2984
rect 3608 2941 3617 2975
rect 3617 2941 3651 2975
rect 3651 2941 3660 2975
rect 3608 2932 3660 2941
rect 2964 2796 3016 2848
rect 4988 2932 5040 2984
rect 4344 2907 4396 2916
rect 4344 2873 4353 2907
rect 4353 2873 4387 2907
rect 4387 2873 4396 2907
rect 4344 2864 4396 2873
rect 5356 2907 5408 2916
rect 5356 2873 5365 2907
rect 5365 2873 5399 2907
rect 5399 2873 5408 2907
rect 5356 2864 5408 2873
rect 4528 2796 4580 2848
rect 5264 2796 5316 2848
rect 7012 2907 7064 2916
rect 7012 2873 7021 2907
rect 7021 2873 7055 2907
rect 7055 2873 7064 2907
rect 7012 2864 7064 2873
rect 7288 2796 7340 2848
rect 9956 3043 10008 3052
rect 9956 3009 9965 3043
rect 9965 3009 9999 3043
rect 9999 3009 10008 3043
rect 9956 3000 10008 3009
rect 10876 3068 10928 3120
rect 17316 3068 17368 3120
rect 11428 2932 11480 2984
rect 12440 2975 12492 2984
rect 12440 2941 12449 2975
rect 12449 2941 12483 2975
rect 12483 2941 12492 2975
rect 12440 2932 12492 2941
rect 13084 2932 13136 2984
rect 15108 3000 15160 3052
rect 16396 3043 16448 3052
rect 16396 3009 16405 3043
rect 16405 3009 16439 3043
rect 16439 3009 16448 3043
rect 16396 3000 16448 3009
rect 16764 3000 16816 3052
rect 13912 2975 13964 2984
rect 13912 2941 13921 2975
rect 13921 2941 13955 2975
rect 13955 2941 13964 2975
rect 13912 2932 13964 2941
rect 17776 2932 17828 2984
rect 9036 2907 9088 2916
rect 9036 2873 9045 2907
rect 9045 2873 9079 2907
rect 9079 2873 9088 2907
rect 9588 2907 9640 2916
rect 9036 2864 9088 2873
rect 9588 2873 9597 2907
rect 9597 2873 9631 2907
rect 9631 2873 9640 2907
rect 9588 2864 9640 2873
rect 10324 2839 10376 2848
rect 10324 2805 10333 2839
rect 10333 2805 10367 2839
rect 10367 2805 10376 2839
rect 10324 2796 10376 2805
rect 12072 2839 12124 2848
rect 12072 2805 12081 2839
rect 12081 2805 12115 2839
rect 12115 2805 12124 2839
rect 12072 2796 12124 2805
rect 13268 2796 13320 2848
rect 13820 2864 13872 2916
rect 15844 2907 15896 2916
rect 15844 2873 15853 2907
rect 15853 2873 15887 2907
rect 15887 2873 15896 2907
rect 15844 2864 15896 2873
rect 18144 2932 18196 2984
rect 20076 2975 20128 2984
rect 20076 2941 20085 2975
rect 20085 2941 20119 2975
rect 20119 2941 20128 2975
rect 20076 2932 20128 2941
rect 19800 2864 19852 2916
rect 17776 2839 17828 2848
rect 17776 2805 17785 2839
rect 17785 2805 17819 2839
rect 17819 2805 17828 2839
rect 17776 2796 17828 2805
rect 18144 2839 18196 2848
rect 18144 2805 18153 2839
rect 18153 2805 18187 2839
rect 18187 2805 18196 2839
rect 18144 2796 18196 2805
rect 8315 2694 8367 2746
rect 8379 2694 8431 2746
rect 8443 2694 8495 2746
rect 8507 2694 8559 2746
rect 15648 2694 15700 2746
rect 15712 2694 15764 2746
rect 15776 2694 15828 2746
rect 15840 2694 15892 2746
rect 1400 2635 1452 2644
rect 1400 2601 1409 2635
rect 1409 2601 1443 2635
rect 1443 2601 1452 2635
rect 1400 2592 1452 2601
rect 3608 2635 3660 2644
rect 3608 2601 3617 2635
rect 3617 2601 3651 2635
rect 3651 2601 3660 2635
rect 3608 2592 3660 2601
rect 4344 2592 4396 2644
rect 3148 2567 3200 2576
rect 3148 2533 3157 2567
rect 3157 2533 3191 2567
rect 3191 2533 3200 2567
rect 3148 2524 3200 2533
rect 2504 2499 2556 2508
rect 2504 2465 2513 2499
rect 2513 2465 2547 2499
rect 2547 2465 2556 2499
rect 2504 2456 2556 2465
rect 2964 2499 3016 2508
rect 2964 2465 2973 2499
rect 2973 2465 3007 2499
rect 3007 2465 3016 2499
rect 2964 2456 3016 2465
rect 4896 2456 4948 2508
rect 5264 2524 5316 2576
rect 7012 2592 7064 2644
rect 7840 2635 7892 2644
rect 7840 2601 7849 2635
rect 7849 2601 7883 2635
rect 7883 2601 7892 2635
rect 7840 2592 7892 2601
rect 6736 2524 6788 2576
rect 7196 2524 7248 2576
rect 9036 2592 9088 2644
rect 10048 2635 10100 2644
rect 10048 2601 10057 2635
rect 10057 2601 10091 2635
rect 10091 2601 10100 2635
rect 10048 2592 10100 2601
rect 11612 2592 11664 2644
rect 12072 2592 12124 2644
rect 6184 2456 6236 2508
rect 7104 2456 7156 2508
rect 10324 2567 10376 2576
rect 10324 2533 10333 2567
rect 10333 2533 10367 2567
rect 10367 2533 10376 2567
rect 10324 2524 10376 2533
rect 13268 2524 13320 2576
rect 13820 2524 13872 2576
rect 13912 2524 13964 2576
rect 11796 2456 11848 2508
rect 13360 2499 13412 2508
rect 13360 2465 13369 2499
rect 13369 2465 13403 2499
rect 13403 2465 13412 2499
rect 13360 2456 13412 2465
rect 15568 2524 15620 2576
rect 17132 2592 17184 2644
rect 17776 2592 17828 2644
rect 18420 2635 18472 2644
rect 6828 2388 6880 2440
rect 17040 2456 17092 2508
rect 18420 2601 18429 2635
rect 18429 2601 18463 2635
rect 18463 2601 18472 2635
rect 18420 2592 18472 2601
rect 18788 2524 18840 2576
rect 6092 2320 6144 2372
rect 4528 2252 4580 2304
rect 4988 2252 5040 2304
rect 6368 2295 6420 2304
rect 6368 2261 6377 2295
rect 6377 2261 6411 2295
rect 6411 2261 6420 2295
rect 6368 2252 6420 2261
rect 7288 2252 7340 2304
rect 15200 2295 15252 2304
rect 15200 2261 15209 2295
rect 15209 2261 15243 2295
rect 15243 2261 15252 2295
rect 15660 2388 15712 2440
rect 15936 2388 15988 2440
rect 20076 2388 20128 2440
rect 21456 2320 21508 2372
rect 15200 2252 15252 2261
rect 4648 2150 4700 2202
rect 4712 2150 4764 2202
rect 4776 2150 4828 2202
rect 4840 2150 4892 2202
rect 11982 2150 12034 2202
rect 12046 2150 12098 2202
rect 12110 2150 12162 2202
rect 12174 2150 12226 2202
rect 19315 2150 19367 2202
rect 19379 2150 19431 2202
rect 19443 2150 19495 2202
rect 19507 2150 19559 2202
rect 9772 76 9824 128
rect 10508 76 10560 128
<< metal2 >>
rect 1766 21570 1822 22000
rect 5354 21570 5410 22000
rect 9034 21570 9090 22000
rect 12714 21570 12770 22000
rect 16394 21570 16450 22000
rect 20074 21570 20130 22000
rect 1766 21542 2084 21570
rect 1766 21520 1822 21542
rect 110 21448 166 21457
rect 110 21383 166 21392
rect 124 18290 152 21383
rect 1306 19816 1362 19825
rect 1306 19751 1362 19760
rect 112 18284 164 18290
rect 112 18226 164 18232
rect 1320 17814 1348 19751
rect 1400 18760 1452 18766
rect 1400 18702 1452 18708
rect 1582 18728 1638 18737
rect 1308 17808 1360 17814
rect 1308 17750 1360 17756
rect 202 16688 258 16697
rect 124 16646 202 16674
rect 124 16017 152 16646
rect 202 16623 258 16632
rect 110 16008 166 16017
rect 1412 15978 1440 18702
rect 1582 18663 1638 18672
rect 1596 18426 1624 18663
rect 1860 18624 1912 18630
rect 1860 18566 1912 18572
rect 1584 18420 1636 18426
rect 1584 18362 1636 18368
rect 1492 18216 1544 18222
rect 1492 18158 1544 18164
rect 1504 17610 1532 18158
rect 1872 17746 1900 18566
rect 2056 18358 2084 21542
rect 5354 21542 5488 21570
rect 5354 21520 5410 21542
rect 4622 19612 4918 19632
rect 4678 19610 4702 19612
rect 4758 19610 4782 19612
rect 4838 19610 4862 19612
rect 4700 19558 4702 19610
rect 4764 19558 4776 19610
rect 4838 19558 4840 19610
rect 4678 19556 4702 19558
rect 4758 19556 4782 19558
rect 4838 19556 4862 19558
rect 4622 19536 4918 19556
rect 4252 19508 4304 19514
rect 4252 19450 4304 19456
rect 4160 19372 4212 19378
rect 4160 19314 4212 19320
rect 2136 19304 2188 19310
rect 4068 19304 4120 19310
rect 2136 19246 2188 19252
rect 3422 19272 3478 19281
rect 2044 18352 2096 18358
rect 2044 18294 2096 18300
rect 1860 17740 1912 17746
rect 1860 17682 1912 17688
rect 1582 17640 1638 17649
rect 1492 17604 1544 17610
rect 1582 17575 1638 17584
rect 1492 17546 1544 17552
rect 1596 17338 1624 17575
rect 1584 17332 1636 17338
rect 1584 17274 1636 17280
rect 1872 16794 1900 17682
rect 1860 16788 1912 16794
rect 1860 16730 1912 16736
rect 1872 16114 1900 16730
rect 1860 16108 1912 16114
rect 1860 16050 1912 16056
rect 110 15943 166 15952
rect 1400 15972 1452 15978
rect 1400 15914 1452 15920
rect 1676 15700 1728 15706
rect 1676 15642 1728 15648
rect 110 14920 166 14929
rect 110 14855 166 14864
rect 124 12782 152 14855
rect 1688 14822 1716 15642
rect 2042 15056 2098 15065
rect 2042 14991 2098 15000
rect 1676 14816 1728 14822
rect 1676 14758 1728 14764
rect 1688 14618 1716 14758
rect 1676 14612 1728 14618
rect 1728 14572 1808 14600
rect 1676 14554 1728 14560
rect 1676 14408 1728 14414
rect 1676 14350 1728 14356
rect 1688 13530 1716 14350
rect 1780 13734 1808 14572
rect 1768 13728 1820 13734
rect 1768 13670 1820 13676
rect 1676 13524 1728 13530
rect 1676 13466 1728 13472
rect 1308 13388 1360 13394
rect 1308 13330 1360 13336
rect 1768 13388 1820 13394
rect 1768 13330 1820 13336
rect 112 12776 164 12782
rect 112 12718 164 12724
rect 20 12640 72 12646
rect 20 12582 72 12588
rect 32 10441 60 12582
rect 112 11892 164 11898
rect 112 11834 164 11840
rect 124 11665 152 11834
rect 110 11656 166 11665
rect 110 11591 166 11600
rect 112 11008 164 11014
rect 112 10950 164 10956
rect 18 10432 74 10441
rect 18 10367 74 10376
rect 124 5001 152 10950
rect 1320 6633 1348 13330
rect 1676 12300 1728 12306
rect 1676 12242 1728 12248
rect 1688 11694 1716 12242
rect 1676 11688 1728 11694
rect 1676 11630 1728 11636
rect 1584 10464 1636 10470
rect 1584 10406 1636 10412
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1412 8838 1440 9998
rect 1596 9518 1624 10406
rect 1584 9512 1636 9518
rect 1584 9454 1636 9460
rect 1584 9172 1636 9178
rect 1584 9114 1636 9120
rect 1400 8832 1452 8838
rect 1400 8774 1452 8780
rect 1412 7002 1440 8774
rect 1596 7954 1624 9114
rect 1780 9042 1808 13330
rect 1952 12640 2004 12646
rect 1952 12582 2004 12588
rect 1860 9376 1912 9382
rect 1860 9318 1912 9324
rect 1768 9036 1820 9042
rect 1768 8978 1820 8984
rect 1780 8634 1808 8978
rect 1768 8628 1820 8634
rect 1768 8570 1820 8576
rect 1872 8022 1900 9318
rect 1964 8673 1992 12582
rect 1950 8664 2006 8673
rect 1950 8599 2006 8608
rect 1952 8356 2004 8362
rect 1952 8298 2004 8304
rect 1964 8022 1992 8298
rect 1860 8016 1912 8022
rect 1860 7958 1912 7964
rect 1952 8016 2004 8022
rect 1952 7958 2004 7964
rect 1584 7948 1636 7954
rect 1584 7890 1636 7896
rect 1596 7002 1624 7890
rect 1400 6996 1452 7002
rect 1400 6938 1452 6944
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 1872 6662 1900 7958
rect 1860 6656 1912 6662
rect 1306 6624 1362 6633
rect 1860 6598 1912 6604
rect 1306 6559 1362 6568
rect 848 6452 900 6458
rect 848 6394 900 6400
rect 110 4992 166 5001
rect 110 4927 166 4936
rect 570 82 626 480
rect 860 82 888 6394
rect 1872 5846 1900 6598
rect 1860 5840 1912 5846
rect 1860 5782 1912 5788
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1412 5370 1440 5646
rect 1400 5364 1452 5370
rect 1400 5306 1452 5312
rect 1768 4548 1820 4554
rect 1768 4490 1820 4496
rect 1780 4282 1808 4490
rect 1872 4486 1900 5782
rect 1860 4480 1912 4486
rect 1860 4422 1912 4428
rect 1768 4276 1820 4282
rect 1768 4218 1820 4224
rect 1768 3460 1820 3466
rect 1768 3402 1820 3408
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 1412 2650 1440 2994
rect 1780 2990 1808 3402
rect 1768 2984 1820 2990
rect 1768 2926 1820 2932
rect 1400 2644 1452 2650
rect 1400 2586 1452 2592
rect 570 54 888 82
rect 1674 82 1730 480
rect 1872 82 1900 4422
rect 2056 4154 2084 14991
rect 2148 14550 2176 19246
rect 2320 19236 2372 19242
rect 4172 19281 4200 19314
rect 4068 19246 4120 19252
rect 4158 19272 4214 19281
rect 3422 19207 3478 19216
rect 2320 19178 2372 19184
rect 2332 18834 2360 19178
rect 3436 19174 3464 19207
rect 4080 19174 4108 19246
rect 4158 19207 4214 19216
rect 2596 19168 2648 19174
rect 2596 19110 2648 19116
rect 2872 19168 2924 19174
rect 2872 19110 2924 19116
rect 3424 19168 3476 19174
rect 3424 19110 3476 19116
rect 4068 19168 4120 19174
rect 4068 19110 4120 19116
rect 2320 18828 2372 18834
rect 2320 18770 2372 18776
rect 2332 18086 2360 18770
rect 2320 18080 2372 18086
rect 2320 18022 2372 18028
rect 2332 17678 2360 18022
rect 2412 17740 2464 17746
rect 2412 17682 2464 17688
rect 2320 17672 2372 17678
rect 2320 17614 2372 17620
rect 2332 16998 2360 17614
rect 2320 16992 2372 16998
rect 2320 16934 2372 16940
rect 2228 16720 2280 16726
rect 2228 16662 2280 16668
rect 2240 16114 2268 16662
rect 2228 16108 2280 16114
rect 2228 16050 2280 16056
rect 2240 15706 2268 16050
rect 2228 15700 2280 15706
rect 2228 15642 2280 15648
rect 2136 14544 2188 14550
rect 2136 14486 2188 14492
rect 2148 14074 2176 14486
rect 2136 14068 2188 14074
rect 2136 14010 2188 14016
rect 2332 13814 2360 16934
rect 2424 16454 2452 17682
rect 2412 16448 2464 16454
rect 2412 16390 2464 16396
rect 2608 15638 2636 19110
rect 2688 18352 2740 18358
rect 2688 18294 2740 18300
rect 2596 15632 2648 15638
rect 2596 15574 2648 15580
rect 2608 14890 2636 15574
rect 2596 14884 2648 14890
rect 2596 14826 2648 14832
rect 2502 14376 2558 14385
rect 2502 14311 2558 14320
rect 2332 13786 2452 13814
rect 2320 13524 2372 13530
rect 2320 13466 2372 13472
rect 2226 13424 2282 13433
rect 2226 13359 2282 13368
rect 2136 12300 2188 12306
rect 2136 12242 2188 12248
rect 2148 11694 2176 12242
rect 2136 11688 2188 11694
rect 2136 11630 2188 11636
rect 2148 11529 2176 11630
rect 2134 11520 2190 11529
rect 2134 11455 2190 11464
rect 2148 10266 2176 11455
rect 2136 10260 2188 10266
rect 2136 10202 2188 10208
rect 2240 7721 2268 13359
rect 2332 12782 2360 13466
rect 2320 12776 2372 12782
rect 2320 12718 2372 12724
rect 2424 12714 2452 13786
rect 2412 12708 2464 12714
rect 2412 12650 2464 12656
rect 2412 12300 2464 12306
rect 2412 12242 2464 12248
rect 2424 11694 2452 12242
rect 2412 11688 2464 11694
rect 2412 11630 2464 11636
rect 2320 10192 2372 10198
rect 2320 10134 2372 10140
rect 2332 9722 2360 10134
rect 2320 9716 2372 9722
rect 2320 9658 2372 9664
rect 2332 9178 2360 9658
rect 2320 9172 2372 9178
rect 2320 9114 2372 9120
rect 2412 8492 2464 8498
rect 2412 8434 2464 8440
rect 2320 8356 2372 8362
rect 2320 8298 2372 8304
rect 2332 7750 2360 8298
rect 2320 7744 2372 7750
rect 2226 7712 2282 7721
rect 2320 7686 2372 7692
rect 2226 7647 2282 7656
rect 2136 7472 2188 7478
rect 2136 7414 2188 7420
rect 2148 7274 2176 7414
rect 2136 7268 2188 7274
rect 2136 7210 2188 7216
rect 2148 5302 2176 7210
rect 2332 7206 2360 7686
rect 2320 7200 2372 7206
rect 2320 7142 2372 7148
rect 2424 6390 2452 8434
rect 2412 6384 2464 6390
rect 2412 6326 2464 6332
rect 2320 6112 2372 6118
rect 2320 6054 2372 6060
rect 2332 5914 2360 6054
rect 2424 5914 2452 6326
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 2412 5908 2464 5914
rect 2412 5850 2464 5856
rect 2136 5296 2188 5302
rect 2136 5238 2188 5244
rect 2148 4826 2176 5238
rect 2228 5092 2280 5098
rect 2332 5080 2360 5850
rect 2516 5846 2544 14311
rect 2596 14000 2648 14006
rect 2596 13942 2648 13948
rect 2608 13870 2636 13942
rect 2596 13864 2648 13870
rect 2596 13806 2648 13812
rect 2608 13394 2636 13806
rect 2596 13388 2648 13394
rect 2596 13330 2648 13336
rect 2596 13184 2648 13190
rect 2596 13126 2648 13132
rect 2608 10538 2636 13126
rect 2700 12986 2728 18294
rect 2884 18222 2912 19110
rect 3148 18760 3200 18766
rect 3148 18702 3200 18708
rect 3160 18426 3188 18702
rect 3148 18420 3200 18426
rect 3148 18362 3200 18368
rect 4080 18222 4108 19110
rect 4264 18816 4292 19450
rect 5460 19378 5488 21542
rect 8680 21542 9090 21570
rect 6736 19440 6788 19446
rect 6736 19382 6788 19388
rect 5448 19372 5500 19378
rect 5448 19314 5500 19320
rect 4344 19304 4396 19310
rect 4344 19246 4396 19252
rect 4988 19304 5040 19310
rect 4988 19246 5040 19252
rect 4356 18834 4384 19246
rect 4172 18788 4292 18816
rect 4344 18828 4396 18834
rect 2872 18216 2924 18222
rect 2872 18158 2924 18164
rect 3608 18216 3660 18222
rect 3608 18158 3660 18164
rect 4068 18216 4120 18222
rect 4068 18158 4120 18164
rect 2778 17232 2834 17241
rect 2778 17167 2834 17176
rect 2792 17134 2820 17167
rect 2780 17128 2832 17134
rect 2780 17070 2832 17076
rect 2792 16522 2820 17070
rect 2780 16516 2832 16522
rect 2780 16458 2832 16464
rect 2884 16402 2912 18158
rect 3240 17060 3292 17066
rect 3240 17002 3292 17008
rect 3056 16584 3108 16590
rect 3056 16526 3108 16532
rect 2792 16374 2912 16402
rect 2688 12980 2740 12986
rect 2688 12922 2740 12928
rect 2700 12782 2728 12922
rect 2792 12918 2820 16374
rect 2872 15496 2924 15502
rect 2872 15438 2924 15444
rect 2780 12912 2832 12918
rect 2780 12854 2832 12860
rect 2688 12776 2740 12782
rect 2688 12718 2740 12724
rect 2700 11694 2728 12718
rect 2792 12442 2820 12854
rect 2780 12436 2832 12442
rect 2780 12378 2832 12384
rect 2884 12374 2912 15438
rect 2964 15360 3016 15366
rect 2964 15302 3016 15308
rect 2976 15026 3004 15302
rect 3068 15094 3096 16526
rect 3148 16516 3200 16522
rect 3148 16458 3200 16464
rect 3056 15088 3108 15094
rect 3056 15030 3108 15036
rect 2964 15020 3016 15026
rect 2964 14962 3016 14968
rect 2964 14612 3016 14618
rect 2964 14554 3016 14560
rect 2976 13190 3004 14554
rect 3068 14550 3096 15030
rect 3056 14544 3108 14550
rect 3056 14486 3108 14492
rect 3056 14272 3108 14278
rect 3056 14214 3108 14220
rect 3068 13938 3096 14214
rect 3056 13932 3108 13938
rect 3056 13874 3108 13880
rect 2964 13184 3016 13190
rect 2964 13126 3016 13132
rect 2964 12776 3016 12782
rect 2964 12718 3016 12724
rect 2872 12368 2924 12374
rect 2872 12310 2924 12316
rect 2688 11688 2740 11694
rect 2688 11630 2740 11636
rect 2700 11354 2728 11630
rect 2688 11348 2740 11354
rect 2688 11290 2740 11296
rect 2872 11212 2924 11218
rect 2872 11154 2924 11160
rect 2596 10532 2648 10538
rect 2596 10474 2648 10480
rect 2608 10130 2636 10474
rect 2596 10124 2648 10130
rect 2596 10066 2648 10072
rect 2504 5840 2556 5846
rect 2504 5782 2556 5788
rect 2516 5234 2544 5782
rect 2504 5228 2556 5234
rect 2504 5170 2556 5176
rect 2280 5052 2360 5080
rect 2228 5034 2280 5040
rect 2608 4978 2636 10066
rect 2884 9722 2912 11154
rect 2872 9716 2924 9722
rect 2872 9658 2924 9664
rect 2884 9042 2912 9658
rect 2872 9036 2924 9042
rect 2872 8978 2924 8984
rect 2884 8634 2912 8978
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2688 6860 2740 6866
rect 2688 6802 2740 6808
rect 2700 6254 2728 6802
rect 2792 6662 2820 7142
rect 2884 6866 2912 8570
rect 2872 6860 2924 6866
rect 2872 6802 2924 6808
rect 2884 6730 2912 6802
rect 2872 6724 2924 6730
rect 2872 6666 2924 6672
rect 2780 6656 2832 6662
rect 2780 6598 2832 6604
rect 2688 6248 2740 6254
rect 2688 6190 2740 6196
rect 2424 4950 2636 4978
rect 2136 4820 2188 4826
rect 2136 4762 2188 4768
rect 2424 4282 2452 4950
rect 2700 4842 2728 6190
rect 2792 5302 2820 6598
rect 2884 6458 2912 6666
rect 2872 6452 2924 6458
rect 2872 6394 2924 6400
rect 2872 5364 2924 5370
rect 2872 5306 2924 5312
rect 2780 5296 2832 5302
rect 2780 5238 2832 5244
rect 2516 4814 2728 4842
rect 2412 4276 2464 4282
rect 2412 4218 2464 4224
rect 1964 4126 2084 4154
rect 1964 3369 1992 4126
rect 2044 3664 2096 3670
rect 2044 3606 2096 3612
rect 1950 3360 2006 3369
rect 1950 3295 2006 3304
rect 2056 2990 2084 3606
rect 2044 2984 2096 2990
rect 2044 2926 2096 2932
rect 2516 2514 2544 4814
rect 2688 4684 2740 4690
rect 2688 4626 2740 4632
rect 2700 4282 2728 4626
rect 2780 4548 2832 4554
rect 2780 4490 2832 4496
rect 2688 4276 2740 4282
rect 2688 4218 2740 4224
rect 2700 3602 2728 4218
rect 2792 4078 2820 4490
rect 2780 4072 2832 4078
rect 2780 4014 2832 4020
rect 2792 3670 2820 4014
rect 2780 3664 2832 3670
rect 2780 3606 2832 3612
rect 2688 3596 2740 3602
rect 2688 3538 2740 3544
rect 2700 3194 2728 3538
rect 2688 3188 2740 3194
rect 2688 3130 2740 3136
rect 2884 2990 2912 5306
rect 2976 4154 3004 12718
rect 3068 11762 3096 13874
rect 3160 12714 3188 16458
rect 3148 12708 3200 12714
rect 3148 12650 3200 12656
rect 3056 11756 3108 11762
rect 3056 11698 3108 11704
rect 3056 11144 3108 11150
rect 3056 11086 3108 11092
rect 3068 8090 3096 11086
rect 3252 10674 3280 17002
rect 3332 16992 3384 16998
rect 3332 16934 3384 16940
rect 3344 14940 3372 16934
rect 3620 16454 3648 18158
rect 3976 17740 4028 17746
rect 3976 17682 4028 17688
rect 3884 17536 3936 17542
rect 3884 17478 3936 17484
rect 3608 16448 3660 16454
rect 3608 16390 3660 16396
rect 3424 15496 3476 15502
rect 3424 15438 3476 15444
rect 3436 15094 3464 15438
rect 3424 15088 3476 15094
rect 3424 15030 3476 15036
rect 3516 14952 3568 14958
rect 3344 14912 3464 14940
rect 3332 14544 3384 14550
rect 3332 14486 3384 14492
rect 3344 12442 3372 14486
rect 3436 13734 3464 14912
rect 3516 14894 3568 14900
rect 3424 13728 3476 13734
rect 3424 13670 3476 13676
rect 3528 13530 3556 14894
rect 3620 14550 3648 16390
rect 3792 15428 3844 15434
rect 3792 15370 3844 15376
rect 3700 14816 3752 14822
rect 3700 14758 3752 14764
rect 3608 14544 3660 14550
rect 3608 14486 3660 14492
rect 3712 14006 3740 14758
rect 3700 14000 3752 14006
rect 3700 13942 3752 13948
rect 3700 13864 3752 13870
rect 3700 13806 3752 13812
rect 3608 13728 3660 13734
rect 3608 13670 3660 13676
rect 3516 13524 3568 13530
rect 3516 13466 3568 13472
rect 3516 12708 3568 12714
rect 3516 12650 3568 12656
rect 3332 12436 3384 12442
rect 3332 12378 3384 12384
rect 3528 12306 3556 12650
rect 3516 12300 3568 12306
rect 3516 12242 3568 12248
rect 3424 11756 3476 11762
rect 3424 11698 3476 11704
rect 3332 11688 3384 11694
rect 3332 11630 3384 11636
rect 3240 10668 3292 10674
rect 3240 10610 3292 10616
rect 3252 10266 3280 10610
rect 3240 10260 3292 10266
rect 3240 10202 3292 10208
rect 3240 9512 3292 9518
rect 3240 9454 3292 9460
rect 3252 9178 3280 9454
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 3344 8090 3372 11630
rect 3436 11626 3464 11698
rect 3424 11620 3476 11626
rect 3424 11562 3476 11568
rect 3436 11354 3464 11562
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 3528 11286 3556 12242
rect 3516 11280 3568 11286
rect 3516 11222 3568 11228
rect 3528 9926 3556 11222
rect 3620 10742 3648 13670
rect 3712 13530 3740 13806
rect 3700 13524 3752 13530
rect 3700 13466 3752 13472
rect 3804 13394 3832 15370
rect 3792 13388 3844 13394
rect 3792 13330 3844 13336
rect 3804 12986 3832 13330
rect 3792 12980 3844 12986
rect 3792 12922 3844 12928
rect 3804 12714 3832 12922
rect 3792 12708 3844 12714
rect 3792 12650 3844 12656
rect 3896 11694 3924 17478
rect 3988 17202 4016 17682
rect 4068 17604 4120 17610
rect 4068 17546 4120 17552
rect 3976 17196 4028 17202
rect 3976 17138 4028 17144
rect 3988 16998 4016 17138
rect 3976 16992 4028 16998
rect 3976 16934 4028 16940
rect 3976 15564 4028 15570
rect 3976 15506 4028 15512
rect 3988 14822 4016 15506
rect 3976 14816 4028 14822
rect 3976 14758 4028 14764
rect 3988 13433 4016 14758
rect 3974 13424 4030 13433
rect 4080 13394 4108 17546
rect 3974 13359 4030 13368
rect 4068 13388 4120 13394
rect 4068 13330 4120 13336
rect 4080 12646 4108 13330
rect 4068 12640 4120 12646
rect 4068 12582 4120 12588
rect 3884 11688 3936 11694
rect 3884 11630 3936 11636
rect 4068 11620 4120 11626
rect 4068 11562 4120 11568
rect 3700 11552 3752 11558
rect 3700 11494 3752 11500
rect 3882 11520 3938 11529
rect 3712 11014 3740 11494
rect 3882 11455 3938 11464
rect 3896 11354 3924 11455
rect 4080 11354 4108 11562
rect 3884 11348 3936 11354
rect 3884 11290 3936 11296
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 4172 11234 4200 18788
rect 4344 18770 4396 18776
rect 4252 18692 4304 18698
rect 4252 18634 4304 18640
rect 4264 18154 4292 18634
rect 4252 18148 4304 18154
rect 4252 18090 4304 18096
rect 4264 17814 4292 18090
rect 4356 17882 4384 18770
rect 4622 18524 4918 18544
rect 4678 18522 4702 18524
rect 4758 18522 4782 18524
rect 4838 18522 4862 18524
rect 4700 18470 4702 18522
rect 4764 18470 4776 18522
rect 4838 18470 4840 18522
rect 4678 18468 4702 18470
rect 4758 18468 4782 18470
rect 4838 18468 4862 18470
rect 4622 18448 4918 18468
rect 4712 18352 4764 18358
rect 4712 18294 4764 18300
rect 4724 18222 4752 18294
rect 4712 18216 4764 18222
rect 4712 18158 4764 18164
rect 4344 17876 4396 17882
rect 4344 17818 4396 17824
rect 4252 17808 4304 17814
rect 4252 17750 4304 17756
rect 5000 17746 5028 19246
rect 5172 19168 5224 19174
rect 5172 19110 5224 19116
rect 5080 18760 5132 18766
rect 5080 18702 5132 18708
rect 4988 17740 5040 17746
rect 4988 17682 5040 17688
rect 4436 17672 4488 17678
rect 5092 17626 5120 18702
rect 4436 17614 4488 17620
rect 4250 16552 4306 16561
rect 4250 16487 4306 16496
rect 4264 15706 4292 16487
rect 4448 16046 4476 17614
rect 5000 17598 5120 17626
rect 4622 17436 4918 17456
rect 4678 17434 4702 17436
rect 4758 17434 4782 17436
rect 4838 17434 4862 17436
rect 4700 17382 4702 17434
rect 4764 17382 4776 17434
rect 4838 17382 4840 17434
rect 4678 17380 4702 17382
rect 4758 17380 4782 17382
rect 4838 17380 4862 17382
rect 4622 17360 4918 17380
rect 5000 16658 5028 17598
rect 5080 17196 5132 17202
rect 5080 17138 5132 17144
rect 4988 16652 5040 16658
rect 4988 16594 5040 16600
rect 5000 16561 5028 16594
rect 4986 16552 5042 16561
rect 4986 16487 5042 16496
rect 4622 16348 4918 16368
rect 4678 16346 4702 16348
rect 4758 16346 4782 16348
rect 4838 16346 4862 16348
rect 4700 16294 4702 16346
rect 4764 16294 4776 16346
rect 4838 16294 4840 16346
rect 4678 16292 4702 16294
rect 4758 16292 4782 16294
rect 4838 16292 4862 16294
rect 4622 16272 4918 16292
rect 4436 16040 4488 16046
rect 4436 15982 4488 15988
rect 4252 15700 4304 15706
rect 4252 15642 4304 15648
rect 4448 14618 4476 15982
rect 5000 15706 5028 16487
rect 4988 15700 5040 15706
rect 4988 15642 5040 15648
rect 4622 15260 4918 15280
rect 4678 15258 4702 15260
rect 4758 15258 4782 15260
rect 4838 15258 4862 15260
rect 4700 15206 4702 15258
rect 4764 15206 4776 15258
rect 4838 15206 4840 15258
rect 4678 15204 4702 15206
rect 4758 15204 4782 15206
rect 4838 15204 4862 15206
rect 4622 15184 4918 15204
rect 4436 14612 4488 14618
rect 4436 14554 4488 14560
rect 4528 14408 4580 14414
rect 4528 14350 4580 14356
rect 4344 13796 4396 13802
rect 4344 13738 4396 13744
rect 4252 12640 4304 12646
rect 4252 12582 4304 12588
rect 4264 11626 4292 12582
rect 4252 11620 4304 11626
rect 4252 11562 4304 11568
rect 4264 11286 4292 11562
rect 3896 11206 4200 11234
rect 4252 11280 4304 11286
rect 4252 11222 4304 11228
rect 3700 11008 3752 11014
rect 3700 10950 3752 10956
rect 3608 10736 3660 10742
rect 3608 10678 3660 10684
rect 3516 9920 3568 9926
rect 3516 9862 3568 9868
rect 3712 9042 3740 10950
rect 3792 10532 3844 10538
rect 3792 10474 3844 10480
rect 3804 9586 3832 10474
rect 3792 9580 3844 9586
rect 3792 9522 3844 9528
rect 3804 9178 3832 9522
rect 3792 9172 3844 9178
rect 3792 9114 3844 9120
rect 3700 9036 3752 9042
rect 3700 8978 3752 8984
rect 3056 8084 3108 8090
rect 3056 8026 3108 8032
rect 3332 8084 3384 8090
rect 3332 8026 3384 8032
rect 3068 7410 3096 8026
rect 3344 7546 3372 8026
rect 3332 7540 3384 7546
rect 3332 7482 3384 7488
rect 3056 7404 3108 7410
rect 3056 7346 3108 7352
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 3056 6316 3108 6322
rect 3056 6258 3108 6264
rect 3068 5778 3096 6258
rect 3160 5778 3188 6734
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 3056 5772 3108 5778
rect 3056 5714 3108 5720
rect 3148 5772 3200 5778
rect 3148 5714 3200 5720
rect 3068 5681 3096 5714
rect 3054 5672 3110 5681
rect 3054 5607 3110 5616
rect 3148 5160 3200 5166
rect 3148 5102 3200 5108
rect 3160 4690 3188 5102
rect 3148 4684 3200 4690
rect 3148 4626 3200 4632
rect 3252 4554 3280 6394
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 3436 5914 3464 6258
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 3700 5840 3752 5846
rect 3700 5782 3752 5788
rect 3712 5302 3740 5782
rect 3792 5568 3844 5574
rect 3792 5510 3844 5516
rect 3700 5296 3752 5302
rect 3700 5238 3752 5244
rect 3712 5098 3740 5238
rect 3804 5166 3832 5510
rect 3792 5160 3844 5166
rect 3792 5102 3844 5108
rect 3700 5092 3752 5098
rect 3700 5034 3752 5040
rect 3712 4758 3740 5034
rect 3700 4752 3752 4758
rect 3700 4694 3752 4700
rect 3240 4548 3292 4554
rect 3240 4490 3292 4496
rect 3712 4154 3740 4694
rect 2976 4126 3096 4154
rect 2964 3596 3016 3602
rect 2964 3538 3016 3544
rect 2872 2984 2924 2990
rect 2872 2926 2924 2932
rect 2976 2854 3004 3538
rect 2964 2848 3016 2854
rect 2964 2790 3016 2796
rect 2976 2514 3004 2790
rect 2504 2508 2556 2514
rect 2504 2450 2556 2456
rect 2964 2508 3016 2514
rect 2964 2450 3016 2456
rect 1674 54 1900 82
rect 2870 82 2926 480
rect 3068 82 3096 4126
rect 3516 4140 3568 4146
rect 3712 4126 3832 4154
rect 3516 4082 3568 4088
rect 3424 4004 3476 4010
rect 3424 3946 3476 3952
rect 3436 3670 3464 3946
rect 3424 3664 3476 3670
rect 3424 3606 3476 3612
rect 3332 3528 3384 3534
rect 3384 3505 3464 3516
rect 3384 3496 3478 3505
rect 3384 3488 3422 3496
rect 3332 3470 3384 3476
rect 3422 3431 3478 3440
rect 3528 2972 3556 4082
rect 3608 3936 3660 3942
rect 3608 3878 3660 3884
rect 3620 3738 3648 3878
rect 3608 3732 3660 3738
rect 3608 3674 3660 3680
rect 3804 3670 3832 4126
rect 3792 3664 3844 3670
rect 3792 3606 3844 3612
rect 3608 2984 3660 2990
rect 3528 2944 3608 2972
rect 3608 2926 3660 2932
rect 3146 2680 3202 2689
rect 3620 2650 3648 2926
rect 3146 2615 3202 2624
rect 3608 2644 3660 2650
rect 3160 2582 3188 2615
rect 3608 2586 3660 2592
rect 3148 2576 3200 2582
rect 3148 2518 3200 2524
rect 2870 54 3096 82
rect 3896 82 3924 11206
rect 4068 11076 4120 11082
rect 4068 11018 4120 11024
rect 4080 9926 4108 11018
rect 4264 10810 4292 11222
rect 4356 11150 4384 13738
rect 4540 13462 4568 14350
rect 4622 14172 4918 14192
rect 4678 14170 4702 14172
rect 4758 14170 4782 14172
rect 4838 14170 4862 14172
rect 4700 14118 4702 14170
rect 4764 14118 4776 14170
rect 4838 14118 4840 14170
rect 4678 14116 4702 14118
rect 4758 14116 4782 14118
rect 4838 14116 4862 14118
rect 4622 14096 4918 14116
rect 4528 13456 4580 13462
rect 4528 13398 4580 13404
rect 4622 13084 4918 13104
rect 4678 13082 4702 13084
rect 4758 13082 4782 13084
rect 4838 13082 4862 13084
rect 4700 13030 4702 13082
rect 4764 13030 4776 13082
rect 4838 13030 4840 13082
rect 4678 13028 4702 13030
rect 4758 13028 4782 13030
rect 4838 13028 4862 13030
rect 4622 13008 4918 13028
rect 4436 12300 4488 12306
rect 4436 12242 4488 12248
rect 4448 11898 4476 12242
rect 4622 11996 4918 12016
rect 4678 11994 4702 11996
rect 4758 11994 4782 11996
rect 4838 11994 4862 11996
rect 4700 11942 4702 11994
rect 4764 11942 4776 11994
rect 4838 11942 4840 11994
rect 4678 11940 4702 11942
rect 4758 11940 4782 11942
rect 4838 11940 4862 11942
rect 4622 11920 4918 11940
rect 4436 11892 4488 11898
rect 4436 11834 4488 11840
rect 4804 11756 4856 11762
rect 4804 11698 4856 11704
rect 4434 11520 4490 11529
rect 4434 11455 4490 11464
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 4448 10996 4476 11455
rect 4816 11218 4844 11698
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 4528 11076 4580 11082
rect 4528 11018 4580 11024
rect 4356 10968 4476 10996
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 4264 10266 4292 10746
rect 4252 10260 4304 10266
rect 4252 10202 4304 10208
rect 4068 9920 4120 9926
rect 4068 9862 4120 9868
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 4080 8634 4108 8910
rect 4250 8800 4306 8809
rect 4250 8735 4306 8744
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 4068 8288 4120 8294
rect 4068 8230 4120 8236
rect 4160 8288 4212 8294
rect 4160 8230 4212 8236
rect 4080 7274 4108 8230
rect 4172 7954 4200 8230
rect 4264 8090 4292 8735
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4356 7970 4384 10968
rect 4540 10282 4568 11018
rect 4622 10908 4918 10928
rect 4678 10906 4702 10908
rect 4758 10906 4782 10908
rect 4838 10906 4862 10908
rect 4700 10854 4702 10906
rect 4764 10854 4776 10906
rect 4838 10854 4840 10906
rect 4678 10852 4702 10854
rect 4758 10852 4782 10854
rect 4838 10852 4862 10854
rect 4622 10832 4918 10852
rect 5000 10606 5028 15642
rect 5092 13326 5120 17138
rect 5080 13320 5132 13326
rect 5080 13262 5132 13268
rect 5080 12708 5132 12714
rect 5080 12650 5132 12656
rect 5092 12306 5120 12650
rect 5080 12300 5132 12306
rect 5080 12242 5132 12248
rect 5092 11558 5120 12242
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 4988 10600 5040 10606
rect 4988 10542 5040 10548
rect 4540 10254 4660 10282
rect 4528 10192 4580 10198
rect 4528 10134 4580 10140
rect 4540 9722 4568 10134
rect 4632 10062 4660 10254
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 4988 9988 5040 9994
rect 4988 9930 5040 9936
rect 4622 9820 4918 9840
rect 4678 9818 4702 9820
rect 4758 9818 4782 9820
rect 4838 9818 4862 9820
rect 4700 9766 4702 9818
rect 4764 9766 4776 9818
rect 4838 9766 4840 9818
rect 4678 9764 4702 9766
rect 4758 9764 4782 9766
rect 4838 9764 4862 9766
rect 4622 9744 4918 9764
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 4436 9444 4488 9450
rect 4436 9386 4488 9392
rect 4448 9178 4476 9386
rect 4436 9172 4488 9178
rect 4436 9114 4488 9120
rect 4528 8832 4580 8838
rect 4528 8774 4580 8780
rect 4540 8498 4568 8774
rect 4622 8732 4918 8752
rect 4678 8730 4702 8732
rect 4758 8730 4782 8732
rect 4838 8730 4862 8732
rect 4700 8678 4702 8730
rect 4764 8678 4776 8730
rect 4838 8678 4840 8730
rect 4678 8676 4702 8678
rect 4758 8676 4782 8678
rect 4838 8676 4862 8678
rect 4622 8656 4918 8676
rect 5000 8566 5028 9930
rect 4988 8560 5040 8566
rect 5092 8537 5120 11494
rect 4988 8502 5040 8508
rect 5078 8528 5134 8537
rect 4528 8492 4580 8498
rect 5078 8463 5134 8472
rect 4528 8434 4580 8440
rect 4540 8362 4568 8434
rect 4436 8356 4488 8362
rect 4436 8298 4488 8304
rect 4528 8356 4580 8362
rect 4528 8298 4580 8304
rect 4448 8090 4476 8298
rect 4436 8084 4488 8090
rect 4436 8026 4488 8032
rect 4160 7948 4212 7954
rect 4356 7942 4476 7970
rect 4160 7890 4212 7896
rect 4172 7546 4200 7890
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 4252 7336 4304 7342
rect 4252 7278 4304 7284
rect 4068 7268 4120 7274
rect 4068 7210 4120 7216
rect 4264 6934 4292 7278
rect 4252 6928 4304 6934
rect 4252 6870 4304 6876
rect 4264 6458 4292 6870
rect 4344 6724 4396 6730
rect 4344 6666 4396 6672
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 4356 6322 4384 6666
rect 4448 6662 4476 7942
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 4622 7644 4918 7664
rect 4678 7642 4702 7644
rect 4758 7642 4782 7644
rect 4838 7642 4862 7644
rect 4700 7590 4702 7642
rect 4764 7590 4776 7642
rect 4838 7590 4840 7642
rect 4678 7588 4702 7590
rect 4758 7588 4782 7590
rect 4838 7588 4862 7590
rect 4622 7568 4918 7588
rect 5000 7410 5028 7822
rect 4988 7404 5040 7410
rect 4988 7346 5040 7352
rect 4436 6656 4488 6662
rect 4436 6598 4488 6604
rect 4622 6556 4918 6576
rect 4678 6554 4702 6556
rect 4758 6554 4782 6556
rect 4838 6554 4862 6556
rect 4700 6502 4702 6554
rect 4764 6502 4776 6554
rect 4838 6502 4840 6554
rect 4678 6500 4702 6502
rect 4758 6500 4782 6502
rect 4838 6500 4862 6502
rect 4622 6480 4918 6500
rect 4344 6316 4396 6322
rect 4344 6258 4396 6264
rect 4988 6316 5040 6322
rect 4988 6258 5040 6264
rect 3976 6248 4028 6254
rect 3976 6190 4028 6196
rect 3988 5642 4016 6190
rect 4252 6180 4304 6186
rect 4252 6122 4304 6128
rect 4264 5914 4292 6122
rect 4252 5908 4304 5914
rect 4252 5850 4304 5856
rect 4068 5772 4120 5778
rect 4068 5714 4120 5720
rect 3976 5636 4028 5642
rect 3976 5578 4028 5584
rect 4080 5370 4108 5714
rect 4622 5468 4918 5488
rect 4678 5466 4702 5468
rect 4758 5466 4782 5468
rect 4838 5466 4862 5468
rect 4700 5414 4702 5466
rect 4764 5414 4776 5466
rect 4838 5414 4840 5466
rect 4678 5412 4702 5414
rect 4758 5412 4782 5414
rect 4838 5412 4862 5414
rect 4622 5392 4918 5412
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4724 4758 4752 4966
rect 5000 4758 5028 6258
rect 4528 4752 4580 4758
rect 4528 4694 4580 4700
rect 4712 4752 4764 4758
rect 4712 4694 4764 4700
rect 4988 4752 5040 4758
rect 4988 4694 5040 4700
rect 4540 4282 4568 4694
rect 4622 4380 4918 4400
rect 4678 4378 4702 4380
rect 4758 4378 4782 4380
rect 4838 4378 4862 4380
rect 4700 4326 4702 4378
rect 4764 4326 4776 4378
rect 4838 4326 4840 4378
rect 4678 4324 4702 4326
rect 4758 4324 4782 4326
rect 4838 4324 4862 4326
rect 4622 4304 4918 4324
rect 4528 4276 4580 4282
rect 4528 4218 4580 4224
rect 5000 4146 5028 4694
rect 5184 4185 5212 19110
rect 5356 18896 5408 18902
rect 5356 18838 5408 18844
rect 5368 18426 5396 18838
rect 5460 18766 5488 19314
rect 5540 19304 5592 19310
rect 5540 19246 5592 19252
rect 6460 19304 6512 19310
rect 6460 19246 6512 19252
rect 5448 18760 5500 18766
rect 5448 18702 5500 18708
rect 5356 18420 5408 18426
rect 5356 18362 5408 18368
rect 5264 17128 5316 17134
rect 5264 17070 5316 17076
rect 5276 16658 5304 17070
rect 5264 16652 5316 16658
rect 5264 16594 5316 16600
rect 5276 16250 5304 16594
rect 5448 16584 5500 16590
rect 5448 16526 5500 16532
rect 5264 16244 5316 16250
rect 5264 16186 5316 16192
rect 5276 16046 5304 16186
rect 5264 16040 5316 16046
rect 5264 15982 5316 15988
rect 5276 15706 5304 15982
rect 5264 15700 5316 15706
rect 5264 15642 5316 15648
rect 5276 15434 5304 15642
rect 5460 15570 5488 16526
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 5264 15428 5316 15434
rect 5264 15370 5316 15376
rect 5264 14884 5316 14890
rect 5264 14826 5316 14832
rect 5276 14618 5304 14826
rect 5460 14618 5488 15506
rect 5264 14612 5316 14618
rect 5264 14554 5316 14560
rect 5448 14612 5500 14618
rect 5448 14554 5500 14560
rect 5264 14476 5316 14482
rect 5264 14418 5316 14424
rect 5276 14074 5304 14418
rect 5264 14068 5316 14074
rect 5264 14010 5316 14016
rect 5356 14068 5408 14074
rect 5356 14010 5408 14016
rect 5276 13462 5304 14010
rect 5264 13456 5316 13462
rect 5264 13398 5316 13404
rect 5276 12986 5304 13398
rect 5264 12980 5316 12986
rect 5264 12922 5316 12928
rect 5264 12640 5316 12646
rect 5264 12582 5316 12588
rect 5276 12442 5304 12582
rect 5264 12436 5316 12442
rect 5264 12378 5316 12384
rect 5368 11354 5396 14010
rect 5552 13814 5580 19246
rect 6184 19236 6236 19242
rect 6184 19178 6236 19184
rect 5816 18964 5868 18970
rect 5816 18906 5868 18912
rect 5632 18828 5684 18834
rect 5632 18770 5684 18776
rect 5644 18426 5672 18770
rect 5632 18420 5684 18426
rect 5632 18362 5684 18368
rect 5644 18222 5672 18362
rect 5632 18216 5684 18222
rect 5632 18158 5684 18164
rect 5632 17740 5684 17746
rect 5632 17682 5684 17688
rect 5644 17270 5672 17682
rect 5632 17264 5684 17270
rect 5632 17206 5684 17212
rect 5644 16658 5672 17206
rect 5724 17128 5776 17134
rect 5724 17070 5776 17076
rect 5632 16652 5684 16658
rect 5632 16594 5684 16600
rect 5632 14884 5684 14890
rect 5632 14826 5684 14832
rect 5644 14482 5672 14826
rect 5632 14476 5684 14482
rect 5632 14418 5684 14424
rect 5736 14278 5764 17070
rect 5724 14272 5776 14278
rect 5644 14232 5724 14260
rect 5644 13977 5672 14232
rect 5724 14214 5776 14220
rect 5630 13968 5686 13977
rect 5630 13903 5686 13912
rect 5644 13870 5672 13903
rect 5460 13786 5580 13814
rect 5632 13864 5684 13870
rect 5632 13806 5684 13812
rect 5356 11348 5408 11354
rect 5356 11290 5408 11296
rect 5354 11248 5410 11257
rect 5354 11183 5410 11192
rect 5368 10146 5396 11183
rect 5460 10198 5488 13786
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5552 12442 5580 13262
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 5736 12374 5764 12922
rect 5724 12368 5776 12374
rect 5724 12310 5776 12316
rect 5724 12232 5776 12238
rect 5724 12174 5776 12180
rect 5632 11688 5684 11694
rect 5538 11656 5594 11665
rect 5632 11630 5684 11636
rect 5538 11591 5594 11600
rect 5276 10118 5396 10146
rect 5448 10192 5500 10198
rect 5448 10134 5500 10140
rect 5276 8022 5304 10118
rect 5356 10056 5408 10062
rect 5356 9998 5408 10004
rect 5368 9722 5396 9998
rect 5356 9716 5408 9722
rect 5356 9658 5408 9664
rect 5264 8016 5316 8022
rect 5264 7958 5316 7964
rect 5448 7948 5500 7954
rect 5368 7908 5448 7936
rect 5368 6662 5396 7908
rect 5448 7890 5500 7896
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 5170 4176 5226 4185
rect 4988 4140 5040 4146
rect 5170 4111 5226 4120
rect 4988 4082 5040 4088
rect 4160 4004 4212 4010
rect 4160 3946 4212 3952
rect 4172 3602 4200 3946
rect 5276 3738 5304 5170
rect 5368 4146 5396 6598
rect 5552 6440 5580 11591
rect 5460 6412 5580 6440
rect 5460 6322 5488 6412
rect 5448 6316 5500 6322
rect 5448 6258 5500 6264
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5448 6180 5500 6186
rect 5448 6122 5500 6128
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 5264 3732 5316 3738
rect 5264 3674 5316 3680
rect 4528 3664 4580 3670
rect 4528 3606 4580 3612
rect 4160 3596 4212 3602
rect 4160 3538 4212 3544
rect 4540 3126 4568 3606
rect 5172 3460 5224 3466
rect 5172 3402 5224 3408
rect 5184 3369 5212 3402
rect 5170 3360 5226 3369
rect 4622 3292 4918 3312
rect 5170 3295 5226 3304
rect 4678 3290 4702 3292
rect 4758 3290 4782 3292
rect 4838 3290 4862 3292
rect 4700 3238 4702 3290
rect 4764 3238 4776 3290
rect 4838 3238 4840 3290
rect 4678 3236 4702 3238
rect 4758 3236 4782 3238
rect 4838 3236 4862 3238
rect 4622 3216 4918 3236
rect 5078 3224 5134 3233
rect 5078 3159 5134 3168
rect 4528 3120 4580 3126
rect 4528 3062 4580 3068
rect 4344 2916 4396 2922
rect 4344 2858 4396 2864
rect 4356 2650 4384 2858
rect 4540 2854 4568 3062
rect 4988 2984 5040 2990
rect 5092 2972 5120 3159
rect 5276 3058 5304 3674
rect 5368 3641 5396 4082
rect 5354 3632 5410 3641
rect 5354 3567 5410 3576
rect 5356 3460 5408 3466
rect 5356 3402 5408 3408
rect 5264 3052 5316 3058
rect 5264 2994 5316 3000
rect 5040 2944 5120 2972
rect 4988 2926 5040 2932
rect 5368 2922 5396 3402
rect 5356 2916 5408 2922
rect 5356 2858 5408 2864
rect 4528 2848 4580 2854
rect 4528 2790 4580 2796
rect 5264 2848 5316 2854
rect 5264 2790 5316 2796
rect 4344 2644 4396 2650
rect 4344 2586 4396 2592
rect 4540 2310 4568 2790
rect 5276 2582 5304 2790
rect 5264 2576 5316 2582
rect 5264 2518 5316 2524
rect 4896 2508 4948 2514
rect 4948 2468 5028 2496
rect 4896 2450 4948 2456
rect 5000 2310 5028 2468
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 4988 2304 5040 2310
rect 4988 2246 5040 2252
rect 4622 2204 4918 2224
rect 4678 2202 4702 2204
rect 4758 2202 4782 2204
rect 4838 2202 4862 2204
rect 4700 2150 4702 2202
rect 4764 2150 4776 2202
rect 4838 2150 4840 2202
rect 4678 2148 4702 2150
rect 4758 2148 4782 2150
rect 4838 2148 4862 2150
rect 4622 2128 4918 2148
rect 5460 1193 5488 6122
rect 5552 5914 5580 6258
rect 5644 6254 5672 11630
rect 5736 11354 5764 12174
rect 5724 11348 5776 11354
rect 5724 11290 5776 11296
rect 5828 11014 5856 18906
rect 6000 18760 6052 18766
rect 6000 18702 6052 18708
rect 6012 18426 6040 18702
rect 6000 18420 6052 18426
rect 6000 18362 6052 18368
rect 6000 17876 6052 17882
rect 6000 17818 6052 17824
rect 5908 17740 5960 17746
rect 5908 17682 5960 17688
rect 5920 17066 5948 17682
rect 5908 17060 5960 17066
rect 5908 17002 5960 17008
rect 5908 15156 5960 15162
rect 5908 15098 5960 15104
rect 5920 14482 5948 15098
rect 5908 14476 5960 14482
rect 5908 14418 5960 14424
rect 5908 12708 5960 12714
rect 5908 12650 5960 12656
rect 5920 12170 5948 12650
rect 5908 12164 5960 12170
rect 5908 12106 5960 12112
rect 5816 11008 5868 11014
rect 5816 10950 5868 10956
rect 5828 10266 5856 10950
rect 5816 10260 5868 10266
rect 5816 10202 5868 10208
rect 5816 9104 5868 9110
rect 5816 9046 5868 9052
rect 5908 9104 5960 9110
rect 5908 9046 5960 9052
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 5736 8514 5764 8978
rect 5828 8838 5856 9046
rect 5816 8832 5868 8838
rect 5816 8774 5868 8780
rect 5920 8634 5948 9046
rect 6012 8634 6040 17818
rect 6092 16992 6144 16998
rect 6092 16934 6144 16940
rect 6104 16522 6132 16934
rect 6092 16516 6144 16522
rect 6092 16458 6144 16464
rect 6092 15428 6144 15434
rect 6092 15370 6144 15376
rect 6104 14074 6132 15370
rect 6092 14068 6144 14074
rect 6092 14010 6144 14016
rect 6092 13184 6144 13190
rect 6092 13126 6144 13132
rect 6104 12850 6132 13126
rect 6092 12844 6144 12850
rect 6092 12786 6144 12792
rect 6090 11928 6146 11937
rect 6090 11863 6146 11872
rect 6104 11830 6132 11863
rect 6092 11824 6144 11830
rect 6092 11766 6144 11772
rect 6092 11348 6144 11354
rect 6092 11290 6144 11296
rect 6104 10810 6132 11290
rect 6092 10804 6144 10810
rect 6092 10746 6144 10752
rect 6092 8968 6144 8974
rect 6092 8910 6144 8916
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 5736 8486 5948 8514
rect 5816 7948 5868 7954
rect 5736 7908 5816 7936
rect 5736 6866 5764 7908
rect 5816 7890 5868 7896
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 5736 6458 5764 6802
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 5632 6248 5684 6254
rect 5632 6190 5684 6196
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5632 5704 5684 5710
rect 5632 5646 5684 5652
rect 5644 5030 5672 5646
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 5552 2009 5580 4558
rect 5538 2000 5594 2009
rect 5538 1935 5594 1944
rect 5644 1737 5672 4966
rect 5828 4010 5856 7482
rect 5920 7410 5948 8486
rect 6012 8022 6040 8570
rect 6104 8498 6132 8910
rect 6092 8492 6144 8498
rect 6092 8434 6144 8440
rect 6000 8016 6052 8022
rect 6000 7958 6052 7964
rect 6012 7546 6040 7958
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 5920 6866 5948 7346
rect 6000 6928 6052 6934
rect 6000 6870 6052 6876
rect 5908 6860 5960 6866
rect 5908 6802 5960 6808
rect 5908 6656 5960 6662
rect 5908 6598 5960 6604
rect 5920 6118 5948 6598
rect 5908 6112 5960 6118
rect 5908 6054 5960 6060
rect 6012 4154 6040 6870
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 5920 4146 6040 4154
rect 5908 4140 6040 4146
rect 5960 4126 6040 4140
rect 5908 4082 5960 4088
rect 6104 4049 6132 4966
rect 6090 4040 6146 4049
rect 5816 4004 5868 4010
rect 6090 3975 6146 3984
rect 5816 3946 5868 3952
rect 6196 2514 6224 19178
rect 6472 19174 6500 19246
rect 6460 19168 6512 19174
rect 6460 19110 6512 19116
rect 6276 18760 6328 18766
rect 6276 18702 6328 18708
rect 6288 13938 6316 18702
rect 6368 17332 6420 17338
rect 6368 17274 6420 17280
rect 6276 13932 6328 13938
rect 6276 13874 6328 13880
rect 6276 13456 6328 13462
rect 6276 13398 6328 13404
rect 6288 12986 6316 13398
rect 6276 12980 6328 12986
rect 6276 12922 6328 12928
rect 6288 12646 6316 12922
rect 6276 12640 6328 12646
rect 6276 12582 6328 12588
rect 6276 12368 6328 12374
rect 6276 12310 6328 12316
rect 6288 11898 6316 12310
rect 6276 11892 6328 11898
rect 6276 11834 6328 11840
rect 6288 11354 6316 11834
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 6276 11144 6328 11150
rect 6276 11086 6328 11092
rect 6288 10810 6316 11086
rect 6276 10804 6328 10810
rect 6276 10746 6328 10752
rect 6276 8968 6328 8974
rect 6276 8910 6328 8916
rect 6288 8566 6316 8910
rect 6276 8560 6328 8566
rect 6276 8502 6328 8508
rect 6380 7002 6408 17274
rect 6472 15978 6500 19110
rect 6644 18828 6696 18834
rect 6644 18770 6696 18776
rect 6656 18426 6684 18770
rect 6644 18420 6696 18426
rect 6644 18362 6696 18368
rect 6748 17762 6776 19382
rect 7012 19372 7064 19378
rect 7012 19314 7064 19320
rect 6828 18760 6880 18766
rect 6828 18702 6880 18708
rect 6656 17734 6776 17762
rect 6552 16788 6604 16794
rect 6552 16730 6604 16736
rect 6460 15972 6512 15978
rect 6460 15914 6512 15920
rect 6460 15360 6512 15366
rect 6460 15302 6512 15308
rect 6472 15162 6500 15302
rect 6460 15156 6512 15162
rect 6460 15098 6512 15104
rect 6564 15042 6592 16730
rect 6472 15014 6592 15042
rect 6472 11529 6500 15014
rect 6656 14940 6684 17734
rect 6736 17672 6788 17678
rect 6736 17614 6788 17620
rect 6564 14912 6684 14940
rect 6564 11762 6592 14912
rect 6644 14476 6696 14482
rect 6644 14418 6696 14424
rect 6656 14113 6684 14418
rect 6642 14104 6698 14113
rect 6642 14039 6644 14048
rect 6696 14039 6698 14048
rect 6644 14010 6696 14016
rect 6656 13979 6684 14010
rect 6644 13932 6696 13938
rect 6644 13874 6696 13880
rect 6656 13841 6684 13874
rect 6642 13832 6698 13841
rect 6642 13767 6698 13776
rect 6552 11756 6604 11762
rect 6552 11698 6604 11704
rect 6458 11520 6514 11529
rect 6458 11455 6514 11464
rect 6644 11144 6696 11150
rect 6644 11086 6696 11092
rect 6656 10266 6684 11086
rect 6748 10266 6776 17614
rect 6840 17270 6868 18702
rect 6920 18080 6972 18086
rect 6920 18022 6972 18028
rect 6828 17264 6880 17270
rect 6828 17206 6880 17212
rect 6840 17134 6868 17206
rect 6828 17128 6880 17134
rect 6828 17070 6880 17076
rect 6932 16726 6960 18022
rect 6920 16720 6972 16726
rect 6920 16662 6972 16668
rect 6828 16584 6880 16590
rect 6828 16526 6880 16532
rect 6840 16114 6868 16526
rect 6932 16250 6960 16662
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 6828 16108 6880 16114
rect 6828 16050 6880 16056
rect 7024 15994 7052 19314
rect 7288 19304 7340 19310
rect 7288 19246 7340 19252
rect 7104 19236 7156 19242
rect 7104 19178 7156 19184
rect 7116 17610 7144 19178
rect 7196 18624 7248 18630
rect 7300 18612 7328 19246
rect 8289 19068 8585 19088
rect 8345 19066 8369 19068
rect 8425 19066 8449 19068
rect 8505 19066 8529 19068
rect 8367 19014 8369 19066
rect 8431 19014 8443 19066
rect 8505 19014 8507 19066
rect 8345 19012 8369 19014
rect 8425 19012 8449 19014
rect 8505 19012 8529 19014
rect 8289 18992 8585 19012
rect 7472 18828 7524 18834
rect 7472 18770 7524 18776
rect 7380 18692 7432 18698
rect 7380 18634 7432 18640
rect 7248 18584 7328 18612
rect 7196 18566 7248 18572
rect 7104 17604 7156 17610
rect 7104 17546 7156 17552
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 7208 17134 7236 17478
rect 7196 17128 7248 17134
rect 7196 17070 7248 17076
rect 6840 15966 7052 15994
rect 6644 10260 6696 10266
rect 6644 10202 6696 10208
rect 6736 10260 6788 10266
rect 6736 10202 6788 10208
rect 6552 10124 6604 10130
rect 6552 10066 6604 10072
rect 6564 9382 6592 10066
rect 6748 9586 6776 10202
rect 6840 10062 6868 15966
rect 7104 15904 7156 15910
rect 7104 15846 7156 15852
rect 7116 15638 7144 15846
rect 7104 15632 7156 15638
rect 7104 15574 7156 15580
rect 7116 14890 7144 15574
rect 7104 14884 7156 14890
rect 7104 14826 7156 14832
rect 7196 14884 7248 14890
rect 7196 14826 7248 14832
rect 7012 14816 7064 14822
rect 7012 14758 7064 14764
rect 7024 14618 7052 14758
rect 7012 14612 7064 14618
rect 7012 14554 7064 14560
rect 6920 14340 6972 14346
rect 6920 14282 6972 14288
rect 6932 12850 6960 14282
rect 7024 13802 7052 14554
rect 7116 14550 7144 14826
rect 7104 14544 7156 14550
rect 7104 14486 7156 14492
rect 7208 14346 7236 14826
rect 7196 14340 7248 14346
rect 7196 14282 7248 14288
rect 7208 13802 7236 14282
rect 7012 13796 7064 13802
rect 7012 13738 7064 13744
rect 7196 13796 7248 13802
rect 7196 13738 7248 13744
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 6932 12442 6960 12786
rect 7012 12708 7064 12714
rect 7012 12650 7064 12656
rect 6920 12436 6972 12442
rect 6920 12378 6972 12384
rect 7024 12374 7052 12650
rect 7012 12368 7064 12374
rect 7012 12310 7064 12316
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 7024 11626 7052 12038
rect 7104 11756 7156 11762
rect 7104 11698 7156 11704
rect 7012 11620 7064 11626
rect 7012 11562 7064 11568
rect 6920 11552 6972 11558
rect 6920 11494 6972 11500
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 6460 7948 6512 7954
rect 6460 7890 6512 7896
rect 6472 7206 6500 7890
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 6368 6996 6420 7002
rect 6368 6938 6420 6944
rect 6276 6860 6328 6866
rect 6276 6802 6328 6808
rect 6288 6186 6316 6802
rect 6472 6390 6500 7142
rect 6564 6730 6592 9318
rect 6932 9042 6960 11494
rect 7024 11354 7052 11562
rect 7116 11354 7144 11698
rect 7012 11348 7064 11354
rect 7012 11290 7064 11296
rect 7104 11348 7156 11354
rect 7104 11290 7156 11296
rect 7024 10810 7052 11290
rect 7196 11280 7248 11286
rect 7196 11222 7248 11228
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 7024 10470 7052 10746
rect 7208 10538 7236 11222
rect 7196 10532 7248 10538
rect 7196 10474 7248 10480
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 7300 10146 7328 18584
rect 7392 18426 7420 18634
rect 7484 18426 7512 18770
rect 8208 18624 8260 18630
rect 8208 18566 8260 18572
rect 7380 18420 7432 18426
rect 7380 18362 7432 18368
rect 7472 18420 7524 18426
rect 7472 18362 7524 18368
rect 7564 18352 7616 18358
rect 7564 18294 7616 18300
rect 7576 17610 7604 18294
rect 8220 18222 8248 18566
rect 7932 18216 7984 18222
rect 7932 18158 7984 18164
rect 8208 18216 8260 18222
rect 8208 18158 8260 18164
rect 7838 17776 7894 17785
rect 7656 17740 7708 17746
rect 7838 17711 7894 17720
rect 7656 17682 7708 17688
rect 7564 17604 7616 17610
rect 7564 17546 7616 17552
rect 7380 16992 7432 16998
rect 7380 16934 7432 16940
rect 7392 14482 7420 16934
rect 7576 16794 7604 17546
rect 7668 17066 7696 17682
rect 7656 17060 7708 17066
rect 7656 17002 7708 17008
rect 7564 16788 7616 16794
rect 7564 16730 7616 16736
rect 7472 15632 7524 15638
rect 7472 15574 7524 15580
rect 7484 15162 7512 15574
rect 7564 15496 7616 15502
rect 7564 15438 7616 15444
rect 7472 15156 7524 15162
rect 7472 15098 7524 15104
rect 7576 14958 7604 15438
rect 7564 14952 7616 14958
rect 7564 14894 7616 14900
rect 7380 14476 7432 14482
rect 7380 14418 7432 14424
rect 7472 14408 7524 14414
rect 7208 10118 7328 10146
rect 7392 14356 7472 14362
rect 7392 14350 7524 14356
rect 7392 14334 7512 14350
rect 6920 9036 6972 9042
rect 6920 8978 6972 8984
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 6840 7750 6868 8502
rect 6932 8090 6960 8978
rect 7104 8424 7156 8430
rect 7104 8366 7156 8372
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 7116 7818 7144 8366
rect 7104 7812 7156 7818
rect 7104 7754 7156 7760
rect 6828 7744 6880 7750
rect 6828 7686 6880 7692
rect 6552 6724 6604 6730
rect 6552 6666 6604 6672
rect 6460 6384 6512 6390
rect 6460 6326 6512 6332
rect 6552 6384 6604 6390
rect 6552 6326 6604 6332
rect 6276 6180 6328 6186
rect 6276 6122 6328 6128
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 6288 3097 6316 4966
rect 6472 4593 6500 6326
rect 6564 4622 6592 6326
rect 6644 5840 6696 5846
rect 6644 5782 6696 5788
rect 6656 5370 6684 5782
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 6840 5273 6868 7686
rect 7116 7342 7144 7754
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 7104 7336 7156 7342
rect 7104 7278 7156 7284
rect 6932 7002 6960 7278
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 7208 6866 7236 10118
rect 7288 10056 7340 10062
rect 7288 9998 7340 10004
rect 7300 9178 7328 9998
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 7196 6860 7248 6866
rect 7196 6802 7248 6808
rect 7208 6186 7236 6802
rect 7012 6180 7064 6186
rect 7012 6122 7064 6128
rect 7196 6180 7248 6186
rect 7196 6122 7248 6128
rect 7024 5574 7052 6122
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 6826 5264 6882 5273
rect 6826 5199 6882 5208
rect 7024 5098 7052 5510
rect 6920 5092 6972 5098
rect 6920 5034 6972 5040
rect 7012 5092 7064 5098
rect 7012 5034 7064 5040
rect 6644 4752 6696 4758
rect 6644 4694 6696 4700
rect 6552 4616 6604 4622
rect 6458 4584 6514 4593
rect 6552 4558 6604 4564
rect 6458 4519 6514 4528
rect 6656 3942 6684 4694
rect 6932 4554 6960 5034
rect 7024 4826 7052 5034
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 7300 4758 7328 7482
rect 7288 4752 7340 4758
rect 7288 4694 7340 4700
rect 6920 4548 6972 4554
rect 6920 4490 6972 4496
rect 6552 3936 6604 3942
rect 6552 3878 6604 3884
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 6564 3670 6592 3878
rect 6656 3738 6684 3878
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 6552 3664 6604 3670
rect 6552 3606 6604 3612
rect 6368 3528 6420 3534
rect 6368 3470 6420 3476
rect 6274 3088 6330 3097
rect 6274 3023 6330 3032
rect 6184 2508 6236 2514
rect 6184 2450 6236 2456
rect 6380 2417 6408 3470
rect 7104 3392 7156 3398
rect 7104 3334 7156 3340
rect 7116 3058 7144 3334
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 7012 2916 7064 2922
rect 7012 2858 7064 2864
rect 7024 2650 7052 2858
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 6736 2576 6788 2582
rect 6736 2518 6788 2524
rect 6748 2428 6776 2518
rect 7116 2514 7144 2994
rect 7300 2854 7328 4694
rect 7392 4554 7420 14334
rect 7472 14272 7524 14278
rect 7472 14214 7524 14220
rect 7484 14074 7512 14214
rect 7472 14068 7524 14074
rect 7472 14010 7524 14016
rect 7576 13954 7604 14894
rect 7484 13926 7604 13954
rect 7484 13258 7512 13926
rect 7564 13796 7616 13802
rect 7564 13738 7616 13744
rect 7472 13252 7524 13258
rect 7472 13194 7524 13200
rect 7484 12918 7512 13194
rect 7472 12912 7524 12918
rect 7472 12854 7524 12860
rect 7472 12436 7524 12442
rect 7472 12378 7524 12384
rect 7484 11218 7512 12378
rect 7576 12102 7604 13738
rect 7564 12096 7616 12102
rect 7564 12038 7616 12044
rect 7472 11212 7524 11218
rect 7472 11154 7524 11160
rect 7484 10810 7512 11154
rect 7668 11014 7696 17002
rect 7748 16720 7800 16726
rect 7748 16662 7800 16668
rect 7760 15910 7788 16662
rect 7748 15904 7800 15910
rect 7748 15846 7800 15852
rect 7760 15706 7788 15846
rect 7748 15700 7800 15706
rect 7748 15642 7800 15648
rect 7748 14000 7800 14006
rect 7748 13942 7800 13948
rect 7760 12782 7788 13942
rect 7748 12776 7800 12782
rect 7748 12718 7800 12724
rect 7852 12458 7880 17711
rect 7944 14006 7972 18158
rect 8220 17746 8248 18158
rect 8289 17980 8585 18000
rect 8345 17978 8369 17980
rect 8425 17978 8449 17980
rect 8505 17978 8529 17980
rect 8367 17926 8369 17978
rect 8431 17926 8443 17978
rect 8505 17926 8507 17978
rect 8345 17924 8369 17926
rect 8425 17924 8449 17926
rect 8505 17924 8529 17926
rect 8289 17904 8585 17924
rect 8208 17740 8260 17746
rect 8208 17682 8260 17688
rect 8220 17066 8248 17682
rect 8208 17060 8260 17066
rect 8208 17002 8260 17008
rect 8289 16892 8585 16912
rect 8345 16890 8369 16892
rect 8425 16890 8449 16892
rect 8505 16890 8529 16892
rect 8367 16838 8369 16890
rect 8431 16838 8443 16890
rect 8505 16838 8507 16890
rect 8345 16836 8369 16838
rect 8425 16836 8449 16838
rect 8505 16836 8529 16838
rect 8289 16816 8585 16836
rect 8024 16652 8076 16658
rect 8024 16594 8076 16600
rect 8116 16652 8168 16658
rect 8116 16594 8168 16600
rect 8036 15638 8064 16594
rect 8128 16561 8156 16594
rect 8114 16552 8170 16561
rect 8114 16487 8170 16496
rect 8208 16040 8260 16046
rect 8208 15982 8260 15988
rect 8116 15904 8168 15910
rect 8116 15846 8168 15852
rect 8024 15632 8076 15638
rect 8024 15574 8076 15580
rect 8036 15502 8064 15574
rect 8024 15496 8076 15502
rect 8024 15438 8076 15444
rect 8036 15026 8064 15438
rect 8024 15020 8076 15026
rect 8024 14962 8076 14968
rect 8024 14884 8076 14890
rect 8024 14826 8076 14832
rect 7932 14000 7984 14006
rect 7932 13942 7984 13948
rect 7932 13388 7984 13394
rect 7932 13330 7984 13336
rect 7944 12481 7972 13330
rect 7760 12430 7880 12458
rect 7930 12472 7986 12481
rect 7760 11778 7788 12430
rect 7930 12407 7986 12416
rect 7944 12374 7972 12407
rect 7840 12368 7892 12374
rect 7840 12310 7892 12316
rect 7932 12368 7984 12374
rect 7932 12310 7984 12316
rect 7852 11898 7880 12310
rect 7840 11892 7892 11898
rect 7840 11834 7892 11840
rect 7760 11750 7972 11778
rect 7656 11008 7708 11014
rect 7656 10950 7708 10956
rect 7840 11008 7892 11014
rect 7840 10950 7892 10956
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7748 10804 7800 10810
rect 7748 10746 7800 10752
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7484 9178 7512 10610
rect 7576 10062 7604 10610
rect 7656 10192 7708 10198
rect 7656 10134 7708 10140
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7668 9382 7696 10134
rect 7656 9376 7708 9382
rect 7656 9318 7708 9324
rect 7472 9172 7524 9178
rect 7472 9114 7524 9120
rect 7668 9110 7696 9318
rect 7656 9104 7708 9110
rect 7656 9046 7708 9052
rect 7472 9036 7524 9042
rect 7472 8978 7524 8984
rect 7484 8090 7512 8978
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7472 7948 7524 7954
rect 7472 7890 7524 7896
rect 7484 7313 7512 7890
rect 7576 7478 7604 8570
rect 7760 8430 7788 10746
rect 7852 9110 7880 10950
rect 7840 9104 7892 9110
rect 7840 9046 7892 9052
rect 7840 8900 7892 8906
rect 7840 8842 7892 8848
rect 7852 8634 7880 8842
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 7748 8424 7800 8430
rect 7748 8366 7800 8372
rect 7564 7472 7616 7478
rect 7944 7426 7972 11750
rect 8036 7546 8064 14826
rect 8128 13841 8156 15846
rect 8220 15706 8248 15982
rect 8289 15804 8585 15824
rect 8345 15802 8369 15804
rect 8425 15802 8449 15804
rect 8505 15802 8529 15804
rect 8367 15750 8369 15802
rect 8431 15750 8443 15802
rect 8505 15750 8507 15802
rect 8345 15748 8369 15750
rect 8425 15748 8449 15750
rect 8505 15748 8529 15750
rect 8289 15728 8585 15748
rect 8208 15700 8260 15706
rect 8208 15642 8260 15648
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 8220 14618 8248 14758
rect 8289 14716 8585 14736
rect 8345 14714 8369 14716
rect 8425 14714 8449 14716
rect 8505 14714 8529 14716
rect 8367 14662 8369 14714
rect 8431 14662 8443 14714
rect 8505 14662 8507 14714
rect 8345 14660 8369 14662
rect 8425 14660 8449 14662
rect 8505 14660 8529 14662
rect 8289 14640 8585 14660
rect 8208 14612 8260 14618
rect 8208 14554 8260 14560
rect 8300 14544 8352 14550
rect 8300 14486 8352 14492
rect 8208 14476 8260 14482
rect 8208 14418 8260 14424
rect 8220 14006 8248 14418
rect 8208 14000 8260 14006
rect 8208 13942 8260 13948
rect 8312 13870 8340 14486
rect 8300 13864 8352 13870
rect 8114 13832 8170 13841
rect 8300 13806 8352 13812
rect 8114 13767 8170 13776
rect 8208 13796 8260 13802
rect 8128 11354 8156 13767
rect 8208 13738 8260 13744
rect 8220 13530 8248 13738
rect 8289 13628 8585 13648
rect 8345 13626 8369 13628
rect 8425 13626 8449 13628
rect 8505 13626 8529 13628
rect 8367 13574 8369 13626
rect 8431 13574 8443 13626
rect 8505 13574 8507 13626
rect 8345 13572 8369 13574
rect 8425 13572 8449 13574
rect 8505 13572 8529 13574
rect 8289 13552 8585 13572
rect 8208 13524 8260 13530
rect 8208 13466 8260 13472
rect 8208 12776 8260 12782
rect 8208 12718 8260 12724
rect 8220 12442 8248 12718
rect 8680 12646 8708 21542
rect 9034 21520 9090 21542
rect 12544 21542 12770 21570
rect 11956 19612 12252 19632
rect 12012 19610 12036 19612
rect 12092 19610 12116 19612
rect 12172 19610 12196 19612
rect 12034 19558 12036 19610
rect 12098 19558 12110 19610
rect 12172 19558 12174 19610
rect 12012 19556 12036 19558
rect 12092 19556 12116 19558
rect 12172 19556 12196 19558
rect 11956 19536 12252 19556
rect 10324 19304 10376 19310
rect 10324 19246 10376 19252
rect 11704 19304 11756 19310
rect 11704 19246 11756 19252
rect 8944 19168 8996 19174
rect 8944 19110 8996 19116
rect 9496 19168 9548 19174
rect 9496 19110 9548 19116
rect 8852 17060 8904 17066
rect 8852 17002 8904 17008
rect 8760 16992 8812 16998
rect 8760 16934 8812 16940
rect 8772 15978 8800 16934
rect 8760 15972 8812 15978
rect 8760 15914 8812 15920
rect 8668 12640 8720 12646
rect 8668 12582 8720 12588
rect 8289 12540 8585 12560
rect 8345 12538 8369 12540
rect 8425 12538 8449 12540
rect 8505 12538 8529 12540
rect 8367 12486 8369 12538
rect 8431 12486 8443 12538
rect 8505 12486 8507 12538
rect 8345 12484 8369 12486
rect 8425 12484 8449 12486
rect 8505 12484 8529 12486
rect 8289 12464 8585 12484
rect 8208 12436 8260 12442
rect 8208 12378 8260 12384
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 8220 11898 8248 12174
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 8289 11452 8585 11472
rect 8345 11450 8369 11452
rect 8425 11450 8449 11452
rect 8505 11450 8529 11452
rect 8367 11398 8369 11450
rect 8431 11398 8443 11450
rect 8505 11398 8507 11450
rect 8345 11396 8369 11398
rect 8425 11396 8449 11398
rect 8505 11396 8529 11398
rect 8289 11376 8585 11396
rect 8116 11348 8168 11354
rect 8116 11290 8168 11296
rect 8128 9722 8156 11290
rect 8208 11212 8260 11218
rect 8208 11154 8260 11160
rect 8220 9926 8248 11154
rect 8680 11082 8708 12582
rect 8864 11218 8892 17002
rect 8852 11212 8904 11218
rect 8852 11154 8904 11160
rect 8668 11076 8720 11082
rect 8668 11018 8720 11024
rect 8680 10470 8708 11018
rect 8668 10464 8720 10470
rect 8668 10406 8720 10412
rect 8760 10464 8812 10470
rect 8760 10406 8812 10412
rect 8289 10364 8585 10384
rect 8345 10362 8369 10364
rect 8425 10362 8449 10364
rect 8505 10362 8529 10364
rect 8367 10310 8369 10362
rect 8431 10310 8443 10362
rect 8505 10310 8507 10362
rect 8345 10308 8369 10310
rect 8425 10308 8449 10310
rect 8505 10308 8529 10310
rect 8289 10288 8585 10308
rect 8208 9920 8260 9926
rect 8208 9862 8260 9868
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 8220 9602 8248 9862
rect 8128 9574 8248 9602
rect 8128 9042 8156 9574
rect 8680 9353 8708 10406
rect 8772 9994 8800 10406
rect 8760 9988 8812 9994
rect 8760 9930 8812 9936
rect 8956 9674 8984 19110
rect 9404 18760 9456 18766
rect 9404 18702 9456 18708
rect 9128 18624 9180 18630
rect 9128 18566 9180 18572
rect 9036 17604 9088 17610
rect 9036 17546 9088 17552
rect 9048 15065 9076 17546
rect 9034 15056 9090 15065
rect 9034 14991 9090 15000
rect 9140 13954 9168 18566
rect 9312 17740 9364 17746
rect 9312 17682 9364 17688
rect 9324 17241 9352 17682
rect 9310 17232 9366 17241
rect 9310 17167 9366 17176
rect 9220 16992 9272 16998
rect 9220 16934 9272 16940
rect 9232 14074 9260 16934
rect 9324 16794 9352 17167
rect 9312 16788 9364 16794
rect 9312 16730 9364 16736
rect 9312 15972 9364 15978
rect 9312 15914 9364 15920
rect 9324 15570 9352 15914
rect 9312 15564 9364 15570
rect 9312 15506 9364 15512
rect 9324 15162 9352 15506
rect 9312 15156 9364 15162
rect 9312 15098 9364 15104
rect 9220 14068 9272 14074
rect 9220 14010 9272 14016
rect 9140 13926 9352 13954
rect 9036 13796 9088 13802
rect 9036 13738 9088 13744
rect 9048 13705 9076 13738
rect 9034 13696 9090 13705
rect 9034 13631 9090 13640
rect 9220 12096 9272 12102
rect 9220 12038 9272 12044
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 9048 10033 9076 11494
rect 9126 10704 9182 10713
rect 9126 10639 9182 10648
rect 9034 10024 9090 10033
rect 9034 9959 9090 9968
rect 8864 9646 8984 9674
rect 8760 9512 8812 9518
rect 8760 9454 8812 9460
rect 8666 9344 8722 9353
rect 8289 9276 8585 9296
rect 8666 9279 8722 9288
rect 8345 9274 8369 9276
rect 8425 9274 8449 9276
rect 8505 9274 8529 9276
rect 8367 9222 8369 9274
rect 8431 9222 8443 9274
rect 8505 9222 8507 9274
rect 8345 9220 8369 9222
rect 8425 9220 8449 9222
rect 8505 9220 8529 9222
rect 8289 9200 8585 9220
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 8116 9036 8168 9042
rect 8116 8978 8168 8984
rect 8128 8090 8156 8978
rect 8220 8634 8248 9114
rect 8680 8906 8708 9279
rect 8668 8900 8720 8906
rect 8668 8842 8720 8848
rect 8666 8664 8722 8673
rect 8208 8628 8260 8634
rect 8666 8599 8722 8608
rect 8208 8570 8260 8576
rect 8220 8362 8248 8570
rect 8680 8430 8708 8599
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8208 8356 8260 8362
rect 8208 8298 8260 8304
rect 8289 8188 8585 8208
rect 8345 8186 8369 8188
rect 8425 8186 8449 8188
rect 8505 8186 8529 8188
rect 8367 8134 8369 8186
rect 8431 8134 8443 8186
rect 8505 8134 8507 8186
rect 8345 8132 8369 8134
rect 8425 8132 8449 8134
rect 8505 8132 8529 8134
rect 8289 8112 8585 8132
rect 8680 8090 8708 8366
rect 8116 8084 8168 8090
rect 8116 8026 8168 8032
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 8392 7812 8444 7818
rect 8392 7754 8444 7760
rect 8116 7744 8168 7750
rect 8116 7686 8168 7692
rect 8024 7540 8076 7546
rect 8024 7482 8076 7488
rect 7564 7414 7616 7420
rect 7668 7398 7972 7426
rect 7470 7304 7526 7313
rect 7470 7239 7526 7248
rect 7484 7206 7512 7239
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 7484 7002 7512 7142
rect 7472 6996 7524 7002
rect 7472 6938 7524 6944
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 7484 5914 7512 6802
rect 7668 6322 7696 7398
rect 7840 7336 7892 7342
rect 7840 7278 7892 7284
rect 7852 6322 7880 7278
rect 8128 6866 8156 7686
rect 8404 7546 8432 7754
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8668 7336 8720 7342
rect 8668 7278 8720 7284
rect 8680 7177 8708 7278
rect 8666 7168 8722 7177
rect 8289 7100 8585 7120
rect 8666 7103 8722 7112
rect 8345 7098 8369 7100
rect 8425 7098 8449 7100
rect 8505 7098 8529 7100
rect 8367 7046 8369 7098
rect 8431 7046 8443 7098
rect 8505 7046 8507 7098
rect 8345 7044 8369 7046
rect 8425 7044 8449 7046
rect 8505 7044 8529 7046
rect 8289 7024 8585 7044
rect 8116 6860 8168 6866
rect 8116 6802 8168 6808
rect 8484 6860 8536 6866
rect 8484 6802 8536 6808
rect 7932 6792 7984 6798
rect 7932 6734 7984 6740
rect 7656 6316 7708 6322
rect 7656 6258 7708 6264
rect 7840 6316 7892 6322
rect 7840 6258 7892 6264
rect 7472 5908 7524 5914
rect 7472 5850 7524 5856
rect 7944 5778 7972 6734
rect 8128 6662 8156 6802
rect 8496 6769 8524 6802
rect 8772 6798 8800 9454
rect 8760 6792 8812 6798
rect 8482 6760 8538 6769
rect 8760 6734 8812 6740
rect 8482 6695 8538 6704
rect 8116 6656 8168 6662
rect 8116 6598 8168 6604
rect 8760 6180 8812 6186
rect 8760 6122 8812 6128
rect 8289 6012 8585 6032
rect 8345 6010 8369 6012
rect 8425 6010 8449 6012
rect 8505 6010 8529 6012
rect 8367 5958 8369 6010
rect 8431 5958 8443 6010
rect 8505 5958 8507 6010
rect 8345 5956 8369 5958
rect 8425 5956 8449 5958
rect 8505 5956 8529 5958
rect 8289 5936 8585 5956
rect 7932 5772 7984 5778
rect 7932 5714 7984 5720
rect 7944 4826 7972 5714
rect 8772 5574 8800 6122
rect 8760 5568 8812 5574
rect 8760 5510 8812 5516
rect 8668 5228 8720 5234
rect 8668 5170 8720 5176
rect 8116 5092 8168 5098
rect 8116 5034 8168 5040
rect 8128 4826 8156 5034
rect 8289 4924 8585 4944
rect 8345 4922 8369 4924
rect 8425 4922 8449 4924
rect 8505 4922 8529 4924
rect 8367 4870 8369 4922
rect 8431 4870 8443 4922
rect 8505 4870 8507 4922
rect 8345 4868 8369 4870
rect 8425 4868 8449 4870
rect 8505 4868 8529 4870
rect 8289 4848 8585 4868
rect 7932 4820 7984 4826
rect 7932 4762 7984 4768
rect 8116 4820 8168 4826
rect 8116 4762 8168 4768
rect 8208 4752 8260 4758
rect 8208 4694 8260 4700
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 7380 4548 7432 4554
rect 7380 4490 7432 4496
rect 7484 3534 7512 4558
rect 8116 4480 8168 4486
rect 8116 4422 8168 4428
rect 7564 4072 7616 4078
rect 7564 4014 7616 4020
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7576 3398 7604 4014
rect 7840 4004 7892 4010
rect 7840 3946 7892 3952
rect 7564 3392 7616 3398
rect 7564 3334 7616 3340
rect 7288 2848 7340 2854
rect 7288 2790 7340 2796
rect 7194 2680 7250 2689
rect 7194 2615 7250 2624
rect 7208 2582 7236 2615
rect 7196 2576 7248 2582
rect 7196 2518 7248 2524
rect 7104 2508 7156 2514
rect 7104 2450 7156 2456
rect 6828 2440 6880 2446
rect 6366 2408 6422 2417
rect 6092 2372 6144 2378
rect 6748 2400 6828 2428
rect 6828 2382 6880 2388
rect 6366 2343 6422 2352
rect 6092 2314 6144 2320
rect 5630 1728 5686 1737
rect 5630 1663 5686 1672
rect 5446 1184 5502 1193
rect 5446 1119 5502 1128
rect 3974 82 4030 480
rect 3896 54 4030 82
rect 570 0 626 54
rect 1674 0 1730 54
rect 2870 0 2926 54
rect 3974 0 4030 54
rect 5170 96 5226 480
rect 6104 82 6132 2314
rect 6380 2310 6408 2343
rect 6368 2304 6420 2310
rect 6368 2246 6420 2252
rect 7288 2304 7340 2310
rect 7288 2246 7340 2252
rect 6274 82 6330 480
rect 6104 54 6330 82
rect 7300 82 7328 2246
rect 7576 1601 7604 3334
rect 7852 2650 7880 3946
rect 8128 3738 8156 4422
rect 8220 4282 8248 4694
rect 8680 4554 8708 5170
rect 8772 5098 8800 5510
rect 8760 5092 8812 5098
rect 8760 5034 8812 5040
rect 8760 4684 8812 4690
rect 8760 4626 8812 4632
rect 8668 4548 8720 4554
rect 8668 4490 8720 4496
rect 8208 4276 8260 4282
rect 8208 4218 8260 4224
rect 8116 3732 8168 3738
rect 8116 3674 8168 3680
rect 8220 3670 8248 4218
rect 8772 4214 8800 4626
rect 8760 4208 8812 4214
rect 8760 4150 8812 4156
rect 8289 3836 8585 3856
rect 8345 3834 8369 3836
rect 8425 3834 8449 3836
rect 8505 3834 8529 3836
rect 8367 3782 8369 3834
rect 8431 3782 8443 3834
rect 8505 3782 8507 3834
rect 8345 3780 8369 3782
rect 8425 3780 8449 3782
rect 8505 3780 8529 3782
rect 8289 3760 8585 3780
rect 8208 3664 8260 3670
rect 8208 3606 8260 3612
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 8128 3398 8156 3470
rect 8116 3392 8168 3398
rect 8116 3334 8168 3340
rect 8220 3194 8248 3606
rect 8864 3194 8892 9646
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 9048 8838 9076 9454
rect 9036 8832 9088 8838
rect 9036 8774 9088 8780
rect 8944 8628 8996 8634
rect 8944 8570 8996 8576
rect 8956 6934 8984 8570
rect 9140 7970 9168 10639
rect 9048 7942 9168 7970
rect 9232 7954 9260 12038
rect 9220 7948 9272 7954
rect 9048 7818 9076 7942
rect 9220 7890 9272 7896
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9036 7812 9088 7818
rect 9036 7754 9088 7760
rect 9036 7336 9088 7342
rect 9036 7278 9088 7284
rect 9048 7002 9076 7278
rect 9036 6996 9088 7002
rect 9036 6938 9088 6944
rect 8944 6928 8996 6934
rect 8944 6870 8996 6876
rect 8942 4856 8998 4865
rect 8942 4791 8998 4800
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 8852 3188 8904 3194
rect 8852 3130 8904 3136
rect 8289 2748 8585 2768
rect 8345 2746 8369 2748
rect 8425 2746 8449 2748
rect 8505 2746 8529 2748
rect 8367 2694 8369 2746
rect 8431 2694 8443 2746
rect 8505 2694 8507 2746
rect 8345 2692 8369 2694
rect 8425 2692 8449 2694
rect 8505 2692 8529 2694
rect 8289 2672 8585 2692
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 7562 1592 7618 1601
rect 7562 1527 7618 1536
rect 7470 82 7526 480
rect 7300 54 7526 82
rect 5170 0 5226 40
rect 6274 0 6330 54
rect 7470 0 7526 54
rect 8666 82 8722 480
rect 8956 82 8984 4791
rect 9036 4072 9088 4078
rect 9036 4014 9088 4020
rect 9048 3738 9076 4014
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 9034 3496 9090 3505
rect 9034 3431 9090 3440
rect 9140 3482 9168 7822
rect 9220 7472 9272 7478
rect 9220 7414 9272 7420
rect 9232 7206 9260 7414
rect 9220 7200 9272 7206
rect 9220 7142 9272 7148
rect 9232 5846 9260 7142
rect 9324 7002 9352 13926
rect 9416 10742 9444 18702
rect 9508 15337 9536 19110
rect 9680 18148 9732 18154
rect 9680 18090 9732 18096
rect 9588 16788 9640 16794
rect 9588 16730 9640 16736
rect 9494 15328 9550 15337
rect 9494 15263 9550 15272
rect 9496 14816 9548 14822
rect 9496 14758 9548 14764
rect 9508 14550 9536 14758
rect 9496 14544 9548 14550
rect 9496 14486 9548 14492
rect 9508 14074 9536 14486
rect 9496 14068 9548 14074
rect 9496 14010 9548 14016
rect 9600 12918 9628 16730
rect 9692 16561 9720 18090
rect 9864 18080 9916 18086
rect 9864 18022 9916 18028
rect 9772 17196 9824 17202
rect 9772 17138 9824 17144
rect 9678 16552 9734 16561
rect 9678 16487 9734 16496
rect 9784 16454 9812 17138
rect 9772 16448 9824 16454
rect 9772 16390 9824 16396
rect 9680 16176 9732 16182
rect 9680 16118 9732 16124
rect 9692 14414 9720 16118
rect 9784 15881 9812 16390
rect 9770 15872 9826 15881
rect 9770 15807 9826 15816
rect 9772 15632 9824 15638
rect 9772 15574 9824 15580
rect 9784 15162 9812 15574
rect 9772 15156 9824 15162
rect 9772 15098 9824 15104
rect 9784 14822 9812 15098
rect 9772 14816 9824 14822
rect 9772 14758 9824 14764
rect 9876 14634 9904 18022
rect 10140 17740 10192 17746
rect 10140 17682 10192 17688
rect 10048 17672 10100 17678
rect 10048 17614 10100 17620
rect 9956 16652 10008 16658
rect 9956 16594 10008 16600
rect 9968 16250 9996 16594
rect 9956 16244 10008 16250
rect 9956 16186 10008 16192
rect 9956 15972 10008 15978
rect 9956 15914 10008 15920
rect 9968 15366 9996 15914
rect 9956 15360 10008 15366
rect 9956 15302 10008 15308
rect 9784 14606 9904 14634
rect 9968 14618 9996 15302
rect 9956 14612 10008 14618
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 9680 13728 9732 13734
rect 9784 13705 9812 14606
rect 9956 14554 10008 14560
rect 10060 14498 10088 17614
rect 10152 17134 10180 17682
rect 10232 17196 10284 17202
rect 10232 17138 10284 17144
rect 10140 17128 10192 17134
rect 10140 17070 10192 17076
rect 10152 16658 10180 17070
rect 10244 16794 10272 17138
rect 10232 16788 10284 16794
rect 10232 16730 10284 16736
rect 10140 16652 10192 16658
rect 10140 16594 10192 16600
rect 10232 16584 10284 16590
rect 10232 16526 10284 16532
rect 10244 15026 10272 16526
rect 10336 16096 10364 19246
rect 11244 19236 11296 19242
rect 11244 19178 11296 19184
rect 11256 18970 11284 19178
rect 11244 18964 11296 18970
rect 11244 18906 11296 18912
rect 11152 18828 11204 18834
rect 11152 18770 11204 18776
rect 11520 18828 11572 18834
rect 11520 18770 11572 18776
rect 10600 18692 10652 18698
rect 10600 18634 10652 18640
rect 10508 18216 10560 18222
rect 10508 18158 10560 18164
rect 10416 17808 10468 17814
rect 10416 17750 10468 17756
rect 10428 17066 10456 17750
rect 10416 17060 10468 17066
rect 10416 17002 10468 17008
rect 10428 16969 10456 17002
rect 10414 16960 10470 16969
rect 10414 16895 10470 16904
rect 10336 16068 10456 16096
rect 10324 15972 10376 15978
rect 10324 15914 10376 15920
rect 10336 15706 10364 15914
rect 10324 15700 10376 15706
rect 10324 15642 10376 15648
rect 10428 15026 10456 16068
rect 10520 15978 10548 18158
rect 10508 15972 10560 15978
rect 10508 15914 10560 15920
rect 10232 15020 10284 15026
rect 10232 14962 10284 14968
rect 10416 15020 10468 15026
rect 10416 14962 10468 14968
rect 10140 14816 10192 14822
rect 10140 14758 10192 14764
rect 9968 14470 10088 14498
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 9876 13802 9904 14010
rect 9864 13796 9916 13802
rect 9864 13738 9916 13744
rect 9680 13670 9732 13676
rect 9770 13696 9826 13705
rect 9692 13394 9720 13670
rect 9770 13631 9826 13640
rect 9770 13560 9826 13569
rect 9770 13495 9826 13504
rect 9680 13388 9732 13394
rect 9680 13330 9732 13336
rect 9692 12986 9720 13330
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9588 12912 9640 12918
rect 9588 12854 9640 12860
rect 9588 12776 9640 12782
rect 9588 12718 9640 12724
rect 9496 11688 9548 11694
rect 9496 11630 9548 11636
rect 9508 11014 9536 11630
rect 9496 11008 9548 11014
rect 9496 10950 9548 10956
rect 9404 10736 9456 10742
rect 9404 10678 9456 10684
rect 9404 9988 9456 9994
rect 9404 9930 9456 9936
rect 9312 6996 9364 7002
rect 9312 6938 9364 6944
rect 9324 6322 9352 6938
rect 9312 6316 9364 6322
rect 9312 6258 9364 6264
rect 9220 5840 9272 5846
rect 9220 5782 9272 5788
rect 9416 3670 9444 9930
rect 9508 9586 9536 10950
rect 9600 10713 9628 12718
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9692 12374 9720 12582
rect 9680 12368 9732 12374
rect 9680 12310 9732 12316
rect 9692 11830 9720 12310
rect 9680 11824 9732 11830
rect 9680 11766 9732 11772
rect 9692 11626 9720 11766
rect 9680 11620 9732 11626
rect 9680 11562 9732 11568
rect 9678 11112 9734 11121
rect 9678 11047 9734 11056
rect 9586 10704 9642 10713
rect 9586 10639 9642 10648
rect 9588 10532 9640 10538
rect 9588 10474 9640 10480
rect 9600 10130 9628 10474
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9496 9580 9548 9586
rect 9496 9522 9548 9528
rect 9588 9104 9640 9110
rect 9588 9046 9640 9052
rect 9600 8294 9628 9046
rect 9588 8288 9640 8294
rect 9588 8230 9640 8236
rect 9600 8129 9628 8230
rect 9586 8120 9642 8129
rect 9496 8084 9548 8090
rect 9586 8055 9642 8064
rect 9496 8026 9548 8032
rect 9508 4690 9536 8026
rect 9692 7342 9720 11047
rect 9680 7336 9732 7342
rect 9680 7278 9732 7284
rect 9784 6882 9812 13495
rect 9876 13462 9904 13738
rect 9864 13456 9916 13462
rect 9864 13398 9916 13404
rect 9864 12912 9916 12918
rect 9864 12854 9916 12860
rect 9876 9625 9904 12854
rect 9968 12306 9996 14470
rect 10048 14408 10100 14414
rect 10048 14350 10100 14356
rect 9956 12300 10008 12306
rect 9956 12242 10008 12248
rect 9968 11898 9996 12242
rect 9956 11892 10008 11898
rect 9956 11834 10008 11840
rect 9956 11620 10008 11626
rect 9956 11562 10008 11568
rect 9968 10266 9996 11562
rect 9956 10260 10008 10266
rect 9956 10202 10008 10208
rect 9956 10056 10008 10062
rect 9956 9998 10008 10004
rect 9862 9616 9918 9625
rect 9862 9551 9918 9560
rect 9876 8906 9904 9551
rect 9968 9178 9996 9998
rect 9956 9172 10008 9178
rect 9956 9114 10008 9120
rect 9864 8900 9916 8906
rect 9864 8842 9916 8848
rect 9876 8634 9904 8842
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9876 6934 9904 7142
rect 9692 6854 9812 6882
rect 9864 6928 9916 6934
rect 9864 6870 9916 6876
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 9496 4684 9548 4690
rect 9496 4626 9548 4632
rect 9404 3664 9456 3670
rect 9404 3606 9456 3612
rect 9218 3496 9274 3505
rect 9140 3454 9218 3482
rect 9048 3126 9076 3431
rect 9140 3233 9168 3454
rect 9218 3431 9274 3440
rect 9416 3398 9444 3606
rect 9600 3602 9628 6054
rect 9692 5681 9720 6854
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 9784 6390 9812 6734
rect 9772 6384 9824 6390
rect 9772 6326 9824 6332
rect 9876 5914 9904 6870
rect 10060 6730 10088 14350
rect 10152 14006 10180 14758
rect 10244 14618 10272 14962
rect 10232 14612 10284 14618
rect 10232 14554 10284 14560
rect 10140 14000 10192 14006
rect 10140 13942 10192 13948
rect 10416 13184 10468 13190
rect 10416 13126 10468 13132
rect 10140 11620 10192 11626
rect 10140 11562 10192 11568
rect 10048 6724 10100 6730
rect 10048 6666 10100 6672
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 9678 5672 9734 5681
rect 9678 5607 9734 5616
rect 10048 5636 10100 5642
rect 10048 5578 10100 5584
rect 10060 5302 10088 5578
rect 10048 5296 10100 5302
rect 10048 5238 10100 5244
rect 10152 4826 10180 11562
rect 10428 11082 10456 13126
rect 10508 12640 10560 12646
rect 10508 12582 10560 12588
rect 10520 11558 10548 12582
rect 10508 11552 10560 11558
rect 10508 11494 10560 11500
rect 10520 11286 10548 11494
rect 10508 11280 10560 11286
rect 10508 11222 10560 11228
rect 10416 11076 10468 11082
rect 10416 11018 10468 11024
rect 10520 10810 10548 11222
rect 10508 10804 10560 10810
rect 10508 10746 10560 10752
rect 10232 10260 10284 10266
rect 10232 10202 10284 10208
rect 10244 9722 10272 10202
rect 10232 9716 10284 9722
rect 10612 9674 10640 18634
rect 11164 18290 11192 18770
rect 11152 18284 11204 18290
rect 11152 18226 11204 18232
rect 10692 18216 10744 18222
rect 10692 18158 10744 18164
rect 10704 17542 10732 18158
rect 10876 18080 10928 18086
rect 10876 18022 10928 18028
rect 10692 17536 10744 17542
rect 10692 17478 10744 17484
rect 10704 17270 10732 17478
rect 10692 17264 10744 17270
rect 10692 17206 10744 17212
rect 10704 14414 10732 17206
rect 10784 16992 10836 16998
rect 10784 16934 10836 16940
rect 10692 14408 10744 14414
rect 10692 14350 10744 14356
rect 10692 11144 10744 11150
rect 10692 11086 10744 11092
rect 10704 10810 10732 11086
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 10692 10600 10744 10606
rect 10692 10542 10744 10548
rect 10232 9658 10284 9664
rect 10428 9646 10640 9674
rect 10324 9172 10376 9178
rect 10324 9114 10376 9120
rect 10336 9081 10364 9114
rect 10322 9072 10378 9081
rect 10322 9007 10378 9016
rect 10428 8974 10456 9646
rect 10416 8968 10468 8974
rect 10416 8910 10468 8916
rect 10600 8900 10652 8906
rect 10600 8842 10652 8848
rect 10232 7948 10284 7954
rect 10232 7890 10284 7896
rect 10244 7546 10272 7890
rect 10508 7744 10560 7750
rect 10508 7686 10560 7692
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 10244 7449 10272 7482
rect 10230 7440 10286 7449
rect 10230 7375 10286 7384
rect 10324 6248 10376 6254
rect 10324 6190 10376 6196
rect 10336 5642 10364 6190
rect 10414 5808 10470 5817
rect 10414 5743 10470 5752
rect 10428 5710 10456 5743
rect 10416 5704 10468 5710
rect 10416 5646 10468 5652
rect 10324 5636 10376 5642
rect 10324 5578 10376 5584
rect 10428 5370 10456 5646
rect 10520 5370 10548 7686
rect 10416 5364 10468 5370
rect 10416 5306 10468 5312
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 10612 5250 10640 8842
rect 10704 8362 10732 10542
rect 10796 10266 10824 16934
rect 10888 11354 10916 18022
rect 11060 17536 11112 17542
rect 11060 17478 11112 17484
rect 11072 14414 11100 17478
rect 11164 15094 11192 18226
rect 11532 18086 11560 18770
rect 11520 18080 11572 18086
rect 11520 18022 11572 18028
rect 11532 17746 11560 18022
rect 11520 17740 11572 17746
rect 11520 17682 11572 17688
rect 11336 17196 11388 17202
rect 11336 17138 11388 17144
rect 11152 15088 11204 15094
rect 11150 15056 11152 15065
rect 11204 15056 11206 15065
rect 11150 14991 11206 15000
rect 11244 15020 11296 15026
rect 11164 14965 11192 14991
rect 11244 14962 11296 14968
rect 11152 14544 11204 14550
rect 11152 14486 11204 14492
rect 11060 14408 11112 14414
rect 11060 14350 11112 14356
rect 10968 14272 11020 14278
rect 10968 14214 11020 14220
rect 10980 13530 11008 14214
rect 11072 14074 11100 14350
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 11164 13734 11192 14486
rect 11152 13728 11204 13734
rect 11152 13670 11204 13676
rect 10968 13524 11020 13530
rect 10968 13466 11020 13472
rect 11152 13524 11204 13530
rect 11152 13466 11204 13472
rect 10980 12850 11008 13466
rect 11058 13288 11114 13297
rect 11058 13223 11114 13232
rect 10968 12844 11020 12850
rect 10968 12786 11020 12792
rect 10968 11688 11020 11694
rect 10968 11630 11020 11636
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 10980 10606 11008 11630
rect 10968 10600 11020 10606
rect 10968 10542 11020 10548
rect 10784 10260 10836 10266
rect 10784 10202 10836 10208
rect 10796 9586 10824 10202
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 10980 9489 11008 9522
rect 10966 9480 11022 9489
rect 10966 9415 11022 9424
rect 10980 9042 11008 9415
rect 10968 9036 11020 9042
rect 10968 8978 11020 8984
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10692 8356 10744 8362
rect 10692 8298 10744 8304
rect 10796 7886 10824 8774
rect 10980 8090 11008 8978
rect 10968 8084 11020 8090
rect 10968 8026 11020 8032
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10796 7342 10824 7822
rect 10876 7472 10928 7478
rect 10876 7414 10928 7420
rect 10784 7336 10836 7342
rect 10784 7278 10836 7284
rect 10796 7002 10824 7278
rect 10888 7206 10916 7414
rect 10876 7200 10928 7206
rect 10876 7142 10928 7148
rect 10784 6996 10836 7002
rect 10784 6938 10836 6944
rect 10888 6186 10916 7142
rect 10876 6180 10928 6186
rect 10876 6122 10928 6128
rect 10888 5846 10916 6122
rect 10876 5840 10928 5846
rect 10876 5782 10928 5788
rect 10520 5222 10640 5250
rect 10782 5264 10838 5273
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 9864 4684 9916 4690
rect 9864 4626 9916 4632
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 9588 3596 9640 3602
rect 9588 3538 9640 3544
rect 9588 3460 9640 3466
rect 9588 3402 9640 3408
rect 9404 3392 9456 3398
rect 9404 3334 9456 3340
rect 9126 3224 9182 3233
rect 9126 3159 9182 3168
rect 9036 3120 9088 3126
rect 9036 3062 9088 3068
rect 9600 2922 9628 3402
rect 9876 3398 9904 4626
rect 9968 4282 9996 4626
rect 9956 4276 10008 4282
rect 9956 4218 10008 4224
rect 10324 4208 10376 4214
rect 10324 4150 10376 4156
rect 10336 3602 10364 4150
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 10048 3596 10100 3602
rect 10048 3538 10100 3544
rect 10324 3596 10376 3602
rect 10324 3538 10376 3544
rect 9864 3392 9916 3398
rect 9864 3334 9916 3340
rect 9968 3058 9996 3538
rect 10060 3369 10088 3538
rect 10046 3360 10102 3369
rect 10046 3295 10102 3304
rect 9956 3052 10008 3058
rect 9956 2994 10008 3000
rect 9968 2961 9996 2994
rect 9954 2952 10010 2961
rect 9036 2916 9088 2922
rect 9036 2858 9088 2864
rect 9588 2916 9640 2922
rect 9954 2887 10010 2896
rect 9588 2858 9640 2864
rect 9048 2650 9076 2858
rect 10060 2650 10088 3295
rect 10324 2848 10376 2854
rect 10324 2790 10376 2796
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 10336 2582 10364 2790
rect 10324 2576 10376 2582
rect 10324 2518 10376 2524
rect 8666 54 8984 82
rect 9770 128 9826 480
rect 10520 134 10548 5222
rect 10888 5234 10916 5782
rect 10782 5199 10838 5208
rect 10876 5228 10928 5234
rect 10796 5166 10824 5199
rect 10876 5170 10928 5176
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 10600 4616 10652 4622
rect 10600 4558 10652 4564
rect 10612 3738 10640 4558
rect 11072 4486 11100 13223
rect 11164 11694 11192 13466
rect 11152 11688 11204 11694
rect 11152 11630 11204 11636
rect 11150 11520 11206 11529
rect 11150 11455 11206 11464
rect 11164 10577 11192 11455
rect 11150 10568 11206 10577
rect 11150 10503 11206 10512
rect 11164 10198 11192 10503
rect 11152 10192 11204 10198
rect 11152 10134 11204 10140
rect 11164 9654 11192 10134
rect 11152 9648 11204 9654
rect 11152 9590 11204 9596
rect 11256 8906 11284 14962
rect 11348 13802 11376 17138
rect 11532 16998 11560 17682
rect 11520 16992 11572 16998
rect 11520 16934 11572 16940
rect 11428 16652 11480 16658
rect 11428 16594 11480 16600
rect 11440 15706 11468 16594
rect 11428 15700 11480 15706
rect 11428 15642 11480 15648
rect 11532 15042 11560 16934
rect 11612 15632 11664 15638
rect 11612 15574 11664 15580
rect 11624 15162 11652 15574
rect 11612 15156 11664 15162
rect 11612 15098 11664 15104
rect 11532 15014 11652 15042
rect 11518 14512 11574 14521
rect 11518 14447 11574 14456
rect 11428 14068 11480 14074
rect 11428 14010 11480 14016
rect 11336 13796 11388 13802
rect 11336 13738 11388 13744
rect 11334 13424 11390 13433
rect 11334 13359 11390 13368
rect 11348 11898 11376 13359
rect 11440 13258 11468 14010
rect 11532 13530 11560 14447
rect 11624 14113 11652 15014
rect 11716 14958 11744 19246
rect 11956 18524 12252 18544
rect 12012 18522 12036 18524
rect 12092 18522 12116 18524
rect 12172 18522 12196 18524
rect 12034 18470 12036 18522
rect 12098 18470 12110 18522
rect 12172 18470 12174 18522
rect 12012 18468 12036 18470
rect 12092 18468 12116 18470
rect 12172 18468 12196 18470
rect 11956 18448 12252 18468
rect 12440 18080 12492 18086
rect 12440 18022 12492 18028
rect 11956 17436 12252 17456
rect 12012 17434 12036 17436
rect 12092 17434 12116 17436
rect 12172 17434 12196 17436
rect 12034 17382 12036 17434
rect 12098 17382 12110 17434
rect 12172 17382 12174 17434
rect 12012 17380 12036 17382
rect 12092 17380 12116 17382
rect 12172 17380 12196 17382
rect 11956 17360 12252 17380
rect 12256 17128 12308 17134
rect 12256 17070 12308 17076
rect 12268 16726 12296 17070
rect 12348 16992 12400 16998
rect 12348 16934 12400 16940
rect 12256 16720 12308 16726
rect 12256 16662 12308 16668
rect 11956 16348 12252 16368
rect 12012 16346 12036 16348
rect 12092 16346 12116 16348
rect 12172 16346 12196 16348
rect 12034 16294 12036 16346
rect 12098 16294 12110 16346
rect 12172 16294 12174 16346
rect 12012 16292 12036 16294
rect 12092 16292 12116 16294
rect 12172 16292 12196 16294
rect 11956 16272 12252 16292
rect 12164 15972 12216 15978
rect 12164 15914 12216 15920
rect 12176 15502 12204 15914
rect 12360 15910 12388 16934
rect 12348 15904 12400 15910
rect 12348 15846 12400 15852
rect 11796 15496 11848 15502
rect 11796 15438 11848 15444
rect 12164 15496 12216 15502
rect 12164 15438 12216 15444
rect 11704 14952 11756 14958
rect 11704 14894 11756 14900
rect 11808 14822 11836 15438
rect 12360 15366 12388 15846
rect 12348 15360 12400 15366
rect 12348 15302 12400 15308
rect 11956 15260 12252 15280
rect 12012 15258 12036 15260
rect 12092 15258 12116 15260
rect 12172 15258 12196 15260
rect 12034 15206 12036 15258
rect 12098 15206 12110 15258
rect 12172 15206 12174 15258
rect 12012 15204 12036 15206
rect 12092 15204 12116 15206
rect 12172 15204 12196 15206
rect 11956 15184 12252 15204
rect 11796 14816 11848 14822
rect 11796 14758 11848 14764
rect 11888 14816 11940 14822
rect 11888 14758 11940 14764
rect 11704 14408 11756 14414
rect 11704 14350 11756 14356
rect 11610 14104 11666 14113
rect 11610 14039 11666 14048
rect 11612 13728 11664 13734
rect 11612 13670 11664 13676
rect 11520 13524 11572 13530
rect 11520 13466 11572 13472
rect 11624 13462 11652 13670
rect 11612 13456 11664 13462
rect 11612 13398 11664 13404
rect 11520 13320 11572 13326
rect 11520 13262 11572 13268
rect 11428 13252 11480 13258
rect 11428 13194 11480 13200
rect 11532 12442 11560 13262
rect 11624 12986 11652 13398
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 11612 12776 11664 12782
rect 11612 12718 11664 12724
rect 11520 12436 11572 12442
rect 11520 12378 11572 12384
rect 11624 12238 11652 12718
rect 11716 12714 11744 14350
rect 11808 13190 11836 14758
rect 11900 13326 11928 14758
rect 11956 14172 12252 14192
rect 12012 14170 12036 14172
rect 12092 14170 12116 14172
rect 12172 14170 12196 14172
rect 12034 14118 12036 14170
rect 12098 14118 12110 14170
rect 12172 14118 12174 14170
rect 12012 14116 12036 14118
rect 12092 14116 12116 14118
rect 12172 14116 12196 14118
rect 11956 14096 12252 14116
rect 11980 13796 12032 13802
rect 11980 13738 12032 13744
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 11796 13184 11848 13190
rect 11992 13172 12020 13738
rect 11796 13126 11848 13132
rect 11900 13144 12020 13172
rect 11796 12912 11848 12918
rect 11796 12854 11848 12860
rect 11704 12708 11756 12714
rect 11704 12650 11756 12656
rect 11808 12238 11836 12854
rect 11900 12782 11928 13144
rect 11956 13084 12252 13104
rect 12012 13082 12036 13084
rect 12092 13082 12116 13084
rect 12172 13082 12196 13084
rect 12034 13030 12036 13082
rect 12098 13030 12110 13082
rect 12172 13030 12174 13082
rect 12012 13028 12036 13030
rect 12092 13028 12116 13030
rect 12172 13028 12196 13030
rect 11956 13008 12252 13028
rect 12360 12986 12388 15302
rect 12348 12980 12400 12986
rect 12348 12922 12400 12928
rect 11888 12776 11940 12782
rect 11888 12718 11940 12724
rect 12072 12708 12124 12714
rect 12072 12650 12124 12656
rect 11888 12640 11940 12646
rect 11888 12582 11940 12588
rect 11900 12374 11928 12582
rect 11888 12368 11940 12374
rect 11888 12310 11940 12316
rect 11612 12232 11664 12238
rect 11612 12174 11664 12180
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 11336 11892 11388 11898
rect 11336 11834 11388 11840
rect 11336 11144 11388 11150
rect 11336 11086 11388 11092
rect 11348 10470 11376 11086
rect 11336 10464 11388 10470
rect 11336 10406 11388 10412
rect 11348 9110 11376 10406
rect 11624 9518 11652 12174
rect 11808 11354 11836 12174
rect 11900 11830 11928 12310
rect 12084 12238 12112 12650
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 11956 11996 12252 12016
rect 12012 11994 12036 11996
rect 12092 11994 12116 11996
rect 12172 11994 12196 11996
rect 12034 11942 12036 11994
rect 12098 11942 12110 11994
rect 12172 11942 12174 11994
rect 12012 11940 12036 11942
rect 12092 11940 12116 11942
rect 12172 11940 12196 11942
rect 11956 11920 12252 11940
rect 12348 11892 12400 11898
rect 12348 11834 12400 11840
rect 11888 11824 11940 11830
rect 11888 11766 11940 11772
rect 11796 11348 11848 11354
rect 11796 11290 11848 11296
rect 12360 11286 12388 11834
rect 12348 11280 12400 11286
rect 12348 11222 12400 11228
rect 11956 10908 12252 10928
rect 12012 10906 12036 10908
rect 12092 10906 12116 10908
rect 12172 10906 12196 10908
rect 12034 10854 12036 10906
rect 12098 10854 12110 10906
rect 12172 10854 12174 10906
rect 12012 10852 12036 10854
rect 12092 10852 12116 10854
rect 12172 10852 12196 10854
rect 11956 10832 12252 10852
rect 12360 10810 12388 11222
rect 12348 10804 12400 10810
rect 12348 10746 12400 10752
rect 12452 10554 12480 18022
rect 12544 17882 12572 21542
rect 12714 21520 12770 21542
rect 16224 21542 16450 21570
rect 13268 19304 13320 19310
rect 13268 19246 13320 19252
rect 12808 18828 12860 18834
rect 12808 18770 12860 18776
rect 12624 18624 12676 18630
rect 12624 18566 12676 18572
rect 12532 17876 12584 17882
rect 12532 17818 12584 17824
rect 12532 16992 12584 16998
rect 12532 16934 12584 16940
rect 12544 13938 12572 16934
rect 12636 15434 12664 18566
rect 12820 18154 12848 18770
rect 13084 18284 13136 18290
rect 13084 18226 13136 18232
rect 12808 18148 12860 18154
rect 12808 18090 12860 18096
rect 12716 18080 12768 18086
rect 12716 18022 12768 18028
rect 12728 17338 12756 18022
rect 12992 17740 13044 17746
rect 12992 17682 13044 17688
rect 12716 17332 12768 17338
rect 12716 17274 12768 17280
rect 13004 17202 13032 17682
rect 12992 17196 13044 17202
rect 12992 17138 13044 17144
rect 12808 16992 12860 16998
rect 12808 16934 12860 16940
rect 12716 16652 12768 16658
rect 12716 16594 12768 16600
rect 12728 16250 12756 16594
rect 12716 16244 12768 16250
rect 12716 16186 12768 16192
rect 12728 15706 12756 16186
rect 12716 15700 12768 15706
rect 12716 15642 12768 15648
rect 12624 15428 12676 15434
rect 12624 15370 12676 15376
rect 12624 15088 12676 15094
rect 12624 15030 12676 15036
rect 12532 13932 12584 13938
rect 12532 13874 12584 13880
rect 12544 13530 12572 13874
rect 12532 13524 12584 13530
rect 12532 13466 12584 13472
rect 12532 12708 12584 12714
rect 12532 12650 12584 12656
rect 12544 12170 12572 12650
rect 12532 12164 12584 12170
rect 12532 12106 12584 12112
rect 12636 12102 12664 15030
rect 12716 14544 12768 14550
rect 12716 14486 12768 14492
rect 12728 14074 12756 14486
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 12820 13814 12848 16934
rect 12992 15496 13044 15502
rect 12992 15438 13044 15444
rect 12900 14816 12952 14822
rect 12900 14758 12952 14764
rect 12912 14550 12940 14758
rect 12900 14544 12952 14550
rect 12900 14486 12952 14492
rect 12728 13786 12848 13814
rect 12912 13802 12940 14486
rect 13004 14414 13032 15438
rect 13096 14521 13124 18226
rect 13176 16652 13228 16658
rect 13176 16594 13228 16600
rect 13188 16046 13216 16594
rect 13176 16040 13228 16046
rect 13176 15982 13228 15988
rect 13280 15892 13308 19246
rect 15622 19068 15918 19088
rect 15678 19066 15702 19068
rect 15758 19066 15782 19068
rect 15838 19066 15862 19068
rect 15700 19014 15702 19066
rect 15764 19014 15776 19066
rect 15838 19014 15840 19066
rect 15678 19012 15702 19014
rect 15758 19012 15782 19014
rect 15838 19012 15862 19014
rect 15622 18992 15918 19012
rect 13728 18828 13780 18834
rect 13728 18770 13780 18776
rect 13740 18290 13768 18770
rect 13728 18284 13780 18290
rect 13728 18226 13780 18232
rect 14556 18216 14608 18222
rect 14556 18158 14608 18164
rect 14740 18216 14792 18222
rect 14740 18158 14792 18164
rect 13728 18148 13780 18154
rect 13728 18090 13780 18096
rect 14372 18148 14424 18154
rect 14372 18090 14424 18096
rect 13636 17196 13688 17202
rect 13636 17138 13688 17144
rect 13360 16720 13412 16726
rect 13360 16662 13412 16668
rect 13188 15864 13308 15892
rect 13082 14512 13138 14521
rect 13082 14447 13138 14456
rect 12992 14408 13044 14414
rect 12992 14350 13044 14356
rect 12900 13796 12952 13802
rect 12624 12096 12676 12102
rect 12624 12038 12676 12044
rect 12728 11665 12756 13786
rect 12900 13738 12952 13744
rect 12900 13252 12952 13258
rect 12900 13194 12952 13200
rect 12808 13184 12860 13190
rect 12808 13126 12860 13132
rect 12820 12850 12848 13126
rect 12808 12844 12860 12850
rect 12808 12786 12860 12792
rect 12714 11656 12770 11665
rect 12714 11591 12770 11600
rect 12624 11076 12676 11082
rect 12624 11018 12676 11024
rect 12360 10526 12480 10554
rect 12532 10532 12584 10538
rect 11796 9920 11848 9926
rect 11796 9862 11848 9868
rect 11612 9512 11664 9518
rect 11612 9454 11664 9460
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11336 9104 11388 9110
rect 11336 9046 11388 9052
rect 11244 8900 11296 8906
rect 11244 8842 11296 8848
rect 11624 8294 11652 9318
rect 11612 8288 11664 8294
rect 11612 8230 11664 8236
rect 11624 8022 11652 8230
rect 11612 8016 11664 8022
rect 11612 7958 11664 7964
rect 11152 7948 11204 7954
rect 11152 7890 11204 7896
rect 11164 7002 11192 7890
rect 11428 7404 11480 7410
rect 11428 7346 11480 7352
rect 11336 7336 11388 7342
rect 11336 7278 11388 7284
rect 11152 6996 11204 7002
rect 11152 6938 11204 6944
rect 11244 6112 11296 6118
rect 11244 6054 11296 6060
rect 11256 5846 11284 6054
rect 11244 5840 11296 5846
rect 11244 5782 11296 5788
rect 11348 5166 11376 7278
rect 11440 6934 11468 7346
rect 11520 7268 11572 7274
rect 11520 7210 11572 7216
rect 11532 7002 11560 7210
rect 11624 7206 11652 7958
rect 11612 7200 11664 7206
rect 11612 7142 11664 7148
rect 11808 7018 11836 9862
rect 11956 9820 12252 9840
rect 12012 9818 12036 9820
rect 12092 9818 12116 9820
rect 12172 9818 12196 9820
rect 12034 9766 12036 9818
rect 12098 9766 12110 9818
rect 12172 9766 12174 9818
rect 12012 9764 12036 9766
rect 12092 9764 12116 9766
rect 12172 9764 12196 9766
rect 11956 9744 12252 9764
rect 12360 9178 12388 10526
rect 12532 10474 12584 10480
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12452 9926 12480 10406
rect 12544 10266 12572 10474
rect 12532 10260 12584 10266
rect 12532 10202 12584 10208
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12452 9722 12480 9862
rect 12440 9716 12492 9722
rect 12440 9658 12492 9664
rect 12440 9512 12492 9518
rect 12440 9454 12492 9460
rect 12348 9172 12400 9178
rect 12348 9114 12400 9120
rect 11956 8732 12252 8752
rect 12012 8730 12036 8732
rect 12092 8730 12116 8732
rect 12172 8730 12196 8732
rect 12034 8678 12036 8730
rect 12098 8678 12110 8730
rect 12172 8678 12174 8730
rect 12012 8676 12036 8678
rect 12092 8676 12116 8678
rect 12172 8676 12196 8678
rect 11956 8656 12252 8676
rect 11888 7812 11940 7818
rect 11888 7754 11940 7760
rect 11900 7478 11928 7754
rect 11956 7644 12252 7664
rect 12012 7642 12036 7644
rect 12092 7642 12116 7644
rect 12172 7642 12196 7644
rect 12034 7590 12036 7642
rect 12098 7590 12110 7642
rect 12172 7590 12174 7642
rect 12012 7588 12036 7590
rect 12092 7588 12116 7590
rect 12172 7588 12196 7590
rect 11956 7568 12252 7588
rect 11888 7472 11940 7478
rect 11888 7414 11940 7420
rect 11520 6996 11572 7002
rect 11808 6990 11928 7018
rect 11520 6938 11572 6944
rect 11428 6928 11480 6934
rect 11428 6870 11480 6876
rect 11796 6928 11848 6934
rect 11796 6870 11848 6876
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 11612 6724 11664 6730
rect 11612 6666 11664 6672
rect 11624 6458 11652 6666
rect 11520 6452 11572 6458
rect 11520 6394 11572 6400
rect 11612 6452 11664 6458
rect 11612 6394 11664 6400
rect 11532 5710 11560 6394
rect 11612 6112 11664 6118
rect 11612 6054 11664 6060
rect 11624 5914 11652 6054
rect 11716 5914 11744 6734
rect 11808 6118 11836 6870
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11612 5908 11664 5914
rect 11612 5850 11664 5856
rect 11704 5908 11756 5914
rect 11704 5850 11756 5856
rect 11520 5704 11572 5710
rect 11520 5646 11572 5652
rect 11520 5228 11572 5234
rect 11520 5170 11572 5176
rect 11336 5160 11388 5166
rect 11336 5102 11388 5108
rect 11244 4820 11296 4826
rect 11348 4808 11376 5102
rect 11428 5092 11480 5098
rect 11428 5034 11480 5040
rect 11296 4780 11376 4808
rect 11244 4762 11296 4768
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 11152 4072 11204 4078
rect 11152 4014 11204 4020
rect 10600 3732 10652 3738
rect 10600 3674 10652 3680
rect 11164 3641 11192 4014
rect 11150 3632 11206 3641
rect 11150 3567 11206 3576
rect 11164 3534 11192 3567
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 10876 3120 10928 3126
rect 10876 3062 10928 3068
rect 9770 76 9772 128
rect 9824 76 9826 128
rect 8666 0 8722 54
rect 9770 0 9826 76
rect 10508 128 10560 134
rect 10508 70 10560 76
rect 10888 82 10916 3062
rect 11440 2990 11468 5034
rect 11532 4758 11560 5170
rect 11520 4752 11572 4758
rect 11520 4694 11572 4700
rect 11704 4752 11756 4758
rect 11704 4694 11756 4700
rect 11716 3942 11744 4694
rect 11796 4140 11848 4146
rect 11796 4082 11848 4088
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 11612 3664 11664 3670
rect 11612 3606 11664 3612
rect 11428 2984 11480 2990
rect 11428 2926 11480 2932
rect 11624 2650 11652 3606
rect 11716 3194 11744 3878
rect 11808 3534 11836 4082
rect 11796 3528 11848 3534
rect 11796 3470 11848 3476
rect 11704 3188 11756 3194
rect 11704 3130 11756 3136
rect 11612 2644 11664 2650
rect 11612 2586 11664 2592
rect 11808 2514 11836 3470
rect 11796 2508 11848 2514
rect 11796 2450 11848 2456
rect 10966 82 11022 480
rect 10888 54 11022 82
rect 11900 82 11928 6990
rect 11956 6556 12252 6576
rect 12012 6554 12036 6556
rect 12092 6554 12116 6556
rect 12172 6554 12196 6556
rect 12034 6502 12036 6554
rect 12098 6502 12110 6554
rect 12172 6502 12174 6554
rect 12012 6500 12036 6502
rect 12092 6500 12116 6502
rect 12172 6500 12196 6502
rect 11956 6480 12252 6500
rect 12348 5840 12400 5846
rect 12348 5782 12400 5788
rect 11956 5468 12252 5488
rect 12012 5466 12036 5468
rect 12092 5466 12116 5468
rect 12172 5466 12196 5468
rect 12034 5414 12036 5466
rect 12098 5414 12110 5466
rect 12172 5414 12174 5466
rect 12012 5412 12036 5414
rect 12092 5412 12116 5414
rect 12172 5412 12196 5414
rect 11956 5392 12252 5412
rect 12360 5370 12388 5782
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12360 5030 12388 5306
rect 12348 5024 12400 5030
rect 12348 4966 12400 4972
rect 12360 4826 12388 4966
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 12348 4616 12400 4622
rect 12348 4558 12400 4564
rect 11956 4380 12252 4400
rect 12012 4378 12036 4380
rect 12092 4378 12116 4380
rect 12172 4378 12196 4380
rect 12034 4326 12036 4378
rect 12098 4326 12110 4378
rect 12172 4326 12174 4378
rect 12012 4324 12036 4326
rect 12092 4324 12116 4326
rect 12172 4324 12196 4326
rect 11956 4304 12252 4324
rect 12360 4154 12388 4558
rect 12268 4126 12388 4154
rect 12268 3670 12296 4126
rect 12346 4040 12402 4049
rect 12346 3975 12348 3984
rect 12400 3975 12402 3984
rect 12348 3946 12400 3952
rect 12360 3670 12388 3946
rect 12256 3664 12308 3670
rect 12256 3606 12308 3612
rect 12348 3664 12400 3670
rect 12348 3606 12400 3612
rect 11956 3292 12252 3312
rect 12012 3290 12036 3292
rect 12092 3290 12116 3292
rect 12172 3290 12196 3292
rect 12034 3238 12036 3290
rect 12098 3238 12110 3290
rect 12172 3238 12174 3290
rect 12012 3236 12036 3238
rect 12092 3236 12116 3238
rect 12172 3236 12196 3238
rect 11956 3216 12252 3236
rect 12452 2990 12480 9454
rect 12544 8974 12572 10202
rect 12636 9110 12664 11018
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 12624 9104 12676 9110
rect 12624 9046 12676 9052
rect 12532 8968 12584 8974
rect 12532 8910 12584 8916
rect 12636 8090 12664 9046
rect 12728 8634 12756 10950
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 12820 9654 12848 9998
rect 12808 9648 12860 9654
rect 12808 9590 12860 9596
rect 12912 8650 12940 13194
rect 13084 11688 13136 11694
rect 13084 11630 13136 11636
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 12716 8628 12768 8634
rect 12716 8570 12768 8576
rect 12820 8622 12940 8650
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12820 7954 12848 8622
rect 12900 8560 12952 8566
rect 12900 8502 12952 8508
rect 12912 8090 12940 8502
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 12808 7948 12860 7954
rect 12808 7890 12860 7896
rect 12624 7472 12676 7478
rect 12624 7414 12676 7420
rect 12636 7274 12664 7414
rect 12532 7268 12584 7274
rect 12532 7210 12584 7216
rect 12624 7268 12676 7274
rect 12624 7210 12676 7216
rect 12544 6730 12572 7210
rect 13004 6934 13032 10610
rect 12992 6928 13044 6934
rect 12992 6870 13044 6876
rect 12808 6792 12860 6798
rect 12808 6734 12860 6740
rect 12532 6724 12584 6730
rect 12532 6666 12584 6672
rect 12716 5704 12768 5710
rect 12716 5646 12768 5652
rect 12728 4826 12756 5646
rect 12820 5234 12848 6734
rect 13004 6390 13032 6870
rect 13096 6798 13124 11630
rect 13188 11370 13216 15864
rect 13268 15632 13320 15638
rect 13268 15574 13320 15580
rect 13280 14822 13308 15574
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 13268 14476 13320 14482
rect 13268 14418 13320 14424
rect 13280 13433 13308 14418
rect 13266 13424 13322 13433
rect 13266 13359 13322 13368
rect 13372 11626 13400 16662
rect 13544 16584 13596 16590
rect 13544 16526 13596 16532
rect 13452 15972 13504 15978
rect 13452 15914 13504 15920
rect 13464 15570 13492 15914
rect 13452 15564 13504 15570
rect 13452 15506 13504 15512
rect 13556 15026 13584 16526
rect 13648 16182 13676 17138
rect 13636 16176 13688 16182
rect 13636 16118 13688 16124
rect 13636 15428 13688 15434
rect 13636 15370 13688 15376
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 13556 14618 13584 14962
rect 13544 14612 13596 14618
rect 13544 14554 13596 14560
rect 13452 14408 13504 14414
rect 13452 14350 13504 14356
rect 13464 13569 13492 14350
rect 13450 13560 13506 13569
rect 13450 13495 13506 13504
rect 13452 13388 13504 13394
rect 13452 13330 13504 13336
rect 13464 12986 13492 13330
rect 13544 13320 13596 13326
rect 13544 13262 13596 13268
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 13556 12442 13584 13262
rect 13544 12436 13596 12442
rect 13544 12378 13596 12384
rect 13556 11762 13584 12378
rect 13544 11756 13596 11762
rect 13544 11698 13596 11704
rect 13452 11688 13504 11694
rect 13452 11630 13504 11636
rect 13360 11620 13412 11626
rect 13360 11562 13412 11568
rect 13188 11342 13400 11370
rect 13268 11280 13320 11286
rect 13268 11222 13320 11228
rect 13280 11082 13308 11222
rect 13268 11076 13320 11082
rect 13268 11018 13320 11024
rect 13280 10810 13308 11018
rect 13268 10804 13320 10810
rect 13268 10746 13320 10752
rect 13268 10192 13320 10198
rect 13268 10134 13320 10140
rect 13176 9376 13228 9382
rect 13280 9364 13308 10134
rect 13228 9336 13308 9364
rect 13176 9318 13228 9324
rect 13372 8498 13400 11342
rect 13464 9994 13492 11630
rect 13648 11257 13676 15370
rect 13740 14482 13768 18090
rect 14188 18080 14240 18086
rect 14188 18022 14240 18028
rect 14200 17785 14228 18022
rect 14186 17776 14242 17785
rect 14096 17740 14148 17746
rect 14186 17711 14242 17720
rect 14096 17682 14148 17688
rect 13820 17536 13872 17542
rect 13820 17478 13872 17484
rect 13832 16130 13860 17478
rect 14108 17338 14136 17682
rect 14188 17536 14240 17542
rect 14188 17478 14240 17484
rect 13912 17332 13964 17338
rect 13912 17274 13964 17280
rect 14096 17332 14148 17338
rect 14096 17274 14148 17280
rect 13924 16250 13952 17274
rect 14108 17066 14136 17274
rect 14096 17060 14148 17066
rect 14096 17002 14148 17008
rect 14004 16992 14056 16998
rect 14004 16934 14056 16940
rect 13912 16244 13964 16250
rect 13912 16186 13964 16192
rect 13832 16102 13952 16130
rect 13728 14476 13780 14482
rect 13728 14418 13780 14424
rect 13726 14240 13782 14249
rect 13726 14175 13782 14184
rect 13740 13462 13768 14175
rect 13924 13530 13952 16102
rect 13912 13524 13964 13530
rect 13912 13466 13964 13472
rect 13728 13456 13780 13462
rect 13728 13398 13780 13404
rect 13912 13388 13964 13394
rect 13912 13330 13964 13336
rect 13728 12980 13780 12986
rect 13728 12922 13780 12928
rect 13634 11248 13690 11257
rect 13634 11183 13690 11192
rect 13636 11144 13688 11150
rect 13636 11086 13688 11092
rect 13544 10736 13596 10742
rect 13544 10678 13596 10684
rect 13452 9988 13504 9994
rect 13452 9930 13504 9936
rect 13556 9654 13584 10678
rect 13648 9994 13676 11086
rect 13740 10810 13768 12922
rect 13924 12850 13952 13330
rect 13912 12844 13964 12850
rect 13912 12786 13964 12792
rect 13924 10849 13952 12786
rect 14016 11354 14044 16934
rect 14094 16552 14150 16561
rect 14094 16487 14150 16496
rect 14108 16182 14136 16487
rect 14096 16176 14148 16182
rect 14096 16118 14148 16124
rect 14096 14476 14148 14482
rect 14096 14418 14148 14424
rect 14108 14074 14136 14418
rect 14096 14068 14148 14074
rect 14096 14010 14148 14016
rect 14096 13796 14148 13802
rect 14096 13738 14148 13744
rect 14108 13462 14136 13738
rect 14096 13456 14148 13462
rect 14096 13398 14148 13404
rect 14108 12374 14136 13398
rect 14096 12368 14148 12374
rect 14096 12310 14148 12316
rect 14108 11898 14136 12310
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 14108 11626 14136 11834
rect 14200 11694 14228 17478
rect 14280 16448 14332 16454
rect 14280 16390 14332 16396
rect 14292 16046 14320 16390
rect 14280 16040 14332 16046
rect 14280 15982 14332 15988
rect 14292 15881 14320 15982
rect 14278 15872 14334 15881
rect 14278 15807 14334 15816
rect 14384 13814 14412 18090
rect 14568 16697 14596 18158
rect 14554 16688 14610 16697
rect 14554 16623 14610 16632
rect 14752 16153 14780 18158
rect 15622 17980 15918 18000
rect 15678 17978 15702 17980
rect 15758 17978 15782 17980
rect 15838 17978 15862 17980
rect 15700 17926 15702 17978
rect 15764 17926 15776 17978
rect 15838 17926 15840 17978
rect 15678 17924 15702 17926
rect 15758 17924 15782 17926
rect 15838 17924 15862 17926
rect 15622 17904 15918 17924
rect 15476 17740 15528 17746
rect 15476 17682 15528 17688
rect 15488 17270 15516 17682
rect 16120 17536 16172 17542
rect 16120 17478 16172 17484
rect 15476 17264 15528 17270
rect 15476 17206 15528 17212
rect 15384 16992 15436 16998
rect 15384 16934 15436 16940
rect 15108 16448 15160 16454
rect 15108 16390 15160 16396
rect 14738 16144 14794 16153
rect 14648 16108 14700 16114
rect 14738 16079 14794 16088
rect 14648 16050 14700 16056
rect 14292 13786 14412 13814
rect 14188 11688 14240 11694
rect 14188 11630 14240 11636
rect 14096 11620 14148 11626
rect 14096 11562 14148 11568
rect 14004 11348 14056 11354
rect 14004 11290 14056 11296
rect 13910 10840 13966 10849
rect 13728 10804 13780 10810
rect 13910 10775 13966 10784
rect 13728 10746 13780 10752
rect 13740 10538 13768 10746
rect 14096 10668 14148 10674
rect 14096 10610 14148 10616
rect 13728 10532 13780 10538
rect 13728 10474 13780 10480
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 13832 9994 13860 10406
rect 13636 9988 13688 9994
rect 13636 9930 13688 9936
rect 13820 9988 13872 9994
rect 13820 9930 13872 9936
rect 13544 9648 13596 9654
rect 13544 9590 13596 9596
rect 13648 9586 13676 9930
rect 14108 9926 14136 10610
rect 13728 9920 13780 9926
rect 13728 9862 13780 9868
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 13636 9580 13688 9586
rect 13636 9522 13688 9528
rect 13648 9178 13676 9522
rect 13740 9450 13768 9862
rect 14108 9625 14136 9862
rect 14094 9616 14150 9625
rect 14094 9551 14150 9560
rect 13728 9444 13780 9450
rect 13728 9386 13780 9392
rect 13636 9172 13688 9178
rect 13636 9114 13688 9120
rect 14096 9036 14148 9042
rect 14096 8978 14148 8984
rect 14108 8945 14136 8978
rect 14094 8936 14150 8945
rect 14094 8871 14150 8880
rect 14108 8634 14136 8871
rect 14096 8628 14148 8634
rect 14096 8570 14148 8576
rect 14292 8498 14320 13786
rect 14372 13524 14424 13530
rect 14372 13466 14424 13472
rect 14384 12850 14412 13466
rect 14372 12844 14424 12850
rect 14372 12786 14424 12792
rect 14464 12708 14516 12714
rect 14464 12650 14516 12656
rect 14476 12442 14504 12650
rect 14464 12436 14516 12442
rect 14464 12378 14516 12384
rect 14476 11898 14504 12378
rect 14556 12232 14608 12238
rect 14556 12174 14608 12180
rect 14464 11892 14516 11898
rect 14464 11834 14516 11840
rect 14568 11558 14596 12174
rect 14660 11558 14688 16050
rect 14752 13569 14780 16079
rect 14924 15972 14976 15978
rect 14924 15914 14976 15920
rect 14738 13560 14794 13569
rect 14738 13495 14794 13504
rect 14556 11552 14608 11558
rect 14556 11494 14608 11500
rect 14648 11552 14700 11558
rect 14648 11494 14700 11500
rect 14372 10736 14424 10742
rect 14372 10678 14424 10684
rect 14384 9722 14412 10678
rect 14568 10674 14596 11494
rect 14556 10668 14608 10674
rect 14556 10610 14608 10616
rect 14556 10192 14608 10198
rect 14556 10134 14608 10140
rect 14568 9722 14596 10134
rect 14372 9716 14424 9722
rect 14372 9658 14424 9664
rect 14556 9716 14608 9722
rect 14556 9658 14608 9664
rect 13360 8492 13412 8498
rect 13360 8434 13412 8440
rect 14280 8492 14332 8498
rect 14280 8434 14332 8440
rect 13176 7880 13228 7886
rect 13176 7822 13228 7828
rect 13188 7546 13216 7822
rect 13176 7540 13228 7546
rect 13176 7482 13228 7488
rect 13372 7410 13400 8434
rect 13544 8288 13596 8294
rect 13544 8230 13596 8236
rect 13556 7750 13584 8230
rect 14292 8090 14320 8434
rect 14752 8430 14780 13495
rect 14936 12186 14964 15914
rect 15016 14408 15068 14414
rect 15016 14350 15068 14356
rect 15028 13190 15056 14350
rect 15016 13184 15068 13190
rect 15016 13126 15068 13132
rect 15028 12850 15056 13126
rect 15016 12844 15068 12850
rect 15016 12786 15068 12792
rect 14936 12158 15056 12186
rect 14924 12096 14976 12102
rect 14924 12038 14976 12044
rect 14936 11830 14964 12038
rect 14924 11824 14976 11830
rect 14924 11766 14976 11772
rect 14740 8424 14792 8430
rect 14740 8366 14792 8372
rect 14280 8084 14332 8090
rect 14280 8026 14332 8032
rect 14004 8016 14056 8022
rect 14004 7958 14056 7964
rect 13544 7744 13596 7750
rect 13544 7686 13596 7692
rect 13452 7472 13504 7478
rect 13452 7414 13504 7420
rect 13360 7404 13412 7410
rect 13360 7346 13412 7352
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 12992 6384 13044 6390
rect 12992 6326 13044 6332
rect 12900 6316 12952 6322
rect 12900 6258 12952 6264
rect 12912 5710 12940 6258
rect 13096 5846 13124 6734
rect 13084 5840 13136 5846
rect 13084 5782 13136 5788
rect 12900 5704 12952 5710
rect 12900 5646 12952 5652
rect 12808 5228 12860 5234
rect 12808 5170 12860 5176
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 12912 4146 12940 5646
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 13268 4752 13320 4758
rect 13268 4694 13320 4700
rect 13084 4616 13136 4622
rect 13084 4558 13136 4564
rect 13096 4214 13124 4558
rect 13084 4208 13136 4214
rect 13084 4150 13136 4156
rect 12900 4140 12952 4146
rect 12900 4082 12952 4088
rect 13280 3942 13308 4694
rect 13372 4622 13400 5170
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13268 3936 13320 3942
rect 13268 3878 13320 3884
rect 13360 3460 13412 3466
rect 13360 3402 13412 3408
rect 13082 3360 13138 3369
rect 13082 3295 13138 3304
rect 13096 3194 13124 3295
rect 13084 3188 13136 3194
rect 13084 3130 13136 3136
rect 13096 2990 13124 3130
rect 12440 2984 12492 2990
rect 12440 2926 12492 2932
rect 13084 2984 13136 2990
rect 13084 2926 13136 2932
rect 12072 2848 12124 2854
rect 12072 2790 12124 2796
rect 13268 2848 13320 2854
rect 13268 2790 13320 2796
rect 12084 2650 12112 2790
rect 12072 2644 12124 2650
rect 12072 2586 12124 2592
rect 13280 2582 13308 2790
rect 13268 2576 13320 2582
rect 13268 2518 13320 2524
rect 13372 2514 13400 3402
rect 13360 2508 13412 2514
rect 13360 2450 13412 2456
rect 11956 2204 12252 2224
rect 12012 2202 12036 2204
rect 12092 2202 12116 2204
rect 12172 2202 12196 2204
rect 12034 2150 12036 2202
rect 12098 2150 12110 2202
rect 12172 2150 12174 2202
rect 12012 2148 12036 2150
rect 12092 2148 12116 2150
rect 12172 2148 12196 2150
rect 11956 2128 12252 2148
rect 12070 82 12126 480
rect 11900 54 12126 82
rect 10966 0 11022 54
rect 12070 0 12126 54
rect 13266 82 13322 480
rect 13464 82 13492 7414
rect 13556 6934 13584 7686
rect 14016 7206 14044 7958
rect 14752 7478 14780 8366
rect 15028 7954 15056 12158
rect 15120 11762 15148 16390
rect 15396 15502 15424 16934
rect 15488 16658 15516 17206
rect 16028 17060 16080 17066
rect 16028 17002 16080 17008
rect 15622 16892 15918 16912
rect 15678 16890 15702 16892
rect 15758 16890 15782 16892
rect 15838 16890 15862 16892
rect 15700 16838 15702 16890
rect 15764 16838 15776 16890
rect 15838 16838 15840 16890
rect 15678 16836 15702 16838
rect 15758 16836 15782 16838
rect 15838 16836 15862 16838
rect 15622 16816 15918 16836
rect 15476 16652 15528 16658
rect 15476 16594 15528 16600
rect 15488 16114 15516 16594
rect 16040 16522 16068 17002
rect 16028 16516 16080 16522
rect 16028 16458 16080 16464
rect 15936 16448 15988 16454
rect 15936 16390 15988 16396
rect 15476 16108 15528 16114
rect 15476 16050 15528 16056
rect 15622 15804 15918 15824
rect 15678 15802 15702 15804
rect 15758 15802 15782 15804
rect 15838 15802 15862 15804
rect 15700 15750 15702 15802
rect 15764 15750 15776 15802
rect 15838 15750 15840 15802
rect 15678 15748 15702 15750
rect 15758 15748 15782 15750
rect 15838 15748 15862 15750
rect 15622 15728 15918 15748
rect 15476 15632 15528 15638
rect 15476 15574 15528 15580
rect 15384 15496 15436 15502
rect 15384 15438 15436 15444
rect 15396 15162 15424 15438
rect 15488 15162 15516 15574
rect 15384 15156 15436 15162
rect 15384 15098 15436 15104
rect 15476 15156 15528 15162
rect 15476 15098 15528 15104
rect 15476 15020 15528 15026
rect 15476 14962 15528 14968
rect 15200 14952 15252 14958
rect 15252 14929 15332 14940
rect 15252 14920 15346 14929
rect 15252 14912 15290 14920
rect 15200 14894 15252 14900
rect 15290 14855 15346 14864
rect 15292 14612 15344 14618
rect 15292 14554 15344 14560
rect 15200 14068 15252 14074
rect 15200 14010 15252 14016
rect 15212 13705 15240 14010
rect 15198 13696 15254 13705
rect 15198 13631 15254 13640
rect 15198 13424 15254 13433
rect 15198 13359 15254 13368
rect 15212 13326 15240 13359
rect 15200 13320 15252 13326
rect 15200 13262 15252 13268
rect 15212 12442 15240 13262
rect 15304 12442 15332 14554
rect 15384 14544 15436 14550
rect 15384 14486 15436 14492
rect 15396 14006 15424 14486
rect 15488 14278 15516 14962
rect 15622 14716 15918 14736
rect 15678 14714 15702 14716
rect 15758 14714 15782 14716
rect 15838 14714 15862 14716
rect 15700 14662 15702 14714
rect 15764 14662 15776 14714
rect 15838 14662 15840 14714
rect 15678 14660 15702 14662
rect 15758 14660 15782 14662
rect 15838 14660 15862 14662
rect 15622 14640 15918 14660
rect 15948 14385 15976 16390
rect 16028 16040 16080 16046
rect 16028 15982 16080 15988
rect 16040 15638 16068 15982
rect 16028 15632 16080 15638
rect 16028 15574 16080 15580
rect 16040 15026 16068 15574
rect 16028 15020 16080 15026
rect 16028 14962 16080 14968
rect 16040 14550 16068 14962
rect 16028 14544 16080 14550
rect 16028 14486 16080 14492
rect 15934 14376 15990 14385
rect 15934 14311 15990 14320
rect 15476 14272 15528 14278
rect 15476 14214 15528 14220
rect 15384 14000 15436 14006
rect 15384 13942 15436 13948
rect 15384 13728 15436 13734
rect 15384 13670 15436 13676
rect 15396 13462 15424 13670
rect 15384 13456 15436 13462
rect 15384 13398 15436 13404
rect 15396 12986 15424 13398
rect 15488 13326 15516 14214
rect 16026 13696 16082 13705
rect 15948 13654 16026 13682
rect 15622 13628 15918 13648
rect 15678 13626 15702 13628
rect 15758 13626 15782 13628
rect 15838 13626 15862 13628
rect 15700 13574 15702 13626
rect 15764 13574 15776 13626
rect 15838 13574 15840 13626
rect 15678 13572 15702 13574
rect 15758 13572 15782 13574
rect 15838 13572 15862 13574
rect 15622 13552 15918 13572
rect 15476 13320 15528 13326
rect 15476 13262 15528 13268
rect 15384 12980 15436 12986
rect 15384 12922 15436 12928
rect 15200 12436 15252 12442
rect 15200 12378 15252 12384
rect 15292 12436 15344 12442
rect 15292 12378 15344 12384
rect 15108 11756 15160 11762
rect 15108 11698 15160 11704
rect 15120 11354 15148 11698
rect 15304 11354 15332 12378
rect 15488 12238 15516 13262
rect 15622 12540 15918 12560
rect 15678 12538 15702 12540
rect 15758 12538 15782 12540
rect 15838 12538 15862 12540
rect 15700 12486 15702 12538
rect 15764 12486 15776 12538
rect 15838 12486 15840 12538
rect 15678 12484 15702 12486
rect 15758 12484 15782 12486
rect 15838 12484 15862 12486
rect 15622 12464 15918 12484
rect 15476 12232 15528 12238
rect 15476 12174 15528 12180
rect 15488 11762 15516 12174
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 15622 11452 15918 11472
rect 15678 11450 15702 11452
rect 15758 11450 15782 11452
rect 15838 11450 15862 11452
rect 15700 11398 15702 11450
rect 15764 11398 15776 11450
rect 15838 11398 15840 11450
rect 15678 11396 15702 11398
rect 15758 11396 15782 11398
rect 15838 11396 15862 11398
rect 15622 11376 15918 11396
rect 15108 11348 15160 11354
rect 15108 11290 15160 11296
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15622 10364 15918 10384
rect 15678 10362 15702 10364
rect 15758 10362 15782 10364
rect 15838 10362 15862 10364
rect 15700 10310 15702 10362
rect 15764 10310 15776 10362
rect 15838 10310 15840 10362
rect 15678 10308 15702 10310
rect 15758 10308 15782 10310
rect 15838 10308 15862 10310
rect 15622 10288 15918 10308
rect 15292 10056 15344 10062
rect 15292 9998 15344 10004
rect 15304 9586 15332 9998
rect 15292 9580 15344 9586
rect 15292 9522 15344 9528
rect 15108 9512 15160 9518
rect 15108 9454 15160 9460
rect 15120 9178 15148 9454
rect 15384 9444 15436 9450
rect 15384 9386 15436 9392
rect 15108 9172 15160 9178
rect 15108 9114 15160 9120
rect 15292 8832 15344 8838
rect 15292 8774 15344 8780
rect 14924 7948 14976 7954
rect 14924 7890 14976 7896
rect 15016 7948 15068 7954
rect 15016 7890 15068 7896
rect 14936 7857 14964 7890
rect 14922 7848 14978 7857
rect 14922 7783 14978 7792
rect 15028 7478 15056 7890
rect 15200 7744 15252 7750
rect 15200 7686 15252 7692
rect 14740 7472 14792 7478
rect 14740 7414 14792 7420
rect 15016 7472 15068 7478
rect 15016 7414 15068 7420
rect 14752 7342 14780 7414
rect 14740 7336 14792 7342
rect 14740 7278 14792 7284
rect 15108 7336 15160 7342
rect 15108 7278 15160 7284
rect 14004 7200 14056 7206
rect 14004 7142 14056 7148
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 13544 6928 13596 6934
rect 13544 6870 13596 6876
rect 13556 6458 13584 6870
rect 13544 6452 13596 6458
rect 13544 6394 13596 6400
rect 14016 6168 14044 7142
rect 14096 6996 14148 7002
rect 14096 6938 14148 6944
rect 14108 6322 14136 6938
rect 14096 6316 14148 6322
rect 14096 6258 14148 6264
rect 14096 6180 14148 6186
rect 14016 6140 14096 6168
rect 14096 6122 14148 6128
rect 14108 5098 14136 6122
rect 14200 5778 14228 7142
rect 15120 7002 15148 7278
rect 15212 7177 15240 7686
rect 15198 7168 15254 7177
rect 15198 7103 15254 7112
rect 15108 6996 15160 7002
rect 15108 6938 15160 6944
rect 14648 6724 14700 6730
rect 14648 6666 14700 6672
rect 14188 5772 14240 5778
rect 14188 5714 14240 5720
rect 14200 5370 14228 5714
rect 14280 5568 14332 5574
rect 14280 5510 14332 5516
rect 14188 5364 14240 5370
rect 14188 5306 14240 5312
rect 14096 5092 14148 5098
rect 14096 5034 14148 5040
rect 14108 4486 14136 5034
rect 14200 4865 14228 5306
rect 14186 4856 14242 4865
rect 14186 4791 14242 4800
rect 14292 4729 14320 5510
rect 14278 4720 14334 4729
rect 14278 4655 14334 4664
rect 14096 4480 14148 4486
rect 14096 4422 14148 4428
rect 14108 3942 14136 4422
rect 14188 4004 14240 4010
rect 14188 3946 14240 3952
rect 14096 3936 14148 3942
rect 14096 3878 14148 3884
rect 14200 3738 14228 3946
rect 14188 3732 14240 3738
rect 14188 3674 14240 3680
rect 13820 3664 13872 3670
rect 13820 3606 13872 3612
rect 13832 2922 13860 3606
rect 13912 2984 13964 2990
rect 13912 2926 13964 2932
rect 13820 2916 13872 2922
rect 13820 2858 13872 2864
rect 13832 2582 13860 2858
rect 13924 2582 13952 2926
rect 13820 2576 13872 2582
rect 13820 2518 13872 2524
rect 13912 2576 13964 2582
rect 13912 2518 13964 2524
rect 13266 54 13492 82
rect 14370 82 14426 480
rect 14660 82 14688 6666
rect 15016 6316 15068 6322
rect 15016 6258 15068 6264
rect 14924 6180 14976 6186
rect 14924 6122 14976 6128
rect 14936 5370 14964 6122
rect 15028 5914 15056 6258
rect 15200 6112 15252 6118
rect 15200 6054 15252 6060
rect 15016 5908 15068 5914
rect 15016 5850 15068 5856
rect 15212 5846 15240 6054
rect 15200 5840 15252 5846
rect 15200 5782 15252 5788
rect 15212 5370 15240 5782
rect 14924 5364 14976 5370
rect 14924 5306 14976 5312
rect 15200 5364 15252 5370
rect 15200 5306 15252 5312
rect 15108 5092 15160 5098
rect 15108 5034 15160 5040
rect 15120 4826 15148 5034
rect 15212 5030 15240 5306
rect 15200 5024 15252 5030
rect 15200 4966 15252 4972
rect 15108 4820 15160 4826
rect 15108 4762 15160 4768
rect 15108 4276 15160 4282
rect 15108 4218 15160 4224
rect 14740 4072 14792 4078
rect 14740 4014 14792 4020
rect 14752 3670 14780 4014
rect 15120 3738 15148 4218
rect 15108 3732 15160 3738
rect 15108 3674 15160 3680
rect 14740 3664 14792 3670
rect 14740 3606 14792 3612
rect 15120 3058 15148 3674
rect 15108 3052 15160 3058
rect 15108 2994 15160 3000
rect 15200 2304 15252 2310
rect 15200 2246 15252 2252
rect 15212 2009 15240 2246
rect 15198 2000 15254 2009
rect 15198 1935 15254 1944
rect 14370 54 14688 82
rect 15304 82 15332 8774
rect 15396 8022 15424 9386
rect 15622 9276 15918 9296
rect 15678 9274 15702 9276
rect 15758 9274 15782 9276
rect 15838 9274 15862 9276
rect 15700 9222 15702 9274
rect 15764 9222 15776 9274
rect 15838 9222 15840 9274
rect 15678 9220 15702 9222
rect 15758 9220 15782 9222
rect 15838 9220 15862 9222
rect 15622 9200 15918 9220
rect 15622 8188 15918 8208
rect 15678 8186 15702 8188
rect 15758 8186 15782 8188
rect 15838 8186 15862 8188
rect 15700 8134 15702 8186
rect 15764 8134 15776 8186
rect 15838 8134 15840 8186
rect 15678 8132 15702 8134
rect 15758 8132 15782 8134
rect 15838 8132 15862 8134
rect 15474 8120 15530 8129
rect 15622 8112 15918 8132
rect 15474 8055 15530 8064
rect 15384 8016 15436 8022
rect 15384 7958 15436 7964
rect 15396 7546 15424 7958
rect 15488 7546 15516 8055
rect 15384 7540 15436 7546
rect 15384 7482 15436 7488
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 15396 7274 15424 7482
rect 15948 7342 15976 13654
rect 16026 13631 16082 13640
rect 16028 12708 16080 12714
rect 16028 12650 16080 12656
rect 16040 12374 16068 12650
rect 16028 12368 16080 12374
rect 16028 12310 16080 12316
rect 16040 12170 16068 12310
rect 16028 12164 16080 12170
rect 16028 12106 16080 12112
rect 16040 11898 16068 12106
rect 16028 11892 16080 11898
rect 16028 11834 16080 11840
rect 16028 11348 16080 11354
rect 16028 11290 16080 11296
rect 16040 10130 16068 11290
rect 16028 10124 16080 10130
rect 16028 10066 16080 10072
rect 16132 8362 16160 17478
rect 16224 16794 16252 21542
rect 16394 21520 16450 21542
rect 19720 21542 20130 21570
rect 16394 20496 16450 20505
rect 16394 20431 16450 20440
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 16304 16652 16356 16658
rect 16304 16594 16356 16600
rect 16316 16250 16344 16594
rect 16304 16244 16356 16250
rect 16304 16186 16356 16192
rect 16304 16108 16356 16114
rect 16304 16050 16356 16056
rect 16212 15972 16264 15978
rect 16212 15914 16264 15920
rect 16224 8956 16252 15914
rect 16316 11898 16344 16050
rect 16408 15910 16436 20431
rect 19289 19612 19585 19632
rect 19345 19610 19369 19612
rect 19425 19610 19449 19612
rect 19505 19610 19529 19612
rect 19367 19558 19369 19610
rect 19431 19558 19443 19610
rect 19505 19558 19507 19610
rect 19345 19556 19369 19558
rect 19425 19556 19449 19558
rect 19505 19556 19529 19558
rect 19289 19536 19585 19556
rect 19064 18964 19116 18970
rect 19064 18906 19116 18912
rect 18420 18216 18472 18222
rect 18420 18158 18472 18164
rect 16764 18080 16816 18086
rect 16764 18022 16816 18028
rect 16580 16108 16632 16114
rect 16580 16050 16632 16056
rect 16396 15904 16448 15910
rect 16396 15846 16448 15852
rect 16488 15360 16540 15366
rect 16488 15302 16540 15308
rect 16396 13932 16448 13938
rect 16396 13874 16448 13880
rect 16408 13258 16436 13874
rect 16396 13252 16448 13258
rect 16396 13194 16448 13200
rect 16396 12844 16448 12850
rect 16500 12832 16528 15302
rect 16592 13297 16620 16050
rect 16776 14958 16804 18022
rect 17224 17740 17276 17746
rect 17224 17682 17276 17688
rect 17236 17338 17264 17682
rect 17224 17332 17276 17338
rect 17224 17274 17276 17280
rect 18328 17060 18380 17066
rect 18328 17002 18380 17008
rect 17316 16652 17368 16658
rect 17316 16594 17368 16600
rect 17132 16448 17184 16454
rect 17132 16390 17184 16396
rect 17040 16176 17092 16182
rect 17040 16118 17092 16124
rect 16764 14952 16816 14958
rect 16764 14894 16816 14900
rect 16672 14612 16724 14618
rect 16672 14554 16724 14560
rect 16684 13841 16712 14554
rect 16776 14414 16804 14894
rect 16856 14816 16908 14822
rect 16856 14758 16908 14764
rect 16764 14408 16816 14414
rect 16764 14350 16816 14356
rect 16670 13832 16726 13841
rect 16670 13767 16726 13776
rect 16764 13796 16816 13802
rect 16764 13738 16816 13744
rect 16672 13728 16724 13734
rect 16672 13670 16724 13676
rect 16578 13288 16634 13297
rect 16578 13223 16634 13232
rect 16448 12804 16528 12832
rect 16396 12786 16448 12792
rect 16500 12442 16528 12804
rect 16488 12436 16540 12442
rect 16488 12378 16540 12384
rect 16580 12436 16632 12442
rect 16580 12378 16632 12384
rect 16304 11892 16356 11898
rect 16304 11834 16356 11840
rect 16304 11280 16356 11286
rect 16304 11222 16356 11228
rect 16316 10810 16344 11222
rect 16488 11144 16540 11150
rect 16488 11086 16540 11092
rect 16304 10804 16356 10810
rect 16304 10746 16356 10752
rect 16316 10538 16344 10746
rect 16304 10532 16356 10538
rect 16304 10474 16356 10480
rect 16316 10266 16344 10474
rect 16500 10266 16528 11086
rect 16304 10260 16356 10266
rect 16304 10202 16356 10208
rect 16488 10260 16540 10266
rect 16488 10202 16540 10208
rect 16592 10198 16620 12378
rect 16580 10192 16632 10198
rect 16580 10134 16632 10140
rect 16488 9988 16540 9994
rect 16488 9930 16540 9936
rect 16396 9716 16448 9722
rect 16396 9658 16448 9664
rect 16408 9110 16436 9658
rect 16396 9104 16448 9110
rect 16396 9046 16448 9052
rect 16304 8968 16356 8974
rect 16224 8928 16304 8956
rect 16224 8566 16252 8928
rect 16304 8910 16356 8916
rect 16408 8634 16436 9046
rect 16396 8628 16448 8634
rect 16396 8570 16448 8576
rect 16212 8560 16264 8566
rect 16212 8502 16264 8508
rect 16304 8560 16356 8566
rect 16304 8502 16356 8508
rect 16316 8430 16344 8502
rect 16500 8480 16528 9930
rect 16408 8452 16528 8480
rect 16304 8424 16356 8430
rect 16304 8366 16356 8372
rect 16120 8356 16172 8362
rect 16120 8298 16172 8304
rect 16304 8288 16356 8294
rect 16304 8230 16356 8236
rect 16316 7342 16344 8230
rect 16408 7449 16436 8452
rect 16488 8356 16540 8362
rect 16488 8298 16540 8304
rect 16500 8090 16528 8298
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 16580 8084 16632 8090
rect 16580 8026 16632 8032
rect 16394 7440 16450 7449
rect 16592 7410 16620 8026
rect 16394 7375 16450 7384
rect 16580 7404 16632 7410
rect 15936 7336 15988 7342
rect 15936 7278 15988 7284
rect 16304 7336 16356 7342
rect 16304 7278 16356 7284
rect 15384 7268 15436 7274
rect 15384 7210 15436 7216
rect 15396 7002 15424 7210
rect 15622 7100 15918 7120
rect 15678 7098 15702 7100
rect 15758 7098 15782 7100
rect 15838 7098 15862 7100
rect 15700 7046 15702 7098
rect 15764 7046 15776 7098
rect 15838 7046 15840 7098
rect 15678 7044 15702 7046
rect 15758 7044 15782 7046
rect 15838 7044 15862 7046
rect 15622 7024 15918 7044
rect 15384 6996 15436 7002
rect 15384 6938 15436 6944
rect 15384 6860 15436 6866
rect 15384 6802 15436 6808
rect 15396 6458 15424 6802
rect 15936 6656 15988 6662
rect 15936 6598 15988 6604
rect 16304 6656 16356 6662
rect 16304 6598 16356 6604
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 15948 6186 15976 6598
rect 16028 6384 16080 6390
rect 16028 6326 16080 6332
rect 15936 6180 15988 6186
rect 15936 6122 15988 6128
rect 15622 6012 15918 6032
rect 15678 6010 15702 6012
rect 15758 6010 15782 6012
rect 15838 6010 15862 6012
rect 15700 5958 15702 6010
rect 15764 5958 15776 6010
rect 15838 5958 15840 6010
rect 15678 5956 15702 5958
rect 15758 5956 15782 5958
rect 15838 5956 15862 5958
rect 15622 5936 15918 5956
rect 15844 5568 15896 5574
rect 15844 5510 15896 5516
rect 15856 5098 15884 5510
rect 15948 5370 15976 6122
rect 16040 5710 16068 6326
rect 16028 5704 16080 5710
rect 16028 5646 16080 5652
rect 15936 5364 15988 5370
rect 15936 5306 15988 5312
rect 15844 5092 15896 5098
rect 15844 5034 15896 5040
rect 15622 4924 15918 4944
rect 15678 4922 15702 4924
rect 15758 4922 15782 4924
rect 15838 4922 15862 4924
rect 15700 4870 15702 4922
rect 15764 4870 15776 4922
rect 15838 4870 15840 4922
rect 15678 4868 15702 4870
rect 15758 4868 15782 4870
rect 15838 4868 15862 4870
rect 15622 4848 15918 4868
rect 15476 4752 15528 4758
rect 15476 4694 15528 4700
rect 15488 4010 15516 4694
rect 15936 4548 15988 4554
rect 15936 4490 15988 4496
rect 15476 4004 15528 4010
rect 15476 3946 15528 3952
rect 15384 3936 15436 3942
rect 15384 3878 15436 3884
rect 15396 3534 15424 3878
rect 15622 3836 15918 3856
rect 15678 3834 15702 3836
rect 15758 3834 15782 3836
rect 15838 3834 15862 3836
rect 15700 3782 15702 3834
rect 15764 3782 15776 3834
rect 15838 3782 15840 3834
rect 15678 3780 15702 3782
rect 15758 3780 15782 3782
rect 15838 3780 15862 3782
rect 15622 3760 15918 3780
rect 15476 3664 15528 3670
rect 15476 3606 15528 3612
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 15488 3194 15516 3606
rect 15948 3466 15976 4490
rect 16040 3942 16068 5646
rect 16316 5642 16344 6598
rect 16408 5692 16436 7375
rect 16580 7346 16632 7352
rect 16684 6798 16712 13670
rect 16776 13190 16804 13738
rect 16868 13433 16896 14758
rect 16948 14000 17000 14006
rect 16948 13942 17000 13948
rect 16960 13530 16988 13942
rect 17052 13734 17080 16118
rect 17040 13728 17092 13734
rect 17040 13670 17092 13676
rect 16948 13524 17000 13530
rect 16948 13466 17000 13472
rect 16854 13424 16910 13433
rect 16854 13359 16910 13368
rect 17040 13388 17092 13394
rect 17040 13330 17092 13336
rect 16764 13184 16816 13190
rect 16764 13126 16816 13132
rect 16776 12850 16804 13126
rect 16764 12844 16816 12850
rect 16764 12786 16816 12792
rect 17052 12646 17080 13330
rect 17040 12640 17092 12646
rect 17040 12582 17092 12588
rect 17040 12300 17092 12306
rect 17040 12242 17092 12248
rect 17052 11626 17080 12242
rect 17040 11620 17092 11626
rect 17040 11562 17092 11568
rect 16856 11552 16908 11558
rect 16856 11494 16908 11500
rect 16764 11076 16816 11082
rect 16764 11018 16816 11024
rect 16776 8974 16804 11018
rect 16868 10266 16896 11494
rect 16856 10260 16908 10266
rect 16856 10202 16908 10208
rect 16856 9512 16908 9518
rect 16856 9454 16908 9460
rect 16764 8968 16816 8974
rect 16764 8910 16816 8916
rect 16868 8820 16896 9454
rect 16948 9444 17000 9450
rect 16948 9386 17000 9392
rect 16776 8792 16896 8820
rect 16672 6792 16724 6798
rect 16672 6734 16724 6740
rect 16684 5846 16712 6734
rect 16776 6338 16804 8792
rect 16856 7336 16908 7342
rect 16856 7278 16908 7284
rect 16868 6934 16896 7278
rect 16856 6928 16908 6934
rect 16856 6870 16908 6876
rect 16868 6458 16896 6870
rect 16856 6452 16908 6458
rect 16856 6394 16908 6400
rect 16776 6310 16896 6338
rect 16672 5840 16724 5846
rect 16672 5782 16724 5788
rect 16408 5664 16712 5692
rect 16304 5636 16356 5642
rect 16304 5578 16356 5584
rect 16488 5160 16540 5166
rect 16408 5120 16488 5148
rect 16304 5024 16356 5030
rect 16304 4966 16356 4972
rect 16316 4826 16344 4966
rect 16304 4820 16356 4826
rect 16304 4762 16356 4768
rect 16304 4684 16356 4690
rect 16304 4626 16356 4632
rect 16316 4146 16344 4626
rect 16408 4622 16436 5120
rect 16488 5102 16540 5108
rect 16396 4616 16448 4622
rect 16396 4558 16448 4564
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16028 3936 16080 3942
rect 16026 3904 16028 3913
rect 16080 3904 16082 3913
rect 16026 3839 16082 3848
rect 16040 3813 16068 3839
rect 15936 3460 15988 3466
rect 15936 3402 15988 3408
rect 15476 3188 15528 3194
rect 15476 3130 15528 3136
rect 15844 3188 15896 3194
rect 15844 3130 15896 3136
rect 15856 2922 15884 3130
rect 15844 2916 15896 2922
rect 15844 2858 15896 2864
rect 15622 2748 15918 2768
rect 15678 2746 15702 2748
rect 15758 2746 15782 2748
rect 15838 2746 15862 2748
rect 15700 2694 15702 2746
rect 15764 2694 15776 2746
rect 15838 2694 15840 2746
rect 15678 2692 15702 2694
rect 15758 2692 15782 2694
rect 15838 2692 15862 2694
rect 15622 2672 15918 2692
rect 15568 2576 15620 2582
rect 15568 2518 15620 2524
rect 15580 2428 15608 2518
rect 15948 2446 15976 3402
rect 16408 3058 16436 4558
rect 16488 4480 16540 4486
rect 16488 4422 16540 4428
rect 16500 4146 16528 4422
rect 16488 4140 16540 4146
rect 16488 4082 16540 4088
rect 16580 4004 16632 4010
rect 16580 3946 16632 3952
rect 16592 3738 16620 3946
rect 16580 3732 16632 3738
rect 16580 3674 16632 3680
rect 16486 3496 16542 3505
rect 16486 3431 16542 3440
rect 16500 3398 16528 3431
rect 16488 3392 16540 3398
rect 16488 3334 16540 3340
rect 16592 3194 16620 3674
rect 16684 3505 16712 5664
rect 16764 4140 16816 4146
rect 16764 4082 16816 4088
rect 16670 3496 16726 3505
rect 16670 3431 16726 3440
rect 16580 3188 16632 3194
rect 16580 3130 16632 3136
rect 16776 3058 16804 4082
rect 16396 3052 16448 3058
rect 16396 2994 16448 3000
rect 16764 3052 16816 3058
rect 16764 2994 16816 3000
rect 15660 2440 15712 2446
rect 15580 2400 15660 2428
rect 15660 2382 15712 2388
rect 15936 2440 15988 2446
rect 15936 2382 15988 2388
rect 15566 82 15622 480
rect 15304 54 15622 82
rect 13266 0 13322 54
rect 14370 0 14426 54
rect 15566 0 15622 54
rect 16762 82 16818 480
rect 16868 82 16896 6310
rect 16960 5710 16988 9386
rect 17052 6882 17080 11562
rect 17144 8022 17172 16390
rect 17328 15910 17356 16594
rect 18236 16584 18288 16590
rect 18236 16526 18288 16532
rect 17408 16244 17460 16250
rect 17408 16186 17460 16192
rect 17960 16244 18012 16250
rect 17960 16186 18012 16192
rect 17316 15904 17368 15910
rect 17316 15846 17368 15852
rect 17316 15564 17368 15570
rect 17316 15506 17368 15512
rect 17328 15162 17356 15506
rect 17316 15156 17368 15162
rect 17316 15098 17368 15104
rect 17328 15026 17356 15098
rect 17316 15020 17368 15026
rect 17316 14962 17368 14968
rect 17420 14482 17448 16186
rect 17972 16153 18000 16186
rect 17958 16144 18014 16153
rect 17958 16079 18014 16088
rect 17972 16046 18000 16079
rect 17960 16040 18012 16046
rect 17960 15982 18012 15988
rect 18052 15700 18104 15706
rect 18052 15642 18104 15648
rect 17776 15564 17828 15570
rect 17776 15506 17828 15512
rect 17788 15162 17816 15506
rect 17776 15156 17828 15162
rect 17776 15098 17828 15104
rect 17788 15065 17816 15098
rect 17774 15056 17830 15065
rect 17774 14991 17830 15000
rect 17590 14920 17646 14929
rect 17590 14855 17646 14864
rect 17604 14822 17632 14855
rect 17592 14816 17644 14822
rect 17592 14758 17644 14764
rect 17684 14816 17736 14822
rect 17684 14758 17736 14764
rect 17224 14476 17276 14482
rect 17224 14418 17276 14424
rect 17408 14476 17460 14482
rect 17408 14418 17460 14424
rect 17236 13734 17264 14418
rect 17420 14006 17448 14418
rect 17408 14000 17460 14006
rect 17408 13942 17460 13948
rect 17224 13728 17276 13734
rect 17224 13670 17276 13676
rect 17236 13462 17264 13670
rect 17224 13456 17276 13462
rect 17224 13398 17276 13404
rect 17236 12628 17264 13398
rect 17420 12986 17448 13942
rect 17500 13728 17552 13734
rect 17500 13670 17552 13676
rect 17408 12980 17460 12986
rect 17408 12922 17460 12928
rect 17512 12918 17540 13670
rect 17500 12912 17552 12918
rect 17500 12854 17552 12860
rect 17316 12640 17368 12646
rect 17236 12600 17316 12628
rect 17316 12582 17368 12588
rect 17224 11552 17276 11558
rect 17224 11494 17276 11500
rect 17236 11286 17264 11494
rect 17224 11280 17276 11286
rect 17224 11222 17276 11228
rect 17328 10606 17356 12582
rect 17500 12300 17552 12306
rect 17500 12242 17552 12248
rect 17408 11756 17460 11762
rect 17408 11698 17460 11704
rect 17316 10600 17368 10606
rect 17316 10542 17368 10548
rect 17316 10464 17368 10470
rect 17316 10406 17368 10412
rect 17224 10192 17276 10198
rect 17224 10134 17276 10140
rect 17236 9722 17264 10134
rect 17328 10062 17356 10406
rect 17316 10056 17368 10062
rect 17316 9998 17368 10004
rect 17224 9716 17276 9722
rect 17224 9658 17276 9664
rect 17420 9518 17448 11698
rect 17512 11694 17540 12242
rect 17500 11688 17552 11694
rect 17500 11630 17552 11636
rect 17592 11620 17644 11626
rect 17592 11562 17644 11568
rect 17500 11552 17552 11558
rect 17500 11494 17552 11500
rect 17512 10713 17540 11494
rect 17498 10704 17554 10713
rect 17498 10639 17554 10648
rect 17408 9512 17460 9518
rect 17408 9454 17460 9460
rect 17316 9036 17368 9042
rect 17316 8978 17368 8984
rect 17328 8294 17356 8978
rect 17408 8492 17460 8498
rect 17408 8434 17460 8440
rect 17316 8288 17368 8294
rect 17316 8230 17368 8236
rect 17132 8016 17184 8022
rect 17132 7958 17184 7964
rect 17224 8016 17276 8022
rect 17224 7958 17276 7964
rect 17144 7002 17172 7958
rect 17236 7818 17264 7958
rect 17224 7812 17276 7818
rect 17224 7754 17276 7760
rect 17236 7478 17264 7754
rect 17224 7472 17276 7478
rect 17224 7414 17276 7420
rect 17328 7313 17356 8230
rect 17420 7886 17448 8434
rect 17512 7886 17540 10639
rect 17604 9081 17632 11562
rect 17696 11082 17724 14758
rect 17776 14408 17828 14414
rect 17776 14350 17828 14356
rect 17684 11076 17736 11082
rect 17684 11018 17736 11024
rect 17788 9674 17816 14350
rect 18064 12782 18092 15642
rect 18248 13394 18276 16526
rect 18340 13938 18368 17002
rect 18432 14958 18460 18158
rect 18788 17332 18840 17338
rect 18788 17274 18840 17280
rect 18512 16652 18564 16658
rect 18512 16594 18564 16600
rect 18524 15910 18552 16594
rect 18512 15904 18564 15910
rect 18512 15846 18564 15852
rect 18420 14952 18472 14958
rect 18420 14894 18472 14900
rect 18418 14512 18474 14521
rect 18418 14447 18420 14456
rect 18472 14447 18474 14456
rect 18420 14418 18472 14424
rect 18432 14006 18460 14418
rect 18420 14000 18472 14006
rect 18420 13942 18472 13948
rect 18328 13932 18380 13938
rect 18328 13874 18380 13880
rect 18236 13388 18288 13394
rect 18236 13330 18288 13336
rect 18248 12918 18276 13330
rect 18236 12912 18288 12918
rect 18236 12854 18288 12860
rect 18248 12789 18276 12854
rect 18052 12776 18104 12782
rect 18052 12718 18104 12724
rect 18064 12442 18092 12718
rect 18144 12640 18196 12646
rect 18144 12582 18196 12588
rect 18052 12436 18104 12442
rect 17880 12396 18052 12424
rect 17880 11218 17908 12396
rect 18052 12378 18104 12384
rect 17960 11688 18012 11694
rect 17960 11630 18012 11636
rect 17972 11218 18000 11630
rect 17868 11212 17920 11218
rect 17868 11154 17920 11160
rect 17960 11212 18012 11218
rect 17960 11154 18012 11160
rect 17880 10690 17908 11154
rect 18156 11014 18184 12582
rect 18236 11212 18288 11218
rect 18236 11154 18288 11160
rect 18144 11008 18196 11014
rect 18144 10950 18196 10956
rect 18248 10742 18276 11154
rect 18236 10736 18288 10742
rect 17880 10662 18000 10690
rect 18236 10678 18288 10684
rect 17868 10464 17920 10470
rect 17868 10406 17920 10412
rect 17696 9646 17816 9674
rect 17590 9072 17646 9081
rect 17590 9007 17646 9016
rect 17604 8974 17632 9007
rect 17592 8968 17644 8974
rect 17592 8910 17644 8916
rect 17408 7880 17460 7886
rect 17408 7822 17460 7828
rect 17500 7880 17552 7886
rect 17500 7822 17552 7828
rect 17500 7404 17552 7410
rect 17500 7346 17552 7352
rect 17314 7304 17370 7313
rect 17314 7239 17370 7248
rect 17132 6996 17184 7002
rect 17132 6938 17184 6944
rect 17052 6854 17172 6882
rect 17040 5840 17092 5846
rect 17040 5782 17092 5788
rect 16948 5704 17000 5710
rect 16948 5646 17000 5652
rect 16960 5030 16988 5646
rect 17052 5302 17080 5782
rect 17040 5296 17092 5302
rect 17040 5238 17092 5244
rect 16948 5024 17000 5030
rect 16948 4966 17000 4972
rect 16948 4820 17000 4826
rect 16948 4762 17000 4768
rect 16960 3670 16988 4762
rect 17144 4154 17172 6854
rect 17316 6180 17368 6186
rect 17316 6122 17368 6128
rect 17224 5704 17276 5710
rect 17224 5646 17276 5652
rect 17236 5166 17264 5646
rect 17224 5160 17276 5166
rect 17224 5102 17276 5108
rect 17328 4690 17356 6122
rect 17512 5574 17540 7346
rect 17696 6798 17724 9646
rect 17880 9586 17908 10406
rect 17972 10266 18000 10662
rect 18236 10600 18288 10606
rect 18236 10542 18288 10548
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 17868 9580 17920 9586
rect 17868 9522 17920 9528
rect 17776 9512 17828 9518
rect 17774 9480 17776 9489
rect 17828 9480 17830 9489
rect 17774 9415 17830 9424
rect 17788 9382 17816 9415
rect 17776 9376 17828 9382
rect 17776 9318 17828 9324
rect 17868 9376 17920 9382
rect 17868 9318 17920 9324
rect 17684 6792 17736 6798
rect 17880 6769 17908 9318
rect 17972 7426 18000 10202
rect 18248 9926 18276 10542
rect 18340 9994 18368 13874
rect 18432 13433 18460 13942
rect 18418 13424 18474 13433
rect 18418 13359 18474 13368
rect 18420 12708 18472 12714
rect 18420 12650 18472 12656
rect 18328 9988 18380 9994
rect 18328 9930 18380 9936
rect 18236 9920 18288 9926
rect 18236 9862 18288 9868
rect 18142 9616 18198 9625
rect 18142 9551 18198 9560
rect 18052 9512 18104 9518
rect 18052 9454 18104 9460
rect 18064 8838 18092 9454
rect 18052 8832 18104 8838
rect 18052 8774 18104 8780
rect 18064 8634 18092 8774
rect 18052 8628 18104 8634
rect 18052 8570 18104 8576
rect 18064 7546 18092 8570
rect 18156 7954 18184 9551
rect 18432 8906 18460 12650
rect 18524 12594 18552 15846
rect 18604 15564 18656 15570
rect 18604 15506 18656 15512
rect 18616 14822 18644 15506
rect 18696 15020 18748 15026
rect 18696 14962 18748 14968
rect 18604 14816 18656 14822
rect 18604 14758 18656 14764
rect 18616 14074 18644 14758
rect 18604 14068 18656 14074
rect 18604 14010 18656 14016
rect 18604 13728 18656 13734
rect 18604 13670 18656 13676
rect 18616 13258 18644 13670
rect 18604 13252 18656 13258
rect 18604 13194 18656 13200
rect 18524 12566 18644 12594
rect 18512 12436 18564 12442
rect 18512 12378 18564 12384
rect 18524 11121 18552 12378
rect 18616 11286 18644 12566
rect 18708 12424 18736 14962
rect 18800 13530 18828 17274
rect 18972 15972 19024 15978
rect 18972 15914 19024 15920
rect 18788 13524 18840 13530
rect 18788 13466 18840 13472
rect 18880 13388 18932 13394
rect 18880 13330 18932 13336
rect 18892 12782 18920 13330
rect 18984 12850 19012 15914
rect 19076 14482 19104 18906
rect 19289 18524 19585 18544
rect 19345 18522 19369 18524
rect 19425 18522 19449 18524
rect 19505 18522 19529 18524
rect 19367 18470 19369 18522
rect 19431 18470 19443 18522
rect 19505 18470 19507 18522
rect 19345 18468 19369 18470
rect 19425 18468 19449 18470
rect 19505 18468 19529 18470
rect 19289 18448 19585 18468
rect 19720 18426 19748 21542
rect 20074 21520 20130 21542
rect 19798 18456 19854 18465
rect 19708 18420 19760 18426
rect 19798 18391 19854 18400
rect 19708 18362 19760 18368
rect 19289 17436 19585 17456
rect 19345 17434 19369 17436
rect 19425 17434 19449 17436
rect 19505 17434 19529 17436
rect 19367 17382 19369 17434
rect 19431 17382 19443 17434
rect 19505 17382 19507 17434
rect 19345 17380 19369 17382
rect 19425 17380 19449 17382
rect 19505 17380 19529 17382
rect 19289 17360 19585 17380
rect 19614 16552 19670 16561
rect 19614 16487 19670 16496
rect 19289 16348 19585 16368
rect 19345 16346 19369 16348
rect 19425 16346 19449 16348
rect 19505 16346 19529 16348
rect 19367 16294 19369 16346
rect 19431 16294 19443 16346
rect 19505 16294 19507 16346
rect 19345 16292 19369 16294
rect 19425 16292 19449 16294
rect 19505 16292 19529 16294
rect 19289 16272 19585 16292
rect 19156 16040 19208 16046
rect 19156 15982 19208 15988
rect 19064 14476 19116 14482
rect 19064 14418 19116 14424
rect 18972 12844 19024 12850
rect 18972 12786 19024 12792
rect 18880 12776 18932 12782
rect 18880 12718 18932 12724
rect 18708 12396 18828 12424
rect 18696 12300 18748 12306
rect 18696 12242 18748 12248
rect 18708 11354 18736 12242
rect 18696 11348 18748 11354
rect 18696 11290 18748 11296
rect 18604 11280 18656 11286
rect 18604 11222 18656 11228
rect 18510 11112 18566 11121
rect 18510 11047 18566 11056
rect 18602 10840 18658 10849
rect 18602 10775 18658 10784
rect 18512 10736 18564 10742
rect 18512 10678 18564 10684
rect 18524 10606 18552 10678
rect 18512 10600 18564 10606
rect 18512 10542 18564 10548
rect 18524 10198 18552 10542
rect 18512 10192 18564 10198
rect 18512 10134 18564 10140
rect 18616 10130 18644 10775
rect 18696 10260 18748 10266
rect 18696 10202 18748 10208
rect 18604 10124 18656 10130
rect 18604 10066 18656 10072
rect 18616 9586 18644 10066
rect 18604 9580 18656 9586
rect 18604 9522 18656 9528
rect 18512 9512 18564 9518
rect 18512 9454 18564 9460
rect 18420 8900 18472 8906
rect 18420 8842 18472 8848
rect 18236 8832 18288 8838
rect 18236 8774 18288 8780
rect 18328 8832 18380 8838
rect 18328 8774 18380 8780
rect 18248 8537 18276 8774
rect 18234 8528 18290 8537
rect 18234 8463 18290 8472
rect 18340 8362 18368 8774
rect 18432 8498 18460 8842
rect 18420 8492 18472 8498
rect 18420 8434 18472 8440
rect 18328 8356 18380 8362
rect 18328 8298 18380 8304
rect 18420 8356 18472 8362
rect 18420 8298 18472 8304
rect 18340 8022 18368 8298
rect 18328 8016 18380 8022
rect 18328 7958 18380 7964
rect 18144 7948 18196 7954
rect 18196 7908 18276 7936
rect 18144 7890 18196 7896
rect 18052 7540 18104 7546
rect 18052 7482 18104 7488
rect 17972 7398 18092 7426
rect 17684 6734 17736 6740
rect 17866 6760 17922 6769
rect 17866 6695 17922 6704
rect 17592 6384 17644 6390
rect 17592 6326 17644 6332
rect 17500 5568 17552 5574
rect 17500 5510 17552 5516
rect 17316 4684 17368 4690
rect 17316 4626 17368 4632
rect 17144 4126 17264 4154
rect 17132 4004 17184 4010
rect 17132 3946 17184 3952
rect 17144 3913 17172 3946
rect 17130 3904 17186 3913
rect 17130 3839 17186 3848
rect 16948 3664 17000 3670
rect 16948 3606 17000 3612
rect 17038 3088 17094 3097
rect 17038 3023 17094 3032
rect 17052 2514 17080 3023
rect 17144 2650 17172 3839
rect 17236 3602 17264 4126
rect 17328 3942 17356 4626
rect 17316 3936 17368 3942
rect 17316 3878 17368 3884
rect 17328 3602 17356 3878
rect 17224 3596 17276 3602
rect 17224 3538 17276 3544
rect 17316 3596 17368 3602
rect 17316 3538 17368 3544
rect 17236 3194 17264 3538
rect 17224 3188 17276 3194
rect 17224 3130 17276 3136
rect 17328 3126 17356 3538
rect 17316 3120 17368 3126
rect 17316 3062 17368 3068
rect 17132 2644 17184 2650
rect 17132 2586 17184 2592
rect 17040 2508 17092 2514
rect 17040 2450 17092 2456
rect 16762 54 16896 82
rect 17604 82 17632 6326
rect 17868 6112 17920 6118
rect 17868 6054 17920 6060
rect 17684 5568 17736 5574
rect 17684 5510 17736 5516
rect 17696 3942 17724 5510
rect 17880 5234 17908 6054
rect 18064 5273 18092 7398
rect 18144 6996 18196 7002
rect 18144 6938 18196 6944
rect 18156 5817 18184 6938
rect 18248 6866 18276 7908
rect 18328 7880 18380 7886
rect 18328 7822 18380 7828
rect 18340 7342 18368 7822
rect 18328 7336 18380 7342
rect 18328 7278 18380 7284
rect 18236 6860 18288 6866
rect 18236 6802 18288 6808
rect 18248 6458 18276 6802
rect 18236 6452 18288 6458
rect 18236 6394 18288 6400
rect 18248 6254 18276 6394
rect 18236 6248 18288 6254
rect 18236 6190 18288 6196
rect 18142 5808 18198 5817
rect 18142 5743 18198 5752
rect 18050 5264 18106 5273
rect 17868 5228 17920 5234
rect 18050 5199 18106 5208
rect 17868 5170 17920 5176
rect 17776 5160 17828 5166
rect 17774 5128 17776 5137
rect 17828 5128 17830 5137
rect 17774 5063 17830 5072
rect 18052 5092 18104 5098
rect 17788 5030 17816 5063
rect 18052 5034 18104 5040
rect 17776 5024 17828 5030
rect 17776 4966 17828 4972
rect 18064 4049 18092 5034
rect 18144 4616 18196 4622
rect 18144 4558 18196 4564
rect 18156 4078 18184 4558
rect 18432 4282 18460 8298
rect 18524 7206 18552 9454
rect 18708 9178 18736 10202
rect 18800 10033 18828 12396
rect 18892 12306 18920 12718
rect 18880 12300 18932 12306
rect 18880 12242 18932 12248
rect 18892 11694 18920 12242
rect 18880 11688 18932 11694
rect 18880 11630 18932 11636
rect 19064 11688 19116 11694
rect 19064 11630 19116 11636
rect 18972 10192 19024 10198
rect 18972 10134 19024 10140
rect 18786 10024 18842 10033
rect 18786 9959 18842 9968
rect 18696 9172 18748 9178
rect 18696 9114 18748 9120
rect 18800 9042 18828 9959
rect 18984 9722 19012 10134
rect 18972 9716 19024 9722
rect 18972 9658 19024 9664
rect 18880 9580 18932 9586
rect 18880 9522 18932 9528
rect 18696 9036 18748 9042
rect 18696 8978 18748 8984
rect 18788 9036 18840 9042
rect 18788 8978 18840 8984
rect 18604 8492 18656 8498
rect 18604 8434 18656 8440
rect 18512 7200 18564 7206
rect 18512 7142 18564 7148
rect 18616 6934 18644 8434
rect 18708 7750 18736 8978
rect 18800 8634 18828 8978
rect 18788 8628 18840 8634
rect 18788 8570 18840 8576
rect 18696 7744 18748 7750
rect 18696 7686 18748 7692
rect 18604 6928 18656 6934
rect 18604 6870 18656 6876
rect 18512 6860 18564 6866
rect 18512 6802 18564 6808
rect 18524 5710 18552 6802
rect 18604 5772 18656 5778
rect 18604 5714 18656 5720
rect 18512 5704 18564 5710
rect 18512 5646 18564 5652
rect 18512 4684 18564 4690
rect 18512 4626 18564 4632
rect 18524 4593 18552 4626
rect 18510 4584 18566 4593
rect 18510 4519 18566 4528
rect 18524 4282 18552 4519
rect 18616 4486 18644 5714
rect 18708 4826 18736 7686
rect 18788 7268 18840 7274
rect 18788 7210 18840 7216
rect 18696 4820 18748 4826
rect 18696 4762 18748 4768
rect 18604 4480 18656 4486
rect 18604 4422 18656 4428
rect 18420 4276 18472 4282
rect 18420 4218 18472 4224
rect 18512 4276 18564 4282
rect 18512 4218 18564 4224
rect 18144 4072 18196 4078
rect 18050 4040 18106 4049
rect 18144 4014 18196 4020
rect 18604 4072 18656 4078
rect 18604 4014 18656 4020
rect 18050 3975 18106 3984
rect 17684 3936 17736 3942
rect 17684 3878 17736 3884
rect 18144 3936 18196 3942
rect 18144 3878 18196 3884
rect 17696 3398 17724 3878
rect 18156 3641 18184 3878
rect 18512 3732 18564 3738
rect 18512 3674 18564 3680
rect 18142 3632 18198 3641
rect 17776 3596 17828 3602
rect 18142 3567 18198 3576
rect 17776 3538 17828 3544
rect 17684 3392 17736 3398
rect 17684 3334 17736 3340
rect 17788 2990 17816 3538
rect 18144 3392 18196 3398
rect 18144 3334 18196 3340
rect 18156 2990 18184 3334
rect 17776 2984 17828 2990
rect 17774 2952 17776 2961
rect 18144 2984 18196 2990
rect 17828 2952 17830 2961
rect 18144 2926 18196 2932
rect 17774 2887 17830 2896
rect 17788 2854 17816 2887
rect 17776 2848 17828 2854
rect 17776 2790 17828 2796
rect 18144 2848 18196 2854
rect 18144 2790 18196 2796
rect 17788 2650 17816 2790
rect 17776 2644 17828 2650
rect 17776 2586 17828 2592
rect 18156 2417 18184 2790
rect 18420 2644 18472 2650
rect 18420 2586 18472 2592
rect 18142 2408 18198 2417
rect 18142 2343 18198 2352
rect 18432 1601 18460 2586
rect 18524 1737 18552 3674
rect 18616 3369 18644 4014
rect 18800 3602 18828 7210
rect 18892 4758 18920 9522
rect 19076 7954 19104 11630
rect 19168 9518 19196 15982
rect 19628 15706 19656 16487
rect 19616 15700 19668 15706
rect 19616 15642 19668 15648
rect 19289 15260 19585 15280
rect 19345 15258 19369 15260
rect 19425 15258 19449 15260
rect 19505 15258 19529 15260
rect 19367 15206 19369 15258
rect 19431 15206 19443 15258
rect 19505 15206 19507 15258
rect 19345 15204 19369 15206
rect 19425 15204 19449 15206
rect 19505 15204 19529 15206
rect 19289 15184 19585 15204
rect 19289 14172 19585 14192
rect 19345 14170 19369 14172
rect 19425 14170 19449 14172
rect 19505 14170 19529 14172
rect 19367 14118 19369 14170
rect 19431 14118 19443 14170
rect 19505 14118 19507 14170
rect 19345 14116 19369 14118
rect 19425 14116 19449 14118
rect 19505 14116 19529 14118
rect 19289 14096 19585 14116
rect 19812 13814 19840 18391
rect 20166 15056 20222 15065
rect 20166 14991 20222 15000
rect 19892 14476 19944 14482
rect 19892 14418 19944 14424
rect 19904 14074 19932 14418
rect 19892 14068 19944 14074
rect 19892 14010 19944 14016
rect 19720 13786 19840 13814
rect 19289 13084 19585 13104
rect 19345 13082 19369 13084
rect 19425 13082 19449 13084
rect 19505 13082 19529 13084
rect 19367 13030 19369 13082
rect 19431 13030 19443 13082
rect 19505 13030 19507 13082
rect 19345 13028 19369 13030
rect 19425 13028 19449 13030
rect 19505 13028 19529 13030
rect 19289 13008 19585 13028
rect 19289 11996 19585 12016
rect 19345 11994 19369 11996
rect 19425 11994 19449 11996
rect 19505 11994 19529 11996
rect 19367 11942 19369 11994
rect 19431 11942 19443 11994
rect 19505 11942 19507 11994
rect 19345 11940 19369 11942
rect 19425 11940 19449 11942
rect 19505 11940 19529 11942
rect 19289 11920 19585 11940
rect 19720 11354 19748 13786
rect 20180 13530 20208 14991
rect 20168 13524 20220 13530
rect 20168 13466 20220 13472
rect 20076 12640 20128 12646
rect 20076 12582 20128 12588
rect 20088 11694 20116 12582
rect 20076 11688 20128 11694
rect 20076 11630 20128 11636
rect 19708 11348 19760 11354
rect 19708 11290 19760 11296
rect 19616 11212 19668 11218
rect 19616 11154 19668 11160
rect 19289 10908 19585 10928
rect 19345 10906 19369 10908
rect 19425 10906 19449 10908
rect 19505 10906 19529 10908
rect 19367 10854 19369 10906
rect 19431 10854 19443 10906
rect 19505 10854 19507 10906
rect 19345 10852 19369 10854
rect 19425 10852 19449 10854
rect 19505 10852 19529 10854
rect 19289 10832 19585 10852
rect 19628 10470 19656 11154
rect 20180 10810 20208 13466
rect 21640 11892 21692 11898
rect 21640 11834 21692 11840
rect 20168 10804 20220 10810
rect 20168 10746 20220 10752
rect 20180 10606 20208 10746
rect 20168 10600 20220 10606
rect 20168 10542 20220 10548
rect 19616 10464 19668 10470
rect 19616 10406 19668 10412
rect 19289 9820 19585 9840
rect 19345 9818 19369 9820
rect 19425 9818 19449 9820
rect 19505 9818 19529 9820
rect 19367 9766 19369 9818
rect 19431 9766 19443 9818
rect 19505 9766 19507 9818
rect 19345 9764 19369 9766
rect 19425 9764 19449 9766
rect 19505 9764 19529 9766
rect 19289 9744 19585 9764
rect 19156 9512 19208 9518
rect 19156 9454 19208 9460
rect 19156 8832 19208 8838
rect 19156 8774 19208 8780
rect 19064 7948 19116 7954
rect 19064 7890 19116 7896
rect 19076 7546 19104 7890
rect 19064 7540 19116 7546
rect 19064 7482 19116 7488
rect 19064 7200 19116 7206
rect 19064 7142 19116 7148
rect 19076 6458 19104 7142
rect 19064 6452 19116 6458
rect 19064 6394 19116 6400
rect 19064 5704 19116 5710
rect 19064 5646 19116 5652
rect 19076 5370 19104 5646
rect 19064 5364 19116 5370
rect 19064 5306 19116 5312
rect 18880 4752 18932 4758
rect 18880 4694 18932 4700
rect 18788 3596 18840 3602
rect 18788 3538 18840 3544
rect 18972 3596 19024 3602
rect 18972 3538 19024 3544
rect 18602 3360 18658 3369
rect 18602 3295 18658 3304
rect 18984 3194 19012 3538
rect 18972 3188 19024 3194
rect 18972 3130 19024 3136
rect 18786 2680 18842 2689
rect 18786 2615 18842 2624
rect 18800 2582 18828 2615
rect 18788 2576 18840 2582
rect 18788 2518 18840 2524
rect 18510 1728 18566 1737
rect 18510 1663 18566 1672
rect 18418 1592 18474 1601
rect 18418 1527 18474 1536
rect 17866 82 17922 480
rect 17604 54 17922 82
rect 16762 0 16818 54
rect 17866 0 17922 54
rect 19062 82 19118 480
rect 19168 82 19196 8774
rect 19289 8732 19585 8752
rect 19345 8730 19369 8732
rect 19425 8730 19449 8732
rect 19505 8730 19529 8732
rect 19367 8678 19369 8730
rect 19431 8678 19443 8730
rect 19505 8678 19507 8730
rect 19345 8676 19369 8678
rect 19425 8676 19449 8678
rect 19505 8676 19529 8678
rect 19289 8656 19585 8676
rect 19289 7644 19585 7664
rect 19345 7642 19369 7644
rect 19425 7642 19449 7644
rect 19505 7642 19529 7644
rect 19367 7590 19369 7642
rect 19431 7590 19443 7642
rect 19505 7590 19507 7642
rect 19345 7588 19369 7590
rect 19425 7588 19449 7590
rect 19505 7588 19529 7590
rect 19289 7568 19585 7588
rect 19628 7342 19656 10406
rect 19708 9920 19760 9926
rect 19708 9862 19760 9868
rect 19720 7857 19748 9862
rect 20180 9674 20208 10542
rect 20088 9646 20208 9674
rect 21548 9648 21600 9654
rect 20088 8945 20116 9646
rect 21548 9590 21600 9596
rect 21560 8945 21588 9590
rect 20074 8936 20130 8945
rect 20074 8871 20130 8880
rect 21546 8936 21602 8945
rect 21546 8871 21602 8880
rect 19984 8628 20036 8634
rect 19984 8570 20036 8576
rect 19706 7848 19762 7857
rect 19706 7783 19762 7792
rect 19616 7336 19668 7342
rect 19616 7278 19668 7284
rect 19289 6556 19585 6576
rect 19345 6554 19369 6556
rect 19425 6554 19449 6556
rect 19505 6554 19529 6556
rect 19367 6502 19369 6554
rect 19431 6502 19443 6554
rect 19505 6502 19507 6554
rect 19345 6500 19369 6502
rect 19425 6500 19449 6502
rect 19505 6500 19529 6502
rect 19289 6480 19585 6500
rect 19289 5468 19585 5488
rect 19345 5466 19369 5468
rect 19425 5466 19449 5468
rect 19505 5466 19529 5468
rect 19367 5414 19369 5466
rect 19431 5414 19443 5466
rect 19505 5414 19507 5466
rect 19345 5412 19369 5414
rect 19425 5412 19449 5414
rect 19505 5412 19529 5414
rect 19289 5392 19585 5412
rect 19720 5030 19748 7783
rect 19800 6996 19852 7002
rect 19800 6938 19852 6944
rect 19708 5024 19760 5030
rect 19708 4966 19760 4972
rect 19720 4486 19748 4966
rect 19708 4480 19760 4486
rect 19708 4422 19760 4428
rect 19289 4380 19585 4400
rect 19345 4378 19369 4380
rect 19425 4378 19449 4380
rect 19505 4378 19529 4380
rect 19367 4326 19369 4378
rect 19431 4326 19443 4378
rect 19505 4326 19507 4378
rect 19345 4324 19369 4326
rect 19425 4324 19449 4326
rect 19505 4324 19529 4326
rect 19289 4304 19585 4324
rect 19289 3292 19585 3312
rect 19345 3290 19369 3292
rect 19425 3290 19449 3292
rect 19505 3290 19529 3292
rect 19367 3238 19369 3290
rect 19431 3238 19443 3290
rect 19505 3238 19507 3290
rect 19345 3236 19369 3238
rect 19425 3236 19449 3238
rect 19505 3236 19529 3238
rect 19289 3216 19585 3236
rect 19720 3194 19748 4422
rect 19708 3188 19760 3194
rect 19708 3130 19760 3136
rect 19812 2922 19840 6938
rect 19996 6254 20024 8570
rect 19984 6248 20036 6254
rect 19984 6190 20036 6196
rect 19890 4720 19946 4729
rect 19890 4655 19946 4664
rect 19800 2916 19852 2922
rect 19800 2858 19852 2864
rect 19289 2204 19585 2224
rect 19345 2202 19369 2204
rect 19425 2202 19449 2204
rect 19505 2202 19529 2204
rect 19367 2150 19369 2202
rect 19431 2150 19443 2202
rect 19505 2150 19507 2202
rect 19345 2148 19369 2150
rect 19425 2148 19449 2150
rect 19505 2148 19529 2150
rect 19289 2128 19585 2148
rect 19062 54 19196 82
rect 19904 82 19932 4655
rect 19996 1601 20024 6190
rect 20088 5166 20116 8871
rect 20168 7200 20220 7206
rect 20168 7142 20220 7148
rect 20180 5545 20208 7142
rect 21652 7041 21680 11834
rect 21638 7032 21694 7041
rect 21638 6967 21640 6976
rect 21692 6967 21694 6976
rect 21640 6938 21692 6944
rect 21652 6907 21680 6938
rect 20444 6792 20496 6798
rect 20444 6734 20496 6740
rect 20456 6458 20484 6734
rect 20444 6452 20496 6458
rect 20444 6394 20496 6400
rect 20166 5536 20222 5545
rect 20166 5471 20222 5480
rect 20076 5160 20128 5166
rect 20076 5102 20128 5108
rect 20076 2984 20128 2990
rect 20076 2926 20128 2932
rect 20088 2446 20116 2926
rect 20076 2440 20128 2446
rect 20076 2382 20128 2388
rect 21456 2372 21508 2378
rect 21456 2314 21508 2320
rect 19982 1592 20038 1601
rect 19982 1527 20038 1536
rect 20166 82 20222 480
rect 19904 54 20222 82
rect 19062 0 19118 54
rect 20166 0 20222 54
rect 21362 82 21418 480
rect 21468 82 21496 2314
rect 21362 54 21496 82
rect 21362 0 21418 54
<< via2 >>
rect 110 21392 166 21448
rect 1306 19760 1362 19816
rect 202 16632 258 16688
rect 110 15952 166 16008
rect 1582 18672 1638 18728
rect 4622 19610 4678 19612
rect 4702 19610 4758 19612
rect 4782 19610 4838 19612
rect 4862 19610 4918 19612
rect 4622 19558 4648 19610
rect 4648 19558 4678 19610
rect 4702 19558 4712 19610
rect 4712 19558 4758 19610
rect 4782 19558 4828 19610
rect 4828 19558 4838 19610
rect 4862 19558 4892 19610
rect 4892 19558 4918 19610
rect 4622 19556 4678 19558
rect 4702 19556 4758 19558
rect 4782 19556 4838 19558
rect 4862 19556 4918 19558
rect 1582 17584 1638 17640
rect 110 14864 166 14920
rect 2042 15000 2098 15056
rect 110 11600 166 11656
rect 18 10376 74 10432
rect 1950 8608 2006 8664
rect 1306 6568 1362 6624
rect 110 4936 166 4992
rect 3422 19216 3478 19272
rect 4158 19216 4214 19272
rect 2502 14320 2558 14376
rect 2226 13368 2282 13424
rect 2134 11464 2190 11520
rect 2226 7656 2282 7712
rect 2778 17176 2834 17232
rect 1950 3304 2006 3360
rect 3974 13368 4030 13424
rect 3882 11464 3938 11520
rect 4622 18522 4678 18524
rect 4702 18522 4758 18524
rect 4782 18522 4838 18524
rect 4862 18522 4918 18524
rect 4622 18470 4648 18522
rect 4648 18470 4678 18522
rect 4702 18470 4712 18522
rect 4712 18470 4758 18522
rect 4782 18470 4828 18522
rect 4828 18470 4838 18522
rect 4862 18470 4892 18522
rect 4892 18470 4918 18522
rect 4622 18468 4678 18470
rect 4702 18468 4758 18470
rect 4782 18468 4838 18470
rect 4862 18468 4918 18470
rect 4250 16496 4306 16552
rect 4622 17434 4678 17436
rect 4702 17434 4758 17436
rect 4782 17434 4838 17436
rect 4862 17434 4918 17436
rect 4622 17382 4648 17434
rect 4648 17382 4678 17434
rect 4702 17382 4712 17434
rect 4712 17382 4758 17434
rect 4782 17382 4828 17434
rect 4828 17382 4838 17434
rect 4862 17382 4892 17434
rect 4892 17382 4918 17434
rect 4622 17380 4678 17382
rect 4702 17380 4758 17382
rect 4782 17380 4838 17382
rect 4862 17380 4918 17382
rect 4986 16496 5042 16552
rect 4622 16346 4678 16348
rect 4702 16346 4758 16348
rect 4782 16346 4838 16348
rect 4862 16346 4918 16348
rect 4622 16294 4648 16346
rect 4648 16294 4678 16346
rect 4702 16294 4712 16346
rect 4712 16294 4758 16346
rect 4782 16294 4828 16346
rect 4828 16294 4838 16346
rect 4862 16294 4892 16346
rect 4892 16294 4918 16346
rect 4622 16292 4678 16294
rect 4702 16292 4758 16294
rect 4782 16292 4838 16294
rect 4862 16292 4918 16294
rect 4622 15258 4678 15260
rect 4702 15258 4758 15260
rect 4782 15258 4838 15260
rect 4862 15258 4918 15260
rect 4622 15206 4648 15258
rect 4648 15206 4678 15258
rect 4702 15206 4712 15258
rect 4712 15206 4758 15258
rect 4782 15206 4828 15258
rect 4828 15206 4838 15258
rect 4862 15206 4892 15258
rect 4892 15206 4918 15258
rect 4622 15204 4678 15206
rect 4702 15204 4758 15206
rect 4782 15204 4838 15206
rect 4862 15204 4918 15206
rect 3054 5616 3110 5672
rect 3422 3440 3478 3496
rect 3146 2624 3202 2680
rect 4622 14170 4678 14172
rect 4702 14170 4758 14172
rect 4782 14170 4838 14172
rect 4862 14170 4918 14172
rect 4622 14118 4648 14170
rect 4648 14118 4678 14170
rect 4702 14118 4712 14170
rect 4712 14118 4758 14170
rect 4782 14118 4828 14170
rect 4828 14118 4838 14170
rect 4862 14118 4892 14170
rect 4892 14118 4918 14170
rect 4622 14116 4678 14118
rect 4702 14116 4758 14118
rect 4782 14116 4838 14118
rect 4862 14116 4918 14118
rect 4622 13082 4678 13084
rect 4702 13082 4758 13084
rect 4782 13082 4838 13084
rect 4862 13082 4918 13084
rect 4622 13030 4648 13082
rect 4648 13030 4678 13082
rect 4702 13030 4712 13082
rect 4712 13030 4758 13082
rect 4782 13030 4828 13082
rect 4828 13030 4838 13082
rect 4862 13030 4892 13082
rect 4892 13030 4918 13082
rect 4622 13028 4678 13030
rect 4702 13028 4758 13030
rect 4782 13028 4838 13030
rect 4862 13028 4918 13030
rect 4622 11994 4678 11996
rect 4702 11994 4758 11996
rect 4782 11994 4838 11996
rect 4862 11994 4918 11996
rect 4622 11942 4648 11994
rect 4648 11942 4678 11994
rect 4702 11942 4712 11994
rect 4712 11942 4758 11994
rect 4782 11942 4828 11994
rect 4828 11942 4838 11994
rect 4862 11942 4892 11994
rect 4892 11942 4918 11994
rect 4622 11940 4678 11942
rect 4702 11940 4758 11942
rect 4782 11940 4838 11942
rect 4862 11940 4918 11942
rect 4434 11464 4490 11520
rect 4250 8744 4306 8800
rect 4622 10906 4678 10908
rect 4702 10906 4758 10908
rect 4782 10906 4838 10908
rect 4862 10906 4918 10908
rect 4622 10854 4648 10906
rect 4648 10854 4678 10906
rect 4702 10854 4712 10906
rect 4712 10854 4758 10906
rect 4782 10854 4828 10906
rect 4828 10854 4838 10906
rect 4862 10854 4892 10906
rect 4892 10854 4918 10906
rect 4622 10852 4678 10854
rect 4702 10852 4758 10854
rect 4782 10852 4838 10854
rect 4862 10852 4918 10854
rect 4622 9818 4678 9820
rect 4702 9818 4758 9820
rect 4782 9818 4838 9820
rect 4862 9818 4918 9820
rect 4622 9766 4648 9818
rect 4648 9766 4678 9818
rect 4702 9766 4712 9818
rect 4712 9766 4758 9818
rect 4782 9766 4828 9818
rect 4828 9766 4838 9818
rect 4862 9766 4892 9818
rect 4892 9766 4918 9818
rect 4622 9764 4678 9766
rect 4702 9764 4758 9766
rect 4782 9764 4838 9766
rect 4862 9764 4918 9766
rect 4622 8730 4678 8732
rect 4702 8730 4758 8732
rect 4782 8730 4838 8732
rect 4862 8730 4918 8732
rect 4622 8678 4648 8730
rect 4648 8678 4678 8730
rect 4702 8678 4712 8730
rect 4712 8678 4758 8730
rect 4782 8678 4828 8730
rect 4828 8678 4838 8730
rect 4862 8678 4892 8730
rect 4892 8678 4918 8730
rect 4622 8676 4678 8678
rect 4702 8676 4758 8678
rect 4782 8676 4838 8678
rect 4862 8676 4918 8678
rect 5078 8472 5134 8528
rect 4622 7642 4678 7644
rect 4702 7642 4758 7644
rect 4782 7642 4838 7644
rect 4862 7642 4918 7644
rect 4622 7590 4648 7642
rect 4648 7590 4678 7642
rect 4702 7590 4712 7642
rect 4712 7590 4758 7642
rect 4782 7590 4828 7642
rect 4828 7590 4838 7642
rect 4862 7590 4892 7642
rect 4892 7590 4918 7642
rect 4622 7588 4678 7590
rect 4702 7588 4758 7590
rect 4782 7588 4838 7590
rect 4862 7588 4918 7590
rect 4622 6554 4678 6556
rect 4702 6554 4758 6556
rect 4782 6554 4838 6556
rect 4862 6554 4918 6556
rect 4622 6502 4648 6554
rect 4648 6502 4678 6554
rect 4702 6502 4712 6554
rect 4712 6502 4758 6554
rect 4782 6502 4828 6554
rect 4828 6502 4838 6554
rect 4862 6502 4892 6554
rect 4892 6502 4918 6554
rect 4622 6500 4678 6502
rect 4702 6500 4758 6502
rect 4782 6500 4838 6502
rect 4862 6500 4918 6502
rect 4622 5466 4678 5468
rect 4702 5466 4758 5468
rect 4782 5466 4838 5468
rect 4862 5466 4918 5468
rect 4622 5414 4648 5466
rect 4648 5414 4678 5466
rect 4702 5414 4712 5466
rect 4712 5414 4758 5466
rect 4782 5414 4828 5466
rect 4828 5414 4838 5466
rect 4862 5414 4892 5466
rect 4892 5414 4918 5466
rect 4622 5412 4678 5414
rect 4702 5412 4758 5414
rect 4782 5412 4838 5414
rect 4862 5412 4918 5414
rect 4622 4378 4678 4380
rect 4702 4378 4758 4380
rect 4782 4378 4838 4380
rect 4862 4378 4918 4380
rect 4622 4326 4648 4378
rect 4648 4326 4678 4378
rect 4702 4326 4712 4378
rect 4712 4326 4758 4378
rect 4782 4326 4828 4378
rect 4828 4326 4838 4378
rect 4862 4326 4892 4378
rect 4892 4326 4918 4378
rect 4622 4324 4678 4326
rect 4702 4324 4758 4326
rect 4782 4324 4838 4326
rect 4862 4324 4918 4326
rect 5630 13912 5686 13968
rect 5354 11192 5410 11248
rect 5538 11600 5594 11656
rect 5170 4120 5226 4176
rect 5170 3304 5226 3360
rect 4622 3290 4678 3292
rect 4702 3290 4758 3292
rect 4782 3290 4838 3292
rect 4862 3290 4918 3292
rect 4622 3238 4648 3290
rect 4648 3238 4678 3290
rect 4702 3238 4712 3290
rect 4712 3238 4758 3290
rect 4782 3238 4828 3290
rect 4828 3238 4838 3290
rect 4862 3238 4892 3290
rect 4892 3238 4918 3290
rect 4622 3236 4678 3238
rect 4702 3236 4758 3238
rect 4782 3236 4838 3238
rect 4862 3236 4918 3238
rect 5078 3168 5134 3224
rect 5354 3576 5410 3632
rect 4622 2202 4678 2204
rect 4702 2202 4758 2204
rect 4782 2202 4838 2204
rect 4862 2202 4918 2204
rect 4622 2150 4648 2202
rect 4648 2150 4678 2202
rect 4702 2150 4712 2202
rect 4712 2150 4758 2202
rect 4782 2150 4828 2202
rect 4828 2150 4838 2202
rect 4862 2150 4892 2202
rect 4892 2150 4918 2202
rect 4622 2148 4678 2150
rect 4702 2148 4758 2150
rect 4782 2148 4838 2150
rect 4862 2148 4918 2150
rect 6090 11872 6146 11928
rect 5538 1944 5594 2000
rect 6090 3984 6146 4040
rect 6642 14068 6698 14104
rect 6642 14048 6644 14068
rect 6644 14048 6696 14068
rect 6696 14048 6698 14068
rect 6642 13776 6698 13832
rect 6458 11464 6514 11520
rect 8289 19066 8345 19068
rect 8369 19066 8425 19068
rect 8449 19066 8505 19068
rect 8529 19066 8585 19068
rect 8289 19014 8315 19066
rect 8315 19014 8345 19066
rect 8369 19014 8379 19066
rect 8379 19014 8425 19066
rect 8449 19014 8495 19066
rect 8495 19014 8505 19066
rect 8529 19014 8559 19066
rect 8559 19014 8585 19066
rect 8289 19012 8345 19014
rect 8369 19012 8425 19014
rect 8449 19012 8505 19014
rect 8529 19012 8585 19014
rect 7838 17720 7894 17776
rect 6826 5208 6882 5264
rect 6458 4528 6514 4584
rect 6274 3032 6330 3088
rect 8289 17978 8345 17980
rect 8369 17978 8425 17980
rect 8449 17978 8505 17980
rect 8529 17978 8585 17980
rect 8289 17926 8315 17978
rect 8315 17926 8345 17978
rect 8369 17926 8379 17978
rect 8379 17926 8425 17978
rect 8449 17926 8495 17978
rect 8495 17926 8505 17978
rect 8529 17926 8559 17978
rect 8559 17926 8585 17978
rect 8289 17924 8345 17926
rect 8369 17924 8425 17926
rect 8449 17924 8505 17926
rect 8529 17924 8585 17926
rect 8289 16890 8345 16892
rect 8369 16890 8425 16892
rect 8449 16890 8505 16892
rect 8529 16890 8585 16892
rect 8289 16838 8315 16890
rect 8315 16838 8345 16890
rect 8369 16838 8379 16890
rect 8379 16838 8425 16890
rect 8449 16838 8495 16890
rect 8495 16838 8505 16890
rect 8529 16838 8559 16890
rect 8559 16838 8585 16890
rect 8289 16836 8345 16838
rect 8369 16836 8425 16838
rect 8449 16836 8505 16838
rect 8529 16836 8585 16838
rect 8114 16496 8170 16552
rect 7930 12416 7986 12472
rect 8289 15802 8345 15804
rect 8369 15802 8425 15804
rect 8449 15802 8505 15804
rect 8529 15802 8585 15804
rect 8289 15750 8315 15802
rect 8315 15750 8345 15802
rect 8369 15750 8379 15802
rect 8379 15750 8425 15802
rect 8449 15750 8495 15802
rect 8495 15750 8505 15802
rect 8529 15750 8559 15802
rect 8559 15750 8585 15802
rect 8289 15748 8345 15750
rect 8369 15748 8425 15750
rect 8449 15748 8505 15750
rect 8529 15748 8585 15750
rect 8289 14714 8345 14716
rect 8369 14714 8425 14716
rect 8449 14714 8505 14716
rect 8529 14714 8585 14716
rect 8289 14662 8315 14714
rect 8315 14662 8345 14714
rect 8369 14662 8379 14714
rect 8379 14662 8425 14714
rect 8449 14662 8495 14714
rect 8495 14662 8505 14714
rect 8529 14662 8559 14714
rect 8559 14662 8585 14714
rect 8289 14660 8345 14662
rect 8369 14660 8425 14662
rect 8449 14660 8505 14662
rect 8529 14660 8585 14662
rect 8114 13776 8170 13832
rect 8289 13626 8345 13628
rect 8369 13626 8425 13628
rect 8449 13626 8505 13628
rect 8529 13626 8585 13628
rect 8289 13574 8315 13626
rect 8315 13574 8345 13626
rect 8369 13574 8379 13626
rect 8379 13574 8425 13626
rect 8449 13574 8495 13626
rect 8495 13574 8505 13626
rect 8529 13574 8559 13626
rect 8559 13574 8585 13626
rect 8289 13572 8345 13574
rect 8369 13572 8425 13574
rect 8449 13572 8505 13574
rect 8529 13572 8585 13574
rect 11956 19610 12012 19612
rect 12036 19610 12092 19612
rect 12116 19610 12172 19612
rect 12196 19610 12252 19612
rect 11956 19558 11982 19610
rect 11982 19558 12012 19610
rect 12036 19558 12046 19610
rect 12046 19558 12092 19610
rect 12116 19558 12162 19610
rect 12162 19558 12172 19610
rect 12196 19558 12226 19610
rect 12226 19558 12252 19610
rect 11956 19556 12012 19558
rect 12036 19556 12092 19558
rect 12116 19556 12172 19558
rect 12196 19556 12252 19558
rect 8289 12538 8345 12540
rect 8369 12538 8425 12540
rect 8449 12538 8505 12540
rect 8529 12538 8585 12540
rect 8289 12486 8315 12538
rect 8315 12486 8345 12538
rect 8369 12486 8379 12538
rect 8379 12486 8425 12538
rect 8449 12486 8495 12538
rect 8495 12486 8505 12538
rect 8529 12486 8559 12538
rect 8559 12486 8585 12538
rect 8289 12484 8345 12486
rect 8369 12484 8425 12486
rect 8449 12484 8505 12486
rect 8529 12484 8585 12486
rect 8289 11450 8345 11452
rect 8369 11450 8425 11452
rect 8449 11450 8505 11452
rect 8529 11450 8585 11452
rect 8289 11398 8315 11450
rect 8315 11398 8345 11450
rect 8369 11398 8379 11450
rect 8379 11398 8425 11450
rect 8449 11398 8495 11450
rect 8495 11398 8505 11450
rect 8529 11398 8559 11450
rect 8559 11398 8585 11450
rect 8289 11396 8345 11398
rect 8369 11396 8425 11398
rect 8449 11396 8505 11398
rect 8529 11396 8585 11398
rect 8289 10362 8345 10364
rect 8369 10362 8425 10364
rect 8449 10362 8505 10364
rect 8529 10362 8585 10364
rect 8289 10310 8315 10362
rect 8315 10310 8345 10362
rect 8369 10310 8379 10362
rect 8379 10310 8425 10362
rect 8449 10310 8495 10362
rect 8495 10310 8505 10362
rect 8529 10310 8559 10362
rect 8559 10310 8585 10362
rect 8289 10308 8345 10310
rect 8369 10308 8425 10310
rect 8449 10308 8505 10310
rect 8529 10308 8585 10310
rect 9034 15000 9090 15056
rect 9310 17176 9366 17232
rect 9034 13640 9090 13696
rect 9126 10648 9182 10704
rect 9034 9968 9090 10024
rect 8666 9288 8722 9344
rect 8289 9274 8345 9276
rect 8369 9274 8425 9276
rect 8449 9274 8505 9276
rect 8529 9274 8585 9276
rect 8289 9222 8315 9274
rect 8315 9222 8345 9274
rect 8369 9222 8379 9274
rect 8379 9222 8425 9274
rect 8449 9222 8495 9274
rect 8495 9222 8505 9274
rect 8529 9222 8559 9274
rect 8559 9222 8585 9274
rect 8289 9220 8345 9222
rect 8369 9220 8425 9222
rect 8449 9220 8505 9222
rect 8529 9220 8585 9222
rect 8666 8608 8722 8664
rect 8289 8186 8345 8188
rect 8369 8186 8425 8188
rect 8449 8186 8505 8188
rect 8529 8186 8585 8188
rect 8289 8134 8315 8186
rect 8315 8134 8345 8186
rect 8369 8134 8379 8186
rect 8379 8134 8425 8186
rect 8449 8134 8495 8186
rect 8495 8134 8505 8186
rect 8529 8134 8559 8186
rect 8559 8134 8585 8186
rect 8289 8132 8345 8134
rect 8369 8132 8425 8134
rect 8449 8132 8505 8134
rect 8529 8132 8585 8134
rect 7470 7248 7526 7304
rect 8666 7112 8722 7168
rect 8289 7098 8345 7100
rect 8369 7098 8425 7100
rect 8449 7098 8505 7100
rect 8529 7098 8585 7100
rect 8289 7046 8315 7098
rect 8315 7046 8345 7098
rect 8369 7046 8379 7098
rect 8379 7046 8425 7098
rect 8449 7046 8495 7098
rect 8495 7046 8505 7098
rect 8529 7046 8559 7098
rect 8559 7046 8585 7098
rect 8289 7044 8345 7046
rect 8369 7044 8425 7046
rect 8449 7044 8505 7046
rect 8529 7044 8585 7046
rect 8482 6704 8538 6760
rect 8289 6010 8345 6012
rect 8369 6010 8425 6012
rect 8449 6010 8505 6012
rect 8529 6010 8585 6012
rect 8289 5958 8315 6010
rect 8315 5958 8345 6010
rect 8369 5958 8379 6010
rect 8379 5958 8425 6010
rect 8449 5958 8495 6010
rect 8495 5958 8505 6010
rect 8529 5958 8559 6010
rect 8559 5958 8585 6010
rect 8289 5956 8345 5958
rect 8369 5956 8425 5958
rect 8449 5956 8505 5958
rect 8529 5956 8585 5958
rect 8289 4922 8345 4924
rect 8369 4922 8425 4924
rect 8449 4922 8505 4924
rect 8529 4922 8585 4924
rect 8289 4870 8315 4922
rect 8315 4870 8345 4922
rect 8369 4870 8379 4922
rect 8379 4870 8425 4922
rect 8449 4870 8495 4922
rect 8495 4870 8505 4922
rect 8529 4870 8559 4922
rect 8559 4870 8585 4922
rect 8289 4868 8345 4870
rect 8369 4868 8425 4870
rect 8449 4868 8505 4870
rect 8529 4868 8585 4870
rect 7194 2624 7250 2680
rect 6366 2352 6422 2408
rect 5630 1672 5686 1728
rect 5446 1128 5502 1184
rect 5170 40 5226 96
rect 8289 3834 8345 3836
rect 8369 3834 8425 3836
rect 8449 3834 8505 3836
rect 8529 3834 8585 3836
rect 8289 3782 8315 3834
rect 8315 3782 8345 3834
rect 8369 3782 8379 3834
rect 8379 3782 8425 3834
rect 8449 3782 8495 3834
rect 8495 3782 8505 3834
rect 8529 3782 8559 3834
rect 8559 3782 8585 3834
rect 8289 3780 8345 3782
rect 8369 3780 8425 3782
rect 8449 3780 8505 3782
rect 8529 3780 8585 3782
rect 8942 4800 8998 4856
rect 8289 2746 8345 2748
rect 8369 2746 8425 2748
rect 8449 2746 8505 2748
rect 8529 2746 8585 2748
rect 8289 2694 8315 2746
rect 8315 2694 8345 2746
rect 8369 2694 8379 2746
rect 8379 2694 8425 2746
rect 8449 2694 8495 2746
rect 8495 2694 8505 2746
rect 8529 2694 8559 2746
rect 8559 2694 8585 2746
rect 8289 2692 8345 2694
rect 8369 2692 8425 2694
rect 8449 2692 8505 2694
rect 8529 2692 8585 2694
rect 7562 1536 7618 1592
rect 9034 3440 9090 3496
rect 9494 15272 9550 15328
rect 9678 16496 9734 16552
rect 9770 15816 9826 15872
rect 10414 16904 10470 16960
rect 9770 13640 9826 13696
rect 9770 13504 9826 13560
rect 9678 11056 9734 11112
rect 9586 10648 9642 10704
rect 9586 8064 9642 8120
rect 9862 9560 9918 9616
rect 9218 3440 9274 3496
rect 9678 5616 9734 5672
rect 10322 9016 10378 9072
rect 10230 7384 10286 7440
rect 10414 5752 10470 5808
rect 11150 15036 11152 15056
rect 11152 15036 11204 15056
rect 11204 15036 11206 15056
rect 11150 15000 11206 15036
rect 11058 13232 11114 13288
rect 10966 9424 11022 9480
rect 9126 3168 9182 3224
rect 10046 3304 10102 3360
rect 9954 2896 10010 2952
rect 10782 5208 10838 5264
rect 11150 11464 11206 11520
rect 11150 10512 11206 10568
rect 11518 14456 11574 14512
rect 11334 13368 11390 13424
rect 11956 18522 12012 18524
rect 12036 18522 12092 18524
rect 12116 18522 12172 18524
rect 12196 18522 12252 18524
rect 11956 18470 11982 18522
rect 11982 18470 12012 18522
rect 12036 18470 12046 18522
rect 12046 18470 12092 18522
rect 12116 18470 12162 18522
rect 12162 18470 12172 18522
rect 12196 18470 12226 18522
rect 12226 18470 12252 18522
rect 11956 18468 12012 18470
rect 12036 18468 12092 18470
rect 12116 18468 12172 18470
rect 12196 18468 12252 18470
rect 11956 17434 12012 17436
rect 12036 17434 12092 17436
rect 12116 17434 12172 17436
rect 12196 17434 12252 17436
rect 11956 17382 11982 17434
rect 11982 17382 12012 17434
rect 12036 17382 12046 17434
rect 12046 17382 12092 17434
rect 12116 17382 12162 17434
rect 12162 17382 12172 17434
rect 12196 17382 12226 17434
rect 12226 17382 12252 17434
rect 11956 17380 12012 17382
rect 12036 17380 12092 17382
rect 12116 17380 12172 17382
rect 12196 17380 12252 17382
rect 11956 16346 12012 16348
rect 12036 16346 12092 16348
rect 12116 16346 12172 16348
rect 12196 16346 12252 16348
rect 11956 16294 11982 16346
rect 11982 16294 12012 16346
rect 12036 16294 12046 16346
rect 12046 16294 12092 16346
rect 12116 16294 12162 16346
rect 12162 16294 12172 16346
rect 12196 16294 12226 16346
rect 12226 16294 12252 16346
rect 11956 16292 12012 16294
rect 12036 16292 12092 16294
rect 12116 16292 12172 16294
rect 12196 16292 12252 16294
rect 11956 15258 12012 15260
rect 12036 15258 12092 15260
rect 12116 15258 12172 15260
rect 12196 15258 12252 15260
rect 11956 15206 11982 15258
rect 11982 15206 12012 15258
rect 12036 15206 12046 15258
rect 12046 15206 12092 15258
rect 12116 15206 12162 15258
rect 12162 15206 12172 15258
rect 12196 15206 12226 15258
rect 12226 15206 12252 15258
rect 11956 15204 12012 15206
rect 12036 15204 12092 15206
rect 12116 15204 12172 15206
rect 12196 15204 12252 15206
rect 11610 14048 11666 14104
rect 11956 14170 12012 14172
rect 12036 14170 12092 14172
rect 12116 14170 12172 14172
rect 12196 14170 12252 14172
rect 11956 14118 11982 14170
rect 11982 14118 12012 14170
rect 12036 14118 12046 14170
rect 12046 14118 12092 14170
rect 12116 14118 12162 14170
rect 12162 14118 12172 14170
rect 12196 14118 12226 14170
rect 12226 14118 12252 14170
rect 11956 14116 12012 14118
rect 12036 14116 12092 14118
rect 12116 14116 12172 14118
rect 12196 14116 12252 14118
rect 11956 13082 12012 13084
rect 12036 13082 12092 13084
rect 12116 13082 12172 13084
rect 12196 13082 12252 13084
rect 11956 13030 11982 13082
rect 11982 13030 12012 13082
rect 12036 13030 12046 13082
rect 12046 13030 12092 13082
rect 12116 13030 12162 13082
rect 12162 13030 12172 13082
rect 12196 13030 12226 13082
rect 12226 13030 12252 13082
rect 11956 13028 12012 13030
rect 12036 13028 12092 13030
rect 12116 13028 12172 13030
rect 12196 13028 12252 13030
rect 11956 11994 12012 11996
rect 12036 11994 12092 11996
rect 12116 11994 12172 11996
rect 12196 11994 12252 11996
rect 11956 11942 11982 11994
rect 11982 11942 12012 11994
rect 12036 11942 12046 11994
rect 12046 11942 12092 11994
rect 12116 11942 12162 11994
rect 12162 11942 12172 11994
rect 12196 11942 12226 11994
rect 12226 11942 12252 11994
rect 11956 11940 12012 11942
rect 12036 11940 12092 11942
rect 12116 11940 12172 11942
rect 12196 11940 12252 11942
rect 11956 10906 12012 10908
rect 12036 10906 12092 10908
rect 12116 10906 12172 10908
rect 12196 10906 12252 10908
rect 11956 10854 11982 10906
rect 11982 10854 12012 10906
rect 12036 10854 12046 10906
rect 12046 10854 12092 10906
rect 12116 10854 12162 10906
rect 12162 10854 12172 10906
rect 12196 10854 12226 10906
rect 12226 10854 12252 10906
rect 11956 10852 12012 10854
rect 12036 10852 12092 10854
rect 12116 10852 12172 10854
rect 12196 10852 12252 10854
rect 15622 19066 15678 19068
rect 15702 19066 15758 19068
rect 15782 19066 15838 19068
rect 15862 19066 15918 19068
rect 15622 19014 15648 19066
rect 15648 19014 15678 19066
rect 15702 19014 15712 19066
rect 15712 19014 15758 19066
rect 15782 19014 15828 19066
rect 15828 19014 15838 19066
rect 15862 19014 15892 19066
rect 15892 19014 15918 19066
rect 15622 19012 15678 19014
rect 15702 19012 15758 19014
rect 15782 19012 15838 19014
rect 15862 19012 15918 19014
rect 13082 14456 13138 14512
rect 12714 11600 12770 11656
rect 11956 9818 12012 9820
rect 12036 9818 12092 9820
rect 12116 9818 12172 9820
rect 12196 9818 12252 9820
rect 11956 9766 11982 9818
rect 11982 9766 12012 9818
rect 12036 9766 12046 9818
rect 12046 9766 12092 9818
rect 12116 9766 12162 9818
rect 12162 9766 12172 9818
rect 12196 9766 12226 9818
rect 12226 9766 12252 9818
rect 11956 9764 12012 9766
rect 12036 9764 12092 9766
rect 12116 9764 12172 9766
rect 12196 9764 12252 9766
rect 11956 8730 12012 8732
rect 12036 8730 12092 8732
rect 12116 8730 12172 8732
rect 12196 8730 12252 8732
rect 11956 8678 11982 8730
rect 11982 8678 12012 8730
rect 12036 8678 12046 8730
rect 12046 8678 12092 8730
rect 12116 8678 12162 8730
rect 12162 8678 12172 8730
rect 12196 8678 12226 8730
rect 12226 8678 12252 8730
rect 11956 8676 12012 8678
rect 12036 8676 12092 8678
rect 12116 8676 12172 8678
rect 12196 8676 12252 8678
rect 11956 7642 12012 7644
rect 12036 7642 12092 7644
rect 12116 7642 12172 7644
rect 12196 7642 12252 7644
rect 11956 7590 11982 7642
rect 11982 7590 12012 7642
rect 12036 7590 12046 7642
rect 12046 7590 12092 7642
rect 12116 7590 12162 7642
rect 12162 7590 12172 7642
rect 12196 7590 12226 7642
rect 12226 7590 12252 7642
rect 11956 7588 12012 7590
rect 12036 7588 12092 7590
rect 12116 7588 12172 7590
rect 12196 7588 12252 7590
rect 11150 3576 11206 3632
rect 11956 6554 12012 6556
rect 12036 6554 12092 6556
rect 12116 6554 12172 6556
rect 12196 6554 12252 6556
rect 11956 6502 11982 6554
rect 11982 6502 12012 6554
rect 12036 6502 12046 6554
rect 12046 6502 12092 6554
rect 12116 6502 12162 6554
rect 12162 6502 12172 6554
rect 12196 6502 12226 6554
rect 12226 6502 12252 6554
rect 11956 6500 12012 6502
rect 12036 6500 12092 6502
rect 12116 6500 12172 6502
rect 12196 6500 12252 6502
rect 11956 5466 12012 5468
rect 12036 5466 12092 5468
rect 12116 5466 12172 5468
rect 12196 5466 12252 5468
rect 11956 5414 11982 5466
rect 11982 5414 12012 5466
rect 12036 5414 12046 5466
rect 12046 5414 12092 5466
rect 12116 5414 12162 5466
rect 12162 5414 12172 5466
rect 12196 5414 12226 5466
rect 12226 5414 12252 5466
rect 11956 5412 12012 5414
rect 12036 5412 12092 5414
rect 12116 5412 12172 5414
rect 12196 5412 12252 5414
rect 11956 4378 12012 4380
rect 12036 4378 12092 4380
rect 12116 4378 12172 4380
rect 12196 4378 12252 4380
rect 11956 4326 11982 4378
rect 11982 4326 12012 4378
rect 12036 4326 12046 4378
rect 12046 4326 12092 4378
rect 12116 4326 12162 4378
rect 12162 4326 12172 4378
rect 12196 4326 12226 4378
rect 12226 4326 12252 4378
rect 11956 4324 12012 4326
rect 12036 4324 12092 4326
rect 12116 4324 12172 4326
rect 12196 4324 12252 4326
rect 12346 4004 12402 4040
rect 12346 3984 12348 4004
rect 12348 3984 12400 4004
rect 12400 3984 12402 4004
rect 11956 3290 12012 3292
rect 12036 3290 12092 3292
rect 12116 3290 12172 3292
rect 12196 3290 12252 3292
rect 11956 3238 11982 3290
rect 11982 3238 12012 3290
rect 12036 3238 12046 3290
rect 12046 3238 12092 3290
rect 12116 3238 12162 3290
rect 12162 3238 12172 3290
rect 12196 3238 12226 3290
rect 12226 3238 12252 3290
rect 11956 3236 12012 3238
rect 12036 3236 12092 3238
rect 12116 3236 12172 3238
rect 12196 3236 12252 3238
rect 13266 13368 13322 13424
rect 13450 13504 13506 13560
rect 14186 17720 14242 17776
rect 13726 14184 13782 14240
rect 13634 11192 13690 11248
rect 14094 16496 14150 16552
rect 14278 15816 14334 15872
rect 14554 16632 14610 16688
rect 15622 17978 15678 17980
rect 15702 17978 15758 17980
rect 15782 17978 15838 17980
rect 15862 17978 15918 17980
rect 15622 17926 15648 17978
rect 15648 17926 15678 17978
rect 15702 17926 15712 17978
rect 15712 17926 15758 17978
rect 15782 17926 15828 17978
rect 15828 17926 15838 17978
rect 15862 17926 15892 17978
rect 15892 17926 15918 17978
rect 15622 17924 15678 17926
rect 15702 17924 15758 17926
rect 15782 17924 15838 17926
rect 15862 17924 15918 17926
rect 14738 16088 14794 16144
rect 13910 10784 13966 10840
rect 14094 9560 14150 9616
rect 14094 8880 14150 8936
rect 14738 13504 14794 13560
rect 13082 3304 13138 3360
rect 11956 2202 12012 2204
rect 12036 2202 12092 2204
rect 12116 2202 12172 2204
rect 12196 2202 12252 2204
rect 11956 2150 11982 2202
rect 11982 2150 12012 2202
rect 12036 2150 12046 2202
rect 12046 2150 12092 2202
rect 12116 2150 12162 2202
rect 12162 2150 12172 2202
rect 12196 2150 12226 2202
rect 12226 2150 12252 2202
rect 11956 2148 12012 2150
rect 12036 2148 12092 2150
rect 12116 2148 12172 2150
rect 12196 2148 12252 2150
rect 15622 16890 15678 16892
rect 15702 16890 15758 16892
rect 15782 16890 15838 16892
rect 15862 16890 15918 16892
rect 15622 16838 15648 16890
rect 15648 16838 15678 16890
rect 15702 16838 15712 16890
rect 15712 16838 15758 16890
rect 15782 16838 15828 16890
rect 15828 16838 15838 16890
rect 15862 16838 15892 16890
rect 15892 16838 15918 16890
rect 15622 16836 15678 16838
rect 15702 16836 15758 16838
rect 15782 16836 15838 16838
rect 15862 16836 15918 16838
rect 15622 15802 15678 15804
rect 15702 15802 15758 15804
rect 15782 15802 15838 15804
rect 15862 15802 15918 15804
rect 15622 15750 15648 15802
rect 15648 15750 15678 15802
rect 15702 15750 15712 15802
rect 15712 15750 15758 15802
rect 15782 15750 15828 15802
rect 15828 15750 15838 15802
rect 15862 15750 15892 15802
rect 15892 15750 15918 15802
rect 15622 15748 15678 15750
rect 15702 15748 15758 15750
rect 15782 15748 15838 15750
rect 15862 15748 15918 15750
rect 15290 14864 15346 14920
rect 15198 13640 15254 13696
rect 15198 13368 15254 13424
rect 15622 14714 15678 14716
rect 15702 14714 15758 14716
rect 15782 14714 15838 14716
rect 15862 14714 15918 14716
rect 15622 14662 15648 14714
rect 15648 14662 15678 14714
rect 15702 14662 15712 14714
rect 15712 14662 15758 14714
rect 15782 14662 15828 14714
rect 15828 14662 15838 14714
rect 15862 14662 15892 14714
rect 15892 14662 15918 14714
rect 15622 14660 15678 14662
rect 15702 14660 15758 14662
rect 15782 14660 15838 14662
rect 15862 14660 15918 14662
rect 15934 14320 15990 14376
rect 15622 13626 15678 13628
rect 15702 13626 15758 13628
rect 15782 13626 15838 13628
rect 15862 13626 15918 13628
rect 15622 13574 15648 13626
rect 15648 13574 15678 13626
rect 15702 13574 15712 13626
rect 15712 13574 15758 13626
rect 15782 13574 15828 13626
rect 15828 13574 15838 13626
rect 15862 13574 15892 13626
rect 15892 13574 15918 13626
rect 15622 13572 15678 13574
rect 15702 13572 15758 13574
rect 15782 13572 15838 13574
rect 15862 13572 15918 13574
rect 15622 12538 15678 12540
rect 15702 12538 15758 12540
rect 15782 12538 15838 12540
rect 15862 12538 15918 12540
rect 15622 12486 15648 12538
rect 15648 12486 15678 12538
rect 15702 12486 15712 12538
rect 15712 12486 15758 12538
rect 15782 12486 15828 12538
rect 15828 12486 15838 12538
rect 15862 12486 15892 12538
rect 15892 12486 15918 12538
rect 15622 12484 15678 12486
rect 15702 12484 15758 12486
rect 15782 12484 15838 12486
rect 15862 12484 15918 12486
rect 15622 11450 15678 11452
rect 15702 11450 15758 11452
rect 15782 11450 15838 11452
rect 15862 11450 15918 11452
rect 15622 11398 15648 11450
rect 15648 11398 15678 11450
rect 15702 11398 15712 11450
rect 15712 11398 15758 11450
rect 15782 11398 15828 11450
rect 15828 11398 15838 11450
rect 15862 11398 15892 11450
rect 15892 11398 15918 11450
rect 15622 11396 15678 11398
rect 15702 11396 15758 11398
rect 15782 11396 15838 11398
rect 15862 11396 15918 11398
rect 15622 10362 15678 10364
rect 15702 10362 15758 10364
rect 15782 10362 15838 10364
rect 15862 10362 15918 10364
rect 15622 10310 15648 10362
rect 15648 10310 15678 10362
rect 15702 10310 15712 10362
rect 15712 10310 15758 10362
rect 15782 10310 15828 10362
rect 15828 10310 15838 10362
rect 15862 10310 15892 10362
rect 15892 10310 15918 10362
rect 15622 10308 15678 10310
rect 15702 10308 15758 10310
rect 15782 10308 15838 10310
rect 15862 10308 15918 10310
rect 14922 7792 14978 7848
rect 15198 7112 15254 7168
rect 14186 4800 14242 4856
rect 14278 4664 14334 4720
rect 15198 1944 15254 2000
rect 15622 9274 15678 9276
rect 15702 9274 15758 9276
rect 15782 9274 15838 9276
rect 15862 9274 15918 9276
rect 15622 9222 15648 9274
rect 15648 9222 15678 9274
rect 15702 9222 15712 9274
rect 15712 9222 15758 9274
rect 15782 9222 15828 9274
rect 15828 9222 15838 9274
rect 15862 9222 15892 9274
rect 15892 9222 15918 9274
rect 15622 9220 15678 9222
rect 15702 9220 15758 9222
rect 15782 9220 15838 9222
rect 15862 9220 15918 9222
rect 15622 8186 15678 8188
rect 15702 8186 15758 8188
rect 15782 8186 15838 8188
rect 15862 8186 15918 8188
rect 15622 8134 15648 8186
rect 15648 8134 15678 8186
rect 15702 8134 15712 8186
rect 15712 8134 15758 8186
rect 15782 8134 15828 8186
rect 15828 8134 15838 8186
rect 15862 8134 15892 8186
rect 15892 8134 15918 8186
rect 15622 8132 15678 8134
rect 15702 8132 15758 8134
rect 15782 8132 15838 8134
rect 15862 8132 15918 8134
rect 15474 8064 15530 8120
rect 16026 13640 16082 13696
rect 16394 20440 16450 20496
rect 19289 19610 19345 19612
rect 19369 19610 19425 19612
rect 19449 19610 19505 19612
rect 19529 19610 19585 19612
rect 19289 19558 19315 19610
rect 19315 19558 19345 19610
rect 19369 19558 19379 19610
rect 19379 19558 19425 19610
rect 19449 19558 19495 19610
rect 19495 19558 19505 19610
rect 19529 19558 19559 19610
rect 19559 19558 19585 19610
rect 19289 19556 19345 19558
rect 19369 19556 19425 19558
rect 19449 19556 19505 19558
rect 19529 19556 19585 19558
rect 16670 13776 16726 13832
rect 16578 13232 16634 13288
rect 16394 7384 16450 7440
rect 15622 7098 15678 7100
rect 15702 7098 15758 7100
rect 15782 7098 15838 7100
rect 15862 7098 15918 7100
rect 15622 7046 15648 7098
rect 15648 7046 15678 7098
rect 15702 7046 15712 7098
rect 15712 7046 15758 7098
rect 15782 7046 15828 7098
rect 15828 7046 15838 7098
rect 15862 7046 15892 7098
rect 15892 7046 15918 7098
rect 15622 7044 15678 7046
rect 15702 7044 15758 7046
rect 15782 7044 15838 7046
rect 15862 7044 15918 7046
rect 15622 6010 15678 6012
rect 15702 6010 15758 6012
rect 15782 6010 15838 6012
rect 15862 6010 15918 6012
rect 15622 5958 15648 6010
rect 15648 5958 15678 6010
rect 15702 5958 15712 6010
rect 15712 5958 15758 6010
rect 15782 5958 15828 6010
rect 15828 5958 15838 6010
rect 15862 5958 15892 6010
rect 15892 5958 15918 6010
rect 15622 5956 15678 5958
rect 15702 5956 15758 5958
rect 15782 5956 15838 5958
rect 15862 5956 15918 5958
rect 15622 4922 15678 4924
rect 15702 4922 15758 4924
rect 15782 4922 15838 4924
rect 15862 4922 15918 4924
rect 15622 4870 15648 4922
rect 15648 4870 15678 4922
rect 15702 4870 15712 4922
rect 15712 4870 15758 4922
rect 15782 4870 15828 4922
rect 15828 4870 15838 4922
rect 15862 4870 15892 4922
rect 15892 4870 15918 4922
rect 15622 4868 15678 4870
rect 15702 4868 15758 4870
rect 15782 4868 15838 4870
rect 15862 4868 15918 4870
rect 15622 3834 15678 3836
rect 15702 3834 15758 3836
rect 15782 3834 15838 3836
rect 15862 3834 15918 3836
rect 15622 3782 15648 3834
rect 15648 3782 15678 3834
rect 15702 3782 15712 3834
rect 15712 3782 15758 3834
rect 15782 3782 15828 3834
rect 15828 3782 15838 3834
rect 15862 3782 15892 3834
rect 15892 3782 15918 3834
rect 15622 3780 15678 3782
rect 15702 3780 15758 3782
rect 15782 3780 15838 3782
rect 15862 3780 15918 3782
rect 16854 13368 16910 13424
rect 16026 3884 16028 3904
rect 16028 3884 16080 3904
rect 16080 3884 16082 3904
rect 16026 3848 16082 3884
rect 15622 2746 15678 2748
rect 15702 2746 15758 2748
rect 15782 2746 15838 2748
rect 15862 2746 15918 2748
rect 15622 2694 15648 2746
rect 15648 2694 15678 2746
rect 15702 2694 15712 2746
rect 15712 2694 15758 2746
rect 15782 2694 15828 2746
rect 15828 2694 15838 2746
rect 15862 2694 15892 2746
rect 15892 2694 15918 2746
rect 15622 2692 15678 2694
rect 15702 2692 15758 2694
rect 15782 2692 15838 2694
rect 15862 2692 15918 2694
rect 16486 3440 16542 3496
rect 16670 3440 16726 3496
rect 17958 16088 18014 16144
rect 17774 15000 17830 15056
rect 17590 14864 17646 14920
rect 17498 10648 17554 10704
rect 18418 14476 18474 14512
rect 18418 14456 18420 14476
rect 18420 14456 18472 14476
rect 18472 14456 18474 14476
rect 17590 9016 17646 9072
rect 17314 7248 17370 7304
rect 17774 9460 17776 9480
rect 17776 9460 17828 9480
rect 17828 9460 17830 9480
rect 17774 9424 17830 9460
rect 18418 13368 18474 13424
rect 18142 9560 18198 9616
rect 19289 18522 19345 18524
rect 19369 18522 19425 18524
rect 19449 18522 19505 18524
rect 19529 18522 19585 18524
rect 19289 18470 19315 18522
rect 19315 18470 19345 18522
rect 19369 18470 19379 18522
rect 19379 18470 19425 18522
rect 19449 18470 19495 18522
rect 19495 18470 19505 18522
rect 19529 18470 19559 18522
rect 19559 18470 19585 18522
rect 19289 18468 19345 18470
rect 19369 18468 19425 18470
rect 19449 18468 19505 18470
rect 19529 18468 19585 18470
rect 19798 18400 19854 18456
rect 19289 17434 19345 17436
rect 19369 17434 19425 17436
rect 19449 17434 19505 17436
rect 19529 17434 19585 17436
rect 19289 17382 19315 17434
rect 19315 17382 19345 17434
rect 19369 17382 19379 17434
rect 19379 17382 19425 17434
rect 19449 17382 19495 17434
rect 19495 17382 19505 17434
rect 19529 17382 19559 17434
rect 19559 17382 19585 17434
rect 19289 17380 19345 17382
rect 19369 17380 19425 17382
rect 19449 17380 19505 17382
rect 19529 17380 19585 17382
rect 19614 16496 19670 16552
rect 19289 16346 19345 16348
rect 19369 16346 19425 16348
rect 19449 16346 19505 16348
rect 19529 16346 19585 16348
rect 19289 16294 19315 16346
rect 19315 16294 19345 16346
rect 19369 16294 19379 16346
rect 19379 16294 19425 16346
rect 19449 16294 19495 16346
rect 19495 16294 19505 16346
rect 19529 16294 19559 16346
rect 19559 16294 19585 16346
rect 19289 16292 19345 16294
rect 19369 16292 19425 16294
rect 19449 16292 19505 16294
rect 19529 16292 19585 16294
rect 18510 11056 18566 11112
rect 18602 10784 18658 10840
rect 18234 8472 18290 8528
rect 17866 6704 17922 6760
rect 17130 3848 17186 3904
rect 17038 3032 17094 3088
rect 18142 5752 18198 5808
rect 18050 5208 18106 5264
rect 17774 5108 17776 5128
rect 17776 5108 17828 5128
rect 17828 5108 17830 5128
rect 17774 5072 17830 5108
rect 18786 9968 18842 10024
rect 18510 4528 18566 4584
rect 18050 3984 18106 4040
rect 18142 3576 18198 3632
rect 17774 2932 17776 2952
rect 17776 2932 17828 2952
rect 17828 2932 17830 2952
rect 17774 2896 17830 2932
rect 18142 2352 18198 2408
rect 19289 15258 19345 15260
rect 19369 15258 19425 15260
rect 19449 15258 19505 15260
rect 19529 15258 19585 15260
rect 19289 15206 19315 15258
rect 19315 15206 19345 15258
rect 19369 15206 19379 15258
rect 19379 15206 19425 15258
rect 19449 15206 19495 15258
rect 19495 15206 19505 15258
rect 19529 15206 19559 15258
rect 19559 15206 19585 15258
rect 19289 15204 19345 15206
rect 19369 15204 19425 15206
rect 19449 15204 19505 15206
rect 19529 15204 19585 15206
rect 19289 14170 19345 14172
rect 19369 14170 19425 14172
rect 19449 14170 19505 14172
rect 19529 14170 19585 14172
rect 19289 14118 19315 14170
rect 19315 14118 19345 14170
rect 19369 14118 19379 14170
rect 19379 14118 19425 14170
rect 19449 14118 19495 14170
rect 19495 14118 19505 14170
rect 19529 14118 19559 14170
rect 19559 14118 19585 14170
rect 19289 14116 19345 14118
rect 19369 14116 19425 14118
rect 19449 14116 19505 14118
rect 19529 14116 19585 14118
rect 20166 15000 20222 15056
rect 19289 13082 19345 13084
rect 19369 13082 19425 13084
rect 19449 13082 19505 13084
rect 19529 13082 19585 13084
rect 19289 13030 19315 13082
rect 19315 13030 19345 13082
rect 19369 13030 19379 13082
rect 19379 13030 19425 13082
rect 19449 13030 19495 13082
rect 19495 13030 19505 13082
rect 19529 13030 19559 13082
rect 19559 13030 19585 13082
rect 19289 13028 19345 13030
rect 19369 13028 19425 13030
rect 19449 13028 19505 13030
rect 19529 13028 19585 13030
rect 19289 11994 19345 11996
rect 19369 11994 19425 11996
rect 19449 11994 19505 11996
rect 19529 11994 19585 11996
rect 19289 11942 19315 11994
rect 19315 11942 19345 11994
rect 19369 11942 19379 11994
rect 19379 11942 19425 11994
rect 19449 11942 19495 11994
rect 19495 11942 19505 11994
rect 19529 11942 19559 11994
rect 19559 11942 19585 11994
rect 19289 11940 19345 11942
rect 19369 11940 19425 11942
rect 19449 11940 19505 11942
rect 19529 11940 19585 11942
rect 19289 10906 19345 10908
rect 19369 10906 19425 10908
rect 19449 10906 19505 10908
rect 19529 10906 19585 10908
rect 19289 10854 19315 10906
rect 19315 10854 19345 10906
rect 19369 10854 19379 10906
rect 19379 10854 19425 10906
rect 19449 10854 19495 10906
rect 19495 10854 19505 10906
rect 19529 10854 19559 10906
rect 19559 10854 19585 10906
rect 19289 10852 19345 10854
rect 19369 10852 19425 10854
rect 19449 10852 19505 10854
rect 19529 10852 19585 10854
rect 19289 9818 19345 9820
rect 19369 9818 19425 9820
rect 19449 9818 19505 9820
rect 19529 9818 19585 9820
rect 19289 9766 19315 9818
rect 19315 9766 19345 9818
rect 19369 9766 19379 9818
rect 19379 9766 19425 9818
rect 19449 9766 19495 9818
rect 19495 9766 19505 9818
rect 19529 9766 19559 9818
rect 19559 9766 19585 9818
rect 19289 9764 19345 9766
rect 19369 9764 19425 9766
rect 19449 9764 19505 9766
rect 19529 9764 19585 9766
rect 18602 3304 18658 3360
rect 18786 2624 18842 2680
rect 18510 1672 18566 1728
rect 18418 1536 18474 1592
rect 19289 8730 19345 8732
rect 19369 8730 19425 8732
rect 19449 8730 19505 8732
rect 19529 8730 19585 8732
rect 19289 8678 19315 8730
rect 19315 8678 19345 8730
rect 19369 8678 19379 8730
rect 19379 8678 19425 8730
rect 19449 8678 19495 8730
rect 19495 8678 19505 8730
rect 19529 8678 19559 8730
rect 19559 8678 19585 8730
rect 19289 8676 19345 8678
rect 19369 8676 19425 8678
rect 19449 8676 19505 8678
rect 19529 8676 19585 8678
rect 19289 7642 19345 7644
rect 19369 7642 19425 7644
rect 19449 7642 19505 7644
rect 19529 7642 19585 7644
rect 19289 7590 19315 7642
rect 19315 7590 19345 7642
rect 19369 7590 19379 7642
rect 19379 7590 19425 7642
rect 19449 7590 19495 7642
rect 19495 7590 19505 7642
rect 19529 7590 19559 7642
rect 19559 7590 19585 7642
rect 19289 7588 19345 7590
rect 19369 7588 19425 7590
rect 19449 7588 19505 7590
rect 19529 7588 19585 7590
rect 20074 8880 20130 8936
rect 21546 8880 21602 8936
rect 19706 7792 19762 7848
rect 19289 6554 19345 6556
rect 19369 6554 19425 6556
rect 19449 6554 19505 6556
rect 19529 6554 19585 6556
rect 19289 6502 19315 6554
rect 19315 6502 19345 6554
rect 19369 6502 19379 6554
rect 19379 6502 19425 6554
rect 19449 6502 19495 6554
rect 19495 6502 19505 6554
rect 19529 6502 19559 6554
rect 19559 6502 19585 6554
rect 19289 6500 19345 6502
rect 19369 6500 19425 6502
rect 19449 6500 19505 6502
rect 19529 6500 19585 6502
rect 19289 5466 19345 5468
rect 19369 5466 19425 5468
rect 19449 5466 19505 5468
rect 19529 5466 19585 5468
rect 19289 5414 19315 5466
rect 19315 5414 19345 5466
rect 19369 5414 19379 5466
rect 19379 5414 19425 5466
rect 19449 5414 19495 5466
rect 19495 5414 19505 5466
rect 19529 5414 19559 5466
rect 19559 5414 19585 5466
rect 19289 5412 19345 5414
rect 19369 5412 19425 5414
rect 19449 5412 19505 5414
rect 19529 5412 19585 5414
rect 19289 4378 19345 4380
rect 19369 4378 19425 4380
rect 19449 4378 19505 4380
rect 19529 4378 19585 4380
rect 19289 4326 19315 4378
rect 19315 4326 19345 4378
rect 19369 4326 19379 4378
rect 19379 4326 19425 4378
rect 19449 4326 19495 4378
rect 19495 4326 19505 4378
rect 19529 4326 19559 4378
rect 19559 4326 19585 4378
rect 19289 4324 19345 4326
rect 19369 4324 19425 4326
rect 19449 4324 19505 4326
rect 19529 4324 19585 4326
rect 19289 3290 19345 3292
rect 19369 3290 19425 3292
rect 19449 3290 19505 3292
rect 19529 3290 19585 3292
rect 19289 3238 19315 3290
rect 19315 3238 19345 3290
rect 19369 3238 19379 3290
rect 19379 3238 19425 3290
rect 19449 3238 19495 3290
rect 19495 3238 19505 3290
rect 19529 3238 19559 3290
rect 19559 3238 19585 3290
rect 19289 3236 19345 3238
rect 19369 3236 19425 3238
rect 19449 3236 19505 3238
rect 19529 3236 19585 3238
rect 19890 4664 19946 4720
rect 19289 2202 19345 2204
rect 19369 2202 19425 2204
rect 19449 2202 19505 2204
rect 19529 2202 19585 2204
rect 19289 2150 19315 2202
rect 19315 2150 19345 2202
rect 19369 2150 19379 2202
rect 19379 2150 19425 2202
rect 19449 2150 19495 2202
rect 19495 2150 19505 2202
rect 19529 2150 19559 2202
rect 19559 2150 19585 2202
rect 19289 2148 19345 2150
rect 19369 2148 19425 2150
rect 19449 2148 19505 2150
rect 19529 2148 19585 2150
rect 21638 6996 21694 7032
rect 21638 6976 21640 6996
rect 21640 6976 21692 6996
rect 21692 6976 21694 6996
rect 20166 5480 20222 5536
rect 19982 1536 20038 1592
<< metal3 >>
rect 0 21448 480 21480
rect 0 21392 110 21448
rect 166 21392 480 21448
rect 0 21360 480 21392
rect 21520 20952 22000 21072
rect 16389 20498 16455 20501
rect 21590 20498 21650 20952
rect 16389 20496 21650 20498
rect 16389 20440 16394 20496
rect 16450 20440 21650 20496
rect 16389 20438 21650 20440
rect 16389 20435 16455 20438
rect 0 20272 480 20392
rect 62 19818 122 20272
rect 1301 19818 1367 19821
rect 62 19816 1367 19818
rect 62 19760 1306 19816
rect 1362 19760 1367 19816
rect 62 19758 1367 19760
rect 1301 19755 1367 19758
rect 4610 19616 4930 19617
rect 4610 19552 4618 19616
rect 4682 19552 4698 19616
rect 4762 19552 4778 19616
rect 4842 19552 4858 19616
rect 4922 19552 4930 19616
rect 4610 19551 4930 19552
rect 11944 19616 12264 19617
rect 11944 19552 11952 19616
rect 12016 19552 12032 19616
rect 12096 19552 12112 19616
rect 12176 19552 12192 19616
rect 12256 19552 12264 19616
rect 11944 19551 12264 19552
rect 19277 19616 19597 19617
rect 19277 19552 19285 19616
rect 19349 19552 19365 19616
rect 19429 19552 19445 19616
rect 19509 19552 19525 19616
rect 19589 19552 19597 19616
rect 19277 19551 19597 19552
rect 0 19184 480 19304
rect 3417 19274 3483 19277
rect 4153 19274 4219 19277
rect 3417 19272 4219 19274
rect 3417 19216 3422 19272
rect 3478 19216 4158 19272
rect 4214 19216 4219 19272
rect 3417 19214 4219 19216
rect 3417 19211 3483 19214
rect 4153 19211 4219 19214
rect 62 18730 122 19184
rect 8277 19072 8597 19073
rect 8277 19008 8285 19072
rect 8349 19008 8365 19072
rect 8429 19008 8445 19072
rect 8509 19008 8525 19072
rect 8589 19008 8597 19072
rect 8277 19007 8597 19008
rect 15610 19072 15930 19073
rect 15610 19008 15618 19072
rect 15682 19008 15698 19072
rect 15762 19008 15778 19072
rect 15842 19008 15858 19072
rect 15922 19008 15930 19072
rect 15610 19007 15930 19008
rect 21520 18912 22000 19032
rect 1577 18730 1643 18733
rect 62 18728 1643 18730
rect 62 18672 1582 18728
rect 1638 18672 1643 18728
rect 62 18670 1643 18672
rect 1577 18667 1643 18670
rect 4610 18528 4930 18529
rect 4610 18464 4618 18528
rect 4682 18464 4698 18528
rect 4762 18464 4778 18528
rect 4842 18464 4858 18528
rect 4922 18464 4930 18528
rect 4610 18463 4930 18464
rect 11944 18528 12264 18529
rect 11944 18464 11952 18528
rect 12016 18464 12032 18528
rect 12096 18464 12112 18528
rect 12176 18464 12192 18528
rect 12256 18464 12264 18528
rect 11944 18463 12264 18464
rect 19277 18528 19597 18529
rect 19277 18464 19285 18528
rect 19349 18464 19365 18528
rect 19429 18464 19445 18528
rect 19509 18464 19525 18528
rect 19589 18464 19597 18528
rect 19277 18463 19597 18464
rect 19793 18458 19859 18461
rect 21590 18458 21650 18912
rect 19793 18456 21650 18458
rect 19793 18400 19798 18456
rect 19854 18400 21650 18456
rect 19793 18398 21650 18400
rect 19793 18395 19859 18398
rect 0 18096 480 18216
rect 62 17642 122 18096
rect 8277 17984 8597 17985
rect 8277 17920 8285 17984
rect 8349 17920 8365 17984
rect 8429 17920 8445 17984
rect 8509 17920 8525 17984
rect 8589 17920 8597 17984
rect 8277 17919 8597 17920
rect 15610 17984 15930 17985
rect 15610 17920 15618 17984
rect 15682 17920 15698 17984
rect 15762 17920 15778 17984
rect 15842 17920 15858 17984
rect 15922 17920 15930 17984
rect 15610 17919 15930 17920
rect 7833 17778 7899 17781
rect 14181 17778 14247 17781
rect 7833 17776 14247 17778
rect 7833 17720 7838 17776
rect 7894 17720 14186 17776
rect 14242 17720 14247 17776
rect 7833 17718 14247 17720
rect 7833 17715 7899 17718
rect 14181 17715 14247 17718
rect 1577 17642 1643 17645
rect 62 17640 1643 17642
rect 62 17584 1582 17640
rect 1638 17584 1643 17640
rect 62 17582 1643 17584
rect 1577 17579 1643 17582
rect 4610 17440 4930 17441
rect 4610 17376 4618 17440
rect 4682 17376 4698 17440
rect 4762 17376 4778 17440
rect 4842 17376 4858 17440
rect 4922 17376 4930 17440
rect 4610 17375 4930 17376
rect 11944 17440 12264 17441
rect 11944 17376 11952 17440
rect 12016 17376 12032 17440
rect 12096 17376 12112 17440
rect 12176 17376 12192 17440
rect 12256 17376 12264 17440
rect 11944 17375 12264 17376
rect 19277 17440 19597 17441
rect 19277 17376 19285 17440
rect 19349 17376 19365 17440
rect 19429 17376 19445 17440
rect 19509 17376 19525 17440
rect 19589 17376 19597 17440
rect 19277 17375 19597 17376
rect 2773 17234 2839 17237
rect 9305 17234 9371 17237
rect 2773 17232 9371 17234
rect 2773 17176 2778 17232
rect 2834 17176 9310 17232
rect 9366 17176 9371 17232
rect 2773 17174 9371 17176
rect 2773 17171 2839 17174
rect 9305 17171 9371 17174
rect 0 17008 480 17128
rect 62 16554 122 17008
rect 10409 16962 10475 16965
rect 10542 16962 10548 16964
rect 10409 16960 10548 16962
rect 10409 16904 10414 16960
rect 10470 16904 10548 16960
rect 10409 16902 10548 16904
rect 10409 16899 10475 16902
rect 10542 16900 10548 16902
rect 10612 16900 10618 16964
rect 8277 16896 8597 16897
rect 8277 16832 8285 16896
rect 8349 16832 8365 16896
rect 8429 16832 8445 16896
rect 8509 16832 8525 16896
rect 8589 16832 8597 16896
rect 8277 16831 8597 16832
rect 15610 16896 15930 16897
rect 15610 16832 15618 16896
rect 15682 16832 15698 16896
rect 15762 16832 15778 16896
rect 15842 16832 15858 16896
rect 15922 16832 15930 16896
rect 21520 16872 22000 16992
rect 15610 16831 15930 16832
rect 197 16690 263 16693
rect 5942 16690 5948 16692
rect 197 16688 5948 16690
rect 197 16632 202 16688
rect 258 16632 5948 16688
rect 197 16630 5948 16632
rect 197 16627 263 16630
rect 5942 16628 5948 16630
rect 6012 16690 6018 16692
rect 14549 16690 14615 16693
rect 6012 16688 14615 16690
rect 6012 16632 14554 16688
rect 14610 16632 14615 16688
rect 6012 16630 14615 16632
rect 6012 16628 6018 16630
rect 14549 16627 14615 16630
rect 4245 16554 4311 16557
rect 62 16552 4311 16554
rect 62 16496 4250 16552
rect 4306 16496 4311 16552
rect 62 16494 4311 16496
rect 4245 16491 4311 16494
rect 4981 16554 5047 16557
rect 8109 16554 8175 16557
rect 4981 16552 8175 16554
rect 4981 16496 4986 16552
rect 5042 16496 8114 16552
rect 8170 16496 8175 16552
rect 4981 16494 8175 16496
rect 4981 16491 5047 16494
rect 8109 16491 8175 16494
rect 9673 16554 9739 16557
rect 14089 16554 14155 16557
rect 9673 16552 14155 16554
rect 9673 16496 9678 16552
rect 9734 16496 14094 16552
rect 14150 16496 14155 16552
rect 9673 16494 14155 16496
rect 9673 16491 9739 16494
rect 14089 16491 14155 16494
rect 19609 16554 19675 16557
rect 21590 16554 21650 16872
rect 19609 16552 21650 16554
rect 19609 16496 19614 16552
rect 19670 16496 21650 16552
rect 19609 16494 21650 16496
rect 19609 16491 19675 16494
rect 4610 16352 4930 16353
rect 4610 16288 4618 16352
rect 4682 16288 4698 16352
rect 4762 16288 4778 16352
rect 4842 16288 4858 16352
rect 4922 16288 4930 16352
rect 4610 16287 4930 16288
rect 11944 16352 12264 16353
rect 11944 16288 11952 16352
rect 12016 16288 12032 16352
rect 12096 16288 12112 16352
rect 12176 16288 12192 16352
rect 12256 16288 12264 16352
rect 11944 16287 12264 16288
rect 19277 16352 19597 16353
rect 19277 16288 19285 16352
rect 19349 16288 19365 16352
rect 19429 16288 19445 16352
rect 19509 16288 19525 16352
rect 19589 16288 19597 16352
rect 19277 16287 19597 16288
rect 14733 16146 14799 16149
rect 17953 16146 18019 16149
rect 14733 16144 18019 16146
rect 14733 16088 14738 16144
rect 14794 16088 17958 16144
rect 18014 16088 18019 16144
rect 14733 16086 18019 16088
rect 14733 16083 14799 16086
rect 17953 16083 18019 16086
rect 0 16008 480 16040
rect 0 15952 110 16008
rect 166 15952 480 16008
rect 0 15920 480 15952
rect 9765 15874 9831 15877
rect 13486 15874 13492 15876
rect 9765 15872 13492 15874
rect 9765 15816 9770 15872
rect 9826 15816 13492 15872
rect 9765 15814 13492 15816
rect 9765 15811 9831 15814
rect 13486 15812 13492 15814
rect 13556 15874 13562 15876
rect 14273 15874 14339 15877
rect 13556 15872 14339 15874
rect 13556 15816 14278 15872
rect 14334 15816 14339 15872
rect 13556 15814 14339 15816
rect 13556 15812 13562 15814
rect 14273 15811 14339 15814
rect 8277 15808 8597 15809
rect 8277 15744 8285 15808
rect 8349 15744 8365 15808
rect 8429 15744 8445 15808
rect 8509 15744 8525 15808
rect 8589 15744 8597 15808
rect 8277 15743 8597 15744
rect 15610 15808 15930 15809
rect 15610 15744 15618 15808
rect 15682 15744 15698 15808
rect 15762 15744 15778 15808
rect 15842 15744 15858 15808
rect 15922 15744 15930 15808
rect 15610 15743 15930 15744
rect 6126 15268 6132 15332
rect 6196 15330 6202 15332
rect 9489 15330 9555 15333
rect 6196 15328 9555 15330
rect 6196 15272 9494 15328
rect 9550 15272 9555 15328
rect 6196 15270 9555 15272
rect 6196 15268 6202 15270
rect 9489 15267 9555 15270
rect 4610 15264 4930 15265
rect 4610 15200 4618 15264
rect 4682 15200 4698 15264
rect 4762 15200 4778 15264
rect 4842 15200 4858 15264
rect 4922 15200 4930 15264
rect 4610 15199 4930 15200
rect 11944 15264 12264 15265
rect 11944 15200 11952 15264
rect 12016 15200 12032 15264
rect 12096 15200 12112 15264
rect 12176 15200 12192 15264
rect 12256 15200 12264 15264
rect 11944 15199 12264 15200
rect 19277 15264 19597 15265
rect 19277 15200 19285 15264
rect 19349 15200 19365 15264
rect 19429 15200 19445 15264
rect 19509 15200 19525 15264
rect 19589 15200 19597 15264
rect 19277 15199 19597 15200
rect 2037 15058 2103 15061
rect 9029 15058 9095 15061
rect 2037 15056 9095 15058
rect 2037 15000 2042 15056
rect 2098 15000 9034 15056
rect 9090 15000 9095 15056
rect 2037 14998 9095 15000
rect 2037 14995 2103 14998
rect 9029 14995 9095 14998
rect 11145 15058 11211 15061
rect 17769 15058 17835 15061
rect 11145 15056 17835 15058
rect 11145 15000 11150 15056
rect 11206 15000 17774 15056
rect 17830 15000 17835 15056
rect 11145 14998 17835 15000
rect 11145 14995 11211 14998
rect 17769 14995 17835 14998
rect 20161 15058 20227 15061
rect 21520 15058 22000 15088
rect 20161 15056 22000 15058
rect 20161 15000 20166 15056
rect 20222 15000 22000 15056
rect 20161 14998 22000 15000
rect 20161 14995 20227 14998
rect 21520 14968 22000 14998
rect 0 14920 480 14952
rect 0 14864 110 14920
rect 166 14864 480 14920
rect 0 14832 480 14864
rect 15285 14922 15351 14925
rect 17585 14922 17651 14925
rect 15285 14920 17651 14922
rect 15285 14864 15290 14920
rect 15346 14864 17590 14920
rect 17646 14864 17651 14920
rect 15285 14862 17651 14864
rect 15285 14859 15351 14862
rect 17585 14859 17651 14862
rect 8277 14720 8597 14721
rect 8277 14656 8285 14720
rect 8349 14656 8365 14720
rect 8429 14656 8445 14720
rect 8509 14656 8525 14720
rect 8589 14656 8597 14720
rect 8277 14655 8597 14656
rect 15610 14720 15930 14721
rect 15610 14656 15618 14720
rect 15682 14656 15698 14720
rect 15762 14656 15778 14720
rect 15842 14656 15858 14720
rect 15922 14656 15930 14720
rect 15610 14655 15930 14656
rect 11513 14514 11579 14517
rect 13077 14514 13143 14517
rect 18413 14514 18479 14517
rect 11513 14512 18479 14514
rect 11513 14456 11518 14512
rect 11574 14456 13082 14512
rect 13138 14456 18418 14512
rect 18474 14456 18479 14512
rect 11513 14454 18479 14456
rect 11513 14451 11579 14454
rect 13077 14451 13143 14454
rect 18413 14451 18479 14454
rect 2497 14378 2563 14381
rect 15929 14378 15995 14381
rect 2497 14376 15995 14378
rect 2497 14320 2502 14376
rect 2558 14320 15934 14376
rect 15990 14320 15995 14376
rect 2497 14318 15995 14320
rect 2497 14315 2563 14318
rect 15929 14315 15995 14318
rect 13486 14180 13492 14244
rect 13556 14242 13562 14244
rect 13721 14242 13787 14245
rect 13556 14240 13787 14242
rect 13556 14184 13726 14240
rect 13782 14184 13787 14240
rect 13556 14182 13787 14184
rect 13556 14180 13562 14182
rect 13721 14179 13787 14182
rect 4610 14176 4930 14177
rect 4610 14112 4618 14176
rect 4682 14112 4698 14176
rect 4762 14112 4778 14176
rect 4842 14112 4858 14176
rect 4922 14112 4930 14176
rect 4610 14111 4930 14112
rect 11944 14176 12264 14177
rect 11944 14112 11952 14176
rect 12016 14112 12032 14176
rect 12096 14112 12112 14176
rect 12176 14112 12192 14176
rect 12256 14112 12264 14176
rect 11944 14111 12264 14112
rect 19277 14176 19597 14177
rect 19277 14112 19285 14176
rect 19349 14112 19365 14176
rect 19429 14112 19445 14176
rect 19509 14112 19525 14176
rect 19589 14112 19597 14176
rect 19277 14111 19597 14112
rect 6637 14106 6703 14109
rect 9622 14106 9628 14108
rect 6637 14104 9628 14106
rect 6637 14048 6642 14104
rect 6698 14048 9628 14104
rect 6637 14046 9628 14048
rect 6637 14043 6703 14046
rect 9622 14044 9628 14046
rect 9692 14106 9698 14108
rect 11605 14106 11671 14109
rect 9692 14104 11671 14106
rect 9692 14048 11610 14104
rect 11666 14048 11671 14104
rect 9692 14046 11671 14048
rect 9692 14044 9698 14046
rect 11605 14043 11671 14046
rect 5625 13970 5691 13973
rect 9070 13970 9076 13972
rect 5625 13968 9076 13970
rect 5625 13912 5630 13968
rect 5686 13912 9076 13968
rect 5625 13910 9076 13912
rect 5625 13907 5691 13910
rect 9070 13908 9076 13910
rect 9140 13908 9146 13972
rect 0 13836 480 13864
rect 0 13772 60 13836
rect 124 13772 480 13836
rect 0 13744 480 13772
rect 6637 13834 6703 13837
rect 8109 13834 8175 13837
rect 6637 13832 8175 13834
rect 6637 13776 6642 13832
rect 6698 13776 8114 13832
rect 8170 13776 8175 13832
rect 6637 13774 8175 13776
rect 6637 13771 6703 13774
rect 8109 13771 8175 13774
rect 16665 13832 16731 13837
rect 16665 13776 16670 13832
rect 16726 13776 16731 13832
rect 16665 13771 16731 13776
rect 9029 13698 9095 13701
rect 9765 13698 9831 13701
rect 15193 13698 15259 13701
rect 9029 13696 15259 13698
rect 9029 13640 9034 13696
rect 9090 13640 9770 13696
rect 9826 13640 15198 13696
rect 15254 13640 15259 13696
rect 9029 13638 15259 13640
rect 9029 13635 9095 13638
rect 9765 13635 9831 13638
rect 15193 13635 15259 13638
rect 16021 13698 16087 13701
rect 16668 13698 16728 13771
rect 16021 13696 16728 13698
rect 16021 13640 16026 13696
rect 16082 13640 16728 13696
rect 16021 13638 16728 13640
rect 16021 13635 16087 13638
rect 8277 13632 8597 13633
rect 8277 13568 8285 13632
rect 8349 13568 8365 13632
rect 8429 13568 8445 13632
rect 8509 13568 8525 13632
rect 8589 13568 8597 13632
rect 8277 13567 8597 13568
rect 15610 13632 15930 13633
rect 15610 13568 15618 13632
rect 15682 13568 15698 13632
rect 15762 13568 15778 13632
rect 15842 13568 15858 13632
rect 15922 13568 15930 13632
rect 15610 13567 15930 13568
rect 9765 13562 9831 13565
rect 13445 13562 13511 13565
rect 9765 13560 13511 13562
rect 9765 13504 9770 13560
rect 9826 13504 13450 13560
rect 13506 13504 13511 13560
rect 9765 13502 13511 13504
rect 9765 13499 9831 13502
rect 13445 13499 13511 13502
rect 14590 13500 14596 13564
rect 14660 13562 14666 13564
rect 14733 13562 14799 13565
rect 14660 13560 14799 13562
rect 14660 13504 14738 13560
rect 14794 13504 14799 13560
rect 14660 13502 14799 13504
rect 14660 13500 14666 13502
rect 14733 13499 14799 13502
rect 2221 13426 2287 13429
rect 3969 13426 4035 13429
rect 11329 13426 11395 13429
rect 13261 13426 13327 13429
rect 2221 13424 13327 13426
rect 2221 13368 2226 13424
rect 2282 13368 3974 13424
rect 4030 13368 11334 13424
rect 11390 13368 13266 13424
rect 13322 13368 13327 13424
rect 2221 13366 13327 13368
rect 2221 13363 2287 13366
rect 3969 13363 4035 13366
rect 11329 13363 11395 13366
rect 13261 13363 13327 13366
rect 15193 13426 15259 13429
rect 16849 13426 16915 13429
rect 15193 13424 16915 13426
rect 15193 13368 15198 13424
rect 15254 13368 16854 13424
rect 16910 13368 16915 13424
rect 15193 13366 16915 13368
rect 15193 13363 15259 13366
rect 16849 13363 16915 13366
rect 18413 13426 18479 13429
rect 18413 13424 21650 13426
rect 18413 13368 18418 13424
rect 18474 13368 21650 13424
rect 18413 13366 21650 13368
rect 18413 13363 18479 13366
rect 11053 13290 11119 13293
rect 16573 13290 16639 13293
rect 11053 13288 16639 13290
rect 11053 13232 11058 13288
rect 11114 13232 16578 13288
rect 16634 13232 16639 13288
rect 11053 13230 16639 13232
rect 11053 13227 11119 13230
rect 16573 13227 16639 13230
rect 4610 13088 4930 13089
rect 4610 13024 4618 13088
rect 4682 13024 4698 13088
rect 4762 13024 4778 13088
rect 4842 13024 4858 13088
rect 4922 13024 4930 13088
rect 4610 13023 4930 13024
rect 11944 13088 12264 13089
rect 11944 13024 11952 13088
rect 12016 13024 12032 13088
rect 12096 13024 12112 13088
rect 12176 13024 12192 13088
rect 12256 13024 12264 13088
rect 11944 13023 12264 13024
rect 19277 13088 19597 13089
rect 19277 13024 19285 13088
rect 19349 13024 19365 13088
rect 19429 13024 19445 13088
rect 19509 13024 19525 13088
rect 19589 13024 19597 13088
rect 21590 13048 21650 13366
rect 19277 13023 19597 13024
rect 21520 12928 22000 13048
rect 0 12656 480 12776
rect 62 12474 122 12656
rect 8277 12544 8597 12545
rect 8277 12480 8285 12544
rect 8349 12480 8365 12544
rect 8429 12480 8445 12544
rect 8509 12480 8525 12544
rect 8589 12480 8597 12544
rect 8277 12479 8597 12480
rect 15610 12544 15930 12545
rect 15610 12480 15618 12544
rect 15682 12480 15698 12544
rect 15762 12480 15778 12544
rect 15842 12480 15858 12544
rect 15922 12480 15930 12544
rect 15610 12479 15930 12480
rect 7925 12474 7991 12477
rect 62 12472 7991 12474
rect 62 12416 7930 12472
rect 7986 12416 7991 12472
rect 62 12414 7991 12416
rect 7925 12411 7991 12414
rect 4610 12000 4930 12001
rect 4610 11936 4618 12000
rect 4682 11936 4698 12000
rect 4762 11936 4778 12000
rect 4842 11936 4858 12000
rect 4922 11936 4930 12000
rect 4610 11935 4930 11936
rect 11944 12000 12264 12001
rect 11944 11936 11952 12000
rect 12016 11936 12032 12000
rect 12096 11936 12112 12000
rect 12176 11936 12192 12000
rect 12256 11936 12264 12000
rect 11944 11935 12264 11936
rect 19277 12000 19597 12001
rect 19277 11936 19285 12000
rect 19349 11936 19365 12000
rect 19429 11936 19445 12000
rect 19509 11936 19525 12000
rect 19589 11936 19597 12000
rect 19277 11935 19597 11936
rect 5942 11868 5948 11932
rect 6012 11930 6018 11932
rect 6085 11930 6151 11933
rect 6012 11928 6151 11930
rect 6012 11872 6090 11928
rect 6146 11872 6151 11928
rect 6012 11870 6151 11872
rect 6012 11868 6018 11870
rect 6085 11867 6151 11870
rect 0 11656 480 11688
rect 0 11600 110 11656
rect 166 11600 480 11656
rect 0 11568 480 11600
rect 5533 11658 5599 11661
rect 12709 11658 12775 11661
rect 5533 11656 12775 11658
rect 5533 11600 5538 11656
rect 5594 11600 12714 11656
rect 12770 11600 12775 11656
rect 5533 11598 12775 11600
rect 5533 11595 5599 11598
rect 12709 11595 12775 11598
rect 2129 11522 2195 11525
rect 3877 11522 3943 11525
rect 4429 11522 4495 11525
rect 6453 11522 6519 11525
rect 2129 11520 6519 11522
rect 2129 11464 2134 11520
rect 2190 11464 3882 11520
rect 3938 11464 4434 11520
rect 4490 11464 6458 11520
rect 6514 11464 6519 11520
rect 2129 11462 6519 11464
rect 2129 11459 2195 11462
rect 3877 11459 3943 11462
rect 4429 11459 4495 11462
rect 6453 11459 6519 11462
rect 9622 11460 9628 11524
rect 9692 11522 9698 11524
rect 11145 11522 11211 11525
rect 9692 11520 11211 11522
rect 9692 11464 11150 11520
rect 11206 11464 11211 11520
rect 9692 11462 11211 11464
rect 9692 11460 9698 11462
rect 11145 11459 11211 11462
rect 8277 11456 8597 11457
rect 8277 11392 8285 11456
rect 8349 11392 8365 11456
rect 8429 11392 8445 11456
rect 8509 11392 8525 11456
rect 8589 11392 8597 11456
rect 8277 11391 8597 11392
rect 15610 11456 15930 11457
rect 15610 11392 15618 11456
rect 15682 11392 15698 11456
rect 15762 11392 15778 11456
rect 15842 11392 15858 11456
rect 15922 11392 15930 11456
rect 15610 11391 15930 11392
rect 5349 11250 5415 11253
rect 13629 11250 13695 11253
rect 5349 11248 13695 11250
rect 5349 11192 5354 11248
rect 5410 11192 13634 11248
rect 13690 11192 13695 11248
rect 5349 11190 13695 11192
rect 5349 11187 5415 11190
rect 13629 11187 13695 11190
rect 9673 11114 9739 11117
rect 18505 11114 18571 11117
rect 9673 11112 18571 11114
rect 9673 11056 9678 11112
rect 9734 11056 18510 11112
rect 18566 11056 18571 11112
rect 9673 11054 18571 11056
rect 9673 11051 9739 11054
rect 18505 11051 18571 11054
rect 4610 10912 4930 10913
rect 4610 10848 4618 10912
rect 4682 10848 4698 10912
rect 4762 10848 4778 10912
rect 4842 10848 4858 10912
rect 4922 10848 4930 10912
rect 4610 10847 4930 10848
rect 11944 10912 12264 10913
rect 11944 10848 11952 10912
rect 12016 10848 12032 10912
rect 12096 10848 12112 10912
rect 12176 10848 12192 10912
rect 12256 10848 12264 10912
rect 11944 10847 12264 10848
rect 19277 10912 19597 10913
rect 19277 10848 19285 10912
rect 19349 10848 19365 10912
rect 19429 10848 19445 10912
rect 19509 10848 19525 10912
rect 19589 10848 19597 10912
rect 21520 10888 22000 11008
rect 19277 10847 19597 10848
rect 13905 10842 13971 10845
rect 18597 10842 18663 10845
rect 13905 10840 18663 10842
rect 13905 10784 13910 10840
rect 13966 10784 18602 10840
rect 18658 10784 18663 10840
rect 13905 10782 18663 10784
rect 13905 10779 13971 10782
rect 18597 10779 18663 10782
rect 9121 10706 9187 10709
rect 9581 10706 9647 10709
rect 17493 10706 17559 10709
rect 9121 10704 17559 10706
rect 9121 10648 9126 10704
rect 9182 10648 9586 10704
rect 9642 10648 17498 10704
rect 17554 10648 17559 10704
rect 9121 10646 17559 10648
rect 9121 10643 9187 10646
rect 9581 10643 9647 10646
rect 17493 10643 17559 10646
rect 11145 10570 11211 10573
rect 21590 10570 21650 10888
rect 11145 10568 21650 10570
rect 11145 10512 11150 10568
rect 11206 10512 21650 10568
rect 11145 10510 21650 10512
rect 11145 10507 11211 10510
rect 0 10432 480 10464
rect 0 10376 18 10432
rect 74 10376 480 10432
rect 0 10344 480 10376
rect 8277 10368 8597 10369
rect 8277 10304 8285 10368
rect 8349 10304 8365 10368
rect 8429 10304 8445 10368
rect 8509 10304 8525 10368
rect 8589 10304 8597 10368
rect 8277 10303 8597 10304
rect 15610 10368 15930 10369
rect 15610 10304 15618 10368
rect 15682 10304 15698 10368
rect 15762 10304 15778 10368
rect 15842 10304 15858 10368
rect 15922 10304 15930 10368
rect 15610 10303 15930 10304
rect 9029 10026 9095 10029
rect 18781 10026 18847 10029
rect 9029 10024 18847 10026
rect 9029 9968 9034 10024
rect 9090 9968 18786 10024
rect 18842 9968 18847 10024
rect 9029 9966 18847 9968
rect 9029 9963 9095 9966
rect 18781 9963 18847 9966
rect 4610 9824 4930 9825
rect 4610 9760 4618 9824
rect 4682 9760 4698 9824
rect 4762 9760 4778 9824
rect 4842 9760 4858 9824
rect 4922 9760 4930 9824
rect 4610 9759 4930 9760
rect 11944 9824 12264 9825
rect 11944 9760 11952 9824
rect 12016 9760 12032 9824
rect 12096 9760 12112 9824
rect 12176 9760 12192 9824
rect 12256 9760 12264 9824
rect 11944 9759 12264 9760
rect 19277 9824 19597 9825
rect 19277 9760 19285 9824
rect 19349 9760 19365 9824
rect 19429 9760 19445 9824
rect 19509 9760 19525 9824
rect 19589 9760 19597 9824
rect 19277 9759 19597 9760
rect 9857 9618 9923 9621
rect 14089 9618 14155 9621
rect 18137 9618 18203 9621
rect 9857 9616 18203 9618
rect 9857 9560 9862 9616
rect 9918 9560 14094 9616
rect 14150 9560 18142 9616
rect 18198 9560 18203 9616
rect 9857 9558 18203 9560
rect 9857 9555 9923 9558
rect 14089 9555 14155 9558
rect 18137 9555 18203 9558
rect 10542 9420 10548 9484
rect 10612 9482 10618 9484
rect 10961 9482 11027 9485
rect 17769 9482 17835 9485
rect 10612 9480 11027 9482
rect 10612 9424 10966 9480
rect 11022 9424 11027 9480
rect 10612 9422 11027 9424
rect 10612 9420 10618 9422
rect 10961 9419 11027 9422
rect 13770 9480 17835 9482
rect 13770 9424 17774 9480
rect 17830 9424 17835 9480
rect 13770 9422 17835 9424
rect 0 9256 480 9376
rect 8661 9346 8727 9349
rect 13770 9346 13830 9422
rect 17769 9419 17835 9422
rect 8661 9344 13830 9346
rect 8661 9288 8666 9344
rect 8722 9288 13830 9344
rect 8661 9286 13830 9288
rect 8661 9283 8727 9286
rect 8277 9280 8597 9281
rect 62 8802 122 9256
rect 8277 9216 8285 9280
rect 8349 9216 8365 9280
rect 8429 9216 8445 9280
rect 8509 9216 8525 9280
rect 8589 9216 8597 9280
rect 8277 9215 8597 9216
rect 15610 9280 15930 9281
rect 15610 9216 15618 9280
rect 15682 9216 15698 9280
rect 15762 9216 15778 9280
rect 15842 9216 15858 9280
rect 15922 9216 15930 9280
rect 15610 9215 15930 9216
rect 10317 9074 10383 9077
rect 17585 9074 17651 9077
rect 10317 9072 17651 9074
rect 10317 9016 10322 9072
rect 10378 9016 17590 9072
rect 17646 9016 17651 9072
rect 10317 9014 17651 9016
rect 10317 9011 10383 9014
rect 17585 9011 17651 9014
rect 14089 8938 14155 8941
rect 20069 8938 20135 8941
rect 21520 8938 22000 8968
rect 14089 8936 20135 8938
rect 14089 8880 14094 8936
rect 14150 8880 20074 8936
rect 20130 8880 20135 8936
rect 14089 8878 20135 8880
rect 21460 8936 22000 8938
rect 21460 8880 21546 8936
rect 21602 8880 22000 8936
rect 21460 8878 22000 8880
rect 14089 8875 14155 8878
rect 20069 8875 20135 8878
rect 21520 8848 22000 8878
rect 4245 8802 4311 8805
rect 62 8800 4311 8802
rect 62 8744 4250 8800
rect 4306 8744 4311 8800
rect 62 8742 4311 8744
rect 4245 8739 4311 8742
rect 4610 8736 4930 8737
rect 4610 8672 4618 8736
rect 4682 8672 4698 8736
rect 4762 8672 4778 8736
rect 4842 8672 4858 8736
rect 4922 8672 4930 8736
rect 4610 8671 4930 8672
rect 11944 8736 12264 8737
rect 11944 8672 11952 8736
rect 12016 8672 12032 8736
rect 12096 8672 12112 8736
rect 12176 8672 12192 8736
rect 12256 8672 12264 8736
rect 11944 8671 12264 8672
rect 19277 8736 19597 8737
rect 19277 8672 19285 8736
rect 19349 8672 19365 8736
rect 19429 8672 19445 8736
rect 19509 8672 19525 8736
rect 19589 8672 19597 8736
rect 19277 8671 19597 8672
rect 1945 8666 2011 8669
rect 62 8664 2011 8666
rect 62 8608 1950 8664
rect 2006 8608 2011 8664
rect 62 8606 2011 8608
rect 62 8288 122 8606
rect 1945 8603 2011 8606
rect 8661 8666 8727 8669
rect 9070 8666 9076 8668
rect 8661 8664 9076 8666
rect 8661 8608 8666 8664
rect 8722 8608 9076 8664
rect 8661 8606 9076 8608
rect 8661 8603 8727 8606
rect 9070 8604 9076 8606
rect 9140 8604 9146 8668
rect 5073 8530 5139 8533
rect 18229 8530 18295 8533
rect 5073 8528 18295 8530
rect 5073 8472 5078 8528
rect 5134 8472 18234 8528
rect 18290 8472 18295 8528
rect 5073 8470 18295 8472
rect 5073 8467 5139 8470
rect 18229 8467 18295 8470
rect 0 8168 480 8288
rect 8277 8192 8597 8193
rect 8277 8128 8285 8192
rect 8349 8128 8365 8192
rect 8429 8128 8445 8192
rect 8509 8128 8525 8192
rect 8589 8128 8597 8192
rect 8277 8127 8597 8128
rect 15610 8192 15930 8193
rect 15610 8128 15618 8192
rect 15682 8128 15698 8192
rect 15762 8128 15778 8192
rect 15842 8128 15858 8192
rect 15922 8128 15930 8192
rect 15610 8127 15930 8128
rect 9581 8122 9647 8125
rect 15469 8122 15535 8125
rect 9581 8120 15535 8122
rect 9581 8064 9586 8120
rect 9642 8064 15474 8120
rect 15530 8064 15535 8120
rect 9581 8062 15535 8064
rect 9581 8059 9647 8062
rect 15469 8059 15535 8062
rect 14917 7850 14983 7853
rect 19701 7850 19767 7853
rect 14917 7848 19767 7850
rect 14917 7792 14922 7848
rect 14978 7792 19706 7848
rect 19762 7792 19767 7848
rect 14917 7790 19767 7792
rect 14917 7787 14983 7790
rect 19701 7787 19767 7790
rect 2221 7714 2287 7717
rect 62 7712 2287 7714
rect 62 7656 2226 7712
rect 2282 7656 2287 7712
rect 62 7654 2287 7656
rect 62 7200 122 7654
rect 2221 7651 2287 7654
rect 4610 7648 4930 7649
rect 4610 7584 4618 7648
rect 4682 7584 4698 7648
rect 4762 7584 4778 7648
rect 4842 7584 4858 7648
rect 4922 7584 4930 7648
rect 4610 7583 4930 7584
rect 11944 7648 12264 7649
rect 11944 7584 11952 7648
rect 12016 7584 12032 7648
rect 12096 7584 12112 7648
rect 12176 7584 12192 7648
rect 12256 7584 12264 7648
rect 11944 7583 12264 7584
rect 19277 7648 19597 7649
rect 19277 7584 19285 7648
rect 19349 7584 19365 7648
rect 19429 7584 19445 7648
rect 19509 7584 19525 7648
rect 19589 7584 19597 7648
rect 19277 7583 19597 7584
rect 10225 7442 10291 7445
rect 16389 7442 16455 7445
rect 10225 7440 16455 7442
rect 10225 7384 10230 7440
rect 10286 7384 16394 7440
rect 16450 7384 16455 7440
rect 10225 7382 16455 7384
rect 10225 7379 10291 7382
rect 16389 7379 16455 7382
rect 7465 7306 7531 7309
rect 17309 7306 17375 7309
rect 7465 7304 17375 7306
rect 7465 7248 7470 7304
rect 7526 7248 17314 7304
rect 17370 7248 17375 7304
rect 7465 7246 17375 7248
rect 7465 7243 7531 7246
rect 17309 7243 17375 7246
rect 0 7080 480 7200
rect 8661 7170 8727 7173
rect 15193 7170 15259 7173
rect 8661 7168 15259 7170
rect 8661 7112 8666 7168
rect 8722 7112 15198 7168
rect 15254 7112 15259 7168
rect 8661 7110 15259 7112
rect 8661 7107 8727 7110
rect 15193 7107 15259 7110
rect 8277 7104 8597 7105
rect 8277 7040 8285 7104
rect 8349 7040 8365 7104
rect 8429 7040 8445 7104
rect 8509 7040 8525 7104
rect 8589 7040 8597 7104
rect 8277 7039 8597 7040
rect 15610 7104 15930 7105
rect 15610 7040 15618 7104
rect 15682 7040 15698 7104
rect 15762 7040 15778 7104
rect 15842 7040 15858 7104
rect 15922 7040 15930 7104
rect 15610 7039 15930 7040
rect 21520 7032 22000 7064
rect 21520 6976 21638 7032
rect 21694 6976 22000 7032
rect 21520 6944 22000 6976
rect 8477 6762 8543 6765
rect 17861 6762 17927 6765
rect 8477 6760 17927 6762
rect 8477 6704 8482 6760
rect 8538 6704 17866 6760
rect 17922 6704 17927 6760
rect 8477 6702 17927 6704
rect 8477 6699 8543 6702
rect 17861 6699 17927 6702
rect 1301 6626 1367 6629
rect 62 6624 1367 6626
rect 62 6568 1306 6624
rect 1362 6568 1367 6624
rect 62 6566 1367 6568
rect 62 6112 122 6566
rect 1301 6563 1367 6566
rect 4610 6560 4930 6561
rect 4610 6496 4618 6560
rect 4682 6496 4698 6560
rect 4762 6496 4778 6560
rect 4842 6496 4858 6560
rect 4922 6496 4930 6560
rect 4610 6495 4930 6496
rect 11944 6560 12264 6561
rect 11944 6496 11952 6560
rect 12016 6496 12032 6560
rect 12096 6496 12112 6560
rect 12176 6496 12192 6560
rect 12256 6496 12264 6560
rect 11944 6495 12264 6496
rect 19277 6560 19597 6561
rect 19277 6496 19285 6560
rect 19349 6496 19365 6560
rect 19429 6496 19445 6560
rect 19509 6496 19525 6560
rect 19589 6496 19597 6560
rect 19277 6495 19597 6496
rect 0 5992 480 6112
rect 8277 6016 8597 6017
rect 8277 5952 8285 6016
rect 8349 5952 8365 6016
rect 8429 5952 8445 6016
rect 8509 5952 8525 6016
rect 8589 5952 8597 6016
rect 8277 5951 8597 5952
rect 15610 6016 15930 6017
rect 15610 5952 15618 6016
rect 15682 5952 15698 6016
rect 15762 5952 15778 6016
rect 15842 5952 15858 6016
rect 15922 5952 15930 6016
rect 15610 5951 15930 5952
rect 10409 5810 10475 5813
rect 18137 5810 18203 5813
rect 10409 5808 18203 5810
rect 10409 5752 10414 5808
rect 10470 5752 18142 5808
rect 18198 5752 18203 5808
rect 10409 5750 18203 5752
rect 10409 5747 10475 5750
rect 18137 5747 18203 5750
rect 3049 5674 3115 5677
rect 9673 5674 9739 5677
rect 3049 5672 9739 5674
rect 3049 5616 3054 5672
rect 3110 5616 9678 5672
rect 9734 5616 9739 5672
rect 3049 5614 9739 5616
rect 3049 5611 3115 5614
rect 9673 5611 9739 5614
rect 20161 5538 20227 5541
rect 20161 5536 21650 5538
rect 20161 5480 20166 5536
rect 20222 5480 21650 5536
rect 20161 5478 21650 5480
rect 20161 5475 20227 5478
rect 4610 5472 4930 5473
rect 4610 5408 4618 5472
rect 4682 5408 4698 5472
rect 4762 5408 4778 5472
rect 4842 5408 4858 5472
rect 4922 5408 4930 5472
rect 4610 5407 4930 5408
rect 11944 5472 12264 5473
rect 11944 5408 11952 5472
rect 12016 5408 12032 5472
rect 12096 5408 12112 5472
rect 12176 5408 12192 5472
rect 12256 5408 12264 5472
rect 11944 5407 12264 5408
rect 19277 5472 19597 5473
rect 19277 5408 19285 5472
rect 19349 5408 19365 5472
rect 19429 5408 19445 5472
rect 19509 5408 19525 5472
rect 19589 5408 19597 5472
rect 19277 5407 19597 5408
rect 54 5204 60 5268
rect 124 5266 130 5268
rect 6821 5266 6887 5269
rect 10777 5266 10843 5269
rect 18045 5266 18111 5269
rect 18270 5266 18276 5268
rect 124 5264 9690 5266
rect 124 5208 6826 5264
rect 6882 5208 9690 5264
rect 124 5206 9690 5208
rect 124 5204 130 5206
rect 6821 5203 6887 5206
rect 9630 5130 9690 5206
rect 10777 5264 18276 5266
rect 10777 5208 10782 5264
rect 10838 5208 18050 5264
rect 18106 5208 18276 5264
rect 10777 5206 18276 5208
rect 10777 5203 10843 5206
rect 18045 5203 18111 5206
rect 18270 5204 18276 5206
rect 18340 5204 18346 5268
rect 17769 5130 17835 5133
rect 9630 5128 17835 5130
rect 9630 5072 17774 5128
rect 17830 5072 17835 5128
rect 9630 5070 17835 5072
rect 17769 5067 17835 5070
rect 21590 5024 21650 5478
rect 0 4992 480 5024
rect 0 4936 110 4992
rect 166 4936 480 4992
rect 0 4904 480 4936
rect 8277 4928 8597 4929
rect 8277 4864 8285 4928
rect 8349 4864 8365 4928
rect 8429 4864 8445 4928
rect 8509 4864 8525 4928
rect 8589 4864 8597 4928
rect 8277 4863 8597 4864
rect 15610 4928 15930 4929
rect 15610 4864 15618 4928
rect 15682 4864 15698 4928
rect 15762 4864 15778 4928
rect 15842 4864 15858 4928
rect 15922 4864 15930 4928
rect 21520 4904 22000 5024
rect 15610 4863 15930 4864
rect 8937 4858 9003 4861
rect 14181 4858 14247 4861
rect 8937 4856 14247 4858
rect 8937 4800 8942 4856
rect 8998 4800 14186 4856
rect 14242 4800 14247 4856
rect 8937 4798 14247 4800
rect 8937 4795 9003 4798
rect 14181 4795 14247 4798
rect 14273 4722 14339 4725
rect 19885 4722 19951 4725
rect 14273 4720 19951 4722
rect 14273 4664 14278 4720
rect 14334 4664 19890 4720
rect 19946 4664 19951 4720
rect 14273 4662 19951 4664
rect 14273 4659 14339 4662
rect 19885 4659 19951 4662
rect 6453 4586 6519 4589
rect 18505 4586 18571 4589
rect 6453 4584 18571 4586
rect 6453 4528 6458 4584
rect 6514 4528 18510 4584
rect 18566 4528 18571 4584
rect 6453 4526 18571 4528
rect 6453 4523 6519 4526
rect 18505 4523 18571 4526
rect 4610 4384 4930 4385
rect 4610 4320 4618 4384
rect 4682 4320 4698 4384
rect 4762 4320 4778 4384
rect 4842 4320 4858 4384
rect 4922 4320 4930 4384
rect 4610 4319 4930 4320
rect 11944 4384 12264 4385
rect 11944 4320 11952 4384
rect 12016 4320 12032 4384
rect 12096 4320 12112 4384
rect 12176 4320 12192 4384
rect 12256 4320 12264 4384
rect 11944 4319 12264 4320
rect 19277 4384 19597 4385
rect 19277 4320 19285 4384
rect 19349 4320 19365 4384
rect 19429 4320 19445 4384
rect 19509 4320 19525 4384
rect 19589 4320 19597 4384
rect 19277 4319 19597 4320
rect 5165 4178 5231 4181
rect 62 4176 5231 4178
rect 62 4120 5170 4176
rect 5226 4120 5231 4176
rect 62 4118 5231 4120
rect 62 3936 122 4118
rect 5165 4115 5231 4118
rect 6085 4042 6151 4045
rect 12341 4042 12407 4045
rect 18045 4042 18111 4045
rect 6085 4040 12407 4042
rect 6085 3984 6090 4040
rect 6146 3984 12346 4040
rect 12402 3984 12407 4040
rect 6085 3982 12407 3984
rect 6085 3979 6151 3982
rect 12341 3979 12407 3982
rect 13770 4040 18111 4042
rect 13770 3984 18050 4040
rect 18106 3984 18111 4040
rect 13770 3982 18111 3984
rect 0 3816 480 3936
rect 8277 3840 8597 3841
rect 8277 3776 8285 3840
rect 8349 3776 8365 3840
rect 8429 3776 8445 3840
rect 8509 3776 8525 3840
rect 8589 3776 8597 3840
rect 8277 3775 8597 3776
rect 13770 3770 13830 3982
rect 18045 3979 18111 3982
rect 16021 3906 16087 3909
rect 17125 3906 17191 3909
rect 16021 3904 17191 3906
rect 16021 3848 16026 3904
rect 16082 3848 17130 3904
rect 17186 3848 17191 3904
rect 16021 3846 17191 3848
rect 16021 3843 16087 3846
rect 17125 3843 17191 3846
rect 15610 3840 15930 3841
rect 15610 3776 15618 3840
rect 15682 3776 15698 3840
rect 15762 3776 15778 3840
rect 15842 3776 15858 3840
rect 15922 3776 15930 3840
rect 15610 3775 15930 3776
rect 8710 3710 13830 3770
rect 5349 3634 5415 3637
rect 8710 3634 8770 3710
rect 5349 3632 8770 3634
rect 5349 3576 5354 3632
rect 5410 3576 8770 3632
rect 5349 3574 8770 3576
rect 11145 3634 11211 3637
rect 18137 3634 18203 3637
rect 11145 3632 18203 3634
rect 11145 3576 11150 3632
rect 11206 3576 18142 3632
rect 18198 3576 18203 3632
rect 11145 3574 18203 3576
rect 5349 3571 5415 3574
rect 11145 3571 11211 3574
rect 18137 3571 18203 3574
rect 3417 3498 3483 3501
rect 9029 3498 9095 3501
rect 3417 3496 9095 3498
rect 3417 3440 3422 3496
rect 3478 3440 9034 3496
rect 9090 3440 9095 3496
rect 3417 3438 9095 3440
rect 3417 3435 3483 3438
rect 9029 3435 9095 3438
rect 9213 3498 9279 3501
rect 16481 3498 16547 3501
rect 9213 3496 16547 3498
rect 9213 3440 9218 3496
rect 9274 3440 16486 3496
rect 16542 3440 16547 3496
rect 9213 3438 16547 3440
rect 9213 3435 9279 3438
rect 16481 3435 16547 3438
rect 16665 3498 16731 3501
rect 16665 3496 21650 3498
rect 16665 3440 16670 3496
rect 16726 3440 21650 3496
rect 16665 3438 21650 3440
rect 16665 3435 16731 3438
rect 1945 3362 2011 3365
rect 62 3360 2011 3362
rect 62 3304 1950 3360
rect 2006 3304 2011 3360
rect 62 3302 2011 3304
rect 62 2848 122 3302
rect 1945 3299 2011 3302
rect 5165 3362 5231 3365
rect 10041 3362 10107 3365
rect 5165 3360 10107 3362
rect 5165 3304 5170 3360
rect 5226 3304 10046 3360
rect 10102 3304 10107 3360
rect 5165 3302 10107 3304
rect 5165 3299 5231 3302
rect 10041 3299 10107 3302
rect 13077 3362 13143 3365
rect 18597 3362 18663 3365
rect 13077 3360 18663 3362
rect 13077 3304 13082 3360
rect 13138 3304 18602 3360
rect 18658 3304 18663 3360
rect 13077 3302 18663 3304
rect 13077 3299 13143 3302
rect 18597 3299 18663 3302
rect 4610 3296 4930 3297
rect 4610 3232 4618 3296
rect 4682 3232 4698 3296
rect 4762 3232 4778 3296
rect 4842 3232 4858 3296
rect 4922 3232 4930 3296
rect 4610 3231 4930 3232
rect 11944 3296 12264 3297
rect 11944 3232 11952 3296
rect 12016 3232 12032 3296
rect 12096 3232 12112 3296
rect 12176 3232 12192 3296
rect 12256 3232 12264 3296
rect 11944 3231 12264 3232
rect 19277 3296 19597 3297
rect 19277 3232 19285 3296
rect 19349 3232 19365 3296
rect 19429 3232 19445 3296
rect 19509 3232 19525 3296
rect 19589 3232 19597 3296
rect 19277 3231 19597 3232
rect 5073 3226 5139 3229
rect 9121 3226 9187 3229
rect 5073 3224 9187 3226
rect 5073 3168 5078 3224
rect 5134 3168 9126 3224
rect 9182 3168 9187 3224
rect 5073 3166 9187 3168
rect 5073 3163 5139 3166
rect 9121 3163 9187 3166
rect 6269 3090 6335 3093
rect 17033 3090 17099 3093
rect 6269 3088 17099 3090
rect 6269 3032 6274 3088
rect 6330 3032 17038 3088
rect 17094 3032 17099 3088
rect 6269 3030 17099 3032
rect 6269 3027 6335 3030
rect 17033 3027 17099 3030
rect 21590 2984 21650 3438
rect 9949 2954 10015 2957
rect 17769 2954 17835 2957
rect 9949 2952 17835 2954
rect 9949 2896 9954 2952
rect 10010 2896 17774 2952
rect 17830 2896 17835 2952
rect 9949 2894 17835 2896
rect 9949 2891 10015 2894
rect 17769 2891 17835 2894
rect 21520 2864 22000 2984
rect 0 2728 480 2848
rect 8277 2752 8597 2753
rect 8277 2688 8285 2752
rect 8349 2688 8365 2752
rect 8429 2688 8445 2752
rect 8509 2688 8525 2752
rect 8589 2688 8597 2752
rect 8277 2687 8597 2688
rect 15610 2752 15930 2753
rect 15610 2688 15618 2752
rect 15682 2688 15698 2752
rect 15762 2688 15778 2752
rect 15842 2688 15858 2752
rect 15922 2688 15930 2752
rect 15610 2687 15930 2688
rect 3141 2682 3207 2685
rect 7189 2682 7255 2685
rect 3141 2680 7255 2682
rect 3141 2624 3146 2680
rect 3202 2624 7194 2680
rect 7250 2624 7255 2680
rect 3141 2622 7255 2624
rect 3141 2619 3207 2622
rect 7189 2619 7255 2622
rect 18270 2620 18276 2684
rect 18340 2682 18346 2684
rect 18781 2682 18847 2685
rect 18340 2680 18847 2682
rect 18340 2624 18786 2680
rect 18842 2624 18847 2680
rect 18340 2622 18847 2624
rect 18340 2620 18346 2622
rect 18781 2619 18847 2622
rect 6361 2410 6427 2413
rect 18137 2410 18203 2413
rect 6361 2408 18203 2410
rect 6361 2352 6366 2408
rect 6422 2352 18142 2408
rect 18198 2352 18203 2408
rect 6361 2350 18203 2352
rect 6361 2347 6427 2350
rect 18137 2347 18203 2350
rect 4610 2208 4930 2209
rect 4610 2144 4618 2208
rect 4682 2144 4698 2208
rect 4762 2144 4778 2208
rect 4842 2144 4858 2208
rect 4922 2144 4930 2208
rect 4610 2143 4930 2144
rect 11944 2208 12264 2209
rect 11944 2144 11952 2208
rect 12016 2144 12032 2208
rect 12096 2144 12112 2208
rect 12176 2144 12192 2208
rect 12256 2144 12264 2208
rect 11944 2143 12264 2144
rect 19277 2208 19597 2209
rect 19277 2144 19285 2208
rect 19349 2144 19365 2208
rect 19429 2144 19445 2208
rect 19509 2144 19525 2208
rect 19589 2144 19597 2208
rect 19277 2143 19597 2144
rect 5533 2002 5599 2005
rect 15193 2002 15259 2005
rect 5533 2000 15259 2002
rect 5533 1944 5538 2000
rect 5594 1944 15198 2000
rect 15254 1944 15259 2000
rect 5533 1942 15259 1944
rect 5533 1939 5599 1942
rect 15193 1939 15259 1942
rect 0 1732 480 1760
rect 0 1668 60 1732
rect 124 1668 480 1732
rect 0 1640 480 1668
rect 5625 1730 5691 1733
rect 18505 1730 18571 1733
rect 5625 1728 18571 1730
rect 5625 1672 5630 1728
rect 5686 1672 18510 1728
rect 18566 1672 18571 1728
rect 5625 1670 18571 1672
rect 5625 1667 5691 1670
rect 18505 1667 18571 1670
rect 7557 1594 7623 1597
rect 18413 1594 18479 1597
rect 7557 1592 18479 1594
rect 7557 1536 7562 1592
rect 7618 1536 18418 1592
rect 18474 1536 18479 1592
rect 7557 1534 18479 1536
rect 7557 1531 7623 1534
rect 18413 1531 18479 1534
rect 19977 1594 20043 1597
rect 19977 1592 21650 1594
rect 19977 1536 19982 1592
rect 20038 1536 21650 1592
rect 19977 1534 21650 1536
rect 19977 1531 20043 1534
rect 5441 1186 5507 1189
rect 62 1184 5507 1186
rect 62 1128 5446 1184
rect 5502 1128 5507 1184
rect 62 1126 5507 1128
rect 62 672 122 1126
rect 5441 1123 5507 1126
rect 21590 1080 21650 1534
rect 21520 960 22000 1080
rect 0 552 480 672
rect 5165 98 5231 101
rect 6126 98 6132 100
rect 5165 96 6132 98
rect 5165 40 5170 96
rect 5226 40 6132 96
rect 5165 38 6132 40
rect 5165 35 5231 38
rect 6126 36 6132 38
rect 6196 36 6202 100
<< via3 >>
rect 4618 19612 4682 19616
rect 4618 19556 4622 19612
rect 4622 19556 4678 19612
rect 4678 19556 4682 19612
rect 4618 19552 4682 19556
rect 4698 19612 4762 19616
rect 4698 19556 4702 19612
rect 4702 19556 4758 19612
rect 4758 19556 4762 19612
rect 4698 19552 4762 19556
rect 4778 19612 4842 19616
rect 4778 19556 4782 19612
rect 4782 19556 4838 19612
rect 4838 19556 4842 19612
rect 4778 19552 4842 19556
rect 4858 19612 4922 19616
rect 4858 19556 4862 19612
rect 4862 19556 4918 19612
rect 4918 19556 4922 19612
rect 4858 19552 4922 19556
rect 11952 19612 12016 19616
rect 11952 19556 11956 19612
rect 11956 19556 12012 19612
rect 12012 19556 12016 19612
rect 11952 19552 12016 19556
rect 12032 19612 12096 19616
rect 12032 19556 12036 19612
rect 12036 19556 12092 19612
rect 12092 19556 12096 19612
rect 12032 19552 12096 19556
rect 12112 19612 12176 19616
rect 12112 19556 12116 19612
rect 12116 19556 12172 19612
rect 12172 19556 12176 19612
rect 12112 19552 12176 19556
rect 12192 19612 12256 19616
rect 12192 19556 12196 19612
rect 12196 19556 12252 19612
rect 12252 19556 12256 19612
rect 12192 19552 12256 19556
rect 19285 19612 19349 19616
rect 19285 19556 19289 19612
rect 19289 19556 19345 19612
rect 19345 19556 19349 19612
rect 19285 19552 19349 19556
rect 19365 19612 19429 19616
rect 19365 19556 19369 19612
rect 19369 19556 19425 19612
rect 19425 19556 19429 19612
rect 19365 19552 19429 19556
rect 19445 19612 19509 19616
rect 19445 19556 19449 19612
rect 19449 19556 19505 19612
rect 19505 19556 19509 19612
rect 19445 19552 19509 19556
rect 19525 19612 19589 19616
rect 19525 19556 19529 19612
rect 19529 19556 19585 19612
rect 19585 19556 19589 19612
rect 19525 19552 19589 19556
rect 8285 19068 8349 19072
rect 8285 19012 8289 19068
rect 8289 19012 8345 19068
rect 8345 19012 8349 19068
rect 8285 19008 8349 19012
rect 8365 19068 8429 19072
rect 8365 19012 8369 19068
rect 8369 19012 8425 19068
rect 8425 19012 8429 19068
rect 8365 19008 8429 19012
rect 8445 19068 8509 19072
rect 8445 19012 8449 19068
rect 8449 19012 8505 19068
rect 8505 19012 8509 19068
rect 8445 19008 8509 19012
rect 8525 19068 8589 19072
rect 8525 19012 8529 19068
rect 8529 19012 8585 19068
rect 8585 19012 8589 19068
rect 8525 19008 8589 19012
rect 15618 19068 15682 19072
rect 15618 19012 15622 19068
rect 15622 19012 15678 19068
rect 15678 19012 15682 19068
rect 15618 19008 15682 19012
rect 15698 19068 15762 19072
rect 15698 19012 15702 19068
rect 15702 19012 15758 19068
rect 15758 19012 15762 19068
rect 15698 19008 15762 19012
rect 15778 19068 15842 19072
rect 15778 19012 15782 19068
rect 15782 19012 15838 19068
rect 15838 19012 15842 19068
rect 15778 19008 15842 19012
rect 15858 19068 15922 19072
rect 15858 19012 15862 19068
rect 15862 19012 15918 19068
rect 15918 19012 15922 19068
rect 15858 19008 15922 19012
rect 4618 18524 4682 18528
rect 4618 18468 4622 18524
rect 4622 18468 4678 18524
rect 4678 18468 4682 18524
rect 4618 18464 4682 18468
rect 4698 18524 4762 18528
rect 4698 18468 4702 18524
rect 4702 18468 4758 18524
rect 4758 18468 4762 18524
rect 4698 18464 4762 18468
rect 4778 18524 4842 18528
rect 4778 18468 4782 18524
rect 4782 18468 4838 18524
rect 4838 18468 4842 18524
rect 4778 18464 4842 18468
rect 4858 18524 4922 18528
rect 4858 18468 4862 18524
rect 4862 18468 4918 18524
rect 4918 18468 4922 18524
rect 4858 18464 4922 18468
rect 11952 18524 12016 18528
rect 11952 18468 11956 18524
rect 11956 18468 12012 18524
rect 12012 18468 12016 18524
rect 11952 18464 12016 18468
rect 12032 18524 12096 18528
rect 12032 18468 12036 18524
rect 12036 18468 12092 18524
rect 12092 18468 12096 18524
rect 12032 18464 12096 18468
rect 12112 18524 12176 18528
rect 12112 18468 12116 18524
rect 12116 18468 12172 18524
rect 12172 18468 12176 18524
rect 12112 18464 12176 18468
rect 12192 18524 12256 18528
rect 12192 18468 12196 18524
rect 12196 18468 12252 18524
rect 12252 18468 12256 18524
rect 12192 18464 12256 18468
rect 19285 18524 19349 18528
rect 19285 18468 19289 18524
rect 19289 18468 19345 18524
rect 19345 18468 19349 18524
rect 19285 18464 19349 18468
rect 19365 18524 19429 18528
rect 19365 18468 19369 18524
rect 19369 18468 19425 18524
rect 19425 18468 19429 18524
rect 19365 18464 19429 18468
rect 19445 18524 19509 18528
rect 19445 18468 19449 18524
rect 19449 18468 19505 18524
rect 19505 18468 19509 18524
rect 19445 18464 19509 18468
rect 19525 18524 19589 18528
rect 19525 18468 19529 18524
rect 19529 18468 19585 18524
rect 19585 18468 19589 18524
rect 19525 18464 19589 18468
rect 8285 17980 8349 17984
rect 8285 17924 8289 17980
rect 8289 17924 8345 17980
rect 8345 17924 8349 17980
rect 8285 17920 8349 17924
rect 8365 17980 8429 17984
rect 8365 17924 8369 17980
rect 8369 17924 8425 17980
rect 8425 17924 8429 17980
rect 8365 17920 8429 17924
rect 8445 17980 8509 17984
rect 8445 17924 8449 17980
rect 8449 17924 8505 17980
rect 8505 17924 8509 17980
rect 8445 17920 8509 17924
rect 8525 17980 8589 17984
rect 8525 17924 8529 17980
rect 8529 17924 8585 17980
rect 8585 17924 8589 17980
rect 8525 17920 8589 17924
rect 15618 17980 15682 17984
rect 15618 17924 15622 17980
rect 15622 17924 15678 17980
rect 15678 17924 15682 17980
rect 15618 17920 15682 17924
rect 15698 17980 15762 17984
rect 15698 17924 15702 17980
rect 15702 17924 15758 17980
rect 15758 17924 15762 17980
rect 15698 17920 15762 17924
rect 15778 17980 15842 17984
rect 15778 17924 15782 17980
rect 15782 17924 15838 17980
rect 15838 17924 15842 17980
rect 15778 17920 15842 17924
rect 15858 17980 15922 17984
rect 15858 17924 15862 17980
rect 15862 17924 15918 17980
rect 15918 17924 15922 17980
rect 15858 17920 15922 17924
rect 4618 17436 4682 17440
rect 4618 17380 4622 17436
rect 4622 17380 4678 17436
rect 4678 17380 4682 17436
rect 4618 17376 4682 17380
rect 4698 17436 4762 17440
rect 4698 17380 4702 17436
rect 4702 17380 4758 17436
rect 4758 17380 4762 17436
rect 4698 17376 4762 17380
rect 4778 17436 4842 17440
rect 4778 17380 4782 17436
rect 4782 17380 4838 17436
rect 4838 17380 4842 17436
rect 4778 17376 4842 17380
rect 4858 17436 4922 17440
rect 4858 17380 4862 17436
rect 4862 17380 4918 17436
rect 4918 17380 4922 17436
rect 4858 17376 4922 17380
rect 11952 17436 12016 17440
rect 11952 17380 11956 17436
rect 11956 17380 12012 17436
rect 12012 17380 12016 17436
rect 11952 17376 12016 17380
rect 12032 17436 12096 17440
rect 12032 17380 12036 17436
rect 12036 17380 12092 17436
rect 12092 17380 12096 17436
rect 12032 17376 12096 17380
rect 12112 17436 12176 17440
rect 12112 17380 12116 17436
rect 12116 17380 12172 17436
rect 12172 17380 12176 17436
rect 12112 17376 12176 17380
rect 12192 17436 12256 17440
rect 12192 17380 12196 17436
rect 12196 17380 12252 17436
rect 12252 17380 12256 17436
rect 12192 17376 12256 17380
rect 19285 17436 19349 17440
rect 19285 17380 19289 17436
rect 19289 17380 19345 17436
rect 19345 17380 19349 17436
rect 19285 17376 19349 17380
rect 19365 17436 19429 17440
rect 19365 17380 19369 17436
rect 19369 17380 19425 17436
rect 19425 17380 19429 17436
rect 19365 17376 19429 17380
rect 19445 17436 19509 17440
rect 19445 17380 19449 17436
rect 19449 17380 19505 17436
rect 19505 17380 19509 17436
rect 19445 17376 19509 17380
rect 19525 17436 19589 17440
rect 19525 17380 19529 17436
rect 19529 17380 19585 17436
rect 19585 17380 19589 17436
rect 19525 17376 19589 17380
rect 10548 16900 10612 16964
rect 8285 16892 8349 16896
rect 8285 16836 8289 16892
rect 8289 16836 8345 16892
rect 8345 16836 8349 16892
rect 8285 16832 8349 16836
rect 8365 16892 8429 16896
rect 8365 16836 8369 16892
rect 8369 16836 8425 16892
rect 8425 16836 8429 16892
rect 8365 16832 8429 16836
rect 8445 16892 8509 16896
rect 8445 16836 8449 16892
rect 8449 16836 8505 16892
rect 8505 16836 8509 16892
rect 8445 16832 8509 16836
rect 8525 16892 8589 16896
rect 8525 16836 8529 16892
rect 8529 16836 8585 16892
rect 8585 16836 8589 16892
rect 8525 16832 8589 16836
rect 15618 16892 15682 16896
rect 15618 16836 15622 16892
rect 15622 16836 15678 16892
rect 15678 16836 15682 16892
rect 15618 16832 15682 16836
rect 15698 16892 15762 16896
rect 15698 16836 15702 16892
rect 15702 16836 15758 16892
rect 15758 16836 15762 16892
rect 15698 16832 15762 16836
rect 15778 16892 15842 16896
rect 15778 16836 15782 16892
rect 15782 16836 15838 16892
rect 15838 16836 15842 16892
rect 15778 16832 15842 16836
rect 15858 16892 15922 16896
rect 15858 16836 15862 16892
rect 15862 16836 15918 16892
rect 15918 16836 15922 16892
rect 15858 16832 15922 16836
rect 5948 16628 6012 16692
rect 4618 16348 4682 16352
rect 4618 16292 4622 16348
rect 4622 16292 4678 16348
rect 4678 16292 4682 16348
rect 4618 16288 4682 16292
rect 4698 16348 4762 16352
rect 4698 16292 4702 16348
rect 4702 16292 4758 16348
rect 4758 16292 4762 16348
rect 4698 16288 4762 16292
rect 4778 16348 4842 16352
rect 4778 16292 4782 16348
rect 4782 16292 4838 16348
rect 4838 16292 4842 16348
rect 4778 16288 4842 16292
rect 4858 16348 4922 16352
rect 4858 16292 4862 16348
rect 4862 16292 4918 16348
rect 4918 16292 4922 16348
rect 4858 16288 4922 16292
rect 11952 16348 12016 16352
rect 11952 16292 11956 16348
rect 11956 16292 12012 16348
rect 12012 16292 12016 16348
rect 11952 16288 12016 16292
rect 12032 16348 12096 16352
rect 12032 16292 12036 16348
rect 12036 16292 12092 16348
rect 12092 16292 12096 16348
rect 12032 16288 12096 16292
rect 12112 16348 12176 16352
rect 12112 16292 12116 16348
rect 12116 16292 12172 16348
rect 12172 16292 12176 16348
rect 12112 16288 12176 16292
rect 12192 16348 12256 16352
rect 12192 16292 12196 16348
rect 12196 16292 12252 16348
rect 12252 16292 12256 16348
rect 12192 16288 12256 16292
rect 19285 16348 19349 16352
rect 19285 16292 19289 16348
rect 19289 16292 19345 16348
rect 19345 16292 19349 16348
rect 19285 16288 19349 16292
rect 19365 16348 19429 16352
rect 19365 16292 19369 16348
rect 19369 16292 19425 16348
rect 19425 16292 19429 16348
rect 19365 16288 19429 16292
rect 19445 16348 19509 16352
rect 19445 16292 19449 16348
rect 19449 16292 19505 16348
rect 19505 16292 19509 16348
rect 19445 16288 19509 16292
rect 19525 16348 19589 16352
rect 19525 16292 19529 16348
rect 19529 16292 19585 16348
rect 19585 16292 19589 16348
rect 19525 16288 19589 16292
rect 13492 15812 13556 15876
rect 8285 15804 8349 15808
rect 8285 15748 8289 15804
rect 8289 15748 8345 15804
rect 8345 15748 8349 15804
rect 8285 15744 8349 15748
rect 8365 15804 8429 15808
rect 8365 15748 8369 15804
rect 8369 15748 8425 15804
rect 8425 15748 8429 15804
rect 8365 15744 8429 15748
rect 8445 15804 8509 15808
rect 8445 15748 8449 15804
rect 8449 15748 8505 15804
rect 8505 15748 8509 15804
rect 8445 15744 8509 15748
rect 8525 15804 8589 15808
rect 8525 15748 8529 15804
rect 8529 15748 8585 15804
rect 8585 15748 8589 15804
rect 8525 15744 8589 15748
rect 15618 15804 15682 15808
rect 15618 15748 15622 15804
rect 15622 15748 15678 15804
rect 15678 15748 15682 15804
rect 15618 15744 15682 15748
rect 15698 15804 15762 15808
rect 15698 15748 15702 15804
rect 15702 15748 15758 15804
rect 15758 15748 15762 15804
rect 15698 15744 15762 15748
rect 15778 15804 15842 15808
rect 15778 15748 15782 15804
rect 15782 15748 15838 15804
rect 15838 15748 15842 15804
rect 15778 15744 15842 15748
rect 15858 15804 15922 15808
rect 15858 15748 15862 15804
rect 15862 15748 15918 15804
rect 15918 15748 15922 15804
rect 15858 15744 15922 15748
rect 6132 15268 6196 15332
rect 4618 15260 4682 15264
rect 4618 15204 4622 15260
rect 4622 15204 4678 15260
rect 4678 15204 4682 15260
rect 4618 15200 4682 15204
rect 4698 15260 4762 15264
rect 4698 15204 4702 15260
rect 4702 15204 4758 15260
rect 4758 15204 4762 15260
rect 4698 15200 4762 15204
rect 4778 15260 4842 15264
rect 4778 15204 4782 15260
rect 4782 15204 4838 15260
rect 4838 15204 4842 15260
rect 4778 15200 4842 15204
rect 4858 15260 4922 15264
rect 4858 15204 4862 15260
rect 4862 15204 4918 15260
rect 4918 15204 4922 15260
rect 4858 15200 4922 15204
rect 11952 15260 12016 15264
rect 11952 15204 11956 15260
rect 11956 15204 12012 15260
rect 12012 15204 12016 15260
rect 11952 15200 12016 15204
rect 12032 15260 12096 15264
rect 12032 15204 12036 15260
rect 12036 15204 12092 15260
rect 12092 15204 12096 15260
rect 12032 15200 12096 15204
rect 12112 15260 12176 15264
rect 12112 15204 12116 15260
rect 12116 15204 12172 15260
rect 12172 15204 12176 15260
rect 12112 15200 12176 15204
rect 12192 15260 12256 15264
rect 12192 15204 12196 15260
rect 12196 15204 12252 15260
rect 12252 15204 12256 15260
rect 12192 15200 12256 15204
rect 19285 15260 19349 15264
rect 19285 15204 19289 15260
rect 19289 15204 19345 15260
rect 19345 15204 19349 15260
rect 19285 15200 19349 15204
rect 19365 15260 19429 15264
rect 19365 15204 19369 15260
rect 19369 15204 19425 15260
rect 19425 15204 19429 15260
rect 19365 15200 19429 15204
rect 19445 15260 19509 15264
rect 19445 15204 19449 15260
rect 19449 15204 19505 15260
rect 19505 15204 19509 15260
rect 19445 15200 19509 15204
rect 19525 15260 19589 15264
rect 19525 15204 19529 15260
rect 19529 15204 19585 15260
rect 19585 15204 19589 15260
rect 19525 15200 19589 15204
rect 8285 14716 8349 14720
rect 8285 14660 8289 14716
rect 8289 14660 8345 14716
rect 8345 14660 8349 14716
rect 8285 14656 8349 14660
rect 8365 14716 8429 14720
rect 8365 14660 8369 14716
rect 8369 14660 8425 14716
rect 8425 14660 8429 14716
rect 8365 14656 8429 14660
rect 8445 14716 8509 14720
rect 8445 14660 8449 14716
rect 8449 14660 8505 14716
rect 8505 14660 8509 14716
rect 8445 14656 8509 14660
rect 8525 14716 8589 14720
rect 8525 14660 8529 14716
rect 8529 14660 8585 14716
rect 8585 14660 8589 14716
rect 8525 14656 8589 14660
rect 15618 14716 15682 14720
rect 15618 14660 15622 14716
rect 15622 14660 15678 14716
rect 15678 14660 15682 14716
rect 15618 14656 15682 14660
rect 15698 14716 15762 14720
rect 15698 14660 15702 14716
rect 15702 14660 15758 14716
rect 15758 14660 15762 14716
rect 15698 14656 15762 14660
rect 15778 14716 15842 14720
rect 15778 14660 15782 14716
rect 15782 14660 15838 14716
rect 15838 14660 15842 14716
rect 15778 14656 15842 14660
rect 15858 14716 15922 14720
rect 15858 14660 15862 14716
rect 15862 14660 15918 14716
rect 15918 14660 15922 14716
rect 15858 14656 15922 14660
rect 13492 14180 13556 14244
rect 4618 14172 4682 14176
rect 4618 14116 4622 14172
rect 4622 14116 4678 14172
rect 4678 14116 4682 14172
rect 4618 14112 4682 14116
rect 4698 14172 4762 14176
rect 4698 14116 4702 14172
rect 4702 14116 4758 14172
rect 4758 14116 4762 14172
rect 4698 14112 4762 14116
rect 4778 14172 4842 14176
rect 4778 14116 4782 14172
rect 4782 14116 4838 14172
rect 4838 14116 4842 14172
rect 4778 14112 4842 14116
rect 4858 14172 4922 14176
rect 4858 14116 4862 14172
rect 4862 14116 4918 14172
rect 4918 14116 4922 14172
rect 4858 14112 4922 14116
rect 11952 14172 12016 14176
rect 11952 14116 11956 14172
rect 11956 14116 12012 14172
rect 12012 14116 12016 14172
rect 11952 14112 12016 14116
rect 12032 14172 12096 14176
rect 12032 14116 12036 14172
rect 12036 14116 12092 14172
rect 12092 14116 12096 14172
rect 12032 14112 12096 14116
rect 12112 14172 12176 14176
rect 12112 14116 12116 14172
rect 12116 14116 12172 14172
rect 12172 14116 12176 14172
rect 12112 14112 12176 14116
rect 12192 14172 12256 14176
rect 12192 14116 12196 14172
rect 12196 14116 12252 14172
rect 12252 14116 12256 14172
rect 12192 14112 12256 14116
rect 19285 14172 19349 14176
rect 19285 14116 19289 14172
rect 19289 14116 19345 14172
rect 19345 14116 19349 14172
rect 19285 14112 19349 14116
rect 19365 14172 19429 14176
rect 19365 14116 19369 14172
rect 19369 14116 19425 14172
rect 19425 14116 19429 14172
rect 19365 14112 19429 14116
rect 19445 14172 19509 14176
rect 19445 14116 19449 14172
rect 19449 14116 19505 14172
rect 19505 14116 19509 14172
rect 19445 14112 19509 14116
rect 19525 14172 19589 14176
rect 19525 14116 19529 14172
rect 19529 14116 19585 14172
rect 19585 14116 19589 14172
rect 19525 14112 19589 14116
rect 9628 14044 9692 14108
rect 9076 13908 9140 13972
rect 60 13772 124 13836
rect 8285 13628 8349 13632
rect 8285 13572 8289 13628
rect 8289 13572 8345 13628
rect 8345 13572 8349 13628
rect 8285 13568 8349 13572
rect 8365 13628 8429 13632
rect 8365 13572 8369 13628
rect 8369 13572 8425 13628
rect 8425 13572 8429 13628
rect 8365 13568 8429 13572
rect 8445 13628 8509 13632
rect 8445 13572 8449 13628
rect 8449 13572 8505 13628
rect 8505 13572 8509 13628
rect 8445 13568 8509 13572
rect 8525 13628 8589 13632
rect 8525 13572 8529 13628
rect 8529 13572 8585 13628
rect 8585 13572 8589 13628
rect 8525 13568 8589 13572
rect 15618 13628 15682 13632
rect 15618 13572 15622 13628
rect 15622 13572 15678 13628
rect 15678 13572 15682 13628
rect 15618 13568 15682 13572
rect 15698 13628 15762 13632
rect 15698 13572 15702 13628
rect 15702 13572 15758 13628
rect 15758 13572 15762 13628
rect 15698 13568 15762 13572
rect 15778 13628 15842 13632
rect 15778 13572 15782 13628
rect 15782 13572 15838 13628
rect 15838 13572 15842 13628
rect 15778 13568 15842 13572
rect 15858 13628 15922 13632
rect 15858 13572 15862 13628
rect 15862 13572 15918 13628
rect 15918 13572 15922 13628
rect 15858 13568 15922 13572
rect 14596 13500 14660 13564
rect 4618 13084 4682 13088
rect 4618 13028 4622 13084
rect 4622 13028 4678 13084
rect 4678 13028 4682 13084
rect 4618 13024 4682 13028
rect 4698 13084 4762 13088
rect 4698 13028 4702 13084
rect 4702 13028 4758 13084
rect 4758 13028 4762 13084
rect 4698 13024 4762 13028
rect 4778 13084 4842 13088
rect 4778 13028 4782 13084
rect 4782 13028 4838 13084
rect 4838 13028 4842 13084
rect 4778 13024 4842 13028
rect 4858 13084 4922 13088
rect 4858 13028 4862 13084
rect 4862 13028 4918 13084
rect 4918 13028 4922 13084
rect 4858 13024 4922 13028
rect 11952 13084 12016 13088
rect 11952 13028 11956 13084
rect 11956 13028 12012 13084
rect 12012 13028 12016 13084
rect 11952 13024 12016 13028
rect 12032 13084 12096 13088
rect 12032 13028 12036 13084
rect 12036 13028 12092 13084
rect 12092 13028 12096 13084
rect 12032 13024 12096 13028
rect 12112 13084 12176 13088
rect 12112 13028 12116 13084
rect 12116 13028 12172 13084
rect 12172 13028 12176 13084
rect 12112 13024 12176 13028
rect 12192 13084 12256 13088
rect 12192 13028 12196 13084
rect 12196 13028 12252 13084
rect 12252 13028 12256 13084
rect 12192 13024 12256 13028
rect 19285 13084 19349 13088
rect 19285 13028 19289 13084
rect 19289 13028 19345 13084
rect 19345 13028 19349 13084
rect 19285 13024 19349 13028
rect 19365 13084 19429 13088
rect 19365 13028 19369 13084
rect 19369 13028 19425 13084
rect 19425 13028 19429 13084
rect 19365 13024 19429 13028
rect 19445 13084 19509 13088
rect 19445 13028 19449 13084
rect 19449 13028 19505 13084
rect 19505 13028 19509 13084
rect 19445 13024 19509 13028
rect 19525 13084 19589 13088
rect 19525 13028 19529 13084
rect 19529 13028 19585 13084
rect 19585 13028 19589 13084
rect 19525 13024 19589 13028
rect 8285 12540 8349 12544
rect 8285 12484 8289 12540
rect 8289 12484 8345 12540
rect 8345 12484 8349 12540
rect 8285 12480 8349 12484
rect 8365 12540 8429 12544
rect 8365 12484 8369 12540
rect 8369 12484 8425 12540
rect 8425 12484 8429 12540
rect 8365 12480 8429 12484
rect 8445 12540 8509 12544
rect 8445 12484 8449 12540
rect 8449 12484 8505 12540
rect 8505 12484 8509 12540
rect 8445 12480 8509 12484
rect 8525 12540 8589 12544
rect 8525 12484 8529 12540
rect 8529 12484 8585 12540
rect 8585 12484 8589 12540
rect 8525 12480 8589 12484
rect 15618 12540 15682 12544
rect 15618 12484 15622 12540
rect 15622 12484 15678 12540
rect 15678 12484 15682 12540
rect 15618 12480 15682 12484
rect 15698 12540 15762 12544
rect 15698 12484 15702 12540
rect 15702 12484 15758 12540
rect 15758 12484 15762 12540
rect 15698 12480 15762 12484
rect 15778 12540 15842 12544
rect 15778 12484 15782 12540
rect 15782 12484 15838 12540
rect 15838 12484 15842 12540
rect 15778 12480 15842 12484
rect 15858 12540 15922 12544
rect 15858 12484 15862 12540
rect 15862 12484 15918 12540
rect 15918 12484 15922 12540
rect 15858 12480 15922 12484
rect 4618 11996 4682 12000
rect 4618 11940 4622 11996
rect 4622 11940 4678 11996
rect 4678 11940 4682 11996
rect 4618 11936 4682 11940
rect 4698 11996 4762 12000
rect 4698 11940 4702 11996
rect 4702 11940 4758 11996
rect 4758 11940 4762 11996
rect 4698 11936 4762 11940
rect 4778 11996 4842 12000
rect 4778 11940 4782 11996
rect 4782 11940 4838 11996
rect 4838 11940 4842 11996
rect 4778 11936 4842 11940
rect 4858 11996 4922 12000
rect 4858 11940 4862 11996
rect 4862 11940 4918 11996
rect 4918 11940 4922 11996
rect 4858 11936 4922 11940
rect 11952 11996 12016 12000
rect 11952 11940 11956 11996
rect 11956 11940 12012 11996
rect 12012 11940 12016 11996
rect 11952 11936 12016 11940
rect 12032 11996 12096 12000
rect 12032 11940 12036 11996
rect 12036 11940 12092 11996
rect 12092 11940 12096 11996
rect 12032 11936 12096 11940
rect 12112 11996 12176 12000
rect 12112 11940 12116 11996
rect 12116 11940 12172 11996
rect 12172 11940 12176 11996
rect 12112 11936 12176 11940
rect 12192 11996 12256 12000
rect 12192 11940 12196 11996
rect 12196 11940 12252 11996
rect 12252 11940 12256 11996
rect 12192 11936 12256 11940
rect 19285 11996 19349 12000
rect 19285 11940 19289 11996
rect 19289 11940 19345 11996
rect 19345 11940 19349 11996
rect 19285 11936 19349 11940
rect 19365 11996 19429 12000
rect 19365 11940 19369 11996
rect 19369 11940 19425 11996
rect 19425 11940 19429 11996
rect 19365 11936 19429 11940
rect 19445 11996 19509 12000
rect 19445 11940 19449 11996
rect 19449 11940 19505 11996
rect 19505 11940 19509 11996
rect 19445 11936 19509 11940
rect 19525 11996 19589 12000
rect 19525 11940 19529 11996
rect 19529 11940 19585 11996
rect 19585 11940 19589 11996
rect 19525 11936 19589 11940
rect 5948 11868 6012 11932
rect 9628 11460 9692 11524
rect 8285 11452 8349 11456
rect 8285 11396 8289 11452
rect 8289 11396 8345 11452
rect 8345 11396 8349 11452
rect 8285 11392 8349 11396
rect 8365 11452 8429 11456
rect 8365 11396 8369 11452
rect 8369 11396 8425 11452
rect 8425 11396 8429 11452
rect 8365 11392 8429 11396
rect 8445 11452 8509 11456
rect 8445 11396 8449 11452
rect 8449 11396 8505 11452
rect 8505 11396 8509 11452
rect 8445 11392 8509 11396
rect 8525 11452 8589 11456
rect 8525 11396 8529 11452
rect 8529 11396 8585 11452
rect 8585 11396 8589 11452
rect 8525 11392 8589 11396
rect 15618 11452 15682 11456
rect 15618 11396 15622 11452
rect 15622 11396 15678 11452
rect 15678 11396 15682 11452
rect 15618 11392 15682 11396
rect 15698 11452 15762 11456
rect 15698 11396 15702 11452
rect 15702 11396 15758 11452
rect 15758 11396 15762 11452
rect 15698 11392 15762 11396
rect 15778 11452 15842 11456
rect 15778 11396 15782 11452
rect 15782 11396 15838 11452
rect 15838 11396 15842 11452
rect 15778 11392 15842 11396
rect 15858 11452 15922 11456
rect 15858 11396 15862 11452
rect 15862 11396 15918 11452
rect 15918 11396 15922 11452
rect 15858 11392 15922 11396
rect 4618 10908 4682 10912
rect 4618 10852 4622 10908
rect 4622 10852 4678 10908
rect 4678 10852 4682 10908
rect 4618 10848 4682 10852
rect 4698 10908 4762 10912
rect 4698 10852 4702 10908
rect 4702 10852 4758 10908
rect 4758 10852 4762 10908
rect 4698 10848 4762 10852
rect 4778 10908 4842 10912
rect 4778 10852 4782 10908
rect 4782 10852 4838 10908
rect 4838 10852 4842 10908
rect 4778 10848 4842 10852
rect 4858 10908 4922 10912
rect 4858 10852 4862 10908
rect 4862 10852 4918 10908
rect 4918 10852 4922 10908
rect 4858 10848 4922 10852
rect 11952 10908 12016 10912
rect 11952 10852 11956 10908
rect 11956 10852 12012 10908
rect 12012 10852 12016 10908
rect 11952 10848 12016 10852
rect 12032 10908 12096 10912
rect 12032 10852 12036 10908
rect 12036 10852 12092 10908
rect 12092 10852 12096 10908
rect 12032 10848 12096 10852
rect 12112 10908 12176 10912
rect 12112 10852 12116 10908
rect 12116 10852 12172 10908
rect 12172 10852 12176 10908
rect 12112 10848 12176 10852
rect 12192 10908 12256 10912
rect 12192 10852 12196 10908
rect 12196 10852 12252 10908
rect 12252 10852 12256 10908
rect 12192 10848 12256 10852
rect 19285 10908 19349 10912
rect 19285 10852 19289 10908
rect 19289 10852 19345 10908
rect 19345 10852 19349 10908
rect 19285 10848 19349 10852
rect 19365 10908 19429 10912
rect 19365 10852 19369 10908
rect 19369 10852 19425 10908
rect 19425 10852 19429 10908
rect 19365 10848 19429 10852
rect 19445 10908 19509 10912
rect 19445 10852 19449 10908
rect 19449 10852 19505 10908
rect 19505 10852 19509 10908
rect 19445 10848 19509 10852
rect 19525 10908 19589 10912
rect 19525 10852 19529 10908
rect 19529 10852 19585 10908
rect 19585 10852 19589 10908
rect 19525 10848 19589 10852
rect 8285 10364 8349 10368
rect 8285 10308 8289 10364
rect 8289 10308 8345 10364
rect 8345 10308 8349 10364
rect 8285 10304 8349 10308
rect 8365 10364 8429 10368
rect 8365 10308 8369 10364
rect 8369 10308 8425 10364
rect 8425 10308 8429 10364
rect 8365 10304 8429 10308
rect 8445 10364 8509 10368
rect 8445 10308 8449 10364
rect 8449 10308 8505 10364
rect 8505 10308 8509 10364
rect 8445 10304 8509 10308
rect 8525 10364 8589 10368
rect 8525 10308 8529 10364
rect 8529 10308 8585 10364
rect 8585 10308 8589 10364
rect 8525 10304 8589 10308
rect 15618 10364 15682 10368
rect 15618 10308 15622 10364
rect 15622 10308 15678 10364
rect 15678 10308 15682 10364
rect 15618 10304 15682 10308
rect 15698 10364 15762 10368
rect 15698 10308 15702 10364
rect 15702 10308 15758 10364
rect 15758 10308 15762 10364
rect 15698 10304 15762 10308
rect 15778 10364 15842 10368
rect 15778 10308 15782 10364
rect 15782 10308 15838 10364
rect 15838 10308 15842 10364
rect 15778 10304 15842 10308
rect 15858 10364 15922 10368
rect 15858 10308 15862 10364
rect 15862 10308 15918 10364
rect 15918 10308 15922 10364
rect 15858 10304 15922 10308
rect 4618 9820 4682 9824
rect 4618 9764 4622 9820
rect 4622 9764 4678 9820
rect 4678 9764 4682 9820
rect 4618 9760 4682 9764
rect 4698 9820 4762 9824
rect 4698 9764 4702 9820
rect 4702 9764 4758 9820
rect 4758 9764 4762 9820
rect 4698 9760 4762 9764
rect 4778 9820 4842 9824
rect 4778 9764 4782 9820
rect 4782 9764 4838 9820
rect 4838 9764 4842 9820
rect 4778 9760 4842 9764
rect 4858 9820 4922 9824
rect 4858 9764 4862 9820
rect 4862 9764 4918 9820
rect 4918 9764 4922 9820
rect 4858 9760 4922 9764
rect 11952 9820 12016 9824
rect 11952 9764 11956 9820
rect 11956 9764 12012 9820
rect 12012 9764 12016 9820
rect 11952 9760 12016 9764
rect 12032 9820 12096 9824
rect 12032 9764 12036 9820
rect 12036 9764 12092 9820
rect 12092 9764 12096 9820
rect 12032 9760 12096 9764
rect 12112 9820 12176 9824
rect 12112 9764 12116 9820
rect 12116 9764 12172 9820
rect 12172 9764 12176 9820
rect 12112 9760 12176 9764
rect 12192 9820 12256 9824
rect 12192 9764 12196 9820
rect 12196 9764 12252 9820
rect 12252 9764 12256 9820
rect 12192 9760 12256 9764
rect 19285 9820 19349 9824
rect 19285 9764 19289 9820
rect 19289 9764 19345 9820
rect 19345 9764 19349 9820
rect 19285 9760 19349 9764
rect 19365 9820 19429 9824
rect 19365 9764 19369 9820
rect 19369 9764 19425 9820
rect 19425 9764 19429 9820
rect 19365 9760 19429 9764
rect 19445 9820 19509 9824
rect 19445 9764 19449 9820
rect 19449 9764 19505 9820
rect 19505 9764 19509 9820
rect 19445 9760 19509 9764
rect 19525 9820 19589 9824
rect 19525 9764 19529 9820
rect 19529 9764 19585 9820
rect 19585 9764 19589 9820
rect 19525 9760 19589 9764
rect 10548 9420 10612 9484
rect 8285 9276 8349 9280
rect 8285 9220 8289 9276
rect 8289 9220 8345 9276
rect 8345 9220 8349 9276
rect 8285 9216 8349 9220
rect 8365 9276 8429 9280
rect 8365 9220 8369 9276
rect 8369 9220 8425 9276
rect 8425 9220 8429 9276
rect 8365 9216 8429 9220
rect 8445 9276 8509 9280
rect 8445 9220 8449 9276
rect 8449 9220 8505 9276
rect 8505 9220 8509 9276
rect 8445 9216 8509 9220
rect 8525 9276 8589 9280
rect 8525 9220 8529 9276
rect 8529 9220 8585 9276
rect 8585 9220 8589 9276
rect 8525 9216 8589 9220
rect 15618 9276 15682 9280
rect 15618 9220 15622 9276
rect 15622 9220 15678 9276
rect 15678 9220 15682 9276
rect 15618 9216 15682 9220
rect 15698 9276 15762 9280
rect 15698 9220 15702 9276
rect 15702 9220 15758 9276
rect 15758 9220 15762 9276
rect 15698 9216 15762 9220
rect 15778 9276 15842 9280
rect 15778 9220 15782 9276
rect 15782 9220 15838 9276
rect 15838 9220 15842 9276
rect 15778 9216 15842 9220
rect 15858 9276 15922 9280
rect 15858 9220 15862 9276
rect 15862 9220 15918 9276
rect 15918 9220 15922 9276
rect 15858 9216 15922 9220
rect 4618 8732 4682 8736
rect 4618 8676 4622 8732
rect 4622 8676 4678 8732
rect 4678 8676 4682 8732
rect 4618 8672 4682 8676
rect 4698 8732 4762 8736
rect 4698 8676 4702 8732
rect 4702 8676 4758 8732
rect 4758 8676 4762 8732
rect 4698 8672 4762 8676
rect 4778 8732 4842 8736
rect 4778 8676 4782 8732
rect 4782 8676 4838 8732
rect 4838 8676 4842 8732
rect 4778 8672 4842 8676
rect 4858 8732 4922 8736
rect 4858 8676 4862 8732
rect 4862 8676 4918 8732
rect 4918 8676 4922 8732
rect 4858 8672 4922 8676
rect 11952 8732 12016 8736
rect 11952 8676 11956 8732
rect 11956 8676 12012 8732
rect 12012 8676 12016 8732
rect 11952 8672 12016 8676
rect 12032 8732 12096 8736
rect 12032 8676 12036 8732
rect 12036 8676 12092 8732
rect 12092 8676 12096 8732
rect 12032 8672 12096 8676
rect 12112 8732 12176 8736
rect 12112 8676 12116 8732
rect 12116 8676 12172 8732
rect 12172 8676 12176 8732
rect 12112 8672 12176 8676
rect 12192 8732 12256 8736
rect 12192 8676 12196 8732
rect 12196 8676 12252 8732
rect 12252 8676 12256 8732
rect 12192 8672 12256 8676
rect 19285 8732 19349 8736
rect 19285 8676 19289 8732
rect 19289 8676 19345 8732
rect 19345 8676 19349 8732
rect 19285 8672 19349 8676
rect 19365 8732 19429 8736
rect 19365 8676 19369 8732
rect 19369 8676 19425 8732
rect 19425 8676 19429 8732
rect 19365 8672 19429 8676
rect 19445 8732 19509 8736
rect 19445 8676 19449 8732
rect 19449 8676 19505 8732
rect 19505 8676 19509 8732
rect 19445 8672 19509 8676
rect 19525 8732 19589 8736
rect 19525 8676 19529 8732
rect 19529 8676 19585 8732
rect 19585 8676 19589 8732
rect 19525 8672 19589 8676
rect 9076 8604 9140 8668
rect 8285 8188 8349 8192
rect 8285 8132 8289 8188
rect 8289 8132 8345 8188
rect 8345 8132 8349 8188
rect 8285 8128 8349 8132
rect 8365 8188 8429 8192
rect 8365 8132 8369 8188
rect 8369 8132 8425 8188
rect 8425 8132 8429 8188
rect 8365 8128 8429 8132
rect 8445 8188 8509 8192
rect 8445 8132 8449 8188
rect 8449 8132 8505 8188
rect 8505 8132 8509 8188
rect 8445 8128 8509 8132
rect 8525 8188 8589 8192
rect 8525 8132 8529 8188
rect 8529 8132 8585 8188
rect 8585 8132 8589 8188
rect 8525 8128 8589 8132
rect 15618 8188 15682 8192
rect 15618 8132 15622 8188
rect 15622 8132 15678 8188
rect 15678 8132 15682 8188
rect 15618 8128 15682 8132
rect 15698 8188 15762 8192
rect 15698 8132 15702 8188
rect 15702 8132 15758 8188
rect 15758 8132 15762 8188
rect 15698 8128 15762 8132
rect 15778 8188 15842 8192
rect 15778 8132 15782 8188
rect 15782 8132 15838 8188
rect 15838 8132 15842 8188
rect 15778 8128 15842 8132
rect 15858 8188 15922 8192
rect 15858 8132 15862 8188
rect 15862 8132 15918 8188
rect 15918 8132 15922 8188
rect 15858 8128 15922 8132
rect 4618 7644 4682 7648
rect 4618 7588 4622 7644
rect 4622 7588 4678 7644
rect 4678 7588 4682 7644
rect 4618 7584 4682 7588
rect 4698 7644 4762 7648
rect 4698 7588 4702 7644
rect 4702 7588 4758 7644
rect 4758 7588 4762 7644
rect 4698 7584 4762 7588
rect 4778 7644 4842 7648
rect 4778 7588 4782 7644
rect 4782 7588 4838 7644
rect 4838 7588 4842 7644
rect 4778 7584 4842 7588
rect 4858 7644 4922 7648
rect 4858 7588 4862 7644
rect 4862 7588 4918 7644
rect 4918 7588 4922 7644
rect 4858 7584 4922 7588
rect 11952 7644 12016 7648
rect 11952 7588 11956 7644
rect 11956 7588 12012 7644
rect 12012 7588 12016 7644
rect 11952 7584 12016 7588
rect 12032 7644 12096 7648
rect 12032 7588 12036 7644
rect 12036 7588 12092 7644
rect 12092 7588 12096 7644
rect 12032 7584 12096 7588
rect 12112 7644 12176 7648
rect 12112 7588 12116 7644
rect 12116 7588 12172 7644
rect 12172 7588 12176 7644
rect 12112 7584 12176 7588
rect 12192 7644 12256 7648
rect 12192 7588 12196 7644
rect 12196 7588 12252 7644
rect 12252 7588 12256 7644
rect 12192 7584 12256 7588
rect 19285 7644 19349 7648
rect 19285 7588 19289 7644
rect 19289 7588 19345 7644
rect 19345 7588 19349 7644
rect 19285 7584 19349 7588
rect 19365 7644 19429 7648
rect 19365 7588 19369 7644
rect 19369 7588 19425 7644
rect 19425 7588 19429 7644
rect 19365 7584 19429 7588
rect 19445 7644 19509 7648
rect 19445 7588 19449 7644
rect 19449 7588 19505 7644
rect 19505 7588 19509 7644
rect 19445 7584 19509 7588
rect 19525 7644 19589 7648
rect 19525 7588 19529 7644
rect 19529 7588 19585 7644
rect 19585 7588 19589 7644
rect 19525 7584 19589 7588
rect 8285 7100 8349 7104
rect 8285 7044 8289 7100
rect 8289 7044 8345 7100
rect 8345 7044 8349 7100
rect 8285 7040 8349 7044
rect 8365 7100 8429 7104
rect 8365 7044 8369 7100
rect 8369 7044 8425 7100
rect 8425 7044 8429 7100
rect 8365 7040 8429 7044
rect 8445 7100 8509 7104
rect 8445 7044 8449 7100
rect 8449 7044 8505 7100
rect 8505 7044 8509 7100
rect 8445 7040 8509 7044
rect 8525 7100 8589 7104
rect 8525 7044 8529 7100
rect 8529 7044 8585 7100
rect 8585 7044 8589 7100
rect 8525 7040 8589 7044
rect 15618 7100 15682 7104
rect 15618 7044 15622 7100
rect 15622 7044 15678 7100
rect 15678 7044 15682 7100
rect 15618 7040 15682 7044
rect 15698 7100 15762 7104
rect 15698 7044 15702 7100
rect 15702 7044 15758 7100
rect 15758 7044 15762 7100
rect 15698 7040 15762 7044
rect 15778 7100 15842 7104
rect 15778 7044 15782 7100
rect 15782 7044 15838 7100
rect 15838 7044 15842 7100
rect 15778 7040 15842 7044
rect 15858 7100 15922 7104
rect 15858 7044 15862 7100
rect 15862 7044 15918 7100
rect 15918 7044 15922 7100
rect 15858 7040 15922 7044
rect 4618 6556 4682 6560
rect 4618 6500 4622 6556
rect 4622 6500 4678 6556
rect 4678 6500 4682 6556
rect 4618 6496 4682 6500
rect 4698 6556 4762 6560
rect 4698 6500 4702 6556
rect 4702 6500 4758 6556
rect 4758 6500 4762 6556
rect 4698 6496 4762 6500
rect 4778 6556 4842 6560
rect 4778 6500 4782 6556
rect 4782 6500 4838 6556
rect 4838 6500 4842 6556
rect 4778 6496 4842 6500
rect 4858 6556 4922 6560
rect 4858 6500 4862 6556
rect 4862 6500 4918 6556
rect 4918 6500 4922 6556
rect 4858 6496 4922 6500
rect 11952 6556 12016 6560
rect 11952 6500 11956 6556
rect 11956 6500 12012 6556
rect 12012 6500 12016 6556
rect 11952 6496 12016 6500
rect 12032 6556 12096 6560
rect 12032 6500 12036 6556
rect 12036 6500 12092 6556
rect 12092 6500 12096 6556
rect 12032 6496 12096 6500
rect 12112 6556 12176 6560
rect 12112 6500 12116 6556
rect 12116 6500 12172 6556
rect 12172 6500 12176 6556
rect 12112 6496 12176 6500
rect 12192 6556 12256 6560
rect 12192 6500 12196 6556
rect 12196 6500 12252 6556
rect 12252 6500 12256 6556
rect 12192 6496 12256 6500
rect 19285 6556 19349 6560
rect 19285 6500 19289 6556
rect 19289 6500 19345 6556
rect 19345 6500 19349 6556
rect 19285 6496 19349 6500
rect 19365 6556 19429 6560
rect 19365 6500 19369 6556
rect 19369 6500 19425 6556
rect 19425 6500 19429 6556
rect 19365 6496 19429 6500
rect 19445 6556 19509 6560
rect 19445 6500 19449 6556
rect 19449 6500 19505 6556
rect 19505 6500 19509 6556
rect 19445 6496 19509 6500
rect 19525 6556 19589 6560
rect 19525 6500 19529 6556
rect 19529 6500 19585 6556
rect 19585 6500 19589 6556
rect 19525 6496 19589 6500
rect 8285 6012 8349 6016
rect 8285 5956 8289 6012
rect 8289 5956 8345 6012
rect 8345 5956 8349 6012
rect 8285 5952 8349 5956
rect 8365 6012 8429 6016
rect 8365 5956 8369 6012
rect 8369 5956 8425 6012
rect 8425 5956 8429 6012
rect 8365 5952 8429 5956
rect 8445 6012 8509 6016
rect 8445 5956 8449 6012
rect 8449 5956 8505 6012
rect 8505 5956 8509 6012
rect 8445 5952 8509 5956
rect 8525 6012 8589 6016
rect 8525 5956 8529 6012
rect 8529 5956 8585 6012
rect 8585 5956 8589 6012
rect 8525 5952 8589 5956
rect 15618 6012 15682 6016
rect 15618 5956 15622 6012
rect 15622 5956 15678 6012
rect 15678 5956 15682 6012
rect 15618 5952 15682 5956
rect 15698 6012 15762 6016
rect 15698 5956 15702 6012
rect 15702 5956 15758 6012
rect 15758 5956 15762 6012
rect 15698 5952 15762 5956
rect 15778 6012 15842 6016
rect 15778 5956 15782 6012
rect 15782 5956 15838 6012
rect 15838 5956 15842 6012
rect 15778 5952 15842 5956
rect 15858 6012 15922 6016
rect 15858 5956 15862 6012
rect 15862 5956 15918 6012
rect 15918 5956 15922 6012
rect 15858 5952 15922 5956
rect 4618 5468 4682 5472
rect 4618 5412 4622 5468
rect 4622 5412 4678 5468
rect 4678 5412 4682 5468
rect 4618 5408 4682 5412
rect 4698 5468 4762 5472
rect 4698 5412 4702 5468
rect 4702 5412 4758 5468
rect 4758 5412 4762 5468
rect 4698 5408 4762 5412
rect 4778 5468 4842 5472
rect 4778 5412 4782 5468
rect 4782 5412 4838 5468
rect 4838 5412 4842 5468
rect 4778 5408 4842 5412
rect 4858 5468 4922 5472
rect 4858 5412 4862 5468
rect 4862 5412 4918 5468
rect 4918 5412 4922 5468
rect 4858 5408 4922 5412
rect 11952 5468 12016 5472
rect 11952 5412 11956 5468
rect 11956 5412 12012 5468
rect 12012 5412 12016 5468
rect 11952 5408 12016 5412
rect 12032 5468 12096 5472
rect 12032 5412 12036 5468
rect 12036 5412 12092 5468
rect 12092 5412 12096 5468
rect 12032 5408 12096 5412
rect 12112 5468 12176 5472
rect 12112 5412 12116 5468
rect 12116 5412 12172 5468
rect 12172 5412 12176 5468
rect 12112 5408 12176 5412
rect 12192 5468 12256 5472
rect 12192 5412 12196 5468
rect 12196 5412 12252 5468
rect 12252 5412 12256 5468
rect 12192 5408 12256 5412
rect 19285 5468 19349 5472
rect 19285 5412 19289 5468
rect 19289 5412 19345 5468
rect 19345 5412 19349 5468
rect 19285 5408 19349 5412
rect 19365 5468 19429 5472
rect 19365 5412 19369 5468
rect 19369 5412 19425 5468
rect 19425 5412 19429 5468
rect 19365 5408 19429 5412
rect 19445 5468 19509 5472
rect 19445 5412 19449 5468
rect 19449 5412 19505 5468
rect 19505 5412 19509 5468
rect 19445 5408 19509 5412
rect 19525 5468 19589 5472
rect 19525 5412 19529 5468
rect 19529 5412 19585 5468
rect 19585 5412 19589 5468
rect 19525 5408 19589 5412
rect 60 5204 124 5268
rect 18276 5204 18340 5268
rect 8285 4924 8349 4928
rect 8285 4868 8289 4924
rect 8289 4868 8345 4924
rect 8345 4868 8349 4924
rect 8285 4864 8349 4868
rect 8365 4924 8429 4928
rect 8365 4868 8369 4924
rect 8369 4868 8425 4924
rect 8425 4868 8429 4924
rect 8365 4864 8429 4868
rect 8445 4924 8509 4928
rect 8445 4868 8449 4924
rect 8449 4868 8505 4924
rect 8505 4868 8509 4924
rect 8445 4864 8509 4868
rect 8525 4924 8589 4928
rect 8525 4868 8529 4924
rect 8529 4868 8585 4924
rect 8585 4868 8589 4924
rect 8525 4864 8589 4868
rect 15618 4924 15682 4928
rect 15618 4868 15622 4924
rect 15622 4868 15678 4924
rect 15678 4868 15682 4924
rect 15618 4864 15682 4868
rect 15698 4924 15762 4928
rect 15698 4868 15702 4924
rect 15702 4868 15758 4924
rect 15758 4868 15762 4924
rect 15698 4864 15762 4868
rect 15778 4924 15842 4928
rect 15778 4868 15782 4924
rect 15782 4868 15838 4924
rect 15838 4868 15842 4924
rect 15778 4864 15842 4868
rect 15858 4924 15922 4928
rect 15858 4868 15862 4924
rect 15862 4868 15918 4924
rect 15918 4868 15922 4924
rect 15858 4864 15922 4868
rect 4618 4380 4682 4384
rect 4618 4324 4622 4380
rect 4622 4324 4678 4380
rect 4678 4324 4682 4380
rect 4618 4320 4682 4324
rect 4698 4380 4762 4384
rect 4698 4324 4702 4380
rect 4702 4324 4758 4380
rect 4758 4324 4762 4380
rect 4698 4320 4762 4324
rect 4778 4380 4842 4384
rect 4778 4324 4782 4380
rect 4782 4324 4838 4380
rect 4838 4324 4842 4380
rect 4778 4320 4842 4324
rect 4858 4380 4922 4384
rect 4858 4324 4862 4380
rect 4862 4324 4918 4380
rect 4918 4324 4922 4380
rect 4858 4320 4922 4324
rect 11952 4380 12016 4384
rect 11952 4324 11956 4380
rect 11956 4324 12012 4380
rect 12012 4324 12016 4380
rect 11952 4320 12016 4324
rect 12032 4380 12096 4384
rect 12032 4324 12036 4380
rect 12036 4324 12092 4380
rect 12092 4324 12096 4380
rect 12032 4320 12096 4324
rect 12112 4380 12176 4384
rect 12112 4324 12116 4380
rect 12116 4324 12172 4380
rect 12172 4324 12176 4380
rect 12112 4320 12176 4324
rect 12192 4380 12256 4384
rect 12192 4324 12196 4380
rect 12196 4324 12252 4380
rect 12252 4324 12256 4380
rect 12192 4320 12256 4324
rect 19285 4380 19349 4384
rect 19285 4324 19289 4380
rect 19289 4324 19345 4380
rect 19345 4324 19349 4380
rect 19285 4320 19349 4324
rect 19365 4380 19429 4384
rect 19365 4324 19369 4380
rect 19369 4324 19425 4380
rect 19425 4324 19429 4380
rect 19365 4320 19429 4324
rect 19445 4380 19509 4384
rect 19445 4324 19449 4380
rect 19449 4324 19505 4380
rect 19505 4324 19509 4380
rect 19445 4320 19509 4324
rect 19525 4380 19589 4384
rect 19525 4324 19529 4380
rect 19529 4324 19585 4380
rect 19585 4324 19589 4380
rect 19525 4320 19589 4324
rect 8285 3836 8349 3840
rect 8285 3780 8289 3836
rect 8289 3780 8345 3836
rect 8345 3780 8349 3836
rect 8285 3776 8349 3780
rect 8365 3836 8429 3840
rect 8365 3780 8369 3836
rect 8369 3780 8425 3836
rect 8425 3780 8429 3836
rect 8365 3776 8429 3780
rect 8445 3836 8509 3840
rect 8445 3780 8449 3836
rect 8449 3780 8505 3836
rect 8505 3780 8509 3836
rect 8445 3776 8509 3780
rect 8525 3836 8589 3840
rect 8525 3780 8529 3836
rect 8529 3780 8585 3836
rect 8585 3780 8589 3836
rect 8525 3776 8589 3780
rect 15618 3836 15682 3840
rect 15618 3780 15622 3836
rect 15622 3780 15678 3836
rect 15678 3780 15682 3836
rect 15618 3776 15682 3780
rect 15698 3836 15762 3840
rect 15698 3780 15702 3836
rect 15702 3780 15758 3836
rect 15758 3780 15762 3836
rect 15698 3776 15762 3780
rect 15778 3836 15842 3840
rect 15778 3780 15782 3836
rect 15782 3780 15838 3836
rect 15838 3780 15842 3836
rect 15778 3776 15842 3780
rect 15858 3836 15922 3840
rect 15858 3780 15862 3836
rect 15862 3780 15918 3836
rect 15918 3780 15922 3836
rect 15858 3776 15922 3780
rect 4618 3292 4682 3296
rect 4618 3236 4622 3292
rect 4622 3236 4678 3292
rect 4678 3236 4682 3292
rect 4618 3232 4682 3236
rect 4698 3292 4762 3296
rect 4698 3236 4702 3292
rect 4702 3236 4758 3292
rect 4758 3236 4762 3292
rect 4698 3232 4762 3236
rect 4778 3292 4842 3296
rect 4778 3236 4782 3292
rect 4782 3236 4838 3292
rect 4838 3236 4842 3292
rect 4778 3232 4842 3236
rect 4858 3292 4922 3296
rect 4858 3236 4862 3292
rect 4862 3236 4918 3292
rect 4918 3236 4922 3292
rect 4858 3232 4922 3236
rect 11952 3292 12016 3296
rect 11952 3236 11956 3292
rect 11956 3236 12012 3292
rect 12012 3236 12016 3292
rect 11952 3232 12016 3236
rect 12032 3292 12096 3296
rect 12032 3236 12036 3292
rect 12036 3236 12092 3292
rect 12092 3236 12096 3292
rect 12032 3232 12096 3236
rect 12112 3292 12176 3296
rect 12112 3236 12116 3292
rect 12116 3236 12172 3292
rect 12172 3236 12176 3292
rect 12112 3232 12176 3236
rect 12192 3292 12256 3296
rect 12192 3236 12196 3292
rect 12196 3236 12252 3292
rect 12252 3236 12256 3292
rect 12192 3232 12256 3236
rect 19285 3292 19349 3296
rect 19285 3236 19289 3292
rect 19289 3236 19345 3292
rect 19345 3236 19349 3292
rect 19285 3232 19349 3236
rect 19365 3292 19429 3296
rect 19365 3236 19369 3292
rect 19369 3236 19425 3292
rect 19425 3236 19429 3292
rect 19365 3232 19429 3236
rect 19445 3292 19509 3296
rect 19445 3236 19449 3292
rect 19449 3236 19505 3292
rect 19505 3236 19509 3292
rect 19445 3232 19509 3236
rect 19525 3292 19589 3296
rect 19525 3236 19529 3292
rect 19529 3236 19585 3292
rect 19585 3236 19589 3292
rect 19525 3232 19589 3236
rect 8285 2748 8349 2752
rect 8285 2692 8289 2748
rect 8289 2692 8345 2748
rect 8345 2692 8349 2748
rect 8285 2688 8349 2692
rect 8365 2748 8429 2752
rect 8365 2692 8369 2748
rect 8369 2692 8425 2748
rect 8425 2692 8429 2748
rect 8365 2688 8429 2692
rect 8445 2748 8509 2752
rect 8445 2692 8449 2748
rect 8449 2692 8505 2748
rect 8505 2692 8509 2748
rect 8445 2688 8509 2692
rect 8525 2748 8589 2752
rect 8525 2692 8529 2748
rect 8529 2692 8585 2748
rect 8585 2692 8589 2748
rect 8525 2688 8589 2692
rect 15618 2748 15682 2752
rect 15618 2692 15622 2748
rect 15622 2692 15678 2748
rect 15678 2692 15682 2748
rect 15618 2688 15682 2692
rect 15698 2748 15762 2752
rect 15698 2692 15702 2748
rect 15702 2692 15758 2748
rect 15758 2692 15762 2748
rect 15698 2688 15762 2692
rect 15778 2748 15842 2752
rect 15778 2692 15782 2748
rect 15782 2692 15838 2748
rect 15838 2692 15842 2748
rect 15778 2688 15842 2692
rect 15858 2748 15922 2752
rect 15858 2692 15862 2748
rect 15862 2692 15918 2748
rect 15918 2692 15922 2748
rect 15858 2688 15922 2692
rect 18276 2620 18340 2684
rect 4618 2204 4682 2208
rect 4618 2148 4622 2204
rect 4622 2148 4678 2204
rect 4678 2148 4682 2204
rect 4618 2144 4682 2148
rect 4698 2204 4762 2208
rect 4698 2148 4702 2204
rect 4702 2148 4758 2204
rect 4758 2148 4762 2204
rect 4698 2144 4762 2148
rect 4778 2204 4842 2208
rect 4778 2148 4782 2204
rect 4782 2148 4838 2204
rect 4838 2148 4842 2204
rect 4778 2144 4842 2148
rect 4858 2204 4922 2208
rect 4858 2148 4862 2204
rect 4862 2148 4918 2204
rect 4918 2148 4922 2204
rect 4858 2144 4922 2148
rect 11952 2204 12016 2208
rect 11952 2148 11956 2204
rect 11956 2148 12012 2204
rect 12012 2148 12016 2204
rect 11952 2144 12016 2148
rect 12032 2204 12096 2208
rect 12032 2148 12036 2204
rect 12036 2148 12092 2204
rect 12092 2148 12096 2204
rect 12032 2144 12096 2148
rect 12112 2204 12176 2208
rect 12112 2148 12116 2204
rect 12116 2148 12172 2204
rect 12172 2148 12176 2204
rect 12112 2144 12176 2148
rect 12192 2204 12256 2208
rect 12192 2148 12196 2204
rect 12196 2148 12252 2204
rect 12252 2148 12256 2204
rect 12192 2144 12256 2148
rect 19285 2204 19349 2208
rect 19285 2148 19289 2204
rect 19289 2148 19345 2204
rect 19345 2148 19349 2204
rect 19285 2144 19349 2148
rect 19365 2204 19429 2208
rect 19365 2148 19369 2204
rect 19369 2148 19425 2204
rect 19425 2148 19429 2204
rect 19365 2144 19429 2148
rect 19445 2204 19509 2208
rect 19445 2148 19449 2204
rect 19449 2148 19505 2204
rect 19505 2148 19509 2204
rect 19445 2144 19509 2148
rect 19525 2204 19589 2208
rect 19525 2148 19529 2204
rect 19529 2148 19585 2204
rect 19585 2148 19589 2204
rect 19525 2144 19589 2148
rect 60 1668 124 1732
rect 6132 36 6196 100
<< metal4 >>
rect 4610 19616 4931 19632
rect 4610 19552 4618 19616
rect 4682 19552 4698 19616
rect 4762 19552 4778 19616
rect 4842 19552 4858 19616
rect 4922 19552 4931 19616
rect 4610 18528 4931 19552
rect 4610 18464 4618 18528
rect 4682 18464 4698 18528
rect 4762 18464 4778 18528
rect 4842 18464 4858 18528
rect 4922 18464 4931 18528
rect 4610 17440 4931 18464
rect 4610 17376 4618 17440
rect 4682 17376 4698 17440
rect 4762 17376 4778 17440
rect 4842 17376 4858 17440
rect 4922 17376 4931 17440
rect 4610 16352 4931 17376
rect 8277 19072 8597 19632
rect 8277 19008 8285 19072
rect 8349 19008 8365 19072
rect 8429 19008 8445 19072
rect 8509 19008 8525 19072
rect 8589 19008 8597 19072
rect 8277 17984 8597 19008
rect 8277 17920 8285 17984
rect 8349 17920 8365 17984
rect 8429 17920 8445 17984
rect 8509 17920 8525 17984
rect 8589 17920 8597 17984
rect 8277 16896 8597 17920
rect 11944 19616 12264 19632
rect 11944 19552 11952 19616
rect 12016 19552 12032 19616
rect 12096 19552 12112 19616
rect 12176 19552 12192 19616
rect 12256 19552 12264 19616
rect 11944 18528 12264 19552
rect 11944 18464 11952 18528
rect 12016 18464 12032 18528
rect 12096 18464 12112 18528
rect 12176 18464 12192 18528
rect 12256 18464 12264 18528
rect 11944 17440 12264 18464
rect 11944 17376 11952 17440
rect 12016 17376 12032 17440
rect 12096 17376 12112 17440
rect 12176 17376 12192 17440
rect 12256 17376 12264 17440
rect 10547 16964 10613 16965
rect 10547 16900 10548 16964
rect 10612 16900 10613 16964
rect 10547 16899 10613 16900
rect 8277 16832 8285 16896
rect 8349 16832 8365 16896
rect 8429 16832 8445 16896
rect 8509 16832 8525 16896
rect 8589 16832 8597 16896
rect 5947 16692 6013 16693
rect 5947 16628 5948 16692
rect 6012 16628 6013 16692
rect 5947 16627 6013 16628
rect 4610 16288 4618 16352
rect 4682 16288 4698 16352
rect 4762 16288 4778 16352
rect 4842 16288 4858 16352
rect 4922 16288 4931 16352
rect 4610 15264 4931 16288
rect 4610 15200 4618 15264
rect 4682 15200 4698 15264
rect 4762 15200 4778 15264
rect 4842 15200 4858 15264
rect 4922 15200 4931 15264
rect 4610 14176 4931 15200
rect 4610 14112 4618 14176
rect 4682 14112 4698 14176
rect 4762 14112 4778 14176
rect 4842 14112 4858 14176
rect 4922 14112 4931 14176
rect 59 13836 125 13837
rect 59 13772 60 13836
rect 124 13834 125 13836
rect 124 13774 306 13834
rect 124 13772 125 13774
rect 59 13771 125 13772
rect 246 12698 306 13774
rect 4610 13088 4931 14112
rect 4610 13024 4618 13088
rect 4682 13024 4698 13088
rect 4762 13024 4778 13088
rect 4842 13024 4858 13088
rect 4922 13024 4931 13088
rect 4610 12000 4931 13024
rect 4610 11936 4618 12000
rect 4682 11936 4698 12000
rect 4762 11936 4778 12000
rect 4842 11936 4858 12000
rect 4922 11936 4931 12000
rect 4610 10912 4931 11936
rect 5950 11933 6010 16627
rect 8277 15808 8597 16832
rect 8277 15744 8285 15808
rect 8349 15744 8365 15808
rect 8429 15744 8445 15808
rect 8509 15744 8525 15808
rect 8589 15744 8597 15808
rect 6131 15332 6197 15333
rect 6131 15268 6132 15332
rect 6196 15268 6197 15332
rect 6131 15267 6197 15268
rect 5947 11932 6013 11933
rect 5947 11868 5948 11932
rect 6012 11868 6013 11932
rect 5947 11867 6013 11868
rect 4610 10848 4618 10912
rect 4682 10848 4698 10912
rect 4762 10848 4778 10912
rect 4842 10848 4858 10912
rect 4922 10848 4931 10912
rect 4610 9824 4931 10848
rect 4610 9760 4618 9824
rect 4682 9760 4698 9824
rect 4762 9760 4778 9824
rect 4842 9760 4858 9824
rect 4922 9760 4931 9824
rect 4610 8736 4931 9760
rect 4610 8672 4618 8736
rect 4682 8672 4698 8736
rect 4762 8672 4778 8736
rect 4842 8672 4858 8736
rect 4922 8672 4931 8736
rect 4610 7648 4931 8672
rect 4610 7584 4618 7648
rect 4682 7584 4698 7648
rect 4762 7584 4778 7648
rect 4842 7584 4858 7648
rect 4922 7584 4931 7648
rect 4610 6560 4931 7584
rect 4610 6496 4618 6560
rect 4682 6496 4698 6560
rect 4762 6496 4778 6560
rect 4842 6496 4858 6560
rect 4922 6496 4931 6560
rect 4610 5472 4931 6496
rect 4610 5408 4618 5472
rect 4682 5408 4698 5472
rect 4762 5408 4778 5472
rect 4842 5408 4858 5472
rect 4922 5408 4931 5472
rect 59 5268 125 5269
rect 59 5204 60 5268
rect 124 5204 125 5268
rect 59 5203 125 5204
rect 62 1733 122 5203
rect 4610 4384 4931 5408
rect 4610 4320 4618 4384
rect 4682 4320 4698 4384
rect 4762 4320 4778 4384
rect 4842 4320 4858 4384
rect 4922 4320 4931 4384
rect 4610 3296 4931 4320
rect 4610 3232 4618 3296
rect 4682 3232 4698 3296
rect 4762 3232 4778 3296
rect 4842 3232 4858 3296
rect 4922 3232 4931 3296
rect 4610 2208 4931 3232
rect 4610 2144 4618 2208
rect 4682 2144 4698 2208
rect 4762 2144 4778 2208
rect 4842 2144 4858 2208
rect 4922 2144 4931 2208
rect 4610 2128 4931 2144
rect 59 1732 125 1733
rect 59 1668 60 1732
rect 124 1668 125 1732
rect 59 1667 125 1668
rect 6134 101 6194 15267
rect 8277 14720 8597 15744
rect 8277 14656 8285 14720
rect 8349 14656 8365 14720
rect 8429 14656 8445 14720
rect 8509 14656 8525 14720
rect 8589 14656 8597 14720
rect 8277 13632 8597 14656
rect 9627 14108 9693 14109
rect 9627 14044 9628 14108
rect 9692 14044 9693 14108
rect 9627 14043 9693 14044
rect 9075 13972 9141 13973
rect 9075 13908 9076 13972
rect 9140 13908 9141 13972
rect 9075 13907 9141 13908
rect 8277 13568 8285 13632
rect 8349 13568 8365 13632
rect 8429 13568 8445 13632
rect 8509 13568 8525 13632
rect 8589 13568 8597 13632
rect 8277 12544 8597 13568
rect 8277 12480 8285 12544
rect 8349 12480 8365 12544
rect 8429 12480 8445 12544
rect 8509 12480 8525 12544
rect 8589 12480 8597 12544
rect 8277 11456 8597 12480
rect 8277 11392 8285 11456
rect 8349 11392 8365 11456
rect 8429 11392 8445 11456
rect 8509 11392 8525 11456
rect 8589 11392 8597 11456
rect 8277 10368 8597 11392
rect 8277 10304 8285 10368
rect 8349 10304 8365 10368
rect 8429 10304 8445 10368
rect 8509 10304 8525 10368
rect 8589 10304 8597 10368
rect 8277 9280 8597 10304
rect 8277 9216 8285 9280
rect 8349 9216 8365 9280
rect 8429 9216 8445 9280
rect 8509 9216 8525 9280
rect 8589 9216 8597 9280
rect 8277 8192 8597 9216
rect 9078 8669 9138 13907
rect 9630 11525 9690 14043
rect 9627 11524 9693 11525
rect 9627 11460 9628 11524
rect 9692 11460 9693 11524
rect 9627 11459 9693 11460
rect 10550 9485 10610 16899
rect 11944 16352 12264 17376
rect 11944 16288 11952 16352
rect 12016 16288 12032 16352
rect 12096 16288 12112 16352
rect 12176 16288 12192 16352
rect 12256 16288 12264 16352
rect 11944 15264 12264 16288
rect 15610 19072 15930 19632
rect 15610 19008 15618 19072
rect 15682 19008 15698 19072
rect 15762 19008 15778 19072
rect 15842 19008 15858 19072
rect 15922 19008 15930 19072
rect 15610 17984 15930 19008
rect 15610 17920 15618 17984
rect 15682 17920 15698 17984
rect 15762 17920 15778 17984
rect 15842 17920 15858 17984
rect 15922 17920 15930 17984
rect 15610 16896 15930 17920
rect 15610 16832 15618 16896
rect 15682 16832 15698 16896
rect 15762 16832 15778 16896
rect 15842 16832 15858 16896
rect 15922 16832 15930 16896
rect 13491 15876 13557 15877
rect 13491 15812 13492 15876
rect 13556 15812 13557 15876
rect 13491 15811 13557 15812
rect 11944 15200 11952 15264
rect 12016 15200 12032 15264
rect 12096 15200 12112 15264
rect 12176 15200 12192 15264
rect 12256 15200 12264 15264
rect 11944 14176 12264 15200
rect 13494 14245 13554 15811
rect 15610 15808 15930 16832
rect 15610 15744 15618 15808
rect 15682 15744 15698 15808
rect 15762 15744 15778 15808
rect 15842 15744 15858 15808
rect 15922 15744 15930 15808
rect 15610 14720 15930 15744
rect 15610 14656 15618 14720
rect 15682 14656 15698 14720
rect 15762 14656 15778 14720
rect 15842 14656 15858 14720
rect 15922 14656 15930 14720
rect 13491 14244 13557 14245
rect 13491 14180 13492 14244
rect 13556 14180 13557 14244
rect 13491 14179 13557 14180
rect 11944 14112 11952 14176
rect 12016 14112 12032 14176
rect 12096 14112 12112 14176
rect 12176 14112 12192 14176
rect 12256 14112 12264 14176
rect 11944 13088 12264 14112
rect 15610 13632 15930 14656
rect 15610 13568 15618 13632
rect 15682 13568 15698 13632
rect 15762 13568 15778 13632
rect 15842 13568 15858 13632
rect 15922 13568 15930 13632
rect 14595 13564 14661 13565
rect 14595 13500 14596 13564
rect 14660 13500 14661 13564
rect 14595 13499 14661 13500
rect 14598 13378 14658 13499
rect 11944 13024 11952 13088
rect 12016 13024 12032 13088
rect 12096 13024 12112 13088
rect 12176 13024 12192 13088
rect 12256 13024 12264 13088
rect 11944 12000 12264 13024
rect 11944 11936 11952 12000
rect 12016 11936 12032 12000
rect 12096 11936 12112 12000
rect 12176 11936 12192 12000
rect 12256 11936 12264 12000
rect 11944 10912 12264 11936
rect 11944 10848 11952 10912
rect 12016 10848 12032 10912
rect 12096 10848 12112 10912
rect 12176 10848 12192 10912
rect 12256 10848 12264 10912
rect 11944 9824 12264 10848
rect 11944 9760 11952 9824
rect 12016 9760 12032 9824
rect 12096 9760 12112 9824
rect 12176 9760 12192 9824
rect 12256 9760 12264 9824
rect 10547 9484 10613 9485
rect 10547 9420 10548 9484
rect 10612 9420 10613 9484
rect 10547 9419 10613 9420
rect 11944 8736 12264 9760
rect 11944 8672 11952 8736
rect 12016 8672 12032 8736
rect 12096 8672 12112 8736
rect 12176 8672 12192 8736
rect 12256 8672 12264 8736
rect 9075 8668 9141 8669
rect 9075 8604 9076 8668
rect 9140 8604 9141 8668
rect 9075 8603 9141 8604
rect 8277 8128 8285 8192
rect 8349 8128 8365 8192
rect 8429 8128 8445 8192
rect 8509 8128 8525 8192
rect 8589 8128 8597 8192
rect 8277 7104 8597 8128
rect 8277 7040 8285 7104
rect 8349 7040 8365 7104
rect 8429 7040 8445 7104
rect 8509 7040 8525 7104
rect 8589 7040 8597 7104
rect 8277 6016 8597 7040
rect 8277 5952 8285 6016
rect 8349 5952 8365 6016
rect 8429 5952 8445 6016
rect 8509 5952 8525 6016
rect 8589 5952 8597 6016
rect 8277 4928 8597 5952
rect 8277 4864 8285 4928
rect 8349 4864 8365 4928
rect 8429 4864 8445 4928
rect 8509 4864 8525 4928
rect 8589 4864 8597 4928
rect 8277 3840 8597 4864
rect 8277 3776 8285 3840
rect 8349 3776 8365 3840
rect 8429 3776 8445 3840
rect 8509 3776 8525 3840
rect 8589 3776 8597 3840
rect 8277 2752 8597 3776
rect 8277 2688 8285 2752
rect 8349 2688 8365 2752
rect 8429 2688 8445 2752
rect 8509 2688 8525 2752
rect 8589 2688 8597 2752
rect 8277 2128 8597 2688
rect 11944 7648 12264 8672
rect 11944 7584 11952 7648
rect 12016 7584 12032 7648
rect 12096 7584 12112 7648
rect 12176 7584 12192 7648
rect 12256 7584 12264 7648
rect 11944 6560 12264 7584
rect 11944 6496 11952 6560
rect 12016 6496 12032 6560
rect 12096 6496 12112 6560
rect 12176 6496 12192 6560
rect 12256 6496 12264 6560
rect 11944 5472 12264 6496
rect 11944 5408 11952 5472
rect 12016 5408 12032 5472
rect 12096 5408 12112 5472
rect 12176 5408 12192 5472
rect 12256 5408 12264 5472
rect 11944 4384 12264 5408
rect 11944 4320 11952 4384
rect 12016 4320 12032 4384
rect 12096 4320 12112 4384
rect 12176 4320 12192 4384
rect 12256 4320 12264 4384
rect 11944 3296 12264 4320
rect 11944 3232 11952 3296
rect 12016 3232 12032 3296
rect 12096 3232 12112 3296
rect 12176 3232 12192 3296
rect 12256 3232 12264 3296
rect 11944 2208 12264 3232
rect 11944 2144 11952 2208
rect 12016 2144 12032 2208
rect 12096 2144 12112 2208
rect 12176 2144 12192 2208
rect 12256 2144 12264 2208
rect 11944 2128 12264 2144
rect 15610 12544 15930 13568
rect 15610 12480 15618 12544
rect 15682 12480 15698 12544
rect 15762 12480 15778 12544
rect 15842 12480 15858 12544
rect 15922 12480 15930 12544
rect 15610 11456 15930 12480
rect 15610 11392 15618 11456
rect 15682 11392 15698 11456
rect 15762 11392 15778 11456
rect 15842 11392 15858 11456
rect 15922 11392 15930 11456
rect 15610 10368 15930 11392
rect 15610 10304 15618 10368
rect 15682 10304 15698 10368
rect 15762 10304 15778 10368
rect 15842 10304 15858 10368
rect 15922 10304 15930 10368
rect 15610 9280 15930 10304
rect 15610 9216 15618 9280
rect 15682 9216 15698 9280
rect 15762 9216 15778 9280
rect 15842 9216 15858 9280
rect 15922 9216 15930 9280
rect 15610 8192 15930 9216
rect 15610 8128 15618 8192
rect 15682 8128 15698 8192
rect 15762 8128 15778 8192
rect 15842 8128 15858 8192
rect 15922 8128 15930 8192
rect 15610 7104 15930 8128
rect 15610 7040 15618 7104
rect 15682 7040 15698 7104
rect 15762 7040 15778 7104
rect 15842 7040 15858 7104
rect 15922 7040 15930 7104
rect 15610 6016 15930 7040
rect 15610 5952 15618 6016
rect 15682 5952 15698 6016
rect 15762 5952 15778 6016
rect 15842 5952 15858 6016
rect 15922 5952 15930 6016
rect 15610 4928 15930 5952
rect 19277 19616 19597 19632
rect 19277 19552 19285 19616
rect 19349 19552 19365 19616
rect 19429 19552 19445 19616
rect 19509 19552 19525 19616
rect 19589 19552 19597 19616
rect 19277 18528 19597 19552
rect 19277 18464 19285 18528
rect 19349 18464 19365 18528
rect 19429 18464 19445 18528
rect 19509 18464 19525 18528
rect 19589 18464 19597 18528
rect 19277 17440 19597 18464
rect 19277 17376 19285 17440
rect 19349 17376 19365 17440
rect 19429 17376 19445 17440
rect 19509 17376 19525 17440
rect 19589 17376 19597 17440
rect 19277 16352 19597 17376
rect 19277 16288 19285 16352
rect 19349 16288 19365 16352
rect 19429 16288 19445 16352
rect 19509 16288 19525 16352
rect 19589 16288 19597 16352
rect 19277 15264 19597 16288
rect 19277 15200 19285 15264
rect 19349 15200 19365 15264
rect 19429 15200 19445 15264
rect 19509 15200 19525 15264
rect 19589 15200 19597 15264
rect 19277 14176 19597 15200
rect 19277 14112 19285 14176
rect 19349 14112 19365 14176
rect 19429 14112 19445 14176
rect 19509 14112 19525 14176
rect 19589 14112 19597 14176
rect 19277 13088 19597 14112
rect 19277 13024 19285 13088
rect 19349 13024 19365 13088
rect 19429 13024 19445 13088
rect 19509 13024 19525 13088
rect 19589 13024 19597 13088
rect 19277 12000 19597 13024
rect 19277 11936 19285 12000
rect 19349 11936 19365 12000
rect 19429 11936 19445 12000
rect 19509 11936 19525 12000
rect 19589 11936 19597 12000
rect 19277 10912 19597 11936
rect 19277 10848 19285 10912
rect 19349 10848 19365 10912
rect 19429 10848 19445 10912
rect 19509 10848 19525 10912
rect 19589 10848 19597 10912
rect 19277 9824 19597 10848
rect 19277 9760 19285 9824
rect 19349 9760 19365 9824
rect 19429 9760 19445 9824
rect 19509 9760 19525 9824
rect 19589 9760 19597 9824
rect 19277 8736 19597 9760
rect 19277 8672 19285 8736
rect 19349 8672 19365 8736
rect 19429 8672 19445 8736
rect 19509 8672 19525 8736
rect 19589 8672 19597 8736
rect 19277 7648 19597 8672
rect 19277 7584 19285 7648
rect 19349 7584 19365 7648
rect 19429 7584 19445 7648
rect 19509 7584 19525 7648
rect 19589 7584 19597 7648
rect 19277 6560 19597 7584
rect 19277 6496 19285 6560
rect 19349 6496 19365 6560
rect 19429 6496 19445 6560
rect 19509 6496 19525 6560
rect 19589 6496 19597 6560
rect 19277 5472 19597 6496
rect 19277 5408 19285 5472
rect 19349 5408 19365 5472
rect 19429 5408 19445 5472
rect 19509 5408 19525 5472
rect 19589 5408 19597 5472
rect 18275 5268 18341 5269
rect 18275 5204 18276 5268
rect 18340 5204 18341 5268
rect 18275 5203 18341 5204
rect 15610 4864 15618 4928
rect 15682 4864 15698 4928
rect 15762 4864 15778 4928
rect 15842 4864 15858 4928
rect 15922 4864 15930 4928
rect 15610 3840 15930 4864
rect 15610 3776 15618 3840
rect 15682 3776 15698 3840
rect 15762 3776 15778 3840
rect 15842 3776 15858 3840
rect 15922 3776 15930 3840
rect 15610 2752 15930 3776
rect 15610 2688 15618 2752
rect 15682 2688 15698 2752
rect 15762 2688 15778 2752
rect 15842 2688 15858 2752
rect 15922 2688 15930 2752
rect 15610 2128 15930 2688
rect 18278 2685 18338 5203
rect 19277 4384 19597 5408
rect 19277 4320 19285 4384
rect 19349 4320 19365 4384
rect 19429 4320 19445 4384
rect 19509 4320 19525 4384
rect 19589 4320 19597 4384
rect 19277 3296 19597 4320
rect 19277 3232 19285 3296
rect 19349 3232 19365 3296
rect 19429 3232 19445 3296
rect 19509 3232 19525 3296
rect 19589 3232 19597 3296
rect 18275 2684 18341 2685
rect 18275 2620 18276 2684
rect 18340 2620 18341 2684
rect 18275 2619 18341 2620
rect 19277 2208 19597 3232
rect 19277 2144 19285 2208
rect 19349 2144 19365 2208
rect 19429 2144 19445 2208
rect 19509 2144 19525 2208
rect 19589 2144 19597 2208
rect 19277 2128 19597 2144
rect 6131 100 6197 101
rect 6131 36 6132 100
rect 6196 36 6197 100
rect 6131 35 6197 36
<< via4 >>
rect 158 12462 394 12698
rect 14510 13142 14746 13378
<< metal5 >>
rect 9500 13378 14788 13420
rect 9500 13142 14510 13378
rect 14746 13142 14788 13378
rect 9500 13100 14788 13142
rect 9500 12740 9820 13100
rect 116 12698 9820 12740
rect 116 12462 158 12698
rect 394 12462 9820 12698
rect 116 12420 9820 12462
use scs8hd_fill_1  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_6 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_conb_1  _133_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_17
timestamp 1586364061
transform 1 0 2668 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_13
timestamp 1586364061
transform 1 0 2300 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_10
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__B
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 222 592
use scs8hd_nor2_4  _093_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use scs8hd_nor2_4  _067_
timestamp 1586364061
transform 1 0 1472 0 1 2720
box -38 -48 866 592
use scs8hd_decap_4  FILLER_1_21 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3036 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 2852 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__B
timestamp 1586364061
transform 1 0 3404 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_35
timestamp 1586364061
transform 1 0 4324 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_29
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_64 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use scs8hd_nor2_4  _092_
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_40
timestamp 1586364061
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_36
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_39
timestamp 1586364061
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4508 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5152 0 1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_5_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_70
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_65
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_71
timestamp 1586364061
transform 1 0 7636 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_70
timestamp 1586364061
transform 1 0 7544 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_66
timestamp 1586364061
transform 1 0 7176 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7360 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 866 592
use scs8hd_decap_4  FILLER_1_77
timestamp 1586364061
transform 1 0 8188 0 1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_81
timestamp 1586364061
transform 1 0 8556 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8648 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8832 0 1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_6.LATCH_5_.latch
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_1_97
timestamp 1586364061
transform 1 0 10028 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_93
timestamp 1586364061
transform 1 0 9660 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_98
timestamp 1586364061
transform 1 0 10120 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__B
timestamp 1586364061
transform 1 0 9936 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__A
timestamp 1586364061
transform 1 0 9844 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_66
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 10304 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 10304 0 -1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_6.LATCH_4_.latch
timestamp 1586364061
transform 1 0 10488 0 -1 2720
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_6.LATCH_3_.latch
timestamp 1586364061
transform 1 0 10488 0 1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_113
timestamp 1586364061
transform 1 0 11500 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_113
timestamp 1586364061
transform 1 0 11500 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11684 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11684 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_121
timestamp 1586364061
transform 1 0 12236 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_117
timestamp 1586364061
transform 1 0 11868 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_121
timestamp 1586364061
transform 1 0 12236 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_117
timestamp 1586364061
transform 1 0 11868 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12052 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_71
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_67
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _148_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_131
timestamp 1586364061
transform 1 0 13156 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_127
timestamp 1586364061
transform 1 0 12788 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_129
timestamp 1586364061
transform 1 0 12972 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12788 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 13340 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 13156 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 12972 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 13708 0 1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_5.LATCH_5_.latch
timestamp 1586364061
transform 1 0 13340 0 -1 2720
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_5.LATCH_4_.latch
timestamp 1586364061
transform 1 0 13892 0 1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_150
timestamp 1586364061
transform 1 0 14904 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_148
timestamp 1586364061
transform 1 0 14720 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_144
timestamp 1586364061
transform 1 0 14352 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14536 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_154
timestamp 1586364061
transform 1 0 15272 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_152
timestamp 1586364061
transform 1 0 15088 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15088 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15456 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_68
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15640 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_0_165
timestamp 1586364061
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_167
timestamp 1586364061
transform 1 0 16468 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_169
timestamp 1586364061
transform 1 0 16652 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_173
timestamp 1586364061
transform 1 0 17020 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_173
timestamp 1586364061
transform 1 0 17020 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _149_
timestamp 1586364061
transform 1 0 17112 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_1_177
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_178
timestamp 1586364061
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__053__A
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__055__A
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_72
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_69
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_193
timestamp 1586364061
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_196
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__057__A
timestamp 1586364061
transform 1 0 19044 0 1 2720
box -38 -48 222 592
use scs8hd_nor2_4  _055_
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use scs8hd_nor2_4  _053_
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_204
timestamp 1586364061
transform 1 0 19872 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_197
timestamp 1586364061
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__057__B
timestamp 1586364061
transform 1 0 19412 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__053__B
timestamp 1586364061
transform 1 0 19320 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_5.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 20884 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 20884 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_200 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 1142 592
use scs8hd_nor2_4  _094_
timestamp 1586364061
transform 1 0 2392 0 -1 3808
box -38 -48 866 592
use scs8hd_conb_1  _134_
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 1840 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__B
timestamp 1586364061
transform 1 0 2208 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_6
timestamp 1586364061
transform 1 0 1656 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_10
timestamp 1586364061
transform 1 0 2024 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 5888 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5244 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5704 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_43
timestamp 1586364061
transform 1 0 5060 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_47
timestamp 1586364061
transform 1 0 5428 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_63
timestamp 1586364061
transform 1 0 6900 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_67
timestamp 1586364061
transform 1 0 7268 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_71
timestamp 1586364061
transform 1 0 7636 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _059_
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_102
timestamp 1586364061
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_106
timestamp 1586364061
transform 1 0 10856 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11040 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_110
timestamp 1586364061
transform 1 0 11224 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_121
timestamp 1586364061
transform 1 0 12236 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_5.LATCH_3_.latch
timestamp 1586364061
transform 1 0 13248 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13064 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_125
timestamp 1586364061
transform 1 0 12604 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_143
timestamp 1586364061
transform 1 0 14260 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_149
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _085_
timestamp 1586364061
transform 1 0 16836 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_163
timestamp 1586364061
transform 1 0 16100 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_2_168
timestamp 1586364061
transform 1 0 16560 0 -1 3808
box -38 -48 314 592
use scs8hd_nor2_4  _057_
timestamp 1586364061
transform 1 0 18400 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__055__B
timestamp 1586364061
transform 1 0 18032 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_180
timestamp 1586364061
transform 1 0 17664 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_186
timestamp 1586364061
transform 1 0 18216 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 20884 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_197
timestamp 1586364061
transform 1 0 19228 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_2_209
timestamp 1586364061
transform 1 0 20332 0 -1 3808
box -38 -48 314 592
use scs8hd_nor2_4  _063_
timestamp 1586364061
transform 1 0 2208 0 1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__063__A
timestamp 1586364061
transform 1 0 2024 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__065__B
timestamp 1586364061
transform 1 0 1656 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_8
timestamp 1586364061
transform 1 0 1840 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3772 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 3220 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_21
timestamp 1586364061
transform 1 0 3036 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_25
timestamp 1586364061
transform 1 0 3404 0 1 3808
box -38 -48 222 592
use scs8hd_or2_4  _083_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5336 0 1 3808
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_38
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_42
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__083__B
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8556 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_73
timestamp 1586364061
transform 1 0 7820 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_77
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10488 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10304 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__B
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_92
timestamp 1586364061
transform 1 0 9568 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_3_97
timestamp 1586364061
transform 1 0 10028 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11684 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_113
timestamp 1586364061
transform 1 0 11500 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_117
timestamp 1586364061
transform 1 0 11868 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_132
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_136
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_140
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14444 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_144
timestamp 1586364061
transform 1 0 14352 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_158
timestamp 1586364061
transform 1 0 15640 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__089__B
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 16192 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_162
timestamp 1586364061
transform 1 0 16008 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_175
timestamp 1586364061
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _096_
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__044__A
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__B
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_179
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_193
timestamp 1586364061
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 20884 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_197
timestamp 1586364061
transform 1 0 19228 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_204
timestamp 1586364061
transform 1 0 19872 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 406 592
use scs8hd_nor2_4  _065_
timestamp 1586364061
transform 1 0 2392 0 -1 4896
box -38 -48 866 592
use scs8hd_conb_1  _137_
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 1840 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__063__B
timestamp 1586364061
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_6
timestamp 1586364061
transform 1 0 1656 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_10
timestamp 1586364061
transform 1 0 2024 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4140 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5888 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_42 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4968 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_50
timestamp 1586364061
transform 1 0 5704 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6440 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7452 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_54
timestamp 1586364061
transform 1 0 6072 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_67
timestamp 1586364061
transform 1 0 7268 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_71
timestamp 1586364061
transform 1 0 7636 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7820 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_88
timestamp 1586364061
transform 1 0 9200 0 -1 4896
box -38 -48 406 592
use scs8hd_nor2_4  _087_
timestamp 1586364061
transform 1 0 9844 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 10856 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_104
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_108
timestamp 1586364061
transform 1 0 11040 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_121
timestamp 1586364061
transform 1 0 12236 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13984 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_125
timestamp 1586364061
transform 1 0 12604 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_138
timestamp 1586364061
transform 1 0 13800 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_142
timestamp 1586364061
transform 1 0 14168 0 -1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_146
timestamp 1586364061
transform 1 0 14536 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_149
timestamp 1586364061
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _089_
timestamp 1586364061
transform 1 0 16836 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16284 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16652 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_163
timestamp 1586364061
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_167
timestamp 1586364061
transform 1 0 16468 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_8  _044_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 18400 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_180
timestamp 1586364061
transform 1 0 17664 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_186
timestamp 1586364061
transform 1 0 18216 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 20884 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_197
timestamp 1586364061
transform 1 0 19228 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_4_209
timestamp 1586364061
transform 1 0 20332 0 -1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1656 0 1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2668 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 3772 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3036 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_19
timestamp 1586364061
transform 1 0 2852 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_23
timestamp 1586364061
transform 1 0 3220 0 1 4896
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_6.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5520 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_40
timestamp 1586364061
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_44
timestamp 1586364061
transform 1 0 5152 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_71
timestamp 1586364061
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8464 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8280 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_75
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_5_89
timestamp 1586364061
transform 1 0 9292 0 1 4896
box -38 -48 406 592
use scs8hd_nor2_4  _086_
timestamp 1586364061
transform 1 0 10764 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 10028 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9660 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_95
timestamp 1586364061
transform 1 0 9844 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_99
timestamp 1586364061
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_103
timestamp 1586364061
transform 1 0 10580 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13984 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 13800 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_132
timestamp 1586364061
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_136
timestamp 1586364061
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_151
timestamp 1586364061
transform 1 0 14996 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_5_156
timestamp 1586364061
transform 1 0 15456 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_168
timestamp 1586364061
transform 1 0 16560 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_173
timestamp 1586364061
transform 1 0 17020 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_177
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 406 592
use scs8hd_inv_8  _045_
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__045__A
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_193
timestamp 1586364061
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_5.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 20884 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_197
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_204
timestamp 1586364061
transform 1 0 19872 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 866 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2576 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_14
timestamp 1586364061
transform 1 0 2392 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_16
timestamp 1586364061
transform 1 0 2576 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_24
timestamp 1586364061
transform 1 0 3312 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_20
timestamp 1586364061
transform 1 0 2944 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_22
timestamp 1586364061
transform 1 0 3128 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_18
timestamp 1586364061
transform 1 0 2760 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2944 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3496 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__064__B
timestamp 1586364061
transform 1 0 3128 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__064__A
timestamp 1586364061
transform 1 0 2760 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_28
timestamp 1586364061
transform 1 0 3680 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3864 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_7_41
timestamp 1586364061
transform 1 0 4876 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_6_43
timestamp 1586364061
transform 1 0 5060 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__062__C
timestamp 1586364061
transform 1 0 5152 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_46
timestamp 1586364061
transform 1 0 5336 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_49
timestamp 1586364061
transform 1 0 5612 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5428 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5796 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__B
timestamp 1586364061
transform 1 0 5520 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_6.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 5984
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 5980 0 -1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__062__A
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__061__B
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_64
timestamp 1586364061
transform 1 0 6992 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_6_70
timestamp 1586364061
transform 1 0 7544 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_71
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__084__C
timestamp 1586364061
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__061__A
timestamp 1586364061
transform 1 0 8188 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_88
timestamp 1586364061
transform 1 0 9200 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_75
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_79
timestamp 1586364061
transform 1 0 8372 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_95
timestamp 1586364061
transform 1 0 9844 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_7_90
timestamp 1586364061
transform 1 0 9384 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_97
timestamp 1586364061
transform 1 0 10028 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10212 0 -1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_6.LATCH_2_.latch
timestamp 1586364061
transform 1 0 10304 0 1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10396 0 -1 5984
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_7_111
timestamp 1586364061
transform 1 0 11316 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_112
timestamp 1586364061
transform 1 0 11408 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_116
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_6_116
timestamp 1586364061
transform 1 0 11776 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12144 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use scs8hd_buf_2  _154_
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_5.LATCH_2_.latch
timestamp 1586364061
transform 1 0 14076 0 1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 13892 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13340 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_6  FILLER_6_135 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13524 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_132
timestamp 1586364061
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_136
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 15272 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15640 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_152
timestamp 1586364061
transform 1 0 15088 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_156
timestamp 1586364061
transform 1 0 15456 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16836 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_163
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_169
timestamp 1586364061
transform 1 0 16652 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_169
timestamp 1586364061
transform 1 0 16652 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_173
timestamp 1586364061
transform 1 0 17020 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_186
timestamp 1586364061
transform 1 0 18216 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_180
timestamp 1586364061
transform 1 0 17664 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 18032 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__B
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_193
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _095_
timestamp 1586364061
transform 1 0 18400 0 -1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _090_
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_204
timestamp 1586364061
transform 1 0 19872 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_197
timestamp 1586364061
transform 1 0 19228 0 1 5984
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_209
timestamp 1586364061
transform 1 0 20332 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20424 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 20884 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 20884 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_197
timestamp 1586364061
transform 1 0 19228 0 -1 5984
box -38 -48 1142 592
use scs8hd_nor2_4  _064_
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 866 592
use scs8hd_conb_1  _135_
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 1840 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2208 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_6
timestamp 1586364061
transform 1 0 1656 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_10
timestamp 1586364061
transform 1 0 2024 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 590 592
use scs8hd_or3_4  _062_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5612 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__049__B
timestamp 1586364061
transform 1 0 5336 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_41
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_45
timestamp 1586364061
transform 1 0 5244 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_48
timestamp 1586364061
transform 1 0 5520 0 -1 7072
box -38 -48 130 592
use scs8hd_nor2_4  _061_
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__091__D
timestamp 1586364061
transform 1 0 7176 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__C
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_58
timestamp 1586364061
transform 1 0 6440 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_64
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__B
timestamp 1586364061
transform 1 0 8372 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9292 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_77
timestamp 1586364061
transform 1 0 8188 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_81
timestamp 1586364061
transform 1 0 8556 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_87
timestamp 1586364061
transform 1 0 9108 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_91
timestamp 1586364061
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_107
timestamp 1586364061
transform 1 0 10948 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11592 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11132 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_111
timestamp 1586364061
transform 1 0 11316 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_123
timestamp 1586364061
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13340 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12604 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_127
timestamp 1586364061
transform 1 0 12788 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_131
timestamp 1586364061
transform 1 0 13156 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_142
timestamp 1586364061
transform 1 0 14168 0 -1 7072
box -38 -48 222 592
use scs8hd_buf_2  _142_
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15824 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14352 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_146
timestamp 1586364061
transform 1 0 14536 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_150
timestamp 1586364061
transform 1 0 14904 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_158
timestamp 1586364061
transform 1 0 15640 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16468 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16192 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_162
timestamp 1586364061
transform 1 0 16008 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_166
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_176
timestamp 1586364061
transform 1 0 17296 0 -1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _097_
timestamp 1586364061
transform 1 0 18032 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_4  FILLER_8_180
timestamp 1586364061
transform 1 0 17664 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_8  FILLER_8_193
timestamp 1586364061
transform 1 0 18860 0 -1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_5.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 20884 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_204
timestamp 1586364061
transform 1 0 19872 0 -1 7072
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2392 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_12
timestamp 1586364061
transform 1 0 2208 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_16
timestamp 1586364061
transform 1 0 2576 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 2944 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 4140 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2760 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_31
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_35
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__049__C
timestamp 1586364061
transform 1 0 5704 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_48
timestamp 1586364061
transform 1 0 5520 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_52
timestamp 1586364061
transform 1 0 5888 0 1 7072
box -38 -48 222 592
use scs8hd_or4_4  _084_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7360 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__084__B
timestamp 1586364061
transform 1 0 7176 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__049__A
timestamp 1586364061
transform 1 0 6072 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_56
timestamp 1586364061
transform 1 0 6256 0 1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 8924 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 8740 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_77
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_81
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _088_
timestamp 1586364061
transform 1 0 10764 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_96
timestamp 1586364061
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_100
timestamp 1586364061
transform 1 0 10304 0 1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  _145_
timestamp 1586364061
transform 1 0 13984 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_132
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_136
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 15272 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 14536 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 15088 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_144
timestamp 1586364061
transform 1 0 14352 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_148
timestamp 1586364061
transform 1 0 14720 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__050__C
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17020 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16468 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_165
timestamp 1586364061
transform 1 0 16284 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_169
timestamp 1586364061
transform 1 0 16652 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_or3_4  _050_
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__050__B
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_193
timestamp 1586364061
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_5.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 20884 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_197
timestamp 1586364061
transform 1 0 19228 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_204
timestamp 1586364061
transform 1 0 19872 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_208
timestamp 1586364061
transform 1 0 20240 0 1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2576 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_14
timestamp 1586364061
transform 1 0 2392 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_2  _144_
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2944 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3680 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_18
timestamp 1586364061
transform 1 0 2760 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_22
timestamp 1586364061
transform 1 0 3128 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_26
timestamp 1586364061
transform 1 0 3496 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_30
timestamp 1586364061
transform 1 0 3864 0 -1 8160
box -38 -48 130 592
use scs8hd_nand3_4  _049_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5336 0 -1 8160
box -38 -48 1326 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4692 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5060 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_36
timestamp 1586364061
transform 1 0 4416 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_41
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_45
timestamp 1586364061
transform 1 0 5244 0 -1 8160
box -38 -48 130 592
use scs8hd_or4_4  _091_
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 6808 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__D
timestamp 1586364061
transform 1 0 7176 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_60
timestamp 1586364061
transform 1 0 6624 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_64
timestamp 1586364061
transform 1 0 6992 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 8372 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 8740 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_77
timestamp 1586364061
transform 1 0 8188 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_81
timestamp 1586364061
transform 1 0 8556 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_85
timestamp 1586364061
transform 1 0 8924 0 -1 8160
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 10948 0 -1 8160
box -38 -48 1050 592
use scs8hd_inv_1  mux_top_ipin_6.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9936 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__082__B
timestamp 1586364061
transform 1 0 10580 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_91
timestamp 1586364061
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_10_99
timestamp 1586364061
transform 1 0 10212 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_105
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_118
timestamp 1586364061
transform 1 0 11960 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_122
timestamp 1586364061
transform 1 0 12328 0 -1 8160
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13156 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_125
timestamp 1586364061
transform 1 0 12604 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_129
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_142
timestamp 1586364061
transform 1 0 14168 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14352 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_146
timestamp 1586364061
transform 1 0 14536 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_152
timestamp 1586364061
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_165
timestamp 1586364061
transform 1 0 16284 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_169
timestamp 1586364061
transform 1 0 16652 0 -1 8160
box -38 -48 406 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 18584 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__050__A
timestamp 1586364061
transform 1 0 18032 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__C
timestamp 1586364061
transform 1 0 18400 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_182
timestamp 1586364061
transform 1 0 17848 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_186
timestamp 1586364061
transform 1 0 18216 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 20884 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_199
timestamp 1586364061
transform 1 0 19412 0 -1 8160
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_10_211
timestamp 1586364061
transform 1 0 20516 0 -1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1840 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 1564 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_17
timestamp 1586364061
transform 1 0 2668 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4324 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__B
timestamp 1586364061
transform 1 0 2852 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3680 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3312 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_21
timestamp 1586364061
transform 1 0 3036 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_26
timestamp 1586364061
transform 1 0 3496 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_30
timestamp 1586364061
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_34
timestamp 1586364061
transform 1 0 4232 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5428 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_44
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_49
timestamp 1586364061
transform 1 0 5612 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_or3_4  _105_
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__105__C
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_71
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _072_
timestamp 1586364061
transform 1 0 8372 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__069__B
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__B
timestamp 1586364061
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_75
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_88
timestamp 1586364061
transform 1 0 9200 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 10580 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__C
timestamp 1586364061
transform 1 0 9384 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_92
timestamp 1586364061
transform 1 0 9568 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_96
timestamp 1586364061
transform 1 0 9936 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_99
timestamp 1586364061
transform 1 0 10212 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13984 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_132
timestamp 1586364061
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_136
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15456 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_149
timestamp 1586364061
transform 1 0 14812 0 1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_11_155
timestamp 1586364061
transform 1 0 15364 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_158
timestamp 1586364061
transform 1 0 15640 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__098__D
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_162
timestamp 1586364061
transform 1 0 16008 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_175
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_179
timestamp 1586364061
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_193
timestamp 1586364061
transform 1 0 18860 0 1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 20884 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 19320 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_197
timestamp 1586364061
transform 1 0 19228 0 1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_11_200
timestamp 1586364061
transform 1 0 19504 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_204
timestamp 1586364061
transform 1 0 19872 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_208
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 406 592
use scs8hd_nor2_4  _066_
timestamp 1586364061
transform 1 0 1472 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_13
timestamp 1586364061
transform 1 0 2300 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_17
timestamp 1586364061
transform 1 0 2668 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_3.LATCH_3_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2852 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_21
timestamp 1586364061
transform 1 0 3036 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_25
timestamp 1586364061
transform 1 0 3404 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_43
timestamp 1586364061
transform 1 0 5060 0 -1 9248
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6164 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7176 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_64
timestamp 1586364061
transform 1 0 6992 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 406 592
use scs8hd_or3_4  _069_
timestamp 1586364061
transform 1 0 7728 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_81
timestamp 1586364061
transform 1 0 8556 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_6  FILLER_12_86
timestamp 1586364061
transform 1 0 9016 0 -1 9248
box -38 -48 590 592
use scs8hd_nor2_4  _082_
timestamp 1586364061
transform 1 0 10580 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9844 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_97
timestamp 1586364061
transform 1 0 10028 0 -1 9248
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12236 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_112
timestamp 1586364061
transform 1 0 11408 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_120
timestamp 1586364061
transform 1 0 12144 0 -1 9248
box -38 -48 130 592
use scs8hd_buf_2  _141_
timestamp 1586364061
transform 1 0 14076 0 -1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_132
timestamp 1586364061
transform 1 0 13248 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_136
timestamp 1586364061
transform 1 0 13616 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_140
timestamp 1586364061
transform 1 0 13984 0 -1 9248
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15456 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_158
timestamp 1586364061
transform 1 0 15640 0 -1 9248
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16192 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17204 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_173
timestamp 1586364061
transform 1 0 17020 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_177
timestamp 1586364061
transform 1 0 17388 0 -1 9248
box -38 -48 222 592
use scs8hd_or4_4  _098_
timestamp 1586364061
transform 1 0 17756 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 17572 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18768 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_190
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_194
timestamp 1586364061
transform 1 0 18952 0 -1 9248
box -38 -48 406 592
use scs8hd_buf_2  _157_
timestamp 1586364061
transform 1 0 19320 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 20884 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_202
timestamp 1586364061
transform 1 0 19688 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_210
timestamp 1586364061
transform 1 0 20424 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_3.LATCH_5_.latch
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1564 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__B
timestamp 1586364061
transform 1 0 2576 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_14
timestamp 1586364061
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_14
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_26
timestamp 1586364061
transform 1 0 3496 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_22
timestamp 1586364061
transform 1 0 3128 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_18
timestamp 1586364061
transform 1 0 2760 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_26
timestamp 1586364061
transform 1 0 3496 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_22
timestamp 1586364061
transform 1 0 3128 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_18
timestamp 1586364061
transform 1 0 2760 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__B
timestamp 1586364061
transform 1 0 2944 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 3312 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 2944 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_30
timestamp 1586364061
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3680 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4232 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_3.LATCH_4_.latch
timestamp 1586364061
transform 1 0 3772 0 1 9248
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_13_44
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_40
timestamp 1586364061
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_53
timestamp 1586364061
transform 1 0 5980 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_49
timestamp 1586364061
transform 1 0 5612 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_45
timestamp 1586364061
transform 1 0 5244 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_48
timestamp 1586364061
transform 1 0 5520 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5796 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5336 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5428 0 -1 10336
box -38 -48 222 592
use scs8hd_conb_1  _132_
timestamp 1586364061
transform 1 0 5704 0 1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4416 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_4  FILLER_14_58
timestamp 1586364061
transform 1 0 6440 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6164 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_64
timestamp 1586364061
transform 1 0 6992 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7176 0 -1 10336
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_14_79
timestamp 1586364061
transform 1 0 8372 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_75
timestamp 1586364061
transform 1 0 8004 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_77
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_73
timestamp 1586364061
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 8188 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_87
timestamp 1586364061
transform 1 0 9108 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_13_81
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 8648 0 1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 8832 0 1 9248
box -38 -48 866 592
use scs8hd_decap_4  FILLER_13_97
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_93
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_104
timestamp 1586364061
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_4.LATCH_5_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_4.LATCH_3_.latch
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_14_108
timestamp 1586364061
transform 1 0 11040 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_3  FILLER_14_116
timestamp 1586364061
transform 1 0 11776 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_buf_2  _147_
timestamp 1586364061
transform 1 0 11408 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_121
timestamp 1586364061
transform 1 0 12236 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_125
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_129
timestamp 1586364061
transform 1 0 12972 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13156 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 12788 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_142
timestamp 1586364061
transform 1 0 14168 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_138
timestamp 1586364061
transform 1 0 13800 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_142
timestamp 1586364061
transform 1 0 14168 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 13984 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13340 0 1 9248
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_4.LATCH_4_.latch
timestamp 1586364061
transform 1 0 12788 0 -1 10336
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15088 0 1 9248
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_4.LATCH_2_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 14904 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14536 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_148
timestamp 1586364061
transform 1 0 14720 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_150
timestamp 1586364061
transform 1 0 14904 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_169
timestamp 1586364061
transform 1 0 16652 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_165
timestamp 1586364061
transform 1 0 16284 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_167
timestamp 1586364061
transform 1 0 16468 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_163
timestamp 1586364061
transform 1 0 16100 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16284 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16652 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_175
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_buf_2  _146_
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_186
timestamp 1586364061
transform 1 0 18216 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_182
timestamp 1586364061
transform 1 0 17848 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__047__A
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_193
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 18400 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__B
timestamp 1586364061
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _081_
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 866 592
use scs8hd_inv_8  _047_
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_13_204
timestamp 1586364061
transform 1 0 19872 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_197
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 19412 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_211
timestamp 1586364061
transform 1 0 20516 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 20884 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 20884 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_199
timestamp 1586364061
transform 1 0 19412 0 -1 10336
box -38 -48 1142 592
use scs8hd_nor2_4  _070_
timestamp 1586364061
transform 1 0 1472 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__070__B
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_13
timestamp 1586364061
transform 1 0 2300 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_17
timestamp 1586364061
transform 1 0 2668 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 3036 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_32
timestamp 1586364061
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _071_
timestamp 1586364061
transform 1 0 4784 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 5888 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__B
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_36
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_49
timestamp 1586364061
transform 1 0 5612 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6256 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_54
timestamp 1586364061
transform 1 0 6072 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_58
timestamp 1586364061
transform 1 0 6440 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 8280 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__C
timestamp 1586364061
transform 1 0 8648 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9200 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_76
timestamp 1586364061
transform 1 0 8096 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_80
timestamp 1586364061
transform 1 0 8464 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_84
timestamp 1586364061
transform 1 0 8832 0 1 10336
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9384 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10396 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_99
timestamp 1586364061
transform 1 0 10212 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_103
timestamp 1586364061
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_107
timestamp 1586364061
transform 1 0 10948 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use scs8hd_inv_1  mux_top_ipin_6.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11132 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _114_
timestamp 1586364061
transform 1 0 13984 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 13800 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_132
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_136
timestamp 1586364061
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15548 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15180 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_149
timestamp 1586364061
transform 1 0 14812 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_155
timestamp 1586364061
transform 1 0 15364 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_159
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__078__B
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15916 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_172
timestamp 1586364061
transform 1 0 16928 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_176
timestamp 1586364061
transform 1 0 17296 0 1 10336
box -38 -48 130 592
use scs8hd_nor2_4  _080_
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__080__B
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_193
timestamp 1586364061
transform 1 0 18860 0 1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_4.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 20884 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_199
timestamp 1586364061
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_204
timestamp 1586364061
transform 1 0 19872 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 406 592
use scs8hd_nor2_4  _068_
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use scs8hd_inv_1  mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__107__D
timestamp 1586364061
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_6
timestamp 1586364061
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_10
timestamp 1586364061
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__106__C
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_3.LATCH_2_.latch
timestamp 1586364061
transform 1 0 5888 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5704 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5060 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_41
timestamp 1586364061
transform 1 0 4876 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_45
timestamp 1586364061
transform 1 0 5244 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_49
timestamp 1586364061
transform 1 0 5612 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7084 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_63
timestamp 1586364061
transform 1 0 6900 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_67
timestamp 1586364061
transform 1 0 7268 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_71
timestamp 1586364061
transform 1 0 7636 0 -1 11424
box -38 -48 314 592
use scs8hd_or3_4  _115_
timestamp 1586364061
transform 1 0 7912 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_6  FILLER_16_83
timestamp 1586364061
transform 1 0 8740 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_89
timestamp 1586364061
transform 1 0 9292 0 -1 11424
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_103
timestamp 1586364061
transform 1 0 10580 0 -1 11424
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11316 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12512 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_122
timestamp 1586364061
transform 1 0 12328 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13064 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12880 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_126
timestamp 1586364061
transform 1 0 12696 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_139
timestamp 1586364061
transform 1 0 13892 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15456 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_158
timestamp 1586364061
transform 1 0 15640 0 -1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 -1 11424
box -38 -48 866 592
use scs8hd_fill_1  FILLER_16_162
timestamp 1586364061
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_172
timestamp 1586364061
transform 1 0 16928 0 -1 11424
box -38 -48 774 592
use scs8hd_nor2_4  _078_
timestamp 1586364061
transform 1 0 17664 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 18676 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_189
timestamp 1586364061
transform 1 0 18492 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_193
timestamp 1586364061
transform 1 0 18860 0 -1 11424
box -38 -48 406 592
use scs8hd_buf_2  _150_
timestamp 1586364061
transform 1 0 19228 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 20884 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_201
timestamp 1586364061
transform 1 0 19596 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  FILLER_16_209
timestamp 1586364061
transform 1 0 20332 0 -1 11424
box -38 -48 314 592
use scs8hd_nor4_4  _107_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 1602 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3956 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 3128 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__C
timestamp 1586364061
transform 1 0 3496 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_20
timestamp 1586364061
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_24
timestamp 1586364061
transform 1 0 3312 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_28
timestamp 1586364061
transform 1 0 3680 0 1 11424
box -38 -48 314 592
use scs8hd_buf_2  _140_
timestamp 1586364061
transform 1 0 5520 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 4968 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 5336 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_40
timestamp 1586364061
transform 1 0 4784 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_44
timestamp 1586364061
transform 1 0 5152 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_52
timestamp 1586364061
transform 1 0 5888 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 6072 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6440 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_56
timestamp 1586364061
transform 1 0 6256 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_60
timestamp 1586364061
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_71
timestamp 1586364061
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8372 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8832 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_75
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_82
timestamp 1586364061
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9568 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9384 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10764 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_103
timestamp 1586364061
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_107
timestamp 1586364061
transform 1 0 10948 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11132 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13064 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12696 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_128
timestamp 1586364061
transform 1 0 12880 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14996 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14444 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14812 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_143
timestamp 1586364061
transform 1 0 14260 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_147
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_160
timestamp 1586364061
transform 1 0 15824 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_4.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16560 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17020 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__B
timestamp 1586364061
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 16376 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16008 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_164
timestamp 1586364061
transform 1 0 16192 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_171
timestamp 1586364061
transform 1 0 16836 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_175
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use scs8hd_inv_8  _046_
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__046__A
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 19044 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_179
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_193
timestamp 1586364061
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 20884 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_197
timestamp 1586364061
transform 1 0 19228 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_204
timestamp 1586364061
transform 1 0 19872 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_208
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 406 592
use scs8hd_nor4_4  _106_
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1602 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_nor2_4  _104_
timestamp 1586364061
transform 1 0 4140 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__060__B
timestamp 1586364061
transform 1 0 3128 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__D
timestamp 1586364061
transform 1 0 3496 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_20
timestamp 1586364061
transform 1 0 2944 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_24
timestamp 1586364061
transform 1 0 3312 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_28
timestamp 1586364061
transform 1 0 3680 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5704 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5520 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_42
timestamp 1586364061
transform 1 0 4968 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_46
timestamp 1586364061
transform 1 0 5336 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6900 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_61
timestamp 1586364061
transform 1 0 6716 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_65
timestamp 1586364061
transform 1 0 7084 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__C
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_78
timestamp 1586364061
transform 1 0 8280 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_82
timestamp 1586364061
transform 1 0 8648 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_86
timestamp 1586364061
transform 1 0 9016 0 -1 12512
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9936 0 -1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_18_107
timestamp 1586364061
transform 1 0 10948 0 -1 12512
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11684 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11408 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_111
timestamp 1586364061
transform 1 0 11316 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_114
timestamp 1586364061
transform 1 0 11592 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_124
timestamp 1586364061
transform 1 0 12512 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13432 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13248 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12696 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_128
timestamp 1586364061
transform 1 0 12880 0 -1 12512
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_149
timestamp 1586364061
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _077_
timestamp 1586364061
transform 1 0 16836 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_163
timestamp 1586364061
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_167
timestamp 1586364061
transform 1 0 16468 0 -1 12512
box -38 -48 406 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 18400 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 18032 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_180
timestamp 1586364061
transform 1 0 17664 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_186
timestamp 1586364061
transform 1 0 18216 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 20884 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_197
timestamp 1586364061
transform 1 0 19228 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_18_209
timestamp 1586364061
transform 1 0 20332 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_6
timestamp 1586364061
transform 1 0 1656 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use scs8hd_buf_2  _143_
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_10
timestamp 1586364061
transform 1 0 2024 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_13
timestamp 1586364061
transform 1 0 2300 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 2208 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__060__A
timestamp 1586364061
transform 1 0 2116 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__060__C
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _102_
timestamp 1586364061
transform 1 0 2392 0 -1 13600
box -38 -48 866 592
use scs8hd_or3_4  _060_
timestamp 1586364061
transform 1 0 2668 0 1 12512
box -38 -48 866 592
use scs8hd_decap_4  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_26
timestamp 1586364061
transform 1 0 3496 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_29
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_30
timestamp 1586364061
transform 1 0 3864 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 3680 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4048 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_7.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_35
timestamp 1586364061
transform 1 0 4324 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_34
timestamp 1586364061
transform 1 0 4232 0 1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5060 0 -1 13600
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4692 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_38
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_41
timestamp 1586364061
transform 1 0 4876 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_58
timestamp 1586364061
transform 1 0 6440 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_54
timestamp 1586364061
transform 1 0 6072 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6624 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_20_71
timestamp 1586364061
transform 1 0 7636 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_71
timestamp 1586364061
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use scs8hd_or3_4  _108_
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 866 592
use scs8hd_inv_1  mux_top_ipin_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8372 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_75
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_88
timestamp 1586364061
transform 1 0 9200 0 1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_20_82
timestamp 1586364061
transform 1 0 8648 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_20_90
timestamp 1586364061
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_95
timestamp 1586364061
transform 1 0 9844 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_92
timestamp 1586364061
transform 1 0 9568 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10028 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_104
timestamp 1586364061
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_99
timestamp 1586364061
transform 1 0 10212 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_20_108
timestamp 1586364061
transform 1 0 11040 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_112
timestamp 1586364061
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_121
timestamp 1586364061
transform 1 0 12236 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_19_116
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12512 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _113_
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__113__B
timestamp 1586364061
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_132
timestamp 1586364061
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_136
timestamp 1586364061
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_140
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_126
timestamp 1586364061
transform 1 0 12696 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_138
timestamp 1586364061
transform 1 0 13800 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_142
timestamp 1586364061
transform 1 0 14168 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_149
timestamp 1586364061
transform 1 0 14812 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 14260 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_156
timestamp 1586364061
transform 1 0 15456 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_152
timestamp 1586364061
transform 1 0 15088 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15640 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14260 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 16836 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_169
timestamp 1586364061
transform 1 0 16652 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_173
timestamp 1586364061
transform 1 0 17020 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_177
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_163
timestamp 1586364061
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_167
timestamp 1586364061
transform 1 0 16468 0 -1 13600
box -38 -48 406 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 18400 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_193
timestamp 1586364061
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_180
timestamp 1586364061
transform 1 0 17664 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_204
timestamp 1586364061
transform 1 0 19872 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_197
timestamp 1586364061
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_209
timestamp 1586364061
transform 1 0 20332 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 20884 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 20884 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_197
timestamp 1586364061
transform 1 0 19228 0 -1 13600
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 1050 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 2576 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_14
timestamp 1586364061
transform 1 0 2392 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _073_
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__073__B
timestamp 1586364061
transform 1 0 3404 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2944 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_18
timestamp 1586364061
transform 1 0 2760 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_22
timestamp 1586364061
transform 1 0 3128 0 1 13600
box -38 -48 314 592
use scs8hd_nor2_4  _118_
timestamp 1586364061
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_36
timestamp 1586364061
transform 1 0 4416 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_21_41
timestamp 1586364061
transform 1 0 4876 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_71
timestamp 1586364061
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_7.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8372 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8832 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9200 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8188 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_75
timestamp 1586364061
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_82
timestamp 1586364061
transform 1 0 8648 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_86
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9752 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9568 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10948 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_90
timestamp 1586364061
transform 1 0 9384 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_105
timestamp 1586364061
transform 1 0 10764 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 12512 0 1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11316 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_109
timestamp 1586364061
transform 1 0 11132 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_113
timestamp 1586364061
transform 1 0 11500 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14076 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13708 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_135
timestamp 1586364061
transform 1 0 13524 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_139
timestamp 1586364061
transform 1 0 13892 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 14260 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15456 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_154
timestamp 1586364061
transform 1 0 15272 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_158
timestamp 1586364061
transform 1 0 15640 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16008 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 17020 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_171
timestamp 1586364061
transform 1 0 16836 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_175
timestamp 1586364061
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 1 13600
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_179
timestamp 1586364061
transform 1 0 17572 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_187
timestamp 1586364061
transform 1 0 18308 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_191
timestamp 1586364061
transform 1 0 18676 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 20884 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19504 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19872 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_198
timestamp 1586364061
transform 1 0 19320 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_202
timestamp 1586364061
transform 1 0 19688 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_206
timestamp 1586364061
transform 1 0 20056 0 1 13600
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2024 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 1564 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_7
timestamp 1586364061
transform 1 0 1748 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3036 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_19
timestamp 1586364061
transform 1 0 2852 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_23
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_4  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_7.LATCH_2_.latch
timestamp 1586364061
transform 1 0 4692 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 5888 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4508 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_36
timestamp 1586364061
transform 1 0 4416 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_50
timestamp 1586364061
transform 1 0 5704 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_7.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7544 0 -1 14688
box -38 -48 1050 592
use scs8hd_inv_1  mux_top_ipin_7.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6532 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6992 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_54
timestamp 1586364061
transform 1 0 6072 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_58
timestamp 1586364061
transform 1 0 6440 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_62
timestamp 1586364061
transform 1 0 6808 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_66
timestamp 1586364061
transform 1 0 7176 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_81
timestamp 1586364061
transform 1 0 8556 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_85
timestamp 1586364061
transform 1 0 8924 0 -1 14688
box -38 -48 590 592
use scs8hd_conb_1  _131_
timestamp 1586364061
transform 1 0 9936 0 -1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10948 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10396 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_91
timestamp 1586364061
transform 1 0 9476 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_99
timestamp 1586364061
transform 1 0 10212 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_103
timestamp 1586364061
transform 1 0 10580 0 -1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12512 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12328 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_116
timestamp 1586364061
transform 1 0 11776 0 -1 14688
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14076 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 13524 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13892 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_133
timestamp 1586364061
transform 1 0 13340 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_137
timestamp 1586364061
transform 1 0 13708 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_144
timestamp 1586364061
transform 1 0 14352 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_22_150
timestamp 1586364061
transform 1 0 14904 0 -1 14688
box -38 -48 130 592
use scs8hd_nor2_4  _126_
timestamp 1586364061
transform 1 0 16836 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_163
timestamp 1586364061
transform 1 0 16100 0 -1 14688
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18400 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_180
timestamp 1586364061
transform 1 0 17664 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_8  FILLER_22_191
timestamp 1586364061
transform 1 0 18676 0 -1 14688
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19412 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 20884 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_202
timestamp 1586364061
transform 1 0 19688 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_210
timestamp 1586364061
transform 1 0 20424 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2208 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_6
timestamp 1586364061
transform 1 0 1656 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_10
timestamp 1586364061
transform 1 0 2024 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_7.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_23
timestamp 1586364061
transform 1 0 3220 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_36
timestamp 1586364061
transform 1 0 4416 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_40
timestamp 1586364061
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7544 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7176 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_68
timestamp 1586364061
transform 1 0 7360 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7728 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 9292 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_81
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_87
timestamp 1586364061
transform 1 0 9108 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 10028 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_91
timestamp 1586364061
transform 1 0 9476 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_95
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_108
timestamp 1586364061
transform 1 0 11040 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_114
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_118
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 13340 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_126
timestamp 1586364061
transform 1 0 12696 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_130
timestamp 1586364061
transform 1 0 13064 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15088 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14720 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_146
timestamp 1586364061
transform 1 0 14536 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_150
timestamp 1586364061
transform 1 0 14904 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17296 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16652 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16284 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_163
timestamp 1586364061
transform 1 0 16100 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_167
timestamp 1586364061
transform 1 0 16468 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_174
timestamp 1586364061
transform 1 0 17112 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_178
timestamp 1586364061
transform 1 0 17480 0 1 14688
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 1 14688
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_4.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_187
timestamp 1586364061
transform 1 0 18308 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_191
timestamp 1586364061
transform 1 0 18676 0 1 14688
box -38 -48 406 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 20884 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19504 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 19872 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_198
timestamp 1586364061
transform 1 0 19320 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_202
timestamp 1586364061
transform 1 0 19688 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_206
timestamp 1586364061
transform 1 0 20056 0 1 14688
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1050 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2576 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_14
timestamp 1586364061
transform 1 0 2392 0 -1 15776
box -38 -48 222 592
use scs8hd_buf_2  _155_
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__040__A
timestamp 1586364061
transform 1 0 3312 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2944 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_18
timestamp 1586364061
transform 1 0 2760 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_22
timestamp 1586364061
transform 1 0 3128 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_26
timestamp 1586364061
transform 1 0 3496 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_30
timestamp 1586364061
transform 1 0 3864 0 -1 15776
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_7.LATCH_4_.latch
timestamp 1586364061
transform 1 0 5520 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 4692 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_36
timestamp 1586364061
transform 1 0 4416 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_41
timestamp 1586364061
transform 1 0 4876 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_46
timestamp 1586364061
transform 1 0 5336 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6716 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_59
timestamp 1586364061
transform 1 0 6532 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_63
timestamp 1586364061
transform 1 0 6900 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 8556 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_76
timestamp 1586364061
transform 1 0 8096 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_80
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_6  FILLER_24_83
timestamp 1586364061
transform 1 0 8740 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_89
timestamp 1586364061
transform 1 0 9292 0 -1 15776
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_104
timestamp 1586364061
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_108
timestamp 1586364061
transform 1 0 11040 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_121
timestamp 1586364061
transform 1 0 12236 0 -1 15776
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 13432 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 12696 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 13064 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_125
timestamp 1586364061
transform 1 0 12604 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_128
timestamp 1586364061
transform 1 0 12880 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_132
timestamp 1586364061
transform 1 0 13248 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_145
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_163
timestamp 1586364061
transform 1 0 16100 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_8  FILLER_24_174
timestamp 1586364061
transform 1 0 17112 0 -1 15776
box -38 -48 774 592
use scs8hd_buf_2  _156_
timestamp 1586364061
transform 1 0 19044 0 -1 15776
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17848 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_185
timestamp 1586364061
transform 1 0 18124 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_193
timestamp 1586364061
transform 1 0 18860 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 20884 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_199
timestamp 1586364061
transform 1 0 19412 0 -1 15776
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_24_211
timestamp 1586364061
transform 1 0 20516 0 -1 15776
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_16
timestamp 1586364061
transform 1 0 2576 0 1 15776
box -38 -48 222 592
use scs8hd_inv_8  _040_
timestamp 1586364061
transform 1 0 3312 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 4324 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2760 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3128 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_20
timestamp 1586364061
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_33
timestamp 1586364061
transform 1 0 4140 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _099_
timestamp 1586364061
transform 1 0 5152 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__100__B
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_37
timestamp 1586364061
transform 1 0 4508 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_41
timestamp 1586364061
transform 1 0 4876 0 1 15776
box -38 -48 314 592
use scs8hd_decap_6  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_7.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 8556 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 8372 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_73
timestamp 1586364061
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_77
timestamp 1586364061
transform 1 0 8188 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 9660 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_90
timestamp 1586364061
transform 1 0 9384 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_25_95
timestamp 1586364061
transform 1 0 9844 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_107
timestamp 1586364061
transform 1 0 10948 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 11132 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_111
timestamp 1586364061
transform 1 0 11316 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_115
timestamp 1586364061
transform 1 0 11684 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_118
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _109_
timestamp 1586364061
transform 1 0 12604 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 14076 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13616 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_134
timestamp 1586364061
transform 1 0 13432 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_138
timestamp 1586364061
transform 1 0 13800 0 1 15776
box -38 -48 314 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 14260 0 1 15776
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15824 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_152
timestamp 1586364061
transform 1 0 15088 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_156
timestamp 1586364061
transform 1 0 15456 0 1 15776
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17296 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16284 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16652 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_163
timestamp 1586364061
transform 1 0 16100 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_167
timestamp 1586364061
transform 1 0 16468 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_174
timestamp 1586364061
transform 1 0 17112 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_178
timestamp 1586364061
transform 1 0 17480 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 1 15776
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17664 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18860 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_182
timestamp 1586364061
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_187
timestamp 1586364061
transform 1 0 18308 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_191
timestamp 1586364061
transform 1 0 18676 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 20884 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19504 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_198
timestamp 1586364061
transform 1 0 19320 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_202
timestamp 1586364061
transform 1 0 19688 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_25_210
timestamp 1586364061
transform 1 0 20424 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_7
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_7
timestamp 1586364061
transform 1 0 1748 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 1840 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_buf_2  _153_
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_11
timestamp 1586364061
transform 1 0 2116 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__048__A
timestamp 1586364061
transform 1 0 2300 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2024 0 -1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _075_
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_26_19
timestamp 1586364061
transform 1 0 2852 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__048__C
timestamp 1586364061
transform 1 0 3036 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_24
timestamp 1586364061
transform 1 0 3312 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__B
timestamp 1586364061
transform 1 0 3496 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_28
timestamp 1586364061
transform 1 0 3680 0 1 16864
box -38 -48 406 592
use scs8hd_decap_4  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4048 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_27_34
timestamp 1586364061
transform 1 0 4232 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_26_36
timestamp 1586364061
transform 1 0 4416 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__103__B
timestamp 1586364061
transform 1 0 4508 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_50
timestamp 1586364061
transform 1 0 5704 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_46
timestamp 1586364061
transform 1 0 5336 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_52
timestamp 1586364061
transform 1 0 5888 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_26_48
timestamp 1586364061
transform 1 0 5520 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 5704 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__B
timestamp 1586364061
transform 1 0 5520 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _103_
timestamp 1586364061
transform 1 0 4508 0 1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _100_
timestamp 1586364061
transform 1 0 4692 0 -1 16864
box -38 -48 866 592
use scs8hd_decap_3  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_54
timestamp 1586364061
transform 1 0 6072 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_60
timestamp 1586364061
transform 1 0 6624 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__C
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_64
timestamp 1586364061
transform 1 0 6992 0 -1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7176 0 -1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _101_
timestamp 1586364061
transform 1 0 7084 0 1 16864
box -38 -48 866 592
use scs8hd_decap_4  FILLER_27_78
timestamp 1586364061
transform 1 0 8280 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_79
timestamp 1586364061
transform 1 0 8372 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_26_75
timestamp 1586364061
transform 1 0 8004 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__B
timestamp 1586364061
transform 1 0 8188 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 8096 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_82
timestamp 1586364061
transform 1 0 8648 0 1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_26_87
timestamp 1586364061
transform 1 0 9108 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 8924 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 8740 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 8924 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_98
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_94
timestamp 1586364061
transform 1 0 9752 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 9936 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_106
timestamp 1586364061
transform 1 0 10856 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_102
timestamp 1586364061
transform 1 0 10488 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__B
timestamp 1586364061
transform 1 0 10304 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _079_
timestamp 1586364061
transform 1 0 10488 0 1 16864
box -38 -48 866 592
use scs8hd_decap_4  FILLER_27_115
timestamp 1586364061
transform 1 0 11684 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_111
timestamp 1586364061
transform 1 0 11316 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_113
timestamp 1586364061
transform 1 0 11500 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11500 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_27_119
timestamp 1586364061
transform 1 0 12052 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_121
timestamp 1586364061
transform 1 0 12236 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 12420 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _110_
timestamp 1586364061
transform 1 0 12696 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13432 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13892 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_125
timestamp 1586364061
transform 1 0 12604 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_135
timestamp 1586364061
transform 1 0 13524 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_132
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_136
timestamp 1586364061
transform 1 0 13616 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_27_141
timestamp 1586364061
transform 1 0 14076 0 1 16864
box -38 -48 314 592
use scs8hd_decap_8  FILLER_27_147
timestamp 1586364061
transform 1 0 14628 0 1 16864
box -38 -48 774 592
use scs8hd_decap_8  FILLER_26_145
timestamp 1586364061
transform 1 0 14444 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 14260 0 -1 16864
box -38 -48 222 592
use scs8hd_conb_1  _129_
timestamp 1586364061
transform 1 0 14352 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_158
timestamp 1586364061
transform 1 0 15640 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_157
timestamp 1586364061
transform 1 0 15548 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15824 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_4.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15364 0 1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_169
timestamp 1586364061
transform 1 0 16652 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_162
timestamp 1586364061
transform 1 0 16008 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_168
timestamp 1586364061
transform 1 0 16560 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16192 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16284 0 -1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16376 0 1 16864
box -38 -48 314 592
use scs8hd_decap_6  FILLER_27_177
timestamp 1586364061
transform 1 0 17388 0 1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_173
timestamp 1586364061
transform 1 0 17020 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16836 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17296 0 -1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18308 0 -1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_179
timestamp 1586364061
transform 1 0 17572 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_12  FILLER_26_190
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_196
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 20884 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 20884 0 1 16864
box -38 -48 314 592
use scs8hd_decap_8  FILLER_26_202
timestamp 1586364061
transform 1 0 19688 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_26_210
timestamp 1586364061
transform 1 0 20424 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 406 592
use scs8hd_or3_4  _048_
timestamp 1586364061
transform 1 0 2392 0 -1 17952
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 1840 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__048__B
timestamp 1586364061
transform 1 0 2208 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_6
timestamp 1586364061
transform 1 0 1656 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_10
timestamp 1586364061
transform 1 0 2024 0 -1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_35
timestamp 1586364061
transform 1 0 4324 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _074_
timestamp 1586364061
transform 1 0 5428 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__052__A
timestamp 1586364061
transform 1 0 4508 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__052__B
timestamp 1586364061
transform 1 0 4876 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 5244 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_39
timestamp 1586364061
transform 1 0 4692 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_43
timestamp 1586364061
transform 1 0 5060 0 -1 17952
box -38 -48 222 592
use scs8hd_or3_4  _076_
timestamp 1586364061
transform 1 0 7544 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__101__B
timestamp 1586364061
transform 1 0 7084 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_28_64
timestamp 1586364061
transform 1 0 6992 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_28_67
timestamp 1586364061
transform 1 0 7268 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 8556 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_79
timestamp 1586364061
transform 1 0 8372 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_83
timestamp 1586364061
transform 1 0 8740 0 -1 17952
box -38 -48 774 592
use scs8hd_nor2_4  _121_
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10948 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_91
timestamp 1586364061
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_102
timestamp 1586364061
transform 1 0 10488 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_106
timestamp 1586364061
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_28_109
timestamp 1586364061
transform 1 0 11132 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_113
timestamp 1586364061
transform 1 0 11500 0 -1 17952
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12880 0 -1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13892 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_125
timestamp 1586364061
transform 1 0 12604 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_131
timestamp 1586364061
transform 1 0 13156 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_8  FILLER_28_142
timestamp 1586364061
transform 1 0 14168 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_28_150
timestamp 1586364061
transform 1 0 14904 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_157
timestamp 1586364061
transform 1 0 15548 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16284 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_168
timestamp 1586364061
transform 1 0 16560 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_180
timestamp 1586364061
transform 1 0 17664 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_192
timestamp 1586364061
transform 1 0 18768 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 20884 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_204
timestamp 1586364061
transform 1 0 19872 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_8  _043_
timestamp 1586364061
transform 1 0 2668 0 1 17952
box -38 -48 866 592
use scs8hd_buf_2  _152_
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__042__A
timestamp 1586364061
transform 1 0 2392 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__043__A
timestamp 1586364061
transform 1 0 2024 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_7
timestamp 1586364061
transform 1 0 1748 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_12
timestamp 1586364061
transform 1 0 2208 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_16
timestamp 1586364061
transform 1 0 2576 0 1 17952
box -38 -48 130 592
use scs8hd_inv_8  _039_
timestamp 1586364061
transform 1 0 4232 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__052__C
timestamp 1586364061
transform 1 0 4048 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__039__A
timestamp 1586364061
transform 1 0 3680 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_26
timestamp 1586364061
transform 1 0 3496 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_30
timestamp 1586364061
transform 1 0 3864 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__056__C
timestamp 1586364061
transform 1 0 5612 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__056__B
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__056__A
timestamp 1586364061
transform 1 0 5244 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_43
timestamp 1586364061
transform 1 0 5060 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_47
timestamp 1586364061
transform 1 0 5428 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_51
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 222 592
use scs8hd_conb_1  _139_
timestamp 1586364061
transform 1 0 6900 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__054__B
timestamp 1586364061
transform 1 0 7360 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__054__C
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_55
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_66
timestamp 1586364061
transform 1 0 7176 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_70
timestamp 1586364061
transform 1 0 7544 0 1 17952
box -38 -48 222 592
use scs8hd_or3_4  _122_
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__122__C
timestamp 1586364061
transform 1 0 7728 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__054__A
timestamp 1586364061
transform 1 0 8924 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_83
timestamp 1586364061
transform 1 0 8740 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_87
timestamp 1586364061
transform 1 0 9108 0 1 17952
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9936 0 1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_3.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10948 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10672 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9752 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_93
timestamp 1586364061
transform 1 0 9660 0 1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_29_99
timestamp 1586364061
transform 1 0 10212 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_103
timestamp 1586364061
transform 1 0 10580 0 1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_29_106
timestamp 1586364061
transform 1 0 10856 0 1 17952
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11684 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_110
timestamp 1586364061
transform 1 0 11224 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_29_117
timestamp 1586364061
transform 1 0 11868 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_121
timestamp 1586364061
transform 1 0 12236 0 1 17952
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13432 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13892 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_126
timestamp 1586364061
transform 1 0 12696 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_130
timestamp 1586364061
transform 1 0 13064 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_137
timestamp 1586364061
transform 1 0 13708 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_141
timestamp 1586364061
transform 1 0 14076 0 1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15456 0 1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14444 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14260 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14904 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_148
timestamp 1586364061
transform 1 0 14720 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_152
timestamp 1586364061
transform 1 0 15088 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_159
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15916 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_163
timestamp 1586364061
transform 1 0 16100 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_175
timestamp 1586364061
transform 1 0 17204 0 1 17952
box -38 -48 774 592
use scs8hd_buf_2  _151_
timestamp 1586364061
transform 1 0 18492 0 1 17952
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_188
timestamp 1586364061
transform 1 0 18400 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_193
timestamp 1586364061
transform 1 0 18860 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 20884 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_197
timestamp 1586364061
transform 1 0 19228 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_29_209
timestamp 1586364061
transform 1 0 20332 0 1 17952
box -38 -48 314 592
use scs8hd_inv_8  _042_
timestamp 1586364061
transform 1 0 2392 0 -1 19040
box -38 -48 866 592
use scs8hd_conb_1  _130_
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_6
timestamp 1586364061
transform 1 0 1656 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_10
timestamp 1586364061
transform 1 0 2024 0 -1 19040
box -38 -48 406 592
use scs8hd_or3_4  _052_
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_23
timestamp 1586364061
transform 1 0 3220 0 -1 19040
box -38 -48 774 592
use scs8hd_or3_4  _056_
timestamp 1586364061
transform 1 0 5612 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_8  FILLER_30_41
timestamp 1586364061
transform 1 0 4876 0 -1 19040
box -38 -48 774 592
use scs8hd_or3_4  _054_
timestamp 1586364061
transform 1 0 7176 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__051__B
timestamp 1586364061
transform 1 0 6900 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_58
timestamp 1586364061
transform 1 0 6440 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_62
timestamp 1586364061
transform 1 0 6808 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_65
timestamp 1586364061
transform 1 0 7084 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 8188 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_75
timestamp 1586364061
transform 1 0 8004 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_79
timestamp 1586364061
transform 1 0 8372 0 -1 19040
box -38 -48 1142 592
use scs8hd_conb_1  _136_
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_3.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10672 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_91
timestamp 1586364061
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_96
timestamp 1586364061
transform 1 0 9936 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_8  FILLER_30_107
timestamp 1586364061
transform 1 0 10948 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11684 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_118
timestamp 1586364061
transform 1 0 11960 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13708 0 -1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12696 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_129
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_12  FILLER_30_140
timestamp 1586364061
transform 1 0 13984 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_152
timestamp 1586364061
transform 1 0 15088 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_166
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_178
timestamp 1586364061
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_190
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 20884 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_202
timestamp 1586364061
transform 1 0 19688 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_30_210
timestamp 1586364061
transform 1 0 20424 0 -1 19040
box -38 -48 222 592
use scs8hd_inv_8  _041_
timestamp 1586364061
transform 1 0 2024 0 1 19040
box -38 -48 866 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__041__A
timestamp 1586364061
transform 1 0 1840 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_7
timestamp 1586364061
transform 1 0 1748 0 1 19040
box -38 -48 130 592
use scs8hd_or3_4  _058_
timestamp 1586364061
transform 1 0 4048 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 3956 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__058__A
timestamp 1586364061
transform 1 0 3772 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__058__B
timestamp 1586364061
transform 1 0 3404 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_19
timestamp 1586364061
transform 1 0 2852 0 1 19040
box -38 -48 590 592
use scs8hd_fill_2  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5612 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__058__C
timestamp 1586364061
transform 1 0 5060 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_41
timestamp 1586364061
transform 1 0 4876 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_45
timestamp 1586364061
transform 1 0 5244 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_52
timestamp 1586364061
transform 1 0 5888 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _051_
timestamp 1586364061
transform 1 0 6900 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__051__A
timestamp 1586364061
transform 1 0 6624 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6072 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_56
timestamp 1586364061
transform 1 0 6256 0 1 19040
box -38 -48 406 592
use scs8hd_conb_1  _138_
timestamp 1586364061
transform 1 0 8556 0 1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_31_72
timestamp 1586364061
transform 1 0 7728 0 1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_31_80
timestamp 1586364061
transform 1 0 8464 0 1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_31_84
timestamp 1586364061
transform 1 0 8832 0 1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10764 0 1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_3.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9752 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9660 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10212 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_92
timestamp 1586364061
transform 1 0 9568 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_97
timestamp 1586364061
transform 1 0 10028 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_101
timestamp 1586364061
transform 1 0 10396 0 1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 12512 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_108
timestamp 1586364061
transform 1 0 11040 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_112
timestamp 1586364061
transform 1 0 11408 0 1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13616 0 1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12604 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14076 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13064 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_128
timestamp 1586364061
transform 1 0 12880 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_132
timestamp 1586364061
transform 1 0 13248 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_139
timestamp 1586364061
transform 1 0 13892 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 15364 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_143
timestamp 1586364061
transform 1 0 14260 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_156
timestamp 1586364061
transform 1 0 15456 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_168
timestamp 1586364061
transform 1 0 16560 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 18216 0 1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_31_180
timestamp 1586364061
transform 1 0 17664 0 1 19040
box -38 -48 590 592
use scs8hd_decap_12  FILLER_31_187
timestamp 1586364061
transform 1 0 18308 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 20884 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_199
timestamp 1586364061
transform 1 0 19412 0 1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_31_211
timestamp 1586364061
transform 1 0 20516 0 1 19040
box -38 -48 130 592
<< labels >>
rlabel metal2 s 1766 21520 1822 22000 6 address[0]
port 0 nsew default input
rlabel metal2 s 2870 0 2926 480 6 address[1]
port 1 nsew default input
rlabel metal2 s 5354 21520 5410 22000 6 address[2]
port 2 nsew default input
rlabel metal2 s 9034 21520 9090 22000 6 address[3]
port 3 nsew default input
rlabel metal3 s 0 552 480 672 6 address[4]
port 4 nsew default input
rlabel metal2 s 12714 21520 12770 22000 6 address[5]
port 5 nsew default input
rlabel metal3 s 0 1640 480 1760 6 address[6]
port 6 nsew default input
rlabel metal2 s 3974 0 4030 480 6 bottom_grid_pin_0_
port 7 nsew default tristate
rlabel metal2 s 6274 0 6330 480 6 bottom_grid_pin_10_
port 8 nsew default tristate
rlabel metal2 s 7470 0 7526 480 6 bottom_grid_pin_12_
port 9 nsew default tristate
rlabel metal2 s 16394 21520 16450 22000 6 bottom_grid_pin_14_
port 10 nsew default tristate
rlabel metal2 s 5170 0 5226 480 6 bottom_grid_pin_2_
port 11 nsew default tristate
rlabel metal3 s 0 2728 480 2848 6 bottom_grid_pin_4_
port 12 nsew default tristate
rlabel metal3 s 0 3816 480 3936 6 bottom_grid_pin_6_
port 13 nsew default tristate
rlabel metal3 s 0 4904 480 5024 6 bottom_grid_pin_8_
port 14 nsew default tristate
rlabel metal3 s 21520 960 22000 1080 6 chanx_left_in[0]
port 15 nsew default input
rlabel metal3 s 0 5992 480 6112 6 chanx_left_in[1]
port 16 nsew default input
rlabel metal3 s 0 7080 480 7200 6 chanx_left_in[2]
port 17 nsew default input
rlabel metal2 s 8666 0 8722 480 6 chanx_left_in[3]
port 18 nsew default input
rlabel metal3 s 21520 2864 22000 2984 6 chanx_left_in[4]
port 19 nsew default input
rlabel metal3 s 0 8168 480 8288 6 chanx_left_in[5]
port 20 nsew default input
rlabel metal2 s 9770 0 9826 480 6 chanx_left_in[6]
port 21 nsew default input
rlabel metal3 s 21520 4904 22000 5024 6 chanx_left_in[7]
port 22 nsew default input
rlabel metal3 s 21520 6944 22000 7064 6 chanx_left_in[8]
port 23 nsew default input
rlabel metal2 s 10966 0 11022 480 6 chanx_left_out[0]
port 24 nsew default tristate
rlabel metal2 s 12070 0 12126 480 6 chanx_left_out[1]
port 25 nsew default tristate
rlabel metal3 s 21520 8848 22000 8968 6 chanx_left_out[2]
port 26 nsew default tristate
rlabel metal2 s 13266 0 13322 480 6 chanx_left_out[3]
port 27 nsew default tristate
rlabel metal3 s 0 9256 480 9376 6 chanx_left_out[4]
port 28 nsew default tristate
rlabel metal3 s 0 10344 480 10464 6 chanx_left_out[5]
port 29 nsew default tristate
rlabel metal2 s 14370 0 14426 480 6 chanx_left_out[6]
port 30 nsew default tristate
rlabel metal2 s 15566 0 15622 480 6 chanx_left_out[7]
port 31 nsew default tristate
rlabel metal3 s 0 11568 480 11688 6 chanx_left_out[8]
port 32 nsew default tristate
rlabel metal3 s 0 12656 480 12776 6 chanx_right_in[0]
port 33 nsew default input
rlabel metal3 s 21520 10888 22000 11008 6 chanx_right_in[1]
port 34 nsew default input
rlabel metal2 s 16762 0 16818 480 6 chanx_right_in[2]
port 35 nsew default input
rlabel metal3 s 0 13744 480 13864 6 chanx_right_in[3]
port 36 nsew default input
rlabel metal3 s 21520 12928 22000 13048 6 chanx_right_in[4]
port 37 nsew default input
rlabel metal3 s 0 14832 480 14952 6 chanx_right_in[5]
port 38 nsew default input
rlabel metal2 s 17866 0 17922 480 6 chanx_right_in[6]
port 39 nsew default input
rlabel metal3 s 21520 14968 22000 15088 6 chanx_right_in[7]
port 40 nsew default input
rlabel metal3 s 0 15920 480 16040 6 chanx_right_in[8]
port 41 nsew default input
rlabel metal2 s 19062 0 19118 480 6 chanx_right_out[0]
port 42 nsew default tristate
rlabel metal3 s 21520 16872 22000 16992 6 chanx_right_out[1]
port 43 nsew default tristate
rlabel metal3 s 0 17008 480 17128 6 chanx_right_out[2]
port 44 nsew default tristate
rlabel metal2 s 20166 0 20222 480 6 chanx_right_out[3]
port 45 nsew default tristate
rlabel metal3 s 0 18096 480 18216 6 chanx_right_out[4]
port 46 nsew default tristate
rlabel metal3 s 0 19184 480 19304 6 chanx_right_out[5]
port 47 nsew default tristate
rlabel metal2 s 20074 21520 20130 22000 6 chanx_right_out[6]
port 48 nsew default tristate
rlabel metal3 s 21520 18912 22000 19032 6 chanx_right_out[7]
port 49 nsew default tristate
rlabel metal2 s 21362 0 21418 480 6 chanx_right_out[8]
port 50 nsew default tristate
rlabel metal2 s 1674 0 1730 480 6 data_in
port 51 nsew default input
rlabel metal2 s 570 0 626 480 6 enable
port 52 nsew default input
rlabel metal3 s 0 21360 480 21480 6 top_grid_pin_14_
port 53 nsew default tristate
rlabel metal3 s 21520 20952 22000 21072 6 top_grid_pin_2_
port 54 nsew default tristate
rlabel metal3 s 0 20272 480 20392 6 top_grid_pin_6_
port 55 nsew default tristate
rlabel metal4 s 4611 2128 4931 19632 6 vpwr
port 56 nsew default input
rlabel metal4 s 8277 2128 8597 19632 6 vgnd
port 57 nsew default input
<< end >>
